module layer_10_featuremap_16(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd31603),
	.w1(32'h3ccb62fa),
	.w2(32'hbc8ecbfb),
	.w3(32'h3cb2d5cc),
	.w4(32'h3cbdccca),
	.w5(32'h3bf2564d),
	.w6(32'h3c3139fe),
	.w7(32'h3c864c80),
	.w8(32'h3c62e410),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc456836),
	.w1(32'hbc4bdf13),
	.w2(32'hb8bbe9d9),
	.w3(32'hbc845e13),
	.w4(32'hbc17b134),
	.w5(32'h3a7c18c8),
	.w6(32'hbbaf113f),
	.w7(32'hbc2156aa),
	.w8(32'hb8f28994),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd395b),
	.w1(32'hbc7dbcf3),
	.w2(32'h3b3eccf8),
	.w3(32'hb9ad436b),
	.w4(32'hbc359324),
	.w5(32'hb959eb3c),
	.w6(32'hbbe2750c),
	.w7(32'hbc56e582),
	.w8(32'hbad526bb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fbe16),
	.w1(32'h3b88215d),
	.w2(32'hbad076a6),
	.w3(32'h3bf7aab2),
	.w4(32'h3c1afbee),
	.w5(32'hbc3b8aa3),
	.w6(32'hb9e63098),
	.w7(32'hbac0b106),
	.w8(32'hbbd5b39c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33f071),
	.w1(32'h3c702c3b),
	.w2(32'h3ac92f6d),
	.w3(32'hbc25c01f),
	.w4(32'h38fbb269),
	.w5(32'hba866528),
	.w6(32'hbc02c768),
	.w7(32'hbb0a7933),
	.w8(32'hbb7598bc),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf2b65),
	.w1(32'h3b0ceac5),
	.w2(32'h3ba711e0),
	.w3(32'hbb06c718),
	.w4(32'hbc31aa2a),
	.w5(32'h3a88a2b3),
	.w6(32'hbbac49d3),
	.w7(32'h3b6f22fb),
	.w8(32'hbb27fe9d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39daf57d),
	.w1(32'hba32b6e8),
	.w2(32'hbc017fae),
	.w3(32'hbc00a4fe),
	.w4(32'hbbce6a55),
	.w5(32'hbc99f6b8),
	.w6(32'hbc077d34),
	.w7(32'hbb9ea40c),
	.w8(32'hbc19cf5a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa7a72),
	.w1(32'hbba7399e),
	.w2(32'hbc8b3fe1),
	.w3(32'hbc139cc9),
	.w4(32'hbbb633cd),
	.w5(32'hbc96f8df),
	.w6(32'hba85fada),
	.w7(32'h3a96d190),
	.w8(32'hbc35632e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc134d6b),
	.w1(32'hba96c278),
	.w2(32'h3c04fee3),
	.w3(32'hbcc8b103),
	.w4(32'hbc75b99e),
	.w5(32'h3b5e5e11),
	.w6(32'hbca37cc0),
	.w7(32'hbc9d6847),
	.w8(32'h3c7cd9bd),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0091a3),
	.w1(32'hba4452e2),
	.w2(32'h3baf1c15),
	.w3(32'hbaf7d4a4),
	.w4(32'hbb955e8c),
	.w5(32'h3b9335a0),
	.w6(32'hb73731ae),
	.w7(32'hbb5db040),
	.w8(32'hbabc6362),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95aa082),
	.w1(32'hbb270cfa),
	.w2(32'hb96d97cf),
	.w3(32'h3b187776),
	.w4(32'hbb0bbd0b),
	.w5(32'h3aae56bc),
	.w6(32'h3bf806c5),
	.w7(32'h3b8727c2),
	.w8(32'hbbcb4f10),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd09a5c),
	.w1(32'h3ba42d2c),
	.w2(32'h3afdf017),
	.w3(32'h3c7b8f4a),
	.w4(32'h3bb49e7f),
	.w5(32'hbbe2c6c9),
	.w6(32'hbbaffe2a),
	.w7(32'hbb7df2eb),
	.w8(32'hbbcae3b2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c12b3),
	.w1(32'h3b505e44),
	.w2(32'h3c0af2e2),
	.w3(32'hbbb543a7),
	.w4(32'hbb808b11),
	.w5(32'h3c07dbc7),
	.w6(32'hbc40f007),
	.w7(32'hbc07be0c),
	.w8(32'h3aa1dcaf),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c353a14),
	.w1(32'hbba988a9),
	.w2(32'hbbf0f061),
	.w3(32'h3be5e055),
	.w4(32'hbb5a4cbb),
	.w5(32'hbc527d66),
	.w6(32'h3c5938bb),
	.w7(32'hbb1187f8),
	.w8(32'hbb5e62e0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8b895),
	.w1(32'h3b4ff16b),
	.w2(32'hbb7ce2ab),
	.w3(32'hbc7316e7),
	.w4(32'hbb886b21),
	.w5(32'h3b5918b7),
	.w6(32'hbc293c0e),
	.w7(32'hbba9d58d),
	.w8(32'h3b8d9dfa),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3782e5),
	.w1(32'hbc2194d3),
	.w2(32'h3b976f39),
	.w3(32'h3a866ddb),
	.w4(32'hba046e56),
	.w5(32'h3bbb5296),
	.w6(32'h3b98f36d),
	.w7(32'h3b1fe1c7),
	.w8(32'h38cbfd31),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadba58b),
	.w1(32'hbb8ed1b0),
	.w2(32'hbb594008),
	.w3(32'h3af2f027),
	.w4(32'hbb82b1cd),
	.w5(32'h3b5b04ff),
	.w6(32'h3be647d4),
	.w7(32'h3a60ba4b),
	.w8(32'h3c040c1e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7092ea),
	.w1(32'hbbc1b996),
	.w2(32'h39acabc6),
	.w3(32'hbc1c9ff3),
	.w4(32'hbc822ae8),
	.w5(32'hbbcd94bd),
	.w6(32'hbb0fe06b),
	.w7(32'hbc51a784),
	.w8(32'hbc263250),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a5248),
	.w1(32'h3ba69157),
	.w2(32'h3c0ff47e),
	.w3(32'h3c0254b8),
	.w4(32'h3ad27875),
	.w5(32'hbbbd1132),
	.w6(32'hbb777702),
	.w7(32'hbb97ac56),
	.w8(32'hbc612522),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c451429),
	.w1(32'hbb8766b3),
	.w2(32'h3bd45947),
	.w3(32'h3c710638),
	.w4(32'h3b0603c2),
	.w5(32'h3bcd3d47),
	.w6(32'hbc1fdd12),
	.w7(32'h3b2390c1),
	.w8(32'h3a8a0825),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ffba1),
	.w1(32'h3b8f655f),
	.w2(32'h3b191ee3),
	.w3(32'h3c112d7f),
	.w4(32'h3b87e925),
	.w5(32'hba1dce8f),
	.w6(32'hbabfc758),
	.w7(32'hbb389aa1),
	.w8(32'h3a4b00cc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a9177),
	.w1(32'h3c29bb57),
	.w2(32'h3c4551ad),
	.w3(32'h3b391575),
	.w4(32'h3c02aea0),
	.w5(32'h3c3a80cf),
	.w6(32'h3b1c5178),
	.w7(32'hbb14a208),
	.w8(32'hbb550d04),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc01723),
	.w1(32'h3c9505c0),
	.w2(32'h3b25e6d8),
	.w3(32'h3d003352),
	.w4(32'h3cd4ff9e),
	.w5(32'hbc2c3132),
	.w6(32'hbc2d7ae6),
	.w7(32'hbc5fcc64),
	.w8(32'hbcd12420),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd25b4),
	.w1(32'h3bebfef0),
	.w2(32'h3b81b7fb),
	.w3(32'hbb98a059),
	.w4(32'hbb8f9197),
	.w5(32'h3ba8d355),
	.w6(32'hbc3011cf),
	.w7(32'hbc19057c),
	.w8(32'h3a23f404),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf523e),
	.w1(32'h3b3fb8dd),
	.w2(32'hba8f0df6),
	.w3(32'h3bba6ed6),
	.w4(32'h3b962308),
	.w5(32'h3b632ef5),
	.w6(32'hbb0c6804),
	.w7(32'hbb9af6c1),
	.w8(32'hbc6b773b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07041b),
	.w1(32'h3c086702),
	.w2(32'h3bc009ec),
	.w3(32'h3bf879d0),
	.w4(32'h3bd019cf),
	.w5(32'h3b62b144),
	.w6(32'hbc073923),
	.w7(32'hbc026cfb),
	.w8(32'hb9237ac7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c486493),
	.w1(32'h3c984e37),
	.w2(32'h39881e6c),
	.w3(32'h3c8551d4),
	.w4(32'h3cc8fa78),
	.w5(32'hba9787f6),
	.w6(32'h38bc10ca),
	.w7(32'h3c2ca19b),
	.w8(32'h3a49f8dc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c977951),
	.w1(32'hbb02a06b),
	.w2(32'h3bbaca01),
	.w3(32'h3c82c312),
	.w4(32'hbbd2e618),
	.w5(32'hbb7e74ba),
	.w6(32'h3cd1bc09),
	.w7(32'hbafd0500),
	.w8(32'hbb157af9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb650892),
	.w1(32'hba9399da),
	.w2(32'hba56f749),
	.w3(32'hbc249c2f),
	.w4(32'hbbc92ab8),
	.w5(32'h3805db7b),
	.w6(32'hbbdb7611),
	.w7(32'hbb9ad186),
	.w8(32'h3b8a3d97),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfac630),
	.w1(32'hbb9391f8),
	.w2(32'h3b67f472),
	.w3(32'h3c8e6eb7),
	.w4(32'hbab346a2),
	.w5(32'h3b4a96fe),
	.w6(32'h3bb0d20b),
	.w7(32'hbb872f57),
	.w8(32'h382be181),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae383a4),
	.w1(32'hbac6c2ff),
	.w2(32'hbaa2e51a),
	.w3(32'hba6f42e9),
	.w4(32'hbb4d8318),
	.w5(32'h3c691dde),
	.w6(32'h3b503d5e),
	.w7(32'hb9a16a60),
	.w8(32'hbbde05de),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc560d1),
	.w1(32'hbad96d3a),
	.w2(32'h3a42b398),
	.w3(32'h3cbb8d10),
	.w4(32'h3c3e0fb5),
	.w5(32'h3c82070c),
	.w6(32'hba828ea9),
	.w7(32'hba7e5dfb),
	.w8(32'h3bc0e946),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf8ada),
	.w1(32'hbb9967cf),
	.w2(32'hbb4c53de),
	.w3(32'h3caa2ecf),
	.w4(32'h3b933dae),
	.w5(32'hbb63f19f),
	.w6(32'h3baebf5a),
	.w7(32'h3b925357),
	.w8(32'hba3b1c1d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c6ea0),
	.w1(32'hbbcb2e1e),
	.w2(32'h3c3a46bd),
	.w3(32'hbbac21d2),
	.w4(32'hbb7ded81),
	.w5(32'h3afdd109),
	.w6(32'hba7ab0af),
	.w7(32'hbb06279c),
	.w8(32'hbbc5fa6c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a92c6),
	.w1(32'hb8b3ab65),
	.w2(32'hbb0fe494),
	.w3(32'h3b4428f2),
	.w4(32'hbc1616ed),
	.w5(32'hbb20bbce),
	.w6(32'hba805ff5),
	.w7(32'hbb2f1551),
	.w8(32'hba8e1ab5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b125c73),
	.w1(32'h38f3e7e1),
	.w2(32'hbbc06fd7),
	.w3(32'h3b46bee6),
	.w4(32'h3b289fb1),
	.w5(32'hbc1545ed),
	.w6(32'hbb7f9541),
	.w7(32'h3ac5bba6),
	.w8(32'h3ac079a2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc78d9b),
	.w1(32'hbc17b8aa),
	.w2(32'hbca063c4),
	.w3(32'h3c170170),
	.w4(32'h3b597007),
	.w5(32'hbae2db3d),
	.w6(32'hbc1765b1),
	.w7(32'h3bdd9025),
	.w8(32'hbb4372f5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea9727),
	.w1(32'hbbaec9a6),
	.w2(32'hbc329bce),
	.w3(32'h38caa30a),
	.w4(32'hbba7fe61),
	.w5(32'hbc1faa1e),
	.w6(32'h3b9687af),
	.w7(32'hbc1224aa),
	.w8(32'hbb20df8e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca52ed6),
	.w1(32'h395d85c8),
	.w2(32'hbc10a8b3),
	.w3(32'h3b934898),
	.w4(32'hbc55533d),
	.w5(32'hbc93b03b),
	.w6(32'h3cba762e),
	.w7(32'h3975c74b),
	.w8(32'hbc92c34e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bf1ad),
	.w1(32'h3c3f3439),
	.w2(32'hbaf80fc7),
	.w3(32'hbc306c42),
	.w4(32'h3ae13421),
	.w5(32'hbb18acfe),
	.w6(32'hbc3205fa),
	.w7(32'hbbf63f88),
	.w8(32'hbb06aafd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dbba4),
	.w1(32'hbb132907),
	.w2(32'h3ba7d3ad),
	.w3(32'hbb342e4b),
	.w4(32'hbb7075a3),
	.w5(32'h3b3e497e),
	.w6(32'hbb4dbfcf),
	.w7(32'hbbbf92ff),
	.w8(32'h3c1493d3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3dd88),
	.w1(32'h3bc6cc1b),
	.w2(32'h39a27120),
	.w3(32'hbac596b8),
	.w4(32'hba755974),
	.w5(32'hbb3bf49c),
	.w6(32'h3b94195a),
	.w7(32'h3bce2a07),
	.w8(32'h3bb7ef11),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cef50),
	.w1(32'hbb8d989e),
	.w2(32'hbb3b3038),
	.w3(32'h3bae400d),
	.w4(32'hbb418773),
	.w5(32'h3950f444),
	.w6(32'h3b6178e8),
	.w7(32'h3952c36f),
	.w8(32'hbac29c53),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba092f6),
	.w1(32'hba9af20b),
	.w2(32'hbb367736),
	.w3(32'h3bde8268),
	.w4(32'h3bd1caa4),
	.w5(32'hbb227741),
	.w6(32'hbb14522b),
	.w7(32'h3912a66a),
	.w8(32'hbc8369ac),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9adbbd),
	.w1(32'h3b4bafa2),
	.w2(32'h3a58d41f),
	.w3(32'hbc021ab9),
	.w4(32'hbbde8932),
	.w5(32'h3ae2bed7),
	.w6(32'hbc3ba705),
	.w7(32'hbc9bbe27),
	.w8(32'hbb04307b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1052d3),
	.w1(32'h3c1240f2),
	.w2(32'h3c35268d),
	.w3(32'hba078e87),
	.w4(32'hbaba8b13),
	.w5(32'h3c1496d2),
	.w6(32'hbc89eb20),
	.w7(32'hbc56e2d0),
	.w8(32'hbc271ac1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ce369),
	.w1(32'h3b8be538),
	.w2(32'h3ab3abbf),
	.w3(32'hba899b48),
	.w4(32'h3aa84e74),
	.w5(32'hbbca0f1a),
	.w6(32'hbc0b26ee),
	.w7(32'hbc10827b),
	.w8(32'hbcb2896d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb300f),
	.w1(32'hbb12576c),
	.w2(32'hba9e102e),
	.w3(32'hbc242f58),
	.w4(32'hbc3bc461),
	.w5(32'hbc16265d),
	.w6(32'hbd003cc5),
	.w7(32'hbc7d2907),
	.w8(32'hbc8713da),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31cd1b),
	.w1(32'h3a209ac4),
	.w2(32'hb91f36a5),
	.w3(32'h3b071c9e),
	.w4(32'h3b737f5c),
	.w5(32'hbab68243),
	.w6(32'hbb7fd362),
	.w7(32'hb9286a71),
	.w8(32'h3b4914b4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba291de5),
	.w1(32'hbbaa9a9d),
	.w2(32'h3bddb8c9),
	.w3(32'hbbb2f4af),
	.w4(32'h3b9a6091),
	.w5(32'h3be971d9),
	.w6(32'hbab5e878),
	.w7(32'h3b92e599),
	.w8(32'h3b408dff),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83cdff),
	.w1(32'h3aa1ce48),
	.w2(32'hbb1aedb4),
	.w3(32'hbafab0b1),
	.w4(32'h3ba85de3),
	.w5(32'hbaa29934),
	.w6(32'h3b85d928),
	.w7(32'hbb0abab7),
	.w8(32'hbc2e4239),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71bff1),
	.w1(32'h3c529b22),
	.w2(32'h3bda121f),
	.w3(32'h3b872d30),
	.w4(32'hbaa70abf),
	.w5(32'h3b9d9d38),
	.w6(32'hbc2ae8b1),
	.w7(32'hbc93746d),
	.w8(32'hbb11ef56),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5f3e5),
	.w1(32'hba7e400a),
	.w2(32'h3bcef8e3),
	.w3(32'hbb863ccc),
	.w4(32'h3a2c49a3),
	.w5(32'h3c28e911),
	.w6(32'h3b7e24b1),
	.w7(32'hb9e45b52),
	.w8(32'hbbce226c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33e184),
	.w1(32'h3bdeb2db),
	.w2(32'h3bf053ae),
	.w3(32'h3c8cf591),
	.w4(32'h3c437af4),
	.w5(32'h3ad5780a),
	.w6(32'hbc013f79),
	.w7(32'hbb90eda0),
	.w8(32'hbb16f9fa),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c198342),
	.w1(32'h3c23a121),
	.w2(32'h396318c0),
	.w3(32'h3b72dcae),
	.w4(32'h3bc4f1a7),
	.w5(32'hbba39b8d),
	.w6(32'h3ba84edd),
	.w7(32'hb885c103),
	.w8(32'hbc44b2ed),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae984c4),
	.w1(32'h3ad07bb5),
	.w2(32'hba8e9d08),
	.w3(32'h3b27dc1a),
	.w4(32'h3bffa70e),
	.w5(32'h3a8b3854),
	.w6(32'hbc2610b9),
	.w7(32'hbc4c9289),
	.w8(32'hbc186cfc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc528b75),
	.w1(32'hbc455c6a),
	.w2(32'hbb76cf00),
	.w3(32'hbbd3bcc2),
	.w4(32'hbb58108a),
	.w5(32'hbc04216e),
	.w6(32'hbc09ee11),
	.w7(32'hbaeaacc2),
	.w8(32'hbb439c4e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadffd0),
	.w1(32'hbb0297be),
	.w2(32'hbb2d4362),
	.w3(32'hbbd92cf8),
	.w4(32'hbbc9eb9f),
	.w5(32'hba687374),
	.w6(32'hbb6cec2e),
	.w7(32'hbb08aa8e),
	.w8(32'hbad80823),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb380db9),
	.w1(32'h39c1c377),
	.w2(32'h3a8bcd60),
	.w3(32'h3b08bce6),
	.w4(32'h3b4483a0),
	.w5(32'hbc21addc),
	.w6(32'h3b4f09a9),
	.w7(32'h3b1fc06f),
	.w8(32'h3be38908),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd01504),
	.w1(32'h3ba14965),
	.w2(32'h3bcda700),
	.w3(32'hbbeb1210),
	.w4(32'hbbf8e081),
	.w5(32'h3a3d5871),
	.w6(32'h3bd766f8),
	.w7(32'h3bc992ca),
	.w8(32'h399f7b9d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4088a),
	.w1(32'h3b97a24a),
	.w2(32'h3a900adb),
	.w3(32'h3b6a1515),
	.w4(32'hbafbfbdb),
	.w5(32'hbbadef96),
	.w6(32'h3b001dd2),
	.w7(32'h3b7cfc0f),
	.w8(32'hbbcd0de7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba089d71),
	.w1(32'hbb17f16a),
	.w2(32'h3bb0a2fe),
	.w3(32'hba6d0c94),
	.w4(32'h3a7ac848),
	.w5(32'hbb4412af),
	.w6(32'h3bdd7cf7),
	.w7(32'hb7d5b95c),
	.w8(32'hbbad6d57),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc79124),
	.w1(32'h3950dbe8),
	.w2(32'h3b05d1d8),
	.w3(32'hbafe18c3),
	.w4(32'hbbd5ccdc),
	.w5(32'hbad21eea),
	.w6(32'hb88128c6),
	.w7(32'hbb5be15a),
	.w8(32'hbacedcb7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac9cad),
	.w1(32'h3b1a84f7),
	.w2(32'hbb81aaf7),
	.w3(32'hbb0f975f),
	.w4(32'hba9c5b67),
	.w5(32'hbc33915a),
	.w6(32'hba8427e2),
	.w7(32'h39937d95),
	.w8(32'hbba684cf),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb330b34),
	.w1(32'hbb2b2694),
	.w2(32'h3af9c73c),
	.w3(32'h3a0b06ea),
	.w4(32'hbb7fcb61),
	.w5(32'h3c1944fa),
	.w6(32'hbb4da940),
	.w7(32'hbb4b1531),
	.w8(32'h3b6ccdf6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf160bb),
	.w1(32'hb9dc27b6),
	.w2(32'hbb2353b9),
	.w3(32'h3bc30db1),
	.w4(32'h3b68568d),
	.w5(32'h39cc135f),
	.w6(32'h3a58ef89),
	.w7(32'h39dc1d25),
	.w8(32'h3b21b2c5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b40dc),
	.w1(32'hbc1136a7),
	.w2(32'h3b918f70),
	.w3(32'h3b7f7814),
	.w4(32'h3b26b57d),
	.w5(32'h3ae0944c),
	.w6(32'h3bbe4ad2),
	.w7(32'h3a614903),
	.w8(32'hbbe571a5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb381f9),
	.w1(32'h3abf784a),
	.w2(32'h3b0f1dd2),
	.w3(32'hbadbb7e1),
	.w4(32'hbb4fc168),
	.w5(32'hbb38d998),
	.w6(32'hbc6d328d),
	.w7(32'hbc26b786),
	.w8(32'hbc15ea37),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a4e29),
	.w1(32'h39f31c66),
	.w2(32'hbb03e956),
	.w3(32'hbc01f240),
	.w4(32'hbb59cb82),
	.w5(32'hbbc10fa8),
	.w6(32'hbc363a1c),
	.w7(32'hbc25ff2d),
	.w8(32'hbc317b3b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34d117),
	.w1(32'h3b97484f),
	.w2(32'h3a7a6c9c),
	.w3(32'h3a315f7e),
	.w4(32'h3a018ddb),
	.w5(32'hba57756d),
	.w6(32'hbbed54e1),
	.w7(32'hbc545f08),
	.w8(32'hbc8ef14f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb647e7b),
	.w1(32'h3b9d9eea),
	.w2(32'hbb0264d7),
	.w3(32'hbbe103df),
	.w4(32'hbb46e2f9),
	.w5(32'h3b29cba4),
	.w6(32'hbbc5367b),
	.w7(32'hbbf6136d),
	.w8(32'hbbb9d228),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac29e4c),
	.w1(32'h3a99f1a3),
	.w2(32'h3bebb58b),
	.w3(32'h3b9cb8a2),
	.w4(32'h3bf68277),
	.w5(32'hbb6832dc),
	.w6(32'hbc257025),
	.w7(32'hbb57f51e),
	.w8(32'hbbce46eb),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb929ab9),
	.w1(32'hbb11054a),
	.w2(32'hbb7881c3),
	.w3(32'hb9aac31b),
	.w4(32'hbb9b7f08),
	.w5(32'hbacfa8bc),
	.w6(32'h3b0ed0a4),
	.w7(32'hbad9e100),
	.w8(32'h3c02713b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf15fbb),
	.w1(32'h3ad24afc),
	.w2(32'hbbc29cf7),
	.w3(32'h3bdf310b),
	.w4(32'hb7b193de),
	.w5(32'hbbdbdc09),
	.w6(32'h3c41de80),
	.w7(32'h3be04cde),
	.w8(32'hbc063dcd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa84136),
	.w1(32'hbbc74cf1),
	.w2(32'hbb4ef064),
	.w3(32'hba9c0e71),
	.w4(32'hbaf86cc8),
	.w5(32'hbb2e35d7),
	.w6(32'hbba05278),
	.w7(32'hbb8cf39b),
	.w8(32'hbac3f496),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c8856),
	.w1(32'hbb52b374),
	.w2(32'hbbd592bd),
	.w3(32'hbb6514f2),
	.w4(32'hbbc0b1e8),
	.w5(32'hbbc78fcc),
	.w6(32'h372b8448),
	.w7(32'hba2cf9bb),
	.w8(32'hbacf7e45),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc028df4),
	.w1(32'hbbb48558),
	.w2(32'hbc07e1f0),
	.w3(32'hbc25538b),
	.w4(32'hba65713d),
	.w5(32'hbc1f7de5),
	.w6(32'hbc790cdb),
	.w7(32'hbb5dbc72),
	.w8(32'hbc5c0555),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d2e89),
	.w1(32'h3b816eaf),
	.w2(32'h3c2287a4),
	.w3(32'h3b60ebe2),
	.w4(32'h3c1b1f8e),
	.w5(32'h3aaf598e),
	.w6(32'hbc057faa),
	.w7(32'hbb8996c4),
	.w8(32'hbbd6b031),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39774571),
	.w1(32'hbb7d253e),
	.w2(32'h3aa18ea4),
	.w3(32'hbb80debe),
	.w4(32'hbaef47e9),
	.w5(32'hba82fe0f),
	.w6(32'hbc49d6c8),
	.w7(32'hbc51d656),
	.w8(32'hbac609c1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0bc89),
	.w1(32'hbaa4e293),
	.w2(32'hbb81167f),
	.w3(32'h3a43dc07),
	.w4(32'hbb40280d),
	.w5(32'hba749f7c),
	.w6(32'hbb0dca59),
	.w7(32'h3a122359),
	.w8(32'hbc0218c3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4601bc),
	.w1(32'h3a17a56b),
	.w2(32'hbb3dee71),
	.w3(32'hbac55d0c),
	.w4(32'h38abcb61),
	.w5(32'hbad14576),
	.w6(32'hbc01dc9b),
	.w7(32'hbbfa9f8a),
	.w8(32'hba5b2507),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba36bff),
	.w1(32'hbb813687),
	.w2(32'h3ad43b97),
	.w3(32'hbb318554),
	.w4(32'hbbc0ff89),
	.w5(32'hb934e65b),
	.w6(32'hb9dd9f65),
	.w7(32'hbb03e57c),
	.w8(32'hbbd2088d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc024ae8),
	.w1(32'hbc1cc6ad),
	.w2(32'hbaf5cc28),
	.w3(32'hbbec8604),
	.w4(32'hbc2001d1),
	.w5(32'hbbbaf269),
	.w6(32'hbba3fd70),
	.w7(32'hbb9ad88b),
	.w8(32'h3a0a0632),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab84ca),
	.w1(32'h3bc618b7),
	.w2(32'h3b945bf7),
	.w3(32'hbb871771),
	.w4(32'hbb625a03),
	.w5(32'h3b760b3d),
	.w6(32'hbbf7cb84),
	.w7(32'hbc164faf),
	.w8(32'h3a0b2718),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb664a64),
	.w1(32'h3c01b1b5),
	.w2(32'hbc08a552),
	.w3(32'hba021273),
	.w4(32'h3bfff60e),
	.w5(32'hbc1f28e2),
	.w6(32'h3b52839d),
	.w7(32'hbb8085a0),
	.w8(32'hbc19ef3d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9192a2),
	.w1(32'h3b6a5ade),
	.w2(32'h375ec9d7),
	.w3(32'hbc688e04),
	.w4(32'hbb8606fa),
	.w5(32'h3b5adf6c),
	.w6(32'hbc75bf31),
	.w7(32'hbc6f0807),
	.w8(32'hb8ad5aa4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69c6f0),
	.w1(32'h3b3fb7f0),
	.w2(32'h3a53cd27),
	.w3(32'hbad4ee21),
	.w4(32'hb921ff78),
	.w5(32'h3b017605),
	.w6(32'hbbe702c4),
	.w7(32'hbc124cc7),
	.w8(32'hbb00a664),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a230efd),
	.w1(32'h39838745),
	.w2(32'h3ba5cc82),
	.w3(32'h3b3f0016),
	.w4(32'h3a393922),
	.w5(32'h3b0293fe),
	.w6(32'h3b5e63c0),
	.w7(32'h3ab0587e),
	.w8(32'h3b104338),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16b326),
	.w1(32'h3baccdbc),
	.w2(32'hbbb08dfc),
	.w3(32'h3b46d282),
	.w4(32'h3c2c435c),
	.w5(32'hbb988703),
	.w6(32'hbc1ef25a),
	.w7(32'hbbdb613f),
	.w8(32'hba146222),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d181f),
	.w1(32'hbaa8214d),
	.w2(32'hbb74ce5f),
	.w3(32'hbbb03346),
	.w4(32'h3a945303),
	.w5(32'h3adc4481),
	.w6(32'hbc1992ba),
	.w7(32'hbc04db37),
	.w8(32'hbbb76815),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b385d1a),
	.w1(32'hbc1e2a10),
	.w2(32'h3b78c08c),
	.w3(32'h3c781d10),
	.w4(32'h3bcad64c),
	.w5(32'hbac8495d),
	.w6(32'h3c2c235d),
	.w7(32'h3b874948),
	.w8(32'hbbda6e53),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9b539),
	.w1(32'h3bc9893c),
	.w2(32'hbbfa0927),
	.w3(32'h3bb7f036),
	.w4(32'h3bb5bf6b),
	.w5(32'h3b8bf123),
	.w6(32'hbc17306c),
	.w7(32'hbb1c4089),
	.w8(32'hbba16ca8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb693306),
	.w1(32'hbbc11c53),
	.w2(32'h3afd310e),
	.w3(32'hb9c6a8ef),
	.w4(32'hbaef2f2c),
	.w5(32'hbae685d0),
	.w6(32'hbb76ff5e),
	.w7(32'hbb820d60),
	.w8(32'hbbd12f40),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12cb10),
	.w1(32'hbb202561),
	.w2(32'hbb850152),
	.w3(32'hbb60c2fd),
	.w4(32'hbb25cd68),
	.w5(32'hbae7ac51),
	.w6(32'hbc1a6908),
	.w7(32'hbbd1db2b),
	.w8(32'hbc05715a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddeab9),
	.w1(32'hbb4681d5),
	.w2(32'hb927a7f8),
	.w3(32'hbb2caac3),
	.w4(32'h3a7dba23),
	.w5(32'h3b79f6f8),
	.w6(32'hbab45074),
	.w7(32'hbb77cb88),
	.w8(32'hbb85da0a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b400319),
	.w1(32'hbb91d830),
	.w2(32'hbb4c913e),
	.w3(32'h3b62d7e0),
	.w4(32'h3aa56a06),
	.w5(32'h3a75df49),
	.w6(32'h3be49b42),
	.w7(32'hbb32229f),
	.w8(32'hbb9cf09c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14493b),
	.w1(32'hbc04f226),
	.w2(32'hbb80e9f2),
	.w3(32'h3a8f8047),
	.w4(32'h3bc51ebb),
	.w5(32'h3aa3ab9a),
	.w6(32'hba1fb139),
	.w7(32'hbbb333ed),
	.w8(32'h3b4cc364),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba39c50),
	.w1(32'hbaa72e26),
	.w2(32'h3a843dfb),
	.w3(32'hbb356839),
	.w4(32'hbb1dcfd6),
	.w5(32'h3b3e364f),
	.w6(32'hbc0eba1d),
	.w7(32'hbba9ca24),
	.w8(32'hbc221482),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd942c2),
	.w1(32'hbba7f7f3),
	.w2(32'hbc6db91a),
	.w3(32'h3c4496ed),
	.w4(32'hbb0c3e6b),
	.w5(32'hbc2bae47),
	.w6(32'hbbe61b7a),
	.w7(32'hbb7e8fff),
	.w8(32'hbc71aecd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5a20c),
	.w1(32'h3c2839a7),
	.w2(32'hbbf9de3e),
	.w3(32'h3a4ed2c6),
	.w4(32'h3c184774),
	.w5(32'hbbd47138),
	.w6(32'hbc8deef0),
	.w7(32'h3bef77e7),
	.w8(32'hbc0a1308),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0c4a5),
	.w1(32'hbc049195),
	.w2(32'hbbcc3b6a),
	.w3(32'h3c0d6e2b),
	.w4(32'h3b2efe32),
	.w5(32'hbabead07),
	.w6(32'hbb6aaaba),
	.w7(32'hbbcfc83c),
	.w8(32'hbb91e501),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8af7f),
	.w1(32'hbbc573d6),
	.w2(32'hbbde18bc),
	.w3(32'h39d82197),
	.w4(32'hbb831876),
	.w5(32'hbc05aa2d),
	.w6(32'hbc8577cb),
	.w7(32'hbc3daddf),
	.w8(32'hbbc0a252),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3ed26),
	.w1(32'hb9f18254),
	.w2(32'hbb8fad22),
	.w3(32'hbb830f6b),
	.w4(32'hbb680e38),
	.w5(32'h3bc5e139),
	.w6(32'hbb347c60),
	.w7(32'h39b4534e),
	.w8(32'hbc15ce8b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aff9f),
	.w1(32'h39a2d997),
	.w2(32'hb98e21f2),
	.w3(32'h3c36c665),
	.w4(32'h3c1967d5),
	.w5(32'hbb579d75),
	.w6(32'hbb1d64e0),
	.w7(32'hb8f647ad),
	.w8(32'hba50c89a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19bcca),
	.w1(32'hbab7b771),
	.w2(32'hbc598d9d),
	.w3(32'hbc2acdc6),
	.w4(32'hbb9c172e),
	.w5(32'hbc90c397),
	.w6(32'hbc851a43),
	.w7(32'hba70643e),
	.w8(32'hbc3c8244),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fec6b),
	.w1(32'h3b186ed1),
	.w2(32'hbbea29f8),
	.w3(32'hbb5fbef9),
	.w4(32'hbb131af2),
	.w5(32'hbb767de6),
	.w6(32'hbc2341a1),
	.w7(32'hbc3111f2),
	.w8(32'hbbd2ac96),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf727d7),
	.w1(32'hbaa12e82),
	.w2(32'hbb0cea11),
	.w3(32'hbb9fcbef),
	.w4(32'hba337aac),
	.w5(32'hbc250a4e),
	.w6(32'hbc0f48b2),
	.w7(32'hbbc8f060),
	.w8(32'hbaa5a34a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02df0c),
	.w1(32'h3c109044),
	.w2(32'hbb808e79),
	.w3(32'hbbf90503),
	.w4(32'hbaadf496),
	.w5(32'hbb32d716),
	.w6(32'hbb14cc07),
	.w7(32'h3a3241e2),
	.w8(32'hbc02cbf8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b060225),
	.w1(32'h3bc7bb2e),
	.w2(32'h38d5c554),
	.w3(32'h3bacc06e),
	.w4(32'h3c2ac44a),
	.w5(32'h3aa38678),
	.w6(32'hbc3ce14c),
	.w7(32'hbbec6482),
	.w8(32'hbb69b8d5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b877478),
	.w1(32'hbb9b7401),
	.w2(32'hbac7d4f6),
	.w3(32'h3c12ac73),
	.w4(32'h3bb3e072),
	.w5(32'hbb526d34),
	.w6(32'hbbb4cfa4),
	.w7(32'hbab539c4),
	.w8(32'hb8cf7a4b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45d484),
	.w1(32'hbb8a4411),
	.w2(32'h3bc6a328),
	.w3(32'hbb067ee7),
	.w4(32'hbc2a5311),
	.w5(32'h3b92286d),
	.w6(32'h3b85ae0f),
	.w7(32'hbb4539a9),
	.w8(32'hbbadc3ef),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f7ab6),
	.w1(32'h3bc98f8f),
	.w2(32'h38ab2b87),
	.w3(32'h3aa2146f),
	.w4(32'h3b3ff986),
	.w5(32'hbaad0af7),
	.w6(32'h3a57a5ad),
	.w7(32'hbbcbe6ff),
	.w8(32'hbba59c9a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b237a),
	.w1(32'h3bafa07c),
	.w2(32'hb94b487c),
	.w3(32'hbb9e1dec),
	.w4(32'h39a913eb),
	.w5(32'hba593323),
	.w6(32'hbc7e294c),
	.w7(32'hbc5b08a1),
	.w8(32'hbac2fd2f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26e227),
	.w1(32'hbbc7f40f),
	.w2(32'h3bf0764c),
	.w3(32'h3b0f60ca),
	.w4(32'hbacfc7dc),
	.w5(32'hbbb5fcf0),
	.w6(32'hbb564b62),
	.w7(32'hbb840e9c),
	.w8(32'hbbbaadbe),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f5494),
	.w1(32'h3ba605e1),
	.w2(32'hb9ae7e65),
	.w3(32'hbbb3d912),
	.w4(32'hbb87a990),
	.w5(32'hbbd32808),
	.w6(32'hbc05b92a),
	.w7(32'hbc08c4d5),
	.w8(32'hbb35cfd8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a757107),
	.w1(32'h3b9721e5),
	.w2(32'h3b9a85ee),
	.w3(32'hbbdf01ed),
	.w4(32'hbbd0ad44),
	.w5(32'h3c482762),
	.w6(32'hbadec27c),
	.w7(32'hbaa0c6bf),
	.w8(32'hbc2d7990),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03b723),
	.w1(32'h3ba11e49),
	.w2(32'hbbaa9ab9),
	.w3(32'h3caaf69b),
	.w4(32'h3c72ae2e),
	.w5(32'hbc0a4f7c),
	.w6(32'hbc1e06f7),
	.w7(32'hbbd9b5df),
	.w8(32'h3a4ca162),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb779c56),
	.w1(32'hbb33c0ab),
	.w2(32'hbb70268c),
	.w3(32'hbbfb544f),
	.w4(32'hbc124138),
	.w5(32'hbb8ec75b),
	.w6(32'hb917cd01),
	.w7(32'hbb08b382),
	.w8(32'h3be4a69b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c3f60),
	.w1(32'h3b463b8d),
	.w2(32'hbc095bbf),
	.w3(32'h3bb9fdd3),
	.w4(32'h3bd0e5d8),
	.w5(32'hbb08fbf3),
	.w6(32'h3b8697ca),
	.w7(32'h3b953c90),
	.w8(32'hbbb8fc22),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66ba58),
	.w1(32'hbbaf7afe),
	.w2(32'hbb8781c1),
	.w3(32'h3ba0c52f),
	.w4(32'h3b640205),
	.w5(32'hbb1c3e99),
	.w6(32'hbbd804c0),
	.w7(32'hbbb20362),
	.w8(32'hbbb28b5b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb935c15),
	.w1(32'hbb7734d8),
	.w2(32'hb9a02b67),
	.w3(32'hbb2db464),
	.w4(32'hbc00bbc6),
	.w5(32'hba571db2),
	.w6(32'hbb6ee6a9),
	.w7(32'hbb202099),
	.w8(32'hb99442ae),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7d725),
	.w1(32'hbaa5f4f4),
	.w2(32'h3a8c93b5),
	.w3(32'h39650535),
	.w4(32'hbac4d3e1),
	.w5(32'h3946cc10),
	.w6(32'hbb321c0f),
	.w7(32'hb9b731a6),
	.w8(32'hb8493e1b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1f914),
	.w1(32'h3b3b28a6),
	.w2(32'h3b5750eb),
	.w3(32'h3ba90a4c),
	.w4(32'h39f8a1d8),
	.w5(32'h3a996cbe),
	.w6(32'h3ba2addc),
	.w7(32'hbb4bd27c),
	.w8(32'hba82dcd0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2ce73),
	.w1(32'hbc06dcbe),
	.w2(32'h3b3f8040),
	.w3(32'h3b8e5905),
	.w4(32'h3a95350a),
	.w5(32'hbb27cc1d),
	.w6(32'hbbc805b2),
	.w7(32'hbc2949b7),
	.w8(32'hb8cd578b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f0beb),
	.w1(32'hb67b2f77),
	.w2(32'h3b0b790a),
	.w3(32'hbc0d105d),
	.w4(32'hbbe7390f),
	.w5(32'h3ab2d2c4),
	.w6(32'hbb9553dd),
	.w7(32'hbb8b79fc),
	.w8(32'hbb4f1224),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8b9df),
	.w1(32'h3c42b9f2),
	.w2(32'h3bf70e3d),
	.w3(32'hba85137e),
	.w4(32'h3bb2ca52),
	.w5(32'h3b5c0748),
	.w6(32'hbc0d269d),
	.w7(32'hbbbf1495),
	.w8(32'hba2fa1f5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c7dc9),
	.w1(32'h3b947996),
	.w2(32'h3b1aefb9),
	.w3(32'hbb9f4f26),
	.w4(32'h3b2da71b),
	.w5(32'h39a7b982),
	.w6(32'hbb044372),
	.w7(32'hbb83e521),
	.w8(32'hbbd47271),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68eadb),
	.w1(32'hbadf7654),
	.w2(32'h3b2831c3),
	.w3(32'hbaa3dae2),
	.w4(32'hbc556903),
	.w5(32'hbb46a8af),
	.w6(32'hbc3fea26),
	.w7(32'hbbdff501),
	.w8(32'hbc095abd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfd217),
	.w1(32'hb9b12d8d),
	.w2(32'hbb130a80),
	.w3(32'hbaf246cf),
	.w4(32'hbc22ded2),
	.w5(32'hbb984475),
	.w6(32'hbb133233),
	.w7(32'hbc0a1415),
	.w8(32'hbc4ac598),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba863c3f),
	.w1(32'h3b0a9daa),
	.w2(32'h3b198de9),
	.w3(32'h3822b957),
	.w4(32'h3c18ac08),
	.w5(32'h3944091f),
	.w6(32'hbb7b6dd8),
	.w7(32'h3a26a01e),
	.w8(32'h3b88a6a3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c638ad4),
	.w1(32'h3b41a78f),
	.w2(32'h3a899984),
	.w3(32'h3ab213fd),
	.w4(32'hbb21adef),
	.w5(32'h39e0f80e),
	.w6(32'hbb4b5196),
	.w7(32'h3b509910),
	.w8(32'h3b12bd5a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a824a),
	.w1(32'hbb0763ba),
	.w2(32'hbc908ab8),
	.w3(32'h3b971728),
	.w4(32'hbbd4f60f),
	.w5(32'hbba3d098),
	.w6(32'hbaae001e),
	.w7(32'h3b2aac5a),
	.w8(32'h39c29095),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63d348),
	.w1(32'hbb810c1f),
	.w2(32'hbc1568ff),
	.w3(32'hbbc99209),
	.w4(32'hbbdee51b),
	.w5(32'hbbd560bb),
	.w6(32'h3b25fb85),
	.w7(32'hbb58a239),
	.w8(32'hbb2d638b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7095ab),
	.w1(32'hba8627a1),
	.w2(32'hbb00c6f6),
	.w3(32'hbb6397b2),
	.w4(32'h39aa803a),
	.w5(32'h3b06da2d),
	.w6(32'hbbcbbb9f),
	.w7(32'hbbdc6e1c),
	.w8(32'hbae8d057),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86b920),
	.w1(32'hbaff4c27),
	.w2(32'hbb0eab06),
	.w3(32'h3bc16cbb),
	.w4(32'hb8a8d9d8),
	.w5(32'hbc27dada),
	.w6(32'hbb0d8ba1),
	.w7(32'hb965ccba),
	.w8(32'hbc1c6dbd),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96e57e),
	.w1(32'h3a91bf13),
	.w2(32'hbb04f847),
	.w3(32'hbbd97bc0),
	.w4(32'hbc2d3d94),
	.w5(32'h3c0ecf8d),
	.w6(32'hbb9c3f04),
	.w7(32'hbb8bf270),
	.w8(32'h3b2c7f3d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad79445),
	.w1(32'h3b8468bf),
	.w2(32'h39d835d5),
	.w3(32'h3c1f35e5),
	.w4(32'h3c3410dd),
	.w5(32'hbb10eafa),
	.w6(32'hbbf45e74),
	.w7(32'hbb73318d),
	.w8(32'hbc3a8696),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e119e),
	.w1(32'hb9a1a609),
	.w2(32'h3afb4dde),
	.w3(32'hbb33f695),
	.w4(32'hbbb69d45),
	.w5(32'hbb15290e),
	.w6(32'hbc3376c5),
	.w7(32'hbc1e0616),
	.w8(32'hbb771a7e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bdf05),
	.w1(32'h3a5c49da),
	.w2(32'h3b81fcaf),
	.w3(32'hbbad30c9),
	.w4(32'hbb74fb92),
	.w5(32'h3bb246d5),
	.w6(32'hbbff2a31),
	.w7(32'hbbcea3b4),
	.w8(32'hbb494253),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06380d),
	.w1(32'hb7f0178e),
	.w2(32'h3a81aaf1),
	.w3(32'h3b3cc96f),
	.w4(32'hbbc421c0),
	.w5(32'hba00b848),
	.w6(32'hbab3410e),
	.w7(32'hbab8808b),
	.w8(32'hbbc1fa31),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c12b7),
	.w1(32'h3ab6ed05),
	.w2(32'hbbc62234),
	.w3(32'h3b3e6cc3),
	.w4(32'h38a5338a),
	.w5(32'hbb0a22cb),
	.w6(32'hbb42567b),
	.w7(32'hbb4388dd),
	.w8(32'hbbd6ac90),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbbb3ca),
	.w1(32'hba34eed3),
	.w2(32'h3c90dd44),
	.w3(32'h3c20ed10),
	.w4(32'hbbfdc196),
	.w5(32'h3be0be09),
	.w6(32'h3c205d16),
	.w7(32'hbc3e93b1),
	.w8(32'hbbf6036d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49009d),
	.w1(32'h3c254a73),
	.w2(32'hbb8b90a4),
	.w3(32'h3befe565),
	.w4(32'h3c1b03c3),
	.w5(32'hbc3e2154),
	.w6(32'hbc3e3724),
	.w7(32'hbc1bc5e0),
	.w8(32'hba853202),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4142),
	.w1(32'h3b055ccf),
	.w2(32'h3a8491ea),
	.w3(32'hbc0f6e86),
	.w4(32'hbb5d20ed),
	.w5(32'hba34b527),
	.w6(32'h3b377841),
	.w7(32'h3bba2ece),
	.w8(32'hba49d0ba),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a4862),
	.w1(32'hbafc05a1),
	.w2(32'h35171694),
	.w3(32'hbb5ad49f),
	.w4(32'hbba9452e),
	.w5(32'h3b55fcbf),
	.w6(32'hbab41194),
	.w7(32'hbb5e4532),
	.w8(32'hb92433f9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50c91d),
	.w1(32'h3ac07c09),
	.w2(32'hbb6881ff),
	.w3(32'h3c0cd4b0),
	.w4(32'h3c0fb95a),
	.w5(32'hbb6215a3),
	.w6(32'hbad1ff64),
	.w7(32'h3bb3406d),
	.w8(32'hbbb3d834),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8718fd),
	.w1(32'h39e087cb),
	.w2(32'h3c484a8b),
	.w3(32'hba15337c),
	.w4(32'h39fbc34a),
	.w5(32'h3c2c4278),
	.w6(32'hbc208272),
	.w7(32'hbbdcbb7c),
	.w8(32'hbc001c09),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d957f),
	.w1(32'h3aeb3bdc),
	.w2(32'h3b15bad3),
	.w3(32'h3c205025),
	.w4(32'h3c093d7a),
	.w5(32'h3b9c026b),
	.w6(32'hbc422649),
	.w7(32'hbbb42f09),
	.w8(32'hbbc545c0),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a581975),
	.w1(32'h3ad33df0),
	.w2(32'h3a9286dd),
	.w3(32'h3bbada33),
	.w4(32'h3b4d1b80),
	.w5(32'hba3f19d1),
	.w6(32'hba9ca975),
	.w7(32'hbb81c998),
	.w8(32'hb8c254e6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6665458),
	.w1(32'h3ab4ab54),
	.w2(32'hbc07aa83),
	.w3(32'h3bace29b),
	.w4(32'h3b615ba2),
	.w5(32'hbb9858c9),
	.w6(32'hbbcaf41e),
	.w7(32'h3a9c0529),
	.w8(32'hbb9418c3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989293),
	.w1(32'h3b59bca5),
	.w2(32'hbaea4c3b),
	.w3(32'hbb790077),
	.w4(32'hbbae0676),
	.w5(32'hb95ebc15),
	.w6(32'hbb9d089c),
	.w7(32'hbb46d0da),
	.w8(32'hbb388c3e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f2ded),
	.w1(32'hbbd320a2),
	.w2(32'hbbaa35b4),
	.w3(32'hbafe2afd),
	.w4(32'hbb56c0b6),
	.w5(32'hbabcd059),
	.w6(32'hbbb98c6b),
	.w7(32'hbb42258e),
	.w8(32'hbbb5de65),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc463b1),
	.w1(32'h39b3b0a9),
	.w2(32'hbb988918),
	.w3(32'h3be62051),
	.w4(32'hbb85f2a3),
	.w5(32'h3aa77a2a),
	.w6(32'h3b36ef06),
	.w7(32'hbc03645c),
	.w8(32'hbc0f398a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb207f8),
	.w1(32'hbbb92f69),
	.w2(32'hbbac5426),
	.w3(32'h3c141635),
	.w4(32'h3a4eff30),
	.w5(32'h38eb72c4),
	.w6(32'h3b810012),
	.w7(32'h3aebc5f5),
	.w8(32'hbbca4e27),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd20086),
	.w1(32'hbb5e3c44),
	.w2(32'hbc1cb849),
	.w3(32'h3aa2f527),
	.w4(32'h3b7a42b7),
	.w5(32'hb9bb3826),
	.w6(32'hbb095c9e),
	.w7(32'hbaf37d64),
	.w8(32'h3b99daf1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ace4d),
	.w1(32'hbb0a7fe5),
	.w2(32'hbac3bb09),
	.w3(32'h3d49f748),
	.w4(32'h3c4d88f7),
	.w5(32'hbaff63e4),
	.w6(32'h3cd6a7bc),
	.w7(32'h3c0291cc),
	.w8(32'hbb6e014d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb587abb),
	.w1(32'hbc5fc9c5),
	.w2(32'h3b187adc),
	.w3(32'h3b6053a6),
	.w4(32'h3adf910c),
	.w5(32'hbbbfaf73),
	.w6(32'h3bb907e3),
	.w7(32'h3919e901),
	.w8(32'hbac41f3c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabef000),
	.w1(32'hbbc647b6),
	.w2(32'hbb69606b),
	.w3(32'h3b5a4f71),
	.w4(32'h3b89b114),
	.w5(32'hbb9fb33b),
	.w6(32'h3b256787),
	.w7(32'h3b2f6723),
	.w8(32'h3c13aca6),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81eb1b),
	.w1(32'h3b9c8f28),
	.w2(32'hba86ab93),
	.w3(32'h3c481ce4),
	.w4(32'h3c8eb7cb),
	.w5(32'h3aead64d),
	.w6(32'h3ccf0225),
	.w7(32'h3ce13b12),
	.w8(32'hbb848206),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02f97a),
	.w1(32'h3b09230e),
	.w2(32'hbb551c15),
	.w3(32'hbb8e9df8),
	.w4(32'h3ad4dd9e),
	.w5(32'hbb16da44),
	.w6(32'hbb2b120f),
	.w7(32'h3b321778),
	.w8(32'hba9ddb1a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05d413),
	.w1(32'hbb877efb),
	.w2(32'h3ced01c9),
	.w3(32'hba8d4db2),
	.w4(32'hbabf65c6),
	.w5(32'h3a4d5af3),
	.w6(32'hbb96c541),
	.w7(32'hbb913b87),
	.w8(32'hbbe6cb6f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7cfa39),
	.w1(32'h3c8eeb1c),
	.w2(32'hbb3c0a4b),
	.w3(32'hbce4cc41),
	.w4(32'hbc80febe),
	.w5(32'h3a3a0164),
	.w6(32'hbd0c7aa1),
	.w7(32'hbc9210e8),
	.w8(32'hbbe57252),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91e3e9),
	.w1(32'hbb8741ed),
	.w2(32'h3c0ccba8),
	.w3(32'hbbf4741a),
	.w4(32'hbbdc207e),
	.w5(32'hbbaf25a3),
	.w6(32'hbbc93134),
	.w7(32'hbbbc3418),
	.w8(32'hbcba746d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccb29b),
	.w1(32'hbb57e381),
	.w2(32'hb8e974e7),
	.w3(32'hbcca0c5b),
	.w4(32'hbca58289),
	.w5(32'hbbc4be6a),
	.w6(32'hbd112d3b),
	.w7(32'hbd0774a5),
	.w8(32'hbbea4e4b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53d9b9),
	.w1(32'h3b08ab7f),
	.w2(32'h3d3e55d5),
	.w3(32'hb8a2d84d),
	.w4(32'h3b8845f1),
	.w5(32'h3b9e69a4),
	.w6(32'hbaea3359),
	.w7(32'h3979253e),
	.w8(32'hbb9dd424),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9956b8),
	.w1(32'h3c9549ea),
	.w2(32'h3a48c9a2),
	.w3(32'hbcd9b4eb),
	.w4(32'hbc885dea),
	.w5(32'hba545fb9),
	.w6(32'hbd18c8e7),
	.w7(32'hbcb5cd3a),
	.w8(32'h3bb12165),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9efcc1),
	.w1(32'h3b307a5f),
	.w2(32'h3a9b3eb6),
	.w3(32'h3af054a7),
	.w4(32'h3bae2cc9),
	.w5(32'hbb8cab3b),
	.w6(32'h3bdd5067),
	.w7(32'h3befe904),
	.w8(32'hbb5d4770),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d4892),
	.w1(32'hbb380681),
	.w2(32'hba398db5),
	.w3(32'hbb3ee575),
	.w4(32'hbbb96459),
	.w5(32'hb9524154),
	.w6(32'hbb6191f1),
	.w7(32'hbbea4ad0),
	.w8(32'hbb9352f3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ceddb9),
	.w1(32'h3a1a76ca),
	.w2(32'hb99c6cb5),
	.w3(32'hb9272669),
	.w4(32'hb9557f38),
	.w5(32'hbaff2fe3),
	.w6(32'hbc4d00ac),
	.w7(32'hbb024cac),
	.w8(32'hbc31a885),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae694f1),
	.w1(32'h3ab615d5),
	.w2(32'hbb4e2014),
	.w3(32'h3b8dad7a),
	.w4(32'h3bdb71ba),
	.w5(32'h3b6121c4),
	.w6(32'hba88b652),
	.w7(32'h3a470fe2),
	.w8(32'h3b88acbe),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba862e0),
	.w1(32'h3ba8a438),
	.w2(32'hbc8816c6),
	.w3(32'h3b38d16e),
	.w4(32'h3a65d3c0),
	.w5(32'h3ca398a5),
	.w6(32'h3b7b6225),
	.w7(32'hb9d7499f),
	.w8(32'h3c9a6282),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc073610),
	.w1(32'hbc5c3c9b),
	.w2(32'hbb037185),
	.w3(32'h3d85d239),
	.w4(32'h3d38adac),
	.w5(32'h3a944bae),
	.w6(32'h3d923689),
	.w7(32'h3d3a7b00),
	.w8(32'h3b9f8352),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4c843),
	.w1(32'hbbd15689),
	.w2(32'h3a847e88),
	.w3(32'hbb18d853),
	.w4(32'hbbb80009),
	.w5(32'hbc03f77e),
	.w6(32'h3b072e89),
	.w7(32'hbbcbba97),
	.w8(32'hbbf32c84),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fc165),
	.w1(32'hbbe4f4a2),
	.w2(32'hbba5df7c),
	.w3(32'h3983e6f9),
	.w4(32'hbbb838a2),
	.w5(32'hbb3f0d43),
	.w6(32'hbb56d007),
	.w7(32'hbbf97e66),
	.w8(32'hbc088d3d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf45a9),
	.w1(32'hbb29b4bc),
	.w2(32'hbba68ac9),
	.w3(32'h3a89f6a4),
	.w4(32'h3b75c47c),
	.w5(32'hbc398109),
	.w6(32'hbbd481c8),
	.w7(32'hbaae604a),
	.w8(32'hbc147a82),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d6c83),
	.w1(32'hbacd6e8f),
	.w2(32'h3c5fa837),
	.w3(32'hbbbb87f5),
	.w4(32'hb9fd977d),
	.w5(32'h3bb64baa),
	.w6(32'hbb91a91f),
	.w7(32'h3ad6ca4b),
	.w8(32'hbc710ca8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60b3b1),
	.w1(32'h3a945820),
	.w2(32'hbb118767),
	.w3(32'hbca7c2b8),
	.w4(32'hbcab8a2a),
	.w5(32'hba5bcbd6),
	.w6(32'hbd2808c9),
	.w7(32'hbd15e078),
	.w8(32'hbc0ede8b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b394276),
	.w1(32'hb9dbfc09),
	.w2(32'hbb2171fe),
	.w3(32'h3a92faf2),
	.w4(32'h3aa7e5d4),
	.w5(32'hbaf2c0dd),
	.w6(32'hbb6b51c2),
	.w7(32'hb89cf059),
	.w8(32'hbb8adbe1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aac8d),
	.w1(32'hbb0155d6),
	.w2(32'h3b8e9c7f),
	.w3(32'h3b182d74),
	.w4(32'h3b895cf4),
	.w5(32'hbae3663d),
	.w6(32'hbbe9ff61),
	.w7(32'hbb9bfe51),
	.w8(32'hbb6958a3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed6490),
	.w1(32'hbb00e7ac),
	.w2(32'hbbac1350),
	.w3(32'h3a9b1377),
	.w4(32'h394bf38c),
	.w5(32'hbbdcffe6),
	.w6(32'h3a8fe0d9),
	.w7(32'hb9d35910),
	.w8(32'h3968f2da),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1250b1),
	.w1(32'h3a44b548),
	.w2(32'hbb0232be),
	.w3(32'h3b26cc98),
	.w4(32'h3b14c759),
	.w5(32'hbae02f14),
	.w6(32'hbb95b18d),
	.w7(32'hbb0127d4),
	.w8(32'hb9414387),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc88d52),
	.w1(32'hbb687802),
	.w2(32'h3abe6c06),
	.w3(32'hbb8d3249),
	.w4(32'hbaa7d950),
	.w5(32'hbc0d178c),
	.w6(32'h3b92e7fa),
	.w7(32'h3bcaedff),
	.w8(32'h3b981ddc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f673e),
	.w1(32'h3be81488),
	.w2(32'hb9704bce),
	.w3(32'h3a1f143d),
	.w4(32'h3bbb8e8f),
	.w5(32'hbb9bc6ce),
	.w6(32'h3b274627),
	.w7(32'h3b5fbd02),
	.w8(32'hbb788224),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b655ec7),
	.w1(32'hb9d05545),
	.w2(32'hbb477f42),
	.w3(32'h3a6eeec4),
	.w4(32'hbb8f259b),
	.w5(32'h3b403cc3),
	.w6(32'hbae9b612),
	.w7(32'hbb75f7f1),
	.w8(32'hbb9fc85a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1e7d3),
	.w1(32'h39c37b06),
	.w2(32'hbb41d3bc),
	.w3(32'hb92e44d8),
	.w4(32'h3b9cc5cd),
	.w5(32'hbb039424),
	.w6(32'hbbe9a36c),
	.w7(32'hbc05cab3),
	.w8(32'hbbcc938a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bbda2),
	.w1(32'hbbd9635d),
	.w2(32'hbc12a155),
	.w3(32'h3b0399a8),
	.w4(32'h3891a6b0),
	.w5(32'hbc12d005),
	.w6(32'hbb330ae1),
	.w7(32'h397f0f6b),
	.w8(32'h3c968779),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc561288),
	.w1(32'hbb057793),
	.w2(32'hba506d10),
	.w3(32'h3c3a0ee6),
	.w4(32'h3c1cca15),
	.w5(32'hbba49ab4),
	.w6(32'h3ce726e6),
	.w7(32'h3d130382),
	.w8(32'hbb777ee3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7af22d),
	.w1(32'hbb833139),
	.w2(32'hbb6ffd19),
	.w3(32'h3b4dcb88),
	.w4(32'h3b5c8163),
	.w5(32'hbbc51155),
	.w6(32'hbc132a89),
	.w7(32'hbb4481dc),
	.w8(32'hbc51d6e6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b108c0b),
	.w1(32'hbc17f21a),
	.w2(32'hbb5c65ff),
	.w3(32'h3c648994),
	.w4(32'h3bcdf9b9),
	.w5(32'hb991e33b),
	.w6(32'h3c48af83),
	.w7(32'hbb2ae518),
	.w8(32'hbbbe34d5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3dfcb),
	.w1(32'hbb424253),
	.w2(32'hba23acc3),
	.w3(32'hbb64de33),
	.w4(32'hbb400095),
	.w5(32'hba04f030),
	.w6(32'h3b7076d5),
	.w7(32'hba006df4),
	.w8(32'h3b0e5ed6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf5a47),
	.w1(32'hbbd787fe),
	.w2(32'h3b1e30ae),
	.w3(32'h3a640a61),
	.w4(32'h3a7fefd3),
	.w5(32'h3b236cd6),
	.w6(32'h3abc7c7c),
	.w7(32'h3a50e134),
	.w8(32'h3b9d0414),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb4ccf),
	.w1(32'h3a588c3d),
	.w2(32'hbb529023),
	.w3(32'h3bf752ef),
	.w4(32'h3baffa29),
	.w5(32'h3ba159a8),
	.w6(32'h3b9f6361),
	.w7(32'h3bc18bf1),
	.w8(32'hbb2d17d6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5818c1),
	.w1(32'h3a740a5a),
	.w2(32'h3aa2e3d9),
	.w3(32'h3b11b7eb),
	.w4(32'h3b92c9a8),
	.w5(32'h3b5ba5aa),
	.w6(32'h3af2ad7e),
	.w7(32'hbb8e4a7d),
	.w8(32'h39b2108a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b129189),
	.w1(32'h3aecb0b5),
	.w2(32'hbd1e7d20),
	.w3(32'h3af4f777),
	.w4(32'h3a141094),
	.w5(32'h3b17698b),
	.w6(32'hb8f79da3),
	.w7(32'h3a153a9f),
	.w8(32'h3d04acc5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce812bf),
	.w1(32'hbcd21f8c),
	.w2(32'hba89510e),
	.w3(32'h3d95bd42),
	.w4(32'h3d588095),
	.w5(32'hb65bab48),
	.w6(32'h3db7e70a),
	.w7(32'h3d8b1f54),
	.w8(32'hbbd788b6),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c0c19),
	.w1(32'h3b556fec),
	.w2(32'h3b3d827d),
	.w3(32'hbb0be009),
	.w4(32'h3ba2cb48),
	.w5(32'hb88e40ea),
	.w6(32'hbbab74d5),
	.w7(32'hb9475f5d),
	.w8(32'hbb45eef8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b574444),
	.w1(32'hb8628851),
	.w2(32'hbbe37528),
	.w3(32'h39b669d8),
	.w4(32'hbb138a5e),
	.w5(32'hba99b651),
	.w6(32'hbb00f592),
	.w7(32'h3ad29866),
	.w8(32'h3a4ccdc4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a140423),
	.w1(32'hbb84faa1),
	.w2(32'h3ada01d9),
	.w3(32'h3c51cf2d),
	.w4(32'h3b99dbc1),
	.w5(32'hbbb2a7b4),
	.w6(32'h3b85bd2f),
	.w7(32'hbae5b342),
	.w8(32'hbc225b4f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd364b),
	.w1(32'hbbfdd5ff),
	.w2(32'hbc1b7cb4),
	.w3(32'hba8dcdd6),
	.w4(32'h3ba9edb2),
	.w5(32'hbb6728a1),
	.w6(32'hbba7b3c4),
	.w7(32'h3bb5d40d),
	.w8(32'h3ad76feb),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf27a31),
	.w1(32'hbbac909e),
	.w2(32'hba70fa81),
	.w3(32'hbaed83f6),
	.w4(32'hbb625e9f),
	.w5(32'hba3db189),
	.w6(32'h3bbbf0a7),
	.w7(32'h3ac01d5c),
	.w8(32'hba9fec6d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7278c4),
	.w1(32'hbb856e22),
	.w2(32'h3b287687),
	.w3(32'h3ac6b97e),
	.w4(32'hbad04d7c),
	.w5(32'hbb133939),
	.w6(32'h3b9938c2),
	.w7(32'h3b862b0e),
	.w8(32'h3be61acf),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ea65f),
	.w1(32'hbb1fa18c),
	.w2(32'h3aa766dc),
	.w3(32'h3b798397),
	.w4(32'hbbb677f2),
	.w5(32'h3b5ecd76),
	.w6(32'h3beea728),
	.w7(32'h3a81c831),
	.w8(32'hbbedca10),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31e9d1),
	.w1(32'hb894eeb1),
	.w2(32'h3b2d11ec),
	.w3(32'h3c808598),
	.w4(32'h3a6387cd),
	.w5(32'hbb93fc5a),
	.w6(32'hba11aee6),
	.w7(32'hbc84cacb),
	.w8(32'hbc1ca325),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb175a31),
	.w1(32'hbb4bd362),
	.w2(32'hbc05b782),
	.w3(32'hbc2ed893),
	.w4(32'hbb521940),
	.w5(32'hbbc1b13d),
	.w6(32'hbbd655a6),
	.w7(32'hbb85fd13),
	.w8(32'hbc207fdd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cafd1),
	.w1(32'h39801424),
	.w2(32'h380bc82c),
	.w3(32'hbb748ead),
	.w4(32'hbadd0146),
	.w5(32'h3bae925d),
	.w6(32'hbbda586e),
	.w7(32'h3a38e74d),
	.w8(32'hbba589b9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c79ca),
	.w1(32'hbafc7613),
	.w2(32'hbabddb22),
	.w3(32'h3ba81656),
	.w4(32'h3b2f5683),
	.w5(32'hb96628af),
	.w6(32'h3baeda92),
	.w7(32'h3b985162),
	.w8(32'hb939c20f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acca1bf),
	.w1(32'h3b0f65cd),
	.w2(32'hbc6b7c5b),
	.w3(32'h3bd763aa),
	.w4(32'hb945ebc7),
	.w5(32'hbb813ea3),
	.w6(32'h3b8ab2e1),
	.w7(32'hba2cef52),
	.w8(32'h3b1de420),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8956c5),
	.w1(32'hbbe0797b),
	.w2(32'hbb027160),
	.w3(32'h3d855bf2),
	.w4(32'h3c9fcd42),
	.w5(32'hba0ec67a),
	.w6(32'h3d148c7d),
	.w7(32'h3c60a62f),
	.w8(32'hbb5a9f14),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07f108),
	.w1(32'h3bc3e011),
	.w2(32'hbd30924c),
	.w3(32'h3b1275f5),
	.w4(32'h3b995b2a),
	.w5(32'hbc0d033f),
	.w6(32'h3adaa3b9),
	.w7(32'hba42a4f7),
	.w8(32'h3cbb479a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc072ef),
	.w1(32'hbc942006),
	.w2(32'hbb02c500),
	.w3(32'h3daf552d),
	.w4(32'h3d9203cb),
	.w5(32'hb9ba8eaf),
	.w6(32'h3df77685),
	.w7(32'h3db99b0b),
	.w8(32'h399b9379),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e0193),
	.w1(32'h3c15611f),
	.w2(32'hbb2a9e06),
	.w3(32'h3b13fcc1),
	.w4(32'h3b19d842),
	.w5(32'h3b84ec52),
	.w6(32'h3ba77314),
	.w7(32'h3b8ef8f8),
	.w8(32'hba63c4f6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7965dd),
	.w1(32'h3b9f40fc),
	.w2(32'h3af50305),
	.w3(32'h3c1a254c),
	.w4(32'h3b8e8c57),
	.w5(32'h3833bc78),
	.w6(32'hbbb82c04),
	.w7(32'hbb60723b),
	.w8(32'hbbe94cec),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89fde2),
	.w1(32'hbbbc5c26),
	.w2(32'hba8c5365),
	.w3(32'h3abfc763),
	.w4(32'hba19354b),
	.w5(32'h3b149272),
	.w6(32'hbc3a2d0b),
	.w7(32'hbbda28bb),
	.w8(32'hbc1f15ae),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a7039),
	.w1(32'h3a914ccf),
	.w2(32'hbb0dbd26),
	.w3(32'hbafeb2e3),
	.w4(32'h3ba283ae),
	.w5(32'h3b40dea1),
	.w6(32'hbaf17722),
	.w7(32'hbb54acf4),
	.w8(32'hbc039791),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe246b4),
	.w1(32'h3aef194e),
	.w2(32'hbc23cdbe),
	.w3(32'h3baa80ce),
	.w4(32'h3afbbfd4),
	.w5(32'h3bbc5a0c),
	.w6(32'h3b588d04),
	.w7(32'h3b99b6b5),
	.w8(32'h3c10abc2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb529df0),
	.w1(32'hbb04bdd3),
	.w2(32'hba9517d2),
	.w3(32'h3cc54273),
	.w4(32'h3ca9c0be),
	.w5(32'h3b2d04b0),
	.w6(32'h3d0872c1),
	.w7(32'h3cc1af1b),
	.w8(32'hbb99ba36),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fbdb7c),
	.w1(32'hbae0f010),
	.w2(32'hba2ce929),
	.w3(32'hbae8ce55),
	.w4(32'hbba9b6f6),
	.w5(32'hbb417851),
	.w6(32'hbb75e4b1),
	.w7(32'hbb32ede6),
	.w8(32'hbac8faf4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96640b),
	.w1(32'hbbb6bbb5),
	.w2(32'hbbc28e07),
	.w3(32'hbb9105f4),
	.w4(32'hba77265f),
	.w5(32'hbc4515dc),
	.w6(32'hbc5d459b),
	.w7(32'h3b3cf304),
	.w8(32'hbc406601),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23df56),
	.w1(32'hbaca46d3),
	.w2(32'h3bfe6941),
	.w3(32'h3b47376d),
	.w4(32'h3bbee948),
	.w5(32'hbc301c20),
	.w6(32'hbc560bbc),
	.w7(32'hbb1db3f6),
	.w8(32'hbc67a3fe),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a6560),
	.w1(32'hbb67e3a4),
	.w2(32'hba40a62b),
	.w3(32'hbc15cd5a),
	.w4(32'hbb9defb5),
	.w5(32'hbaf8cc23),
	.w6(32'hbca84c4e),
	.w7(32'hbc09d4a0),
	.w8(32'hbb4d5362),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d2ac2),
	.w1(32'hb8d0cab2),
	.w2(32'hbd01a273),
	.w3(32'h3bd874ff),
	.w4(32'h3b2b9929),
	.w5(32'h3c19757e),
	.w6(32'h3b91d2d5),
	.w7(32'hbb082960),
	.w8(32'h3cf4c5b0),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dbdb7),
	.w1(32'hbc565e01),
	.w2(32'h3aed11ae),
	.w3(32'h3d9e3d8e),
	.w4(32'h3d7778be),
	.w5(32'h39d89b77),
	.w6(32'h3dcac8a7),
	.w7(32'h3d8fe3bc),
	.w8(32'hbbc15d00),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac980d7),
	.w1(32'hbae92bb7),
	.w2(32'h3bba9094),
	.w3(32'hbbb930bf),
	.w4(32'hbaedc924),
	.w5(32'h3bea398f),
	.w6(32'hbb250f4d),
	.w7(32'hbb63e492),
	.w8(32'h3b315c62),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af89e07),
	.w1(32'hbadf047e),
	.w2(32'h3b3a4651),
	.w3(32'h3b2d3ac9),
	.w4(32'hbb38338a),
	.w5(32'h3a44dd97),
	.w6(32'hbafa49c9),
	.w7(32'hbbaa273f),
	.w8(32'hbaa8025c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac45519),
	.w1(32'h3bf6269b),
	.w2(32'h3bb2755a),
	.w3(32'h38645c4e),
	.w4(32'h3b90bca0),
	.w5(32'h3b8bc802),
	.w6(32'h39d8d4e9),
	.w7(32'h3b1e3c04),
	.w8(32'h388966b8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24c283),
	.w1(32'h3a7b9d81),
	.w2(32'hbb9a8da0),
	.w3(32'h3acab041),
	.w4(32'hbb34762c),
	.w5(32'hbb82d7b1),
	.w6(32'hba8c8d72),
	.w7(32'hbb5bf390),
	.w8(32'hbb05b91a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb783167),
	.w1(32'hbbb02927),
	.w2(32'hbbe49e70),
	.w3(32'hbb0bfdbe),
	.w4(32'hbba053e0),
	.w5(32'hbb840964),
	.w6(32'hb842f8dd),
	.w7(32'h3a0c6d29),
	.w8(32'h395cc749),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d4ca8),
	.w1(32'hbb982d81),
	.w2(32'hbb8c2d7e),
	.w3(32'hbb55e7e8),
	.w4(32'h3bb2d496),
	.w5(32'h3bb3bf35),
	.w6(32'hbbe4be41),
	.w7(32'h3b8c0f45),
	.w8(32'hbb771308),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c9dea),
	.w1(32'hb99c2648),
	.w2(32'h3b8a74a2),
	.w3(32'h3b6260a9),
	.w4(32'h3bad439d),
	.w5(32'hbb0eef44),
	.w6(32'h3ab3273a),
	.w7(32'hbb6b18ca),
	.w8(32'h3b45ec78),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a2c95),
	.w1(32'h3b117ac3),
	.w2(32'hbb336969),
	.w3(32'h3ac8d92c),
	.w4(32'h3bc2960b),
	.w5(32'hbaf526e8),
	.w6(32'h3b8adc94),
	.w7(32'h3b88e0cf),
	.w8(32'hbafd36a3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36f500),
	.w1(32'h3bae0cac),
	.w2(32'hbb85d6fb),
	.w3(32'h3b67f06d),
	.w4(32'h39356164),
	.w5(32'hbab96245),
	.w6(32'hbbd178f9),
	.w7(32'h3a3b60ad),
	.w8(32'hbb9cd3e1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad74ccf),
	.w1(32'h3b80e535),
	.w2(32'hbb4a8805),
	.w3(32'h3a4279f5),
	.w4(32'h3b131ef7),
	.w5(32'h38066d7c),
	.w6(32'hbbb0c124),
	.w7(32'hbb2500e1),
	.w8(32'hb9c3b98e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bf84a),
	.w1(32'hbb119cea),
	.w2(32'h3ac1b57c),
	.w3(32'h3bab131f),
	.w4(32'h3bc73aa3),
	.w5(32'hbb91bde6),
	.w6(32'h3b9eefc1),
	.w7(32'h39cd8644),
	.w8(32'h3aaff4cc),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeffec7),
	.w1(32'h3a816b62),
	.w2(32'hbae9e79b),
	.w3(32'hbaae4291),
	.w4(32'hbb8c8b13),
	.w5(32'hbb65f287),
	.w6(32'hbba77b9f),
	.w7(32'hbb8c1834),
	.w8(32'hbb5249ad),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb903ac0b),
	.w1(32'hbabc74c9),
	.w2(32'hbb17b0de),
	.w3(32'hb984fc7e),
	.w4(32'hbb19db49),
	.w5(32'h3b4100c1),
	.w6(32'hba81d0c7),
	.w7(32'hbb4a2204),
	.w8(32'h3bf3fd08),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961e673),
	.w1(32'hbb62aff1),
	.w2(32'h3aa22c24),
	.w3(32'hbb73f18d),
	.w4(32'hbb7b892b),
	.w5(32'h3b0b61e1),
	.w6(32'h3bb98293),
	.w7(32'h3ac46081),
	.w8(32'hbacee470),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8bfcb),
	.w1(32'h3b697a8b),
	.w2(32'hbb1d3aed),
	.w3(32'hbb2f1cff),
	.w4(32'h3b85e73f),
	.w5(32'hbb1b09f9),
	.w6(32'h3a7bb952),
	.w7(32'h3b2f8244),
	.w8(32'hbae8ad1d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997bc45),
	.w1(32'hba0beb7f),
	.w2(32'h399a56b5),
	.w3(32'hba9b292f),
	.w4(32'h3a8d7a71),
	.w5(32'h3a515bf4),
	.w6(32'h3b890379),
	.w7(32'h3b51d593),
	.w8(32'hbab12726),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad9e99),
	.w1(32'hbb38ade8),
	.w2(32'hbbbbad77),
	.w3(32'hbad7d8b7),
	.w4(32'hbbde3956),
	.w5(32'h39da06d1),
	.w6(32'h3b430d26),
	.w7(32'hbbb97b23),
	.w8(32'hbb868557),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb862a45),
	.w1(32'hba2ee0d5),
	.w2(32'hba950c99),
	.w3(32'h3bb2083a),
	.w4(32'h3a2dea20),
	.w5(32'h3a5819b6),
	.w6(32'hbafe35a1),
	.w7(32'hbc39b35a),
	.w8(32'hbc33ce58),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b505160),
	.w1(32'hbb0de9dc),
	.w2(32'hbaf61608),
	.w3(32'hbb6fab05),
	.w4(32'hbbbcb8b5),
	.w5(32'hbb5356d4),
	.w6(32'hbc5f133c),
	.w7(32'hbbca7628),
	.w8(32'h3ae539b5),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d718f),
	.w1(32'hba07e140),
	.w2(32'h3b4d263f),
	.w3(32'h3a9b113d),
	.w4(32'h3b0d6eb1),
	.w5(32'h39968831),
	.w6(32'h3ba5c82b),
	.w7(32'h3b2a5cb4),
	.w8(32'hbc1df4eb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b732680),
	.w1(32'h3a617a39),
	.w2(32'h3b86bca4),
	.w3(32'h3b35c55b),
	.w4(32'hbbbe4759),
	.w5(32'h3b876e70),
	.w6(32'hbc0d029a),
	.w7(32'hbb99c52c),
	.w8(32'h3be769fa),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42405f),
	.w1(32'h3b66cb5d),
	.w2(32'h3b98edc4),
	.w3(32'h3ab4fc5c),
	.w4(32'h3b7d58f0),
	.w5(32'hbac16dc2),
	.w6(32'h3c00e11a),
	.w7(32'h3bed328a),
	.w8(32'h3b0ea352),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4658cb),
	.w1(32'hbbec9da8),
	.w2(32'h3a49f425),
	.w3(32'hbc16bddb),
	.w4(32'hbbb003d9),
	.w5(32'h3a12e3c2),
	.w6(32'h3b758431),
	.w7(32'h3b21657f),
	.w8(32'h3bfb62b4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1ad66),
	.w1(32'h3b36984b),
	.w2(32'h3aa92ab1),
	.w3(32'h3ba1642e),
	.w4(32'h3be9c3de),
	.w5(32'hba27795a),
	.w6(32'h3beb5177),
	.w7(32'h3c167329),
	.w8(32'h39ee176c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af659ee),
	.w1(32'h3969e610),
	.w2(32'h3bb9ca3c),
	.w3(32'h3a7d330e),
	.w4(32'h3b908780),
	.w5(32'hbb0e5128),
	.w6(32'hbbc742dd),
	.w7(32'hb9dd27a4),
	.w8(32'hbb6a88dd),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d66fe),
	.w1(32'h3b9a8959),
	.w2(32'h3a145b61),
	.w3(32'h394bb95e),
	.w4(32'hb84eefd5),
	.w5(32'hbb664c8c),
	.w6(32'h3afc6dc5),
	.w7(32'h3bee2be4),
	.w8(32'hbac093d3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c66ac8),
	.w1(32'hba4da44b),
	.w2(32'h3c65277e),
	.w3(32'hb9ec9f4d),
	.w4(32'hb9500aff),
	.w5(32'h3bbba8a1),
	.w6(32'hbabbe3af),
	.w7(32'hba9733ea),
	.w8(32'h3a473791),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82c032),
	.w1(32'h3c77d3ed),
	.w2(32'h3bb28103),
	.w3(32'hbbb353a9),
	.w4(32'hbb102ce7),
	.w5(32'h39974b60),
	.w6(32'hbc257d95),
	.w7(32'hbbb9935b),
	.w8(32'h3b8ae692),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b585374),
	.w1(32'h3b3a2886),
	.w2(32'h3b0bc7b5),
	.w3(32'hbbc39d98),
	.w4(32'h39a7a2f2),
	.w5(32'h3a013090),
	.w6(32'hbb210d5e),
	.w7(32'h3ada5b0f),
	.w8(32'hbb2f7dfa),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba55e22),
	.w1(32'h3a3a2f3d),
	.w2(32'h3afe88c7),
	.w3(32'h3ba3175c),
	.w4(32'hba5d80bd),
	.w5(32'h3b2391be),
	.w6(32'h3b0460a0),
	.w7(32'hbbaabd01),
	.w8(32'h3bf8a5a7),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93663c7),
	.w1(32'h3bc51ce1),
	.w2(32'hbb19c155),
	.w3(32'h3b9cfe9e),
	.w4(32'h3b7d47d8),
	.w5(32'hbbbd9f38),
	.w6(32'h3c1478cd),
	.w7(32'h3be4c319),
	.w8(32'hbb84deba),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad051f),
	.w1(32'hbb8039b4),
	.w2(32'hbb8cbdfb),
	.w3(32'h3b060c35),
	.w4(32'hbb40e7e3),
	.w5(32'h38dcba96),
	.w6(32'h3994105d),
	.w7(32'h3b298dda),
	.w8(32'hbbdc793b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb967674),
	.w1(32'hba11acd0),
	.w2(32'hbc15e5a6),
	.w3(32'h3a91b1e4),
	.w4(32'hbb0706e0),
	.w5(32'hbc026b0b),
	.w6(32'hba6664eb),
	.w7(32'h3b4d4477),
	.w8(32'hbbf06b44),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74993b),
	.w1(32'h3b3b87e7),
	.w2(32'h3aca83f0),
	.w3(32'hbba1c44f),
	.w4(32'h3aa0bcec),
	.w5(32'h3b0e429f),
	.w6(32'hbbe088b1),
	.w7(32'hbb14a1f1),
	.w8(32'h3b25eefa),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule