module layer_10_featuremap_148(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a81604),
	.w1(32'h370b5d69),
	.w2(32'hb7d92dac),
	.w3(32'hb645ef5e),
	.w4(32'h36e62d48),
	.w5(32'hb7feb83f),
	.w6(32'h37a79cc3),
	.w7(32'hb752450b),
	.w8(32'h377edf81),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f52d2),
	.w1(32'h3882c328),
	.w2(32'h38765dc0),
	.w3(32'h38a7a905),
	.w4(32'h38948b90),
	.w5(32'h386473db),
	.w6(32'h38a948c1),
	.w7(32'h389bc603),
	.w8(32'h3870c800),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c1c1f8),
	.w1(32'hb7461ef6),
	.w2(32'hb72d7b25),
	.w3(32'hb6ef3026),
	.w4(32'hb71ddbfa),
	.w5(32'hb73b3385),
	.w6(32'hb73e9216),
	.w7(32'hb71fc938),
	.w8(32'hb620e2cf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72ae124),
	.w1(32'hb7b5677b),
	.w2(32'hb7995a0a),
	.w3(32'hb726e74d),
	.w4(32'hb6a81127),
	.w5(32'h37087ea4),
	.w6(32'hb7b39c1b),
	.w7(32'hb819431a),
	.w8(32'hb80136ba),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eacd3b),
	.w1(32'hb745d5ce),
	.w2(32'h379509df),
	.w3(32'hb6aa40f9),
	.w4(32'hb7833818),
	.w5(32'h37304693),
	.w6(32'hb6b98ee3),
	.w7(32'h378334bc),
	.w8(32'hb7302820),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70154cd),
	.w1(32'hb72a48d4),
	.w2(32'h378e35df),
	.w3(32'hb7433b31),
	.w4(32'hb74ec903),
	.w5(32'h37899a08),
	.w6(32'h35f47135),
	.w7(32'h37cd1bd9),
	.w8(32'hb535762b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7defada),
	.w1(32'h373ce444),
	.w2(32'h380c76d3),
	.w3(32'hb7cb5fb4),
	.w4(32'h36860f62),
	.w5(32'h374296fc),
	.w6(32'h3605a101),
	.w7(32'h37923a6c),
	.w8(32'hb73e5574),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8abf7bd),
	.w1(32'hb85067be),
	.w2(32'hb606a590),
	.w3(32'hb8a7b110),
	.w4(32'hb8ceadc7),
	.w5(32'hb8940775),
	.w6(32'hb92b2c07),
	.w7(32'hb960b989),
	.w8(32'hb95b77f9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cfe1b1),
	.w1(32'h387290ec),
	.w2(32'h38877032),
	.w3(32'h382b76cf),
	.w4(32'h381f300c),
	.w5(32'h3864a3bd),
	.w6(32'h38214380),
	.w7(32'hb7b9605b),
	.w8(32'hb7afe539),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3c8e5),
	.w1(32'h388e4cd6),
	.w2(32'hb86e5a23),
	.w3(32'h38f15160),
	.w4(32'h38dda25e),
	.w5(32'h360030bd),
	.w6(32'h38d8c36f),
	.w7(32'h3886ab85),
	.w8(32'hb747113e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bb01c0),
	.w1(32'hb818d2e3),
	.w2(32'h38b9dfea),
	.w3(32'hb6e85ddf),
	.w4(32'h380ecd7c),
	.w5(32'h38872086),
	.w6(32'hb7d566f9),
	.w7(32'h3821de15),
	.w8(32'h38bd0f45),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b785c9),
	.w1(32'hb8638148),
	.w2(32'h3856a922),
	.w3(32'hb809f1ba),
	.w4(32'hb830e4ca),
	.w5(32'h36974052),
	.w6(32'hb841bdbf),
	.w7(32'hb79edc55),
	.w8(32'hb809533a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a047e7),
	.w1(32'h380da79d),
	.w2(32'hb8a63f99),
	.w3(32'h3808a6f0),
	.w4(32'h386740d8),
	.w5(32'hb89e0750),
	.w6(32'h379f9dbb),
	.w7(32'hb60ae704),
	.w8(32'hb91822cd),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c816e9),
	.w1(32'h37be3b7a),
	.w2(32'h378fcb08),
	.w3(32'h385cb923),
	.w4(32'hb78e310d),
	.w5(32'h37ec0ef4),
	.w6(32'h388a5618),
	.w7(32'h3786e57d),
	.w8(32'h37da25da),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0c351),
	.w1(32'h3855d25e),
	.w2(32'h367dd303),
	.w3(32'h38891f00),
	.w4(32'h382db767),
	.w5(32'h373b8794),
	.w6(32'h38115c00),
	.w7(32'hb87f2b3c),
	.w8(32'hb8a8e66e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e4407f),
	.w1(32'h388f4c75),
	.w2(32'h3754456c),
	.w3(32'h391b970c),
	.w4(32'h381762fc),
	.w5(32'h37335043),
	.w6(32'h382b1a1c),
	.w7(32'hb8923a08),
	.w8(32'hb8864983),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37742b9b),
	.w1(32'h33b5c713),
	.w2(32'h389b5248),
	.w3(32'h39284803),
	.w4(32'h38bd6c62),
	.w5(32'h39304982),
	.w6(32'h38888832),
	.w7(32'h37aa5018),
	.w8(32'h39188bc8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914a292),
	.w1(32'hb901ef69),
	.w2(32'hb92b74fe),
	.w3(32'hb934a3dc),
	.w4(32'hb930f184),
	.w5(32'hb95b149a),
	.w6(32'hb9b6e91b),
	.w7(32'hb9a28013),
	.w8(32'hb9a1fb1c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a51441),
	.w1(32'hb6d96e96),
	.w2(32'hb866780f),
	.w3(32'hb887192c),
	.w4(32'hb81f3806),
	.w5(32'hb8b63c6b),
	.w6(32'hb903f6d3),
	.w7(32'hb8f575a4),
	.w8(32'hb90875a8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3657afd5),
	.w1(32'hb59ea6cd),
	.w2(32'h36dc57ba),
	.w3(32'h34d043c9),
	.w4(32'hb502c41f),
	.w5(32'h36f84574),
	.w6(32'h35c05646),
	.w7(32'h370007f0),
	.w8(32'h370fd297),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dd855d),
	.w1(32'hb73d3a13),
	.w2(32'h37c3f23b),
	.w3(32'h36c22dd2),
	.w4(32'hb766ae60),
	.w5(32'h37a7cd1d),
	.w6(32'hb6c8a1bb),
	.w7(32'h37baac42),
	.w8(32'h369954a2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc0471),
	.w1(32'hb6852723),
	.w2(32'hb6f08169),
	.w3(32'h37ed5270),
	.w4(32'h3735ea73),
	.w5(32'h36095321),
	.w6(32'h378bfad8),
	.w7(32'hb66f90ab),
	.w8(32'h37061a92),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7977653),
	.w1(32'hb93df684),
	.w2(32'hb9137fc7),
	.w3(32'hb8bfab8c),
	.w4(32'hb9276d6b),
	.w5(32'hb8e6939b),
	.w6(32'hb9cad67b),
	.w7(32'hb9d910eb),
	.w8(32'hba218eb4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966a456),
	.w1(32'h3916079d),
	.w2(32'h37ea6478),
	.w3(32'h39908697),
	.w4(32'h3929688c),
	.w5(32'hb74fd729),
	.w6(32'h39275e91),
	.w7(32'h3823dba8),
	.w8(32'hb91272b3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d2bb6),
	.w1(32'hb84d2897),
	.w2(32'hb8dea1a7),
	.w3(32'h391f149f),
	.w4(32'hb8ed69d9),
	.w5(32'hb99dc2d0),
	.w6(32'h38766310),
	.w7(32'hb9258814),
	.w8(32'hb9a136cc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d3ac55),
	.w1(32'h383e90bc),
	.w2(32'h3866e2b4),
	.w3(32'hb6977bac),
	.w4(32'h38572721),
	.w5(32'h3874723f),
	.w6(32'h378a692e),
	.w7(32'h377c45e5),
	.w8(32'h3756623e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3711be9f),
	.w1(32'hb63c6027),
	.w2(32'h378dd984),
	.w3(32'h363c6a02),
	.w4(32'hb706f50c),
	.w5(32'h372f53e2),
	.w6(32'h36eca3de),
	.w7(32'h3764813d),
	.w8(32'h37092253),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389993fc),
	.w1(32'h385945d7),
	.w2(32'hb6e57198),
	.w3(32'h3868a636),
	.w4(32'h3889a7f5),
	.w5(32'h3779edea),
	.w6(32'h3841f5fa),
	.w7(32'h38712cf6),
	.w8(32'h37f53fa6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382a6582),
	.w1(32'h3875d146),
	.w2(32'h391a24f6),
	.w3(32'h38833697),
	.w4(32'hb8edb734),
	.w5(32'h387dfb85),
	.w6(32'hb8a2a85b),
	.w7(32'h36d669bf),
	.w8(32'h3878ffc4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f20e07),
	.w1(32'h39290220),
	.w2(32'h391a00f3),
	.w3(32'h393ab0c7),
	.w4(32'h397e148d),
	.w5(32'h39718d7c),
	.w6(32'h37c7aee5),
	.w7(32'h38a91ff0),
	.w8(32'h38da5c42),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3827d784),
	.w1(32'hb73071bc),
	.w2(32'h37a8efb7),
	.w3(32'h383578f2),
	.w4(32'hb76c9a07),
	.w5(32'h37a27fa7),
	.w6(32'hb6e2d834),
	.w7(32'h37315ef1),
	.w8(32'h370a411c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b8a276),
	.w1(32'h377307dd),
	.w2(32'h3731846c),
	.w3(32'h36c3b7eb),
	.w4(32'hb6f31446),
	.w5(32'h380a48e0),
	.w6(32'hb7203b62),
	.w7(32'h37b1c29f),
	.w8(32'h38206c17),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914a16b),
	.w1(32'h370cdd69),
	.w2(32'hb80b05f7),
	.w3(32'h39222c4b),
	.w4(32'hb7f7e675),
	.w5(32'hb888f439),
	.w6(32'h38ec9c51),
	.w7(32'hb7c89308),
	.w8(32'hb8784928),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f1277),
	.w1(32'hb603addf),
	.w2(32'h385ff55d),
	.w3(32'h382a4892),
	.w4(32'hb78918b9),
	.w5(32'h384a321d),
	.w6(32'h37c3d488),
	.w7(32'h37defd55),
	.w8(32'h376f66d8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812f500),
	.w1(32'hb6d988a9),
	.w2(32'hb59629e0),
	.w3(32'h3829dda5),
	.w4(32'h3650ab2b),
	.w5(32'h369d7f85),
	.w6(32'h363b99d7),
	.w7(32'h35c01e7a),
	.w8(32'h372f7674),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6978720),
	.w1(32'hb715bd90),
	.w2(32'h3724e6e9),
	.w3(32'hb6efb398),
	.w4(32'hb7b9e7b1),
	.w5(32'hb732e315),
	.w6(32'hb8008b43),
	.w7(32'hb8127beb),
	.w8(32'hb85de2d7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fc49a),
	.w1(32'hb8b9fccb),
	.w2(32'h377a5537),
	.w3(32'hb987b194),
	.w4(32'h383dc09a),
	.w5(32'h38ca71c9),
	.w6(32'hb94c2c76),
	.w7(32'hb8b7651e),
	.w8(32'hb81cba78),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90009ad),
	.w1(32'h39ab87c5),
	.w2(32'h3956a2f1),
	.w3(32'h3865764c),
	.w4(32'h399962ad),
	.w5(32'h398bbce4),
	.w6(32'h38e37e3e),
	.w7(32'h396f49af),
	.w8(32'h3925016d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39040324),
	.w1(32'h39a96539),
	.w2(32'h38fb7ee5),
	.w3(32'hb70c00fb),
	.w4(32'h392e23a9),
	.w5(32'h38b92628),
	.w6(32'h38097cb1),
	.w7(32'h388cbfd2),
	.w8(32'hb6345223),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385f4f35),
	.w1(32'h380e9cd7),
	.w2(32'h3785ea94),
	.w3(32'h3883a2df),
	.w4(32'h38241749),
	.w5(32'h3709eea5),
	.w6(32'h387ae76f),
	.w7(32'h3818a826),
	.w8(32'h36a56b0c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e8a63d),
	.w1(32'hb84562d6),
	.w2(32'h38a22cb0),
	.w3(32'h373b9fd9),
	.w4(32'hb70f247f),
	.w5(32'h38c1dde3),
	.w6(32'hb84c722b),
	.w7(32'h3841e5e8),
	.w8(32'h3829805f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a18db7),
	.w1(32'hb75d5bec),
	.w2(32'hb5f7d9a2),
	.w3(32'h383d491c),
	.w4(32'h377b433d),
	.w5(32'h37e02474),
	.w6(32'hb0f8a7d0),
	.w7(32'h37ea5b12),
	.w8(32'h385090f4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cd65bc),
	.w1(32'h384bbed8),
	.w2(32'h38ea49a0),
	.w3(32'hb81cc53d),
	.w4(32'h38351332),
	.w5(32'h38baa960),
	.w6(32'hb87ee435),
	.w7(32'h38b08583),
	.w8(32'h388eb2b4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d08e55),
	.w1(32'h381bf6ec),
	.w2(32'h38b4b185),
	.w3(32'h38c19601),
	.w4(32'h3955a8a5),
	.w5(32'hb822e8e8),
	.w6(32'hb8aa3a7a),
	.w7(32'h389bc1b6),
	.w8(32'hb9a985d2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919da18),
	.w1(32'h39789104),
	.w2(32'h37d4c15a),
	.w3(32'h392cafae),
	.w4(32'h3991e6b7),
	.w5(32'h387fabab),
	.w6(32'h38964875),
	.w7(32'h383e60a2),
	.w8(32'hb87517cb),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919f171),
	.w1(32'h392dc9ec),
	.w2(32'h37b14c46),
	.w3(32'h394c1d69),
	.w4(32'h396c3433),
	.w5(32'h3589ef88),
	.w6(32'h38fd7155),
	.w7(32'h3820d1ac),
	.w8(32'hb91a90f6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac15bb),
	.w1(32'h39c4b2a1),
	.w2(32'h39449eac),
	.w3(32'h39aab8ca),
	.w4(32'h39da4bb7),
	.w5(32'h3969a470),
	.w6(32'h39842ef1),
	.w7(32'h3909bd8b),
	.w8(32'hb86ac811),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7597c04),
	.w1(32'hb81f5bf5),
	.w2(32'hb85d2d07),
	.w3(32'hb7f76763),
	.w4(32'hb8ec2e0f),
	.w5(32'hb89e7a8d),
	.w6(32'hb9a1e546),
	.w7(32'hb9b68285),
	.w8(32'hb9a15eec),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb829a706),
	.w1(32'hb86f6663),
	.w2(32'hb73ea170),
	.w3(32'hb7c56742),
	.w4(32'h381c8449),
	.w5(32'h37f5bca6),
	.w6(32'hb88215d5),
	.w7(32'hb78ecf4a),
	.w8(32'hb72ff05a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b7b22d),
	.w1(32'h38e45d7b),
	.w2(32'h38cc7004),
	.w3(32'h39148021),
	.w4(32'h390fe4c0),
	.w5(32'h386f32aa),
	.w6(32'h3900aea2),
	.w7(32'h37a636e8),
	.w8(32'hb87d7d52),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf24d4),
	.w1(32'h382e51e8),
	.w2(32'h38396194),
	.w3(32'h390df7f4),
	.w4(32'h38bf58eb),
	.w5(32'h381c8c60),
	.w6(32'h3804baa3),
	.w7(32'h37662427),
	.w8(32'h3782ae40),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382aa2d9),
	.w1(32'h3817aa0e),
	.w2(32'hb8128c63),
	.w3(32'h3824eda5),
	.w4(32'h385e7cde),
	.w5(32'hb7da375d),
	.w6(32'h38060f25),
	.w7(32'hb80a2822),
	.w8(32'hb7557b56),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382e184a),
	.w1(32'hb7e5e221),
	.w2(32'hb765fd49),
	.w3(32'h37c1c859),
	.w4(32'hb82c7cfd),
	.w5(32'hb7cc314f),
	.w6(32'hb7c7ad77),
	.w7(32'hb82a3c75),
	.w8(32'hb87c2481),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c80133),
	.w1(32'hb8a50b1a),
	.w2(32'hb8e7b7ed),
	.w3(32'hb8dc9322),
	.w4(32'hb8dd3bc8),
	.w5(32'hb8e11333),
	.w6(32'hb93397b5),
	.w7(32'hb94ec011),
	.w8(32'hb98922c7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3612713c),
	.w1(32'hb793ac12),
	.w2(32'hb6ef842d),
	.w3(32'hb7411f5d),
	.w4(32'hb8023e58),
	.w5(32'hb8024777),
	.w6(32'hb821072f),
	.w7(32'hb8268c74),
	.w8(32'hb86230eb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36271484),
	.w1(32'hb83d6dc5),
	.w2(32'h3817e6b3),
	.w3(32'h361e6ef9),
	.w4(32'hb8097652),
	.w5(32'h3848113c),
	.w6(32'hb85cfccd),
	.w7(32'h37dec128),
	.w8(32'h3723f319),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aa71e3),
	.w1(32'hb6e619f9),
	.w2(32'h37a58a2e),
	.w3(32'h37f6684e),
	.w4(32'h33d5132d),
	.w5(32'h37c5cf8a),
	.w6(32'hb7078a38),
	.w7(32'h378b36b5),
	.w8(32'h37a33699),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380bcc93),
	.w1(32'h36862e74),
	.w2(32'h384d9a6d),
	.w3(32'h3810531e),
	.w4(32'hb73c0a53),
	.w5(32'h380f6e03),
	.w6(32'hb6471c8d),
	.w7(32'h381530da),
	.w8(32'h372a53fa),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378f7d6d),
	.w1(32'h3802938d),
	.w2(32'h38242bb6),
	.w3(32'h37a97d0e),
	.w4(32'h383d7437),
	.w5(32'h3814467a),
	.w6(32'h3725bc9c),
	.w7(32'h37d215bb),
	.w8(32'h3785fc39),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce67cd),
	.w1(32'h373980e5),
	.w2(32'h38802709),
	.w3(32'h37ba59c0),
	.w4(32'h3832f81c),
	.w5(32'h383a8349),
	.w6(32'hb76c2924),
	.w7(32'h37c92b0d),
	.w8(32'h36ab320b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a95dcb),
	.w1(32'h35a31154),
	.w2(32'hb73c7d85),
	.w3(32'h3747d308),
	.w4(32'h3752a14f),
	.w5(32'hb817eb11),
	.w6(32'hb87122fc),
	.w7(32'hb871b3d1),
	.w8(32'hb8ef75f4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80cdfdd),
	.w1(32'hb89de664),
	.w2(32'hb84be740),
	.w3(32'hb8c2ecde),
	.w4(32'hb8625c21),
	.w5(32'hb800723c),
	.w6(32'hb8cc0e3b),
	.w7(32'hb8e58011),
	.w8(32'hb8c22674),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f5311e),
	.w1(32'h37b20a6e),
	.w2(32'hb819abf1),
	.w3(32'hb6cc6501),
	.w4(32'h380fdb8d),
	.w5(32'hb80d9784),
	.w6(32'h3791b0b3),
	.w7(32'hb8183d55),
	.w8(32'h37b7ae41),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787c1b0),
	.w1(32'hb7419c51),
	.w2(32'hb6bfd620),
	.w3(32'h36a4e1ad),
	.w4(32'hb7307956),
	.w5(32'hb6c2bf84),
	.w6(32'hb724eae7),
	.w7(32'hb5e004b4),
	.w8(32'h37263040),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782c004),
	.w1(32'hb6d321f9),
	.w2(32'h368e8a02),
	.w3(32'hb7a4772e),
	.w4(32'hb806149a),
	.w5(32'hb64a4363),
	.w6(32'hb6ca6338),
	.w7(32'hb78cca85),
	.w8(32'hb6e91aed),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fa493f),
	.w1(32'hb7a9a69c),
	.w2(32'h37a22e90),
	.w3(32'hb6d37c50),
	.w4(32'hb7bf795e),
	.w5(32'h37606b48),
	.w6(32'hb6b42014),
	.w7(32'h37e28f28),
	.w8(32'h37a4fb8f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6faa836),
	.w1(32'hb70d5f82),
	.w2(32'hb6e7628b),
	.w3(32'h36772c30),
	.w4(32'h37f78f54),
	.w5(32'h3841f95e),
	.w6(32'hb867b0fc),
	.w7(32'hb8063300),
	.w8(32'hb78d4e6a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39327250),
	.w1(32'h37fc9e1a),
	.w2(32'h38a3be2d),
	.w3(32'h3927d952),
	.w4(32'hb74f7f73),
	.w5(32'hb6a32fe8),
	.w6(32'hb83fbf4f),
	.w7(32'h37868734),
	.w8(32'hb8fb8a39),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899a26d),
	.w1(32'hb8a5b3da),
	.w2(32'hb93aafd5),
	.w3(32'hb73bac8b),
	.w4(32'hb8a73c6f),
	.w5(32'hb943b91f),
	.w6(32'hb93da553),
	.w7(32'hb972ee24),
	.w8(32'hb9a6e924),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971cd43),
	.w1(32'h39775fb9),
	.w2(32'h3790550c),
	.w3(32'h398c80df),
	.w4(32'h395facf1),
	.w5(32'hb783c108),
	.w6(32'h39045e26),
	.w7(32'h388e8636),
	.w8(32'hb8e027c3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73156b0),
	.w1(32'hb6a07974),
	.w2(32'hb71701b3),
	.w3(32'hb73f11ae),
	.w4(32'hb6a2f78f),
	.w5(32'hb7218a18),
	.w6(32'hb5cf2163),
	.w7(32'hb6bd0362),
	.w8(32'h36e0825b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d53f3f),
	.w1(32'hb704ec71),
	.w2(32'h37298a72),
	.w3(32'hb71aabcf),
	.w4(32'hb6c8e794),
	.w5(32'h3759185f),
	.w6(32'h369a44d4),
	.w7(32'h37882bc9),
	.w8(32'h36a1045a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb771cc6a),
	.w1(32'hb6b1d133),
	.w2(32'h369af477),
	.w3(32'hb735bbd5),
	.w4(32'hb6998b0c),
	.w5(32'h3690df37),
	.w6(32'h36b9e398),
	.w7(32'h3768d551),
	.w8(32'h36a7bc1c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370d6639),
	.w1(32'h362a5bd7),
	.w2(32'h380604aa),
	.w3(32'h3733d088),
	.w4(32'hb5acc013),
	.w5(32'h380d017e),
	.w6(32'hb802d2c7),
	.w7(32'hb67594cc),
	.w8(32'h365666ae),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cd01e4),
	.w1(32'h3697a3ee),
	.w2(32'h3781a5dd),
	.w3(32'hb7408531),
	.w4(32'hb710d320),
	.w5(32'h368cf7a7),
	.w6(32'hb670a724),
	.w7(32'h368e7f88),
	.w8(32'h37d1181f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a24c88),
	.w1(32'hb8b56617),
	.w2(32'hb90e033d),
	.w3(32'hb8dcd185),
	.w4(32'hb8b34f14),
	.w5(32'hb8918a18),
	.w6(32'hb91fdc89),
	.w7(32'hb9430204),
	.w8(32'hb92b2d0b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e091df),
	.w1(32'hb946c111),
	.w2(32'hb93122d7),
	.w3(32'hb8fa310b),
	.w4(32'hb989b6be),
	.w5(32'hb94c0fcc),
	.w6(32'hb984bdc8),
	.w7(32'hb9a6841d),
	.w8(32'hb99d837e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d72fce),
	.w1(32'h38e4b2b1),
	.w2(32'h35ba188b),
	.w3(32'h38f59d82),
	.w4(32'h38ef5af4),
	.w5(32'hb800cee2),
	.w6(32'h3890c905),
	.w7(32'hb598bd9c),
	.w8(32'hb881d3be),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b85141),
	.w1(32'hb71f3a82),
	.w2(32'hb7f271db),
	.w3(32'hb7be4dbb),
	.w4(32'hb80a9ee2),
	.w5(32'hb868294e),
	.w6(32'hb88e7a73),
	.w7(32'hb88bbd34),
	.w8(32'hb8e6cb7d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38138d19),
	.w1(32'hb6db9135),
	.w2(32'h361e52d0),
	.w3(32'h38442f1b),
	.w4(32'hb715c742),
	.w5(32'hb73f6512),
	.w6(32'h3703252b),
	.w7(32'h373683e2),
	.w8(32'hb8800dc5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894f9e0),
	.w1(32'hb8a8f64a),
	.w2(32'h3830fe5c),
	.w3(32'h38961f94),
	.w4(32'hb88f9b53),
	.w5(32'h382044c8),
	.w6(32'hb89740f6),
	.w7(32'h381c5814),
	.w8(32'hb79b3728),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72e5b3d),
	.w1(32'hb8afaf87),
	.w2(32'hb8de4735),
	.w3(32'hb7f79730),
	.w4(32'hb8c465ba),
	.w5(32'hb916f701),
	.w6(32'hb90168de),
	.w7(32'hb91bb2d8),
	.w8(32'hb937ac8e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ab51b3),
	.w1(32'hb75c7296),
	.w2(32'h364c3735),
	.w3(32'hb59ce817),
	.w4(32'hb7122849),
	.w5(32'h36e0dbfa),
	.w6(32'hb784a0c3),
	.w7(32'hb51a6d8a),
	.w8(32'h3627a2b2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3695ffc4),
	.w1(32'h37007a69),
	.w2(32'h34b500d2),
	.w3(32'h37044519),
	.w4(32'h37088cd9),
	.w5(32'hb5b4f8f3),
	.w6(32'h36ee8fbb),
	.w7(32'h35466183),
	.w8(32'h36db9057),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374d3df4),
	.w1(32'hb8b676b6),
	.w2(32'h3696aae4),
	.w3(32'h37150070),
	.w4(32'hb89f73cc),
	.w5(32'h370bc05d),
	.w6(32'hb8b97f3c),
	.w7(32'hb707647c),
	.w8(32'h372e22e0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37998ac8),
	.w1(32'h367e8dff),
	.w2(32'h36d3179b),
	.w3(32'h37d5f708),
	.w4(32'h360b143e),
	.w5(32'h35d5fa55),
	.w6(32'h35d88453),
	.w7(32'h37227302),
	.w8(32'h37843464),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f1f1af),
	.w1(32'h38ec7816),
	.w2(32'h38a1b14d),
	.w3(32'h38cb3383),
	.w4(32'h3901c91c),
	.w5(32'h38837d66),
	.w6(32'h38b54f3d),
	.w7(32'h38b1efb9),
	.w8(32'h38cd76a8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c059a5),
	.w1(32'hb717fec1),
	.w2(32'h3744702f),
	.w3(32'h3743837f),
	.w4(32'hb7490260),
	.w5(32'h370ee34e),
	.w6(32'hb790ddff),
	.w7(32'hb52eb915),
	.w8(32'hb72d2e1b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e05f6f),
	.w1(32'h3708a3d5),
	.w2(32'hb8010182),
	.w3(32'h376f54c4),
	.w4(32'hb68e6319),
	.w5(32'hb791b07d),
	.w6(32'h371b98f0),
	.w7(32'hb78099c8),
	.w8(32'hb8678c8e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fb61e),
	.w1(32'hb99f6eae),
	.w2(32'hb967ef4e),
	.w3(32'hb9b1b874),
	.w4(32'hb9b0f6e6),
	.w5(32'hb9401f71),
	.w6(32'hb9f1c543),
	.w7(32'hb9ea41b5),
	.w8(32'hb9aeb3e3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb779ee8b),
	.w1(32'h388ab421),
	.w2(32'h379554a9),
	.w3(32'hb65cc4fa),
	.w4(32'h382b62dd),
	.w5(32'hb788b4bf),
	.w6(32'hb78ee1b2),
	.w7(32'h383dfed4),
	.w8(32'hb71345d2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379487db),
	.w1(32'hb74c8e6b),
	.w2(32'hb6c53383),
	.w3(32'h383d0b3d),
	.w4(32'hb73942ab),
	.w5(32'hb7c480cc),
	.w6(32'h37a04511),
	.w7(32'hb892fd78),
	.w8(32'hb93be7ce),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aeb7c9),
	.w1(32'h37fb4f50),
	.w2(32'hb857a24b),
	.w3(32'h38b4777c),
	.w4(32'h38360baf),
	.w5(32'hb88b8b35),
	.w6(32'h385291bd),
	.w7(32'h388eab74),
	.w8(32'hb822b959),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384d905a),
	.w1(32'hb825c2db),
	.w2(32'h375ba4d7),
	.w3(32'h3890925b),
	.w4(32'hb790a429),
	.w5(32'hb74c69be),
	.w6(32'hb8a68c52),
	.w7(32'hb8543ae9),
	.w8(32'hb9425578),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a63071),
	.w1(32'hb667a886),
	.w2(32'hb771512f),
	.w3(32'h38b00c35),
	.w4(32'hb660eb3b),
	.w5(32'hb7e9ba8b),
	.w6(32'h37b85bc1),
	.w7(32'hb8444b7a),
	.w8(32'hb8956acb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388fe359),
	.w1(32'h38b0e049),
	.w2(32'h37d732e1),
	.w3(32'h38b0dfcd),
	.w4(32'h38a7af80),
	.w5(32'h37c48a48),
	.w6(32'h3888dccf),
	.w7(32'h3873b2dd),
	.w8(32'hb701514a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb836a252),
	.w1(32'hb8b9d4aa),
	.w2(32'hb812649b),
	.w3(32'hb8b62d4d),
	.w4(32'hb89a4d9e),
	.w5(32'hb89d348f),
	.w6(32'hb8a306f6),
	.w7(32'hb8183dca),
	.w8(32'hb912d83f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386fb888),
	.w1(32'h39255891),
	.w2(32'hb942c2d1),
	.w3(32'hb8d166ff),
	.w4(32'h39125a36),
	.w5(32'hb94806b9),
	.w6(32'hb913ff39),
	.w7(32'hb95cba82),
	.w8(32'hb9d5f09f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899c279),
	.w1(32'h39143593),
	.w2(32'hb89ade79),
	.w3(32'h3902ec3c),
	.w4(32'h39ccfb74),
	.w5(32'h38d37189),
	.w6(32'hb6b75fee),
	.w7(32'h38fd1ecd),
	.w8(32'hb9349124),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1aa54),
	.w1(32'hb933548d),
	.w2(32'hb941346c),
	.w3(32'hb8d02a35),
	.w4(32'hb96dc6fd),
	.w5(32'hb93f9f54),
	.w6(32'hb95a776a),
	.w7(32'hb994a364),
	.w8(32'hb9a95c1b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b9aa94),
	.w1(32'h3952fb11),
	.w2(32'h39155a5f),
	.w3(32'h3937915c),
	.w4(32'h3a043dc2),
	.w5(32'h398fb224),
	.w6(32'h394f3179),
	.w7(32'h39197b9f),
	.w8(32'h383ec3ca),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e2621),
	.w1(32'h3959d979),
	.w2(32'h38f704fe),
	.w3(32'h39127992),
	.w4(32'h38b13c41),
	.w5(32'hb64fe10f),
	.w6(32'h39735bcb),
	.w7(32'hb8fec683),
	.w8(32'hb9352613),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8861318),
	.w1(32'h37057916),
	.w2(32'hb7b4c13f),
	.w3(32'hb890c84c),
	.w4(32'h3884389d),
	.w5(32'hb83ed15c),
	.w6(32'hb8f70b75),
	.w7(32'h38a677ac),
	.w8(32'hb97082b1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369bcf47),
	.w1(32'hb94bef7e),
	.w2(32'hb9ab7ece),
	.w3(32'hb8ebac48),
	.w4(32'hb8fd133c),
	.w5(32'hb91fab41),
	.w6(32'hb8b7e073),
	.w7(32'hb8aa8e32),
	.w8(32'hb99704a7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee735a),
	.w1(32'hb973378e),
	.w2(32'hb98ede81),
	.w3(32'hb8c2f3e6),
	.w4(32'hb980980c),
	.w5(32'hb92928a9),
	.w6(32'hb97f049a),
	.w7(32'hb996c980),
	.w8(32'hb9b9ec68),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6e54e),
	.w1(32'h38380be5),
	.w2(32'hb69e87eb),
	.w3(32'h390b2087),
	.w4(32'h37b18474),
	.w5(32'h371fa9d2),
	.w6(32'h38e7da78),
	.w7(32'h37fe0f8a),
	.w8(32'h370ce352),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38198bfb),
	.w1(32'hb70cdeeb),
	.w2(32'hb7a6d8f6),
	.w3(32'h37d5a3b1),
	.w4(32'hb5cf3dbb),
	.w5(32'hb7a8942f),
	.w6(32'hb4b0441b),
	.w7(32'hb7829488),
	.w8(32'hb7b00294),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3800d2d4),
	.w1(32'hb7b62b62),
	.w2(32'h3858211e),
	.w3(32'h37f6374b),
	.w4(32'h383abd88),
	.w5(32'h38d5c8d5),
	.w6(32'h37442bfb),
	.w7(32'h378b6391),
	.w8(32'h38357b77),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc05e0),
	.w1(32'hb8b70566),
	.w2(32'hb91087f6),
	.w3(32'h36b0fd31),
	.w4(32'hb8834c2a),
	.w5(32'hb8e4332d),
	.w6(32'h38365bde),
	.w7(32'hb894c7b5),
	.w8(32'hb96e3850),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904d4f1),
	.w1(32'h3985902f),
	.w2(32'h3927a2de),
	.w3(32'h397ae843),
	.w4(32'h397a19b0),
	.w5(32'hb76b402a),
	.w6(32'h3885d3c6),
	.w7(32'h36e0bec3),
	.w8(32'hb8cff075),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37079489),
	.w1(32'h38da0319),
	.w2(32'h389b9146),
	.w3(32'h389ce3b2),
	.w4(32'h38e20957),
	.w5(32'h3891b93e),
	.w6(32'h38036077),
	.w7(32'hb80a6725),
	.w8(32'hb7f14344),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79183ff),
	.w1(32'h38d1fe22),
	.w2(32'h3814e6ee),
	.w3(32'h381ab8ae),
	.w4(32'h38c1cf7a),
	.w5(32'h38a5c5d9),
	.w6(32'h3858cb15),
	.w7(32'hb8623391),
	.w8(32'h377612a4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71efc63),
	.w1(32'h37151cde),
	.w2(32'h3689f48e),
	.w3(32'hb7b12a0c),
	.w4(32'hb8450029),
	.w5(32'hb868c855),
	.w6(32'hb86954a2),
	.w7(32'hb85f3d69),
	.w8(32'hb8899497),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373a210e),
	.w1(32'h390fc5e5),
	.w2(32'h391ff9cc),
	.w3(32'h38c21da1),
	.w4(32'h391e87a6),
	.w5(32'h390d14f2),
	.w6(32'hb702262e),
	.w7(32'hb80a555c),
	.w8(32'hb788a9ba),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387a63e9),
	.w1(32'h38907089),
	.w2(32'h379a8b84),
	.w3(32'h3888b0b5),
	.w4(32'h38a10f55),
	.w5(32'h3652afef),
	.w6(32'h388105e7),
	.w7(32'h380d61a3),
	.w8(32'hb81cb494),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a5c900),
	.w1(32'hb72e7e2f),
	.w2(32'h37424bc5),
	.w3(32'h372cdae5),
	.w4(32'hb7395e23),
	.w5(32'h372a2606),
	.w6(32'hb52505d3),
	.w7(32'h37a02639),
	.w8(32'hb7488c01),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb743033d),
	.w1(32'hb73ce626),
	.w2(32'h36f47301),
	.w3(32'hb6df06a4),
	.w4(32'hb73c7c31),
	.w5(32'h370552f1),
	.w6(32'hb642a982),
	.w7(32'h3705ce31),
	.w8(32'hb5e4f370),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7109b29),
	.w1(32'hb71dce0d),
	.w2(32'h36c01305),
	.w3(32'hb6667340),
	.w4(32'hb730c75f),
	.w5(32'h36d68503),
	.w6(32'h34e00fea),
	.w7(32'h373b2d19),
	.w8(32'hb5e115f7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6feceb4),
	.w1(32'hb6818966),
	.w2(32'hb6b58743),
	.w3(32'hb6dfebbc),
	.w4(32'hb652bc97),
	.w5(32'hb7332b23),
	.w6(32'h3648e742),
	.w7(32'hb3896d54),
	.w8(32'hb64a5d2f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388fd901),
	.w1(32'h376566be),
	.w2(32'hb79cdc41),
	.w3(32'h38bf8645),
	.w4(32'h3789b6d0),
	.w5(32'hb81d3c44),
	.w6(32'h381520a9),
	.w7(32'h378534ba),
	.w8(32'hb8747724),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37927b4a),
	.w1(32'h374acf24),
	.w2(32'h37df080c),
	.w3(32'h3793f24f),
	.w4(32'h37a08aa7),
	.w5(32'h380b3b79),
	.w6(32'h37427469),
	.w7(32'h37f39e86),
	.w8(32'hb5d7c349),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82195fc),
	.w1(32'hb811c02d),
	.w2(32'hb8104e96),
	.w3(32'hb821c941),
	.w4(32'hb82aeb77),
	.w5(32'hb818c353),
	.w6(32'hb899b3f6),
	.w7(32'hb8c7e5f8),
	.w8(32'hb8bf6ae2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a2968),
	.w1(32'h390a7a6e),
	.w2(32'h38e609dd),
	.w3(32'h39298275),
	.w4(32'h391c7f58),
	.w5(32'h38cfec30),
	.w6(32'h39194e00),
	.w7(32'h3908b14f),
	.w8(32'h388202d4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb716786c),
	.w1(32'h3783a944),
	.w2(32'h36bcdbf3),
	.w3(32'hb6edeaf3),
	.w4(32'h37420c96),
	.w5(32'hb69f2b81),
	.w6(32'h37aeb1a7),
	.w7(32'h3789873a),
	.w8(32'h36e8566a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3683494f),
	.w1(32'hb7871412),
	.w2(32'h36d58f22),
	.w3(32'h374374d1),
	.w4(32'hb788bd8a),
	.w5(32'h376e6fa1),
	.w6(32'hb6f18779),
	.w7(32'h37877fdd),
	.w8(32'hb71f438d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70d21cb),
	.w1(32'hb7b30645),
	.w2(32'h37d64900),
	.w3(32'h36b14eae),
	.w4(32'hb73035b7),
	.w5(32'h37fbcd2a),
	.w6(32'hb766db17),
	.w7(32'h37b8ddb4),
	.w8(32'hb5b9941b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e56cdd),
	.w1(32'hb9a8bf85),
	.w2(32'hb990bd4b),
	.w3(32'h37e4f5ae),
	.w4(32'hb91f02fc),
	.w5(32'hb98a4e0e),
	.w6(32'hb9594da6),
	.w7(32'hb807c17f),
	.w8(32'hb9777f49),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c23c6),
	.w1(32'hb7889721),
	.w2(32'hb95cfb5e),
	.w3(32'hb9746356),
	.w4(32'hb8cfdcb0),
	.w5(32'hb9dcc28d),
	.w6(32'hb7796d3b),
	.w7(32'hb87286f9),
	.w8(32'hb99639d8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4c36b),
	.w1(32'h38ea9c08),
	.w2(32'hb9d62b52),
	.w3(32'hb9d0db2c),
	.w4(32'h3992fb26),
	.w5(32'hb932f717),
	.w6(32'h3958bab5),
	.w7(32'h39a02129),
	.w8(32'hba095f77),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fad37),
	.w1(32'h398ad6da),
	.w2(32'h39a2ea79),
	.w3(32'hbaab5727),
	.w4(32'h38e43176),
	.w5(32'h39aa28af),
	.w6(32'h39b730d1),
	.w7(32'h3998c070),
	.w8(32'h39a5d411),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a912b2),
	.w1(32'hb96a4a28),
	.w2(32'hb90d4855),
	.w3(32'h398dd386),
	.w4(32'h375b86e9),
	.w5(32'hb82d7718),
	.w6(32'hb91d8900),
	.w7(32'hb90f6ef6),
	.w8(32'hb943b265),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9007e0b),
	.w1(32'h3a3bf67d),
	.w2(32'h396fa13c),
	.w3(32'hb928dc19),
	.w4(32'h39b89a97),
	.w5(32'hb90e3ad9),
	.w6(32'h38b3eb4f),
	.w7(32'h38d1f411),
	.w8(32'h3a123312),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972e321),
	.w1(32'h3a5bddc9),
	.w2(32'h389097eb),
	.w3(32'hb940df8f),
	.w4(32'h3a8f6849),
	.w5(32'h390dcc4e),
	.w6(32'h3983f626),
	.w7(32'h397c44e1),
	.w8(32'h3a47289a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a533a03),
	.w1(32'hb827cb41),
	.w2(32'hb8ad5b5e),
	.w3(32'h3986cd09),
	.w4(32'h38d7130d),
	.w5(32'hb906e1db),
	.w6(32'hb808dc55),
	.w7(32'h37b6fc08),
	.w8(32'hb97d1e87),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93942bb),
	.w1(32'h399e1e37),
	.w2(32'h39a96e7f),
	.w3(32'hb9ab8b74),
	.w4(32'h39ad957d),
	.w5(32'h39d00ab7),
	.w6(32'h39c8aa37),
	.w7(32'h39b13e15),
	.w8(32'h39bd46eb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39466f),
	.w1(32'hb9f826f3),
	.w2(32'hba089ee3),
	.w3(32'h3a196da0),
	.w4(32'hb9bbec9f),
	.w5(32'hba1db551),
	.w6(32'hb9d145a6),
	.w7(32'hb9d82bae),
	.w8(32'hba043562),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a369e),
	.w1(32'h388f0fec),
	.w2(32'h38f43a4c),
	.w3(32'hba0d3adf),
	.w4(32'h38327060),
	.w5(32'hb755dd2e),
	.w6(32'h39248dcc),
	.w7(32'h396d3a34),
	.w8(32'hb8aa73f4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb775508b),
	.w1(32'h3a3a65cb),
	.w2(32'h3a0b51e3),
	.w3(32'hb92d1ecc),
	.w4(32'h39d66718),
	.w5(32'h3a1bbc17),
	.w6(32'h3a112f95),
	.w7(32'h3a02086e),
	.w8(32'h3a441c42),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a460e61),
	.w1(32'hb9e419c4),
	.w2(32'hb96646c7),
	.w3(32'h3a4d4365),
	.w4(32'hb83569a9),
	.w5(32'h3881e28e),
	.w6(32'hb962d89c),
	.w7(32'hb9562779),
	.w8(32'hb9821cce),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2444a0),
	.w1(32'hb8f25814),
	.w2(32'hb8e215a1),
	.w3(32'hba011b62),
	.w4(32'hb993dc33),
	.w5(32'hba47ab4d),
	.w6(32'h39854564),
	.w7(32'h3a13077f),
	.w8(32'h39da9cc4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d8fc0),
	.w1(32'hb9ab69e9),
	.w2(32'hb9d5cd2e),
	.w3(32'hb9319f85),
	.w4(32'hb96948d7),
	.w5(32'hb901fd14),
	.w6(32'hb9028f10),
	.w7(32'hb9268907),
	.w8(32'hb9a7ac3b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92aff39),
	.w1(32'hbaa36bb5),
	.w2(32'hba8a541d),
	.w3(32'h393a3a37),
	.w4(32'hba8e41a8),
	.w5(32'hba8034bf),
	.w6(32'hbab61ea0),
	.w7(32'hbaba3695),
	.w8(32'hba825dc8),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89b459),
	.w1(32'h38474cd3),
	.w2(32'hb8f9ccad),
	.w3(32'hba803987),
	.w4(32'h39c20878),
	.w5(32'hba353c7f),
	.w6(32'hb9a50858),
	.w7(32'h398f5e90),
	.w8(32'h3a4bf49e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39dfd4),
	.w1(32'h3928ff03),
	.w2(32'h38d86ae3),
	.w3(32'hba5597d1),
	.w4(32'h388032fa),
	.w5(32'hb9339b1a),
	.w6(32'h399482cf),
	.w7(32'h399510b8),
	.w8(32'h36ad1000),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8334925),
	.w1(32'hba172b52),
	.w2(32'hba029015),
	.w3(32'hb9444a89),
	.w4(32'hb9151ac4),
	.w5(32'h38f7fad0),
	.w6(32'hba205ebd),
	.w7(32'hb9d6655c),
	.w8(32'hb9230b7c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fc2d9),
	.w1(32'h39e9d126),
	.w2(32'h3a344794),
	.w3(32'h3999d1ef),
	.w4(32'h3a0efa1a),
	.w5(32'h3a412420),
	.w6(32'h39b8714f),
	.w7(32'h39fc9e11),
	.w8(32'h3a58de93),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dee4b),
	.w1(32'h3917bb8d),
	.w2(32'h396b0862),
	.w3(32'h3a5e0fae),
	.w4(32'h38f3bf00),
	.w5(32'h38d74e19),
	.w6(32'h383c08b8),
	.w7(32'h39079cae),
	.w8(32'h38a8a32d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39679bdd),
	.w1(32'h38a29621),
	.w2(32'h38186845),
	.w3(32'h3904b5a7),
	.w4(32'h389e15ef),
	.w5(32'hb5537d36),
	.w6(32'h38b93645),
	.w7(32'h38fe749e),
	.w8(32'hb89ba2b0),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f15d3a),
	.w1(32'hba0e7512),
	.w2(32'hba5621ee),
	.w3(32'hb66561bf),
	.w4(32'hb9f1e932),
	.w5(32'hba36f8a9),
	.w6(32'h373bfe75),
	.w7(32'hb95cb6c2),
	.w8(32'hb9ef7a90),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba597331),
	.w1(32'hb9ad1b95),
	.w2(32'hb9b1693f),
	.w3(32'hba255b18),
	.w4(32'h37e76850),
	.w5(32'h3a5ae445),
	.w6(32'hb9e83247),
	.w7(32'hb978fb61),
	.w8(32'hba3b329c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93b8e4),
	.w1(32'hba0863aa),
	.w2(32'h3988d0e9),
	.w3(32'h39df2cb0),
	.w4(32'h38193dec),
	.w5(32'h38f99334),
	.w6(32'hba0869dc),
	.w7(32'hb9351e27),
	.w8(32'hba00def3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8acf981),
	.w1(32'hb9a56457),
	.w2(32'hb9b77203),
	.w3(32'h3985701e),
	.w4(32'hb9a33dfc),
	.w5(32'hba10bfc3),
	.w6(32'hb980ce0a),
	.w7(32'hb99792fa),
	.w8(32'hb9dd971c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb948f),
	.w1(32'h38726493),
	.w2(32'hb7b16bf3),
	.w3(32'hb9ed67d8),
	.w4(32'h393b758f),
	.w5(32'h381a4f3c),
	.w6(32'hb8b673eb),
	.w7(32'h394f36f0),
	.w8(32'h39614fe6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38800650),
	.w1(32'hb89adb74),
	.w2(32'h39fc1921),
	.w3(32'h387bba2f),
	.w4(32'h39d6f3b1),
	.w5(32'h3a13e8e2),
	.w6(32'hba020500),
	.w7(32'hb9813db0),
	.w8(32'h3889f1b5),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990530c),
	.w1(32'hb90961e0),
	.w2(32'hb9eee2d5),
	.w3(32'h3842c7f3),
	.w4(32'hb7970458),
	.w5(32'hb955aed8),
	.w6(32'hb9760d2f),
	.w7(32'hb74da7c4),
	.w8(32'hb92c70c0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fdfd26),
	.w1(32'h39dd5a4d),
	.w2(32'h38e8a0d6),
	.w3(32'h38ec7a93),
	.w4(32'h39a09311),
	.w5(32'hb932e2a8),
	.w6(32'hb85083db),
	.w7(32'h39183c12),
	.w8(32'hb9033e97),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d53d52),
	.w1(32'hba832794),
	.w2(32'hb99f3801),
	.w3(32'hb99dc59d),
	.w4(32'hba29bbe2),
	.w5(32'h39a8966a),
	.w6(32'hba48d3b0),
	.w7(32'hb89025b8),
	.w8(32'hb8e454d0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9943e62),
	.w1(32'hb9af3a9e),
	.w2(32'hb9852d35),
	.w3(32'h3932f551),
	.w4(32'hb9d54754),
	.w5(32'hb8a45faa),
	.w6(32'hb93f1de0),
	.w7(32'hb970d331),
	.w8(32'h388c3192),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb878d951),
	.w1(32'hb996e2db),
	.w2(32'hba0a05bd),
	.w3(32'hb8329762),
	.w4(32'hb9938cdf),
	.w5(32'hb9f17bb6),
	.w6(32'h380c58a2),
	.w7(32'hb9178fd8),
	.w8(32'hb9cc7aba),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba114895),
	.w1(32'hb9806647),
	.w2(32'hb9889992),
	.w3(32'hb9fa4c93),
	.w4(32'hb89062f2),
	.w5(32'hb90b4d6b),
	.w6(32'hb9791428),
	.w7(32'hb9734882),
	.w8(32'hb9bc51bc),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7a4c7),
	.w1(32'h389bcdc3),
	.w2(32'hb972afdc),
	.w3(32'hb9481ad8),
	.w4(32'h39a37b11),
	.w5(32'h389b5aed),
	.w6(32'hb8c33761),
	.w7(32'hb9d013be),
	.w8(32'hb94cb8ec),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a633cf1),
	.w1(32'hb9536af4),
	.w2(32'hb94059a4),
	.w3(32'h39b8afa9),
	.w4(32'hb70a59ff),
	.w5(32'hb923e3ea),
	.w6(32'hb9911350),
	.w7(32'hb9b556ad),
	.w8(32'hba7b0930),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1e279),
	.w1(32'h3a461e4b),
	.w2(32'h3a0ed12f),
	.w3(32'hb99567ba),
	.w4(32'h3a1164ec),
	.w5(32'h39f15191),
	.w6(32'h3a938508),
	.w7(32'h3a84138f),
	.w8(32'h3a5bf3b0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06760c),
	.w1(32'hb989cf64),
	.w2(32'hb9d285cb),
	.w3(32'h39edf185),
	.w4(32'hb89ccc28),
	.w5(32'hb94ab087),
	.w6(32'hb815bea6),
	.w7(32'hb7ccf8fa),
	.w8(32'hb9853ec3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c635c3),
	.w1(32'h393f7137),
	.w2(32'h394b4c1b),
	.w3(32'hb92b5a9a),
	.w4(32'h391fbcd5),
	.w5(32'h3947fe36),
	.w6(32'h3936c603),
	.w7(32'h3925941f),
	.w8(32'h397a425a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ad473),
	.w1(32'h399b1156),
	.w2(32'h39ed8663),
	.w3(32'h3921df76),
	.w4(32'h39daf608),
	.w5(32'h3a19c918),
	.w6(32'h39cc9cc7),
	.w7(32'h39f9d960),
	.w8(32'h3a27fd84),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a334ac5),
	.w1(32'hb72b108d),
	.w2(32'hb9401bda),
	.w3(32'h3a1e2e33),
	.w4(32'hb8b42d57),
	.w5(32'hb9d2141e),
	.w6(32'h38849e9e),
	.w7(32'hb58c2c5a),
	.w8(32'hb93b4e3a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac1fd4),
	.w1(32'h39868be9),
	.w2(32'h3989d647),
	.w3(32'hb9e959f0),
	.w4(32'h3926250f),
	.w5(32'h38f05fca),
	.w6(32'h386a62c5),
	.w7(32'h38e38f08),
	.w8(32'h38dd8130),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397daae5),
	.w1(32'hb947543c),
	.w2(32'hb9a3a397),
	.w3(32'h39171bd9),
	.w4(32'hb99ff007),
	.w5(32'hb8fbe879),
	.w6(32'h3854ce69),
	.w7(32'hb6a7a364),
	.w8(32'hb8d68616),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a3999),
	.w1(32'hba29f8e1),
	.w2(32'hba3dd0f2),
	.w3(32'hb97d046b),
	.w4(32'hba22c527),
	.w5(32'hba52510d),
	.w6(32'hb9a21cfd),
	.w7(32'hba135de5),
	.w8(32'hba293468),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e08f6),
	.w1(32'hb9bb5b1f),
	.w2(32'hb914bf45),
	.w3(32'hba563992),
	.w4(32'h37fb8e73),
	.w5(32'h3958ea1b),
	.w6(32'hb9a6648a),
	.w7(32'hb99d8f3a),
	.w8(32'hb98909d9),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f5b96),
	.w1(32'h3a5e887d),
	.w2(32'h3a3c1332),
	.w3(32'hb8e6d771),
	.w4(32'h39dbde16),
	.w5(32'h3a31ddfb),
	.w6(32'h3a5639f7),
	.w7(32'h3a3fc8dd),
	.w8(32'h3aa8f889),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab69707),
	.w1(32'h3992dd9c),
	.w2(32'h388b6551),
	.w3(32'h3a8a7850),
	.w4(32'h39ba4fcf),
	.w5(32'h398f9570),
	.w6(32'h38a3f189),
	.w7(32'hb909222e),
	.w8(32'h3959fe73),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936b4a1),
	.w1(32'hb6d62e43),
	.w2(32'hb8c45e94),
	.w3(32'h397dfcc7),
	.w4(32'h38c90449),
	.w5(32'h39a5359f),
	.w6(32'h398d3182),
	.w7(32'h39c0c674),
	.w8(32'h37479908),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fdd757),
	.w1(32'h3a8bed78),
	.w2(32'h3a7bc8b1),
	.w3(32'h39a05f09),
	.w4(32'h3a038db9),
	.w5(32'hba2ad55f),
	.w6(32'h3a304f9d),
	.w7(32'h3a2c0c5f),
	.w8(32'h3a40ddac),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b56a99),
	.w1(32'hba8a4ae8),
	.w2(32'hb7cbea69),
	.w3(32'hb9854718),
	.w4(32'hba0ca08a),
	.w5(32'h39e84c64),
	.w6(32'hba896855),
	.w7(32'hb98845e1),
	.w8(32'hba085d7f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a296c2),
	.w1(32'hb990b405),
	.w2(32'hb8b10d51),
	.w3(32'h36b5721b),
	.w4(32'hb7fbd466),
	.w5(32'h39368b85),
	.w6(32'hb9e99148),
	.w7(32'hb9912a73),
	.w8(32'hb99abe8f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8959ce9),
	.w1(32'hba2abcf3),
	.w2(32'hba3bd2fe),
	.w3(32'h38bcf9de),
	.w4(32'hba1e2213),
	.w5(32'hba4e6cb6),
	.w6(32'hba1a0262),
	.w7(32'hba31d070),
	.w8(32'hba1c8c50),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ab634),
	.w1(32'h3913b164),
	.w2(32'h399db1d8),
	.w3(32'hba44ed9d),
	.w4(32'h3815bf75),
	.w5(32'h38968802),
	.w6(32'hb97a4637),
	.w7(32'h392c7014),
	.w8(32'h39f6859f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938820b),
	.w1(32'h3a3f534b),
	.w2(32'h3a37f339),
	.w3(32'hb829fe7a),
	.w4(32'hb981f582),
	.w5(32'hba342d10),
	.w6(32'h3a9a3c1a),
	.w7(32'h3a8b6b2d),
	.w8(32'h38b9c467),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382cd0bf),
	.w1(32'h393c3e6b),
	.w2(32'hb93756c8),
	.w3(32'hb9eeb6b9),
	.w4(32'hb8d560d3),
	.w5(32'hba12176f),
	.w6(32'h3981815c),
	.w7(32'h3984cc45),
	.w8(32'hb955bc12),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4cc28),
	.w1(32'h39b10cbb),
	.w2(32'hba0af7e0),
	.w3(32'hba35b406),
	.w4(32'h39ed067f),
	.w5(32'h3949109e),
	.w6(32'h39e81002),
	.w7(32'h39a312fa),
	.w8(32'h3991c2fc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2967bb),
	.w1(32'hb77c920e),
	.w2(32'h385bc26b),
	.w3(32'h3a351526),
	.w4(32'h38914166),
	.w5(32'h39680372),
	.w6(32'h389672ea),
	.w7(32'h3771a336),
	.w8(32'h399cd7ed),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caf9f6),
	.w1(32'hb9f3eb0c),
	.w2(32'hb983434d),
	.w3(32'h39e9ff11),
	.w4(32'hba1d6f3e),
	.w5(32'hb9883725),
	.w6(32'hb98418cc),
	.w7(32'h39057b3b),
	.w8(32'hb841aaec),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcf8aa),
	.w1(32'hba1e5487),
	.w2(32'hb9ae533c),
	.w3(32'hb9c4cb4a),
	.w4(32'hb969fa04),
	.w5(32'hb8fc64ca),
	.w6(32'hba5bc612),
	.w7(32'hba2bb5a1),
	.w8(32'hb9fe4975),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c7cab),
	.w1(32'h3a1430c8),
	.w2(32'h39231317),
	.w3(32'h38ceb8fc),
	.w4(32'h3a0d4363),
	.w5(32'h395b1810),
	.w6(32'h38add87f),
	.w7(32'h3a05cfb7),
	.w8(32'h3a97286a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5606a5),
	.w1(32'h39b3ee24),
	.w2(32'h39a27537),
	.w3(32'hb84870fd),
	.w4(32'h39944ffa),
	.w5(32'h398e20c7),
	.w6(32'h398edc92),
	.w7(32'h3901e432),
	.w8(32'h392920e7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992bbfd),
	.w1(32'hb8b76b3f),
	.w2(32'hb9b4ae64),
	.w3(32'h38e174b8),
	.w4(32'hb90e4632),
	.w5(32'hba1c7d2a),
	.w6(32'h37ef00c8),
	.w7(32'hb90b0f9b),
	.w8(32'hba0d4598),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954b262),
	.w1(32'h3926aeea),
	.w2(32'h39821f6d),
	.w3(32'hb981faf7),
	.w4(32'h397d88ff),
	.w5(32'h38b7fa89),
	.w6(32'h3766e8f6),
	.w7(32'h39141e93),
	.w8(32'h37dd1a52),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9085dba),
	.w1(32'hb9a3068f),
	.w2(32'hb9c209f8),
	.w3(32'hb975ec25),
	.w4(32'hb9b22574),
	.w5(32'hb9c7aa3e),
	.w6(32'hb97c9f7f),
	.w7(32'hb963795f),
	.w8(32'hb9d557ac),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a0186),
	.w1(32'h39728e4a),
	.w2(32'hb954dc28),
	.w3(32'hba0fe019),
	.w4(32'hb8cb442e),
	.w5(32'hb90f3839),
	.w6(32'h388f048c),
	.w7(32'hb9892aa3),
	.w8(32'hb938f612),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0be8a),
	.w1(32'h3a2a18fe),
	.w2(32'h3a124667),
	.w3(32'hb9a18e8d),
	.w4(32'h39b93d33),
	.w5(32'h3a042461),
	.w6(32'h3a20bf97),
	.w7(32'h3a0edbb0),
	.w8(32'h3a68c5a5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6873e7),
	.w1(32'hb7182a34),
	.w2(32'h39842dbe),
	.w3(32'h3a395189),
	.w4(32'h390da73d),
	.w5(32'h39b5d73d),
	.w6(32'hb760583f),
	.w7(32'h38028913),
	.w8(32'h398380b5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6129b),
	.w1(32'h38995837),
	.w2(32'h39aa4662),
	.w3(32'h39628380),
	.w4(32'hb6d5b4c8),
	.w5(32'h3a08c2d4),
	.w6(32'hb8f242e0),
	.w7(32'h3a106ed4),
	.w8(32'h3a11adf0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a232ac8),
	.w1(32'hb993ff4f),
	.w2(32'hb967d62b),
	.w3(32'h39de1f4a),
	.w4(32'hba337c81),
	.w5(32'hba1a8834),
	.w6(32'h38d7487d),
	.w7(32'hb8c2fb11),
	.w8(32'hb917a34b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d1394),
	.w1(32'hb9a21cb5),
	.w2(32'hb9030a84),
	.w3(32'hb9b0ce57),
	.w4(32'hb96a6b64),
	.w5(32'hb8caf32b),
	.w6(32'h3724e55b),
	.w7(32'h3993a049),
	.w8(32'h387ae3ea),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9152410),
	.w1(32'h38c474ce),
	.w2(32'hb943df41),
	.w3(32'hb85b59e2),
	.w4(32'hb838c194),
	.w5(32'hb9fc2c93),
	.w6(32'h39dcdc5a),
	.w7(32'h392786e8),
	.w8(32'hb933abcf),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f58c7),
	.w1(32'h39535380),
	.w2(32'h3988d9d1),
	.w3(32'hb9b5afa5),
	.w4(32'h390480fb),
	.w5(32'h39bb4eb6),
	.w6(32'hb99b327f),
	.w7(32'h39c7ccf8),
	.w8(32'h3a422343),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b66362),
	.w1(32'h39d90c7b),
	.w2(32'h3a17ff78),
	.w3(32'h39881eb4),
	.w4(32'h39d007ab),
	.w5(32'h3a0a8bb7),
	.w6(32'h39bea16c),
	.w7(32'h39e47d6c),
	.w8(32'h3a055187),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2366c8),
	.w1(32'hb7e4297a),
	.w2(32'hb9796af7),
	.w3(32'h39ef112b),
	.w4(32'hb92a88dc),
	.w5(32'hb9d2010f),
	.w6(32'h391242fc),
	.w7(32'h37c79a51),
	.w8(32'hb93f5e09),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b983c),
	.w1(32'hb856b4ca),
	.w2(32'hb90610e9),
	.w3(32'hb9b2962e),
	.w4(32'hb8f052bc),
	.w5(32'hb9c92f2b),
	.w6(32'h38986039),
	.w7(32'hb799e8fb),
	.w8(32'hb94f15ab),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983164b),
	.w1(32'hb9eed4ee),
	.w2(32'hba17c353),
	.w3(32'hb9a6df39),
	.w4(32'hb92a78d2),
	.w5(32'hb98a662d),
	.w6(32'hb9672cf8),
	.w7(32'hb99deb16),
	.w8(32'hb9fb3ae8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1462b4),
	.w1(32'h3933e41c),
	.w2(32'h3926751d),
	.w3(32'hb97cac4a),
	.w4(32'h38345172),
	.w5(32'hb87e5c7f),
	.w6(32'h37a6bf87),
	.w7(32'h3905a33a),
	.w8(32'hb8372a59),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3751fd9a),
	.w1(32'hb9a3cf52),
	.w2(32'hb899df12),
	.w3(32'hb92ccab0),
	.w4(32'hba78d507),
	.w5(32'hba8b797f),
	.w6(32'h3a15bffd),
	.w7(32'hb91f6199),
	.w8(32'hb89a888f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e503f6),
	.w1(32'hba0364d8),
	.w2(32'hba124807),
	.w3(32'h39558db0),
	.w4(32'hb9f836fa),
	.w5(32'hba305506),
	.w6(32'hba201e2b),
	.w7(32'hba055e61),
	.w8(32'hba0215e7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0326ba),
	.w1(32'hb8110c91),
	.w2(32'hb98aea41),
	.w3(32'hba090329),
	.w4(32'hb97a8c25),
	.w5(32'hb9fc705e),
	.w6(32'hb86ba8e2),
	.w7(32'hb9f07b21),
	.w8(32'hb9812587),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f93218),
	.w1(32'h3854f8be),
	.w2(32'h39d31c03),
	.w3(32'hb9907cef),
	.w4(32'h39a27f28),
	.w5(32'h3a107d09),
	.w6(32'hb98a8136),
	.w7(32'hb90ad393),
	.w8(32'h38ffbd52),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a278eb8),
	.w1(32'hb9b54c80),
	.w2(32'hba26d7af),
	.w3(32'h3a23c089),
	.w4(32'hb92a9e97),
	.w5(32'hba04e643),
	.w6(32'h38ca8e18),
	.w7(32'hb8961026),
	.w8(32'hba0652b3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba235f60),
	.w1(32'hb9af2e86),
	.w2(32'hb9aff7f6),
	.w3(32'hba05819b),
	.w4(32'hba0e1597),
	.w5(32'hba1022a0),
	.w6(32'h390514a3),
	.w7(32'h3965c66e),
	.w8(32'hb98c25eb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e021f1),
	.w1(32'hb9b7cf60),
	.w2(32'hba07bd5a),
	.w3(32'hb9fcd213),
	.w4(32'hba02b161),
	.w5(32'hba434aa0),
	.w6(32'hb93817ff),
	.w7(32'hba12fcc2),
	.w8(32'hba2cb016),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4071c2),
	.w1(32'hb9839a77),
	.w2(32'hb8a59b70),
	.w3(32'hba7f44f8),
	.w4(32'hb94264c9),
	.w5(32'h363ee180),
	.w6(32'hb9929629),
	.w7(32'hb93d021d),
	.w8(32'hb9511d4c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a6f7b5),
	.w1(32'h3785ff01),
	.w2(32'hb7ca56a9),
	.w3(32'h385f38c5),
	.w4(32'hb8a1b8d8),
	.w5(32'hb8045d42),
	.w6(32'h3924bb06),
	.w7(32'hb91c43c2),
	.w8(32'hb9817651),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb792c457),
	.w1(32'hba42cd7f),
	.w2(32'hb7d0091b),
	.w3(32'hb89ae13c),
	.w4(32'hb9f5cc51),
	.w5(32'h3851fcd4),
	.w6(32'hb9e86123),
	.w7(32'hb93bd057),
	.w8(32'hba3ac63e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34e43f94),
	.w1(32'hb985550a),
	.w2(32'hb92f3deb),
	.w3(32'h3952f50b),
	.w4(32'hb9e78136),
	.w5(32'hb9a62453),
	.w6(32'hb95fe989),
	.w7(32'hb96d357f),
	.w8(32'hb984d263),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c7954),
	.w1(32'hba58bed1),
	.w2(32'hb9c54014),
	.w3(32'hb968dfc8),
	.w4(32'hba2661bb),
	.w5(32'hb981d419),
	.w6(32'hba490319),
	.w7(32'hba410cd3),
	.w8(32'hb982605b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807e28f),
	.w1(32'hb9962c02),
	.w2(32'hba11eda4),
	.w3(32'h3912289c),
	.w4(32'hb95a2ae1),
	.w5(32'hb9cc9eab),
	.w6(32'h389cc902),
	.w7(32'hb9026c29),
	.w8(32'hb9b222aa),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba198efd),
	.w1(32'h381be26f),
	.w2(32'hb88233b4),
	.w3(32'hb9cd513c),
	.w4(32'h38abcbc7),
	.w5(32'h38e15383),
	.w6(32'h390fd14b),
	.w7(32'h344fe7b1),
	.w8(32'h395536c9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39293578),
	.w1(32'hb9850264),
	.w2(32'hb9f0b033),
	.w3(32'h3984402b),
	.w4(32'hb952b151),
	.w5(32'hb9fd9e74),
	.w6(32'h38935e3b),
	.w7(32'hb91310ba),
	.w8(32'hb9c81deb),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba308fdf),
	.w1(32'hb9bad3fc),
	.w2(32'hba15f0b3),
	.w3(32'hba2477ea),
	.w4(32'hb9c0c714),
	.w5(32'hba0177a5),
	.w6(32'hb981da87),
	.w7(32'hb9e06308),
	.w8(32'hba1a69df),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15db78),
	.w1(32'h394ccbea),
	.w2(32'h3982ed4c),
	.w3(32'hba050067),
	.w4(32'h39060f7f),
	.w5(32'h39a39ca3),
	.w6(32'h38ce4bc6),
	.w7(32'h394d8d5c),
	.w8(32'h39d126f9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a387dd1),
	.w1(32'h38aabeb5),
	.w2(32'h37172ed3),
	.w3(32'h3a1b9c6d),
	.w4(32'hb8ef4512),
	.w5(32'h374f6a44),
	.w6(32'h38c72d12),
	.w7(32'h37bac40e),
	.w8(32'h38658b30),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a872b7),
	.w1(32'hb9a0b19e),
	.w2(32'hb99f2f89),
	.w3(32'h37f9db7d),
	.w4(32'hb9e2aab1),
	.w5(32'hb9bae51c),
	.w6(32'hb87edcc2),
	.w7(32'h392f6986),
	.w8(32'hb897e99a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad5966),
	.w1(32'hb97479cb),
	.w2(32'hb74469e9),
	.w3(32'hb98216ae),
	.w4(32'h3885b34d),
	.w5(32'h38408afe),
	.w6(32'hb9860e7a),
	.w7(32'hb92fd7d6),
	.w8(32'hb925f105),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972063d),
	.w1(32'hb9c474e8),
	.w2(32'hba0d1428),
	.w3(32'hb95fa73c),
	.w4(32'hb9a40dc9),
	.w5(32'h38444ea9),
	.w6(32'h39189ff6),
	.w7(32'hb9a93e52),
	.w8(32'hba29cfe5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb6619),
	.w1(32'hb9bbb12d),
	.w2(32'h39de8b3b),
	.w3(32'h398503da),
	.w4(32'hb7bbd987),
	.w5(32'hb7ea11cb),
	.w6(32'hba10f8cb),
	.w7(32'hb9d7818f),
	.w8(32'hb5c4d113),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397adbd6),
	.w1(32'hb94cf2c9),
	.w2(32'hb9042b69),
	.w3(32'h392827a4),
	.w4(32'hb50d18aa),
	.w5(32'hb8ec8a80),
	.w6(32'hb8a81af1),
	.w7(32'h398653b9),
	.w8(32'hb93fe5b1),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ca58d),
	.w1(32'hb9616b8f),
	.w2(32'hb985bab2),
	.w3(32'hb980fdc7),
	.w4(32'hb9b98bef),
	.w5(32'hb9de4b7f),
	.w6(32'h390c5301),
	.w7(32'hb922310f),
	.w8(32'hb98fe86d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfb67a),
	.w1(32'h38b3e6ec),
	.w2(32'hb83ecdd1),
	.w3(32'hba0be47c),
	.w4(32'hb8b7b211),
	.w5(32'hb9103c94),
	.w6(32'h397176bb),
	.w7(32'h398a556c),
	.w8(32'h38e3247b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb836babe),
	.w1(32'h3a4253fd),
	.w2(32'h3a614804),
	.w3(32'hb880b9d5),
	.w4(32'h3a826478),
	.w5(32'h3a44fc9f),
	.w6(32'hb9363cbd),
	.w7(32'h3a4c8128),
	.w8(32'h3ad9c10f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4c2b2),
	.w1(32'h3973b82a),
	.w2(32'hba62c42a),
	.w3(32'h3a5dca6b),
	.w4(32'h38f7fdf0),
	.w5(32'hb9d05275),
	.w6(32'h3a70cdc9),
	.w7(32'h3a269083),
	.w8(32'hb96c1f8e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16ffc3),
	.w1(32'hba6d7a84),
	.w2(32'hba6a55b7),
	.w3(32'h3a232555),
	.w4(32'hba6952d0),
	.w5(32'hba896d97),
	.w6(32'hba92e84d),
	.w7(32'hba786df8),
	.w8(32'hba5f2969),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43df4d),
	.w1(32'hb7381520),
	.w2(32'hb944640c),
	.w3(32'hba49c7b6),
	.w4(32'hb898da41),
	.w5(32'hb9d3de51),
	.w6(32'hb7e3e982),
	.w7(32'h3859ab97),
	.w8(32'hb9073d33),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999f9e2),
	.w1(32'hb9d65bbd),
	.w2(32'hb9d5a38e),
	.w3(32'hb9eb0166),
	.w4(32'hb9d11bf6),
	.w5(32'hb9ff0983),
	.w6(32'hb9e90a66),
	.w7(32'hb9ba468f),
	.w8(32'hb99b0dc9),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2db02),
	.w1(32'hb8bf09ce),
	.w2(32'hb89f7023),
	.w3(32'hb9dfd445),
	.w4(32'hb7233f20),
	.w5(32'h378188da),
	.w6(32'hb9750035),
	.w7(32'hb912e162),
	.w8(32'hb968316f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f62c4),
	.w1(32'hb9afff26),
	.w2(32'hb9b5c52c),
	.w3(32'h378c3a5f),
	.w4(32'hb87f8fa3),
	.w5(32'hb966e53f),
	.w6(32'hb8b0f3b8),
	.w7(32'hb93d3bd5),
	.w8(32'hb991011a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1241a4),
	.w1(32'hba0a3de5),
	.w2(32'hba5c2036),
	.w3(32'hba0d4df3),
	.w4(32'hb9e34d7f),
	.w5(32'hba1f34c5),
	.w6(32'hb84bbd59),
	.w7(32'hb9b78690),
	.w8(32'hba235436),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76b15c),
	.w1(32'hb9f76134),
	.w2(32'hb9ec4546),
	.w3(32'hba2c9f50),
	.w4(32'hb9e51cc3),
	.w5(32'hba022ddb),
	.w6(32'hba10e183),
	.w7(32'hb9e20e58),
	.w8(32'hb9b67e0f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d377fc),
	.w1(32'h397d458b),
	.w2(32'h39b08b8b),
	.w3(32'hb9d0cab2),
	.w4(32'hb773ac82),
	.w5(32'h3844d108),
	.w6(32'h343d0ce8),
	.w7(32'hb92b4ac7),
	.w8(32'h399b5c31),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5c13a),
	.w1(32'h390f5b0c),
	.w2(32'hb8113f2b),
	.w3(32'h384884c0),
	.w4(32'hb6acd569),
	.w5(32'hb9d2d935),
	.w6(32'h3992bde8),
	.w7(32'h39af89f1),
	.w8(32'h37d0e5de),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a62e37),
	.w1(32'h39d292d7),
	.w2(32'hb9a8e1ef),
	.w3(32'hb9c0e70f),
	.w4(32'hb9ad90c3),
	.w5(32'hba42ca7e),
	.w6(32'h3a5b565b),
	.w7(32'hb933aeb9),
	.w8(32'hb8bf1acc),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92735b4),
	.w1(32'hb8e11b29),
	.w2(32'hb97b3041),
	.w3(32'hb9945984),
	.w4(32'hb82fd98f),
	.w5(32'hba00b871),
	.w6(32'hb7a9b80b),
	.w7(32'h3869308b),
	.w8(32'hb94652bd),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3ed32),
	.w1(32'hb8063468),
	.w2(32'hb938dd55),
	.w3(32'hba023c89),
	.w4(32'hb918efc6),
	.w5(32'hb9962f33),
	.w6(32'hb92ab485),
	.w7(32'hb919afa0),
	.w8(32'hb8d157a7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f7587),
	.w1(32'hba215c9a),
	.w2(32'hba22e2c9),
	.w3(32'hb9df9d33),
	.w4(32'hb9df5301),
	.w5(32'hb9ee4924),
	.w6(32'hba06c3c3),
	.w7(32'hba29d419),
	.w8(32'hba148015),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06c8c0),
	.w1(32'hba2a3f3c),
	.w2(32'hba22dba7),
	.w3(32'hb98fc688),
	.w4(32'hba214b8f),
	.w5(32'hba3c9d21),
	.w6(32'hba406ca9),
	.w7(32'hba19cff7),
	.w8(32'hb9f88029),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17e60f),
	.w1(32'hb982e77b),
	.w2(32'hb978d659),
	.w3(32'hba187598),
	.w4(32'hb90d5d8a),
	.w5(32'hb9a84ec0),
	.w6(32'hb96a8a7b),
	.w7(32'hb9366404),
	.w8(32'hb97bfeca),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986cd7b),
	.w1(32'hb9889566),
	.w2(32'hb9c8406d),
	.w3(32'hb9983e10),
	.w4(32'hb9649c22),
	.w5(32'hb9e17a34),
	.w6(32'hb94e0c05),
	.w7(32'hb95005ff),
	.w8(32'hb9872e83),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a462e5),
	.w1(32'hba2fe0c5),
	.w2(32'hba4d5f1a),
	.w3(32'hb9a081ca),
	.w4(32'hb7ce296c),
	.w5(32'h38a897d9),
	.w6(32'hb9fe8f69),
	.w7(32'hb9e3795d),
	.w8(32'hba49737c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa45580),
	.w1(32'h39bd1681),
	.w2(32'h3a307cc2),
	.w3(32'hb9907bb0),
	.w4(32'h39d4ab6c),
	.w5(32'h3a19fcee),
	.w6(32'h39778356),
	.w7(32'h39b1651e),
	.w8(32'h39d5e243),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a320ca1),
	.w1(32'h39039214),
	.w2(32'hb90ffa10),
	.w3(32'h398d53cf),
	.w4(32'hb82a88c3),
	.w5(32'hb9976ccb),
	.w6(32'h37e62ba4),
	.w7(32'h38f33ed8),
	.w8(32'hb90fa961),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20dbb7),
	.w1(32'h39b2b33b),
	.w2(32'hb95b865d),
	.w3(32'hba1fa865),
	.w4(32'h381fb1e5),
	.w5(32'hb986439d),
	.w6(32'h399f6ed2),
	.w7(32'h3927027c),
	.w8(32'hb9981a62),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9972166),
	.w1(32'hb98bd2a7),
	.w2(32'hb99f69e6),
	.w3(32'hb9e5f934),
	.w4(32'hb9a311f5),
	.w5(32'hba0bb763),
	.w6(32'hb8ec2079),
	.w7(32'hb92db60c),
	.w8(32'hb9a92434),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f759a4),
	.w1(32'h3a1b1fff),
	.w2(32'hb8bd14e8),
	.w3(32'hba0c935f),
	.w4(32'h3a590e97),
	.w5(32'h3a25c954),
	.w6(32'h3a6b8b5d),
	.w7(32'h3a8ae88b),
	.w8(32'hb8e4f263),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80acd4),
	.w1(32'hb8f4b4dc),
	.w2(32'hb9f885bf),
	.w3(32'h39fb3549),
	.w4(32'hb9928f5f),
	.w5(32'hba0af7b5),
	.w6(32'h385edc75),
	.w7(32'hb8c0e8de),
	.w8(32'hba0c07e2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06e5a9),
	.w1(32'hba0e3c17),
	.w2(32'hba5ebdf7),
	.w3(32'hba4bf00d),
	.w4(32'hba0369ae),
	.w5(32'hba2555e6),
	.w6(32'hb6dac392),
	.w7(32'hb9477d26),
	.w8(32'hba1b0736),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba566563),
	.w1(32'hb7545e5d),
	.w2(32'h38f939d0),
	.w3(32'hba12800f),
	.w4(32'h384e11e6),
	.w5(32'h3917b6f1),
	.w6(32'h3687126e),
	.w7(32'h387d83c0),
	.w8(32'hb65cb61a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7802f5e),
	.w1(32'h39279f69),
	.w2(32'h394ad8ee),
	.w3(32'hb707d68e),
	.w4(32'h38fa8b7b),
	.w5(32'h390c8671),
	.w6(32'h38bb2ffa),
	.w7(32'h38a6570c),
	.w8(32'h38b0c808),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule