module layer_8_featuremap_210(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4b573),
	.w1(32'hbb6b3dd2),
	.w2(32'hbb0dd9ab),
	.w3(32'hbc28cd51),
	.w4(32'h3b448b62),
	.w5(32'hbc35561b),
	.w6(32'h3a577cb5),
	.w7(32'hbbc4dc84),
	.w8(32'hbbd59e6b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe57e1),
	.w1(32'hb90945af),
	.w2(32'hbb47961b),
	.w3(32'hbba85f0f),
	.w4(32'h39c0e082),
	.w5(32'hbb086b06),
	.w6(32'hba2ab07f),
	.w7(32'h3ac07fdb),
	.w8(32'h3b837f42),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88abc89),
	.w1(32'h3c2e9fff),
	.w2(32'h3bdba521),
	.w3(32'hbaf4215e),
	.w4(32'h3c95705c),
	.w5(32'h3bcae395),
	.w6(32'hbab04043),
	.w7(32'hbbaec345),
	.w8(32'hbc910f75),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5375ac),
	.w1(32'h3beccf51),
	.w2(32'hbbc12c29),
	.w3(32'h3b8431d7),
	.w4(32'h3bafad99),
	.w5(32'h3c609d8e),
	.w6(32'hbc2bbc3a),
	.w7(32'hbb95e7b8),
	.w8(32'hbbff0919),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36d1cb),
	.w1(32'h3bdde120),
	.w2(32'h3be3a504),
	.w3(32'h3bd826b0),
	.w4(32'h3a38de76),
	.w5(32'h3a9281fe),
	.w6(32'h3b7ec7b3),
	.w7(32'h39cff2ac),
	.w8(32'hbb55bc4c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4554ee),
	.w1(32'hbc34bc03),
	.w2(32'hbc92592d),
	.w3(32'h3b001f38),
	.w4(32'hbbd33d13),
	.w5(32'hbc1f3cee),
	.w6(32'hbb80b826),
	.w7(32'hba042b65),
	.w8(32'hbb319782),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2b3cd),
	.w1(32'h3acc7274),
	.w2(32'h3a86a493),
	.w3(32'hbc27c3cd),
	.w4(32'hba788776),
	.w5(32'hb969717e),
	.w6(32'h3aebadd8),
	.w7(32'hbb467ea7),
	.w8(32'hbb497061),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b155c),
	.w1(32'hbb660e95),
	.w2(32'h3add1343),
	.w3(32'h3a51ff5e),
	.w4(32'hbb56c797),
	.w5(32'h3c6a11b5),
	.w6(32'hbc3b7c21),
	.w7(32'hbc848f71),
	.w8(32'hbb646066),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8df05),
	.w1(32'h3b57e981),
	.w2(32'h3c1be241),
	.w3(32'h3c0529aa),
	.w4(32'hbbe34a92),
	.w5(32'hb84784bb),
	.w6(32'h3a1611eb),
	.w7(32'hba9959e3),
	.w8(32'hbb956456),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab43a98),
	.w1(32'h3d18163e),
	.w2(32'h3cfb9972),
	.w3(32'hbae7774e),
	.w4(32'h3c9fd3ad),
	.w5(32'h3b36dc48),
	.w6(32'h3c213cd9),
	.w7(32'h3b19a450),
	.w8(32'hbb7dce19),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c597059),
	.w1(32'hbcb702c9),
	.w2(32'hbd010318),
	.w3(32'hbc05d2a1),
	.w4(32'h3c04d5e9),
	.w5(32'hbc827496),
	.w6(32'hbbdfc811),
	.w7(32'h3c07c11d),
	.w8(32'h3c2dcad0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc409f3c),
	.w1(32'h39dac49b),
	.w2(32'hbbb9dfaf),
	.w3(32'hbc07d600),
	.w4(32'h3bdea880),
	.w5(32'h3bd59316),
	.w6(32'hb92bc6b5),
	.w7(32'h3a62c406),
	.w8(32'h3c5e7924),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c003a98),
	.w1(32'h3a9aa2bb),
	.w2(32'hbc84fc33),
	.w3(32'h3b85f4c2),
	.w4(32'h3cb3017c),
	.w5(32'h3c766271),
	.w6(32'hbb8fac63),
	.w7(32'hbbcacf72),
	.w8(32'hbbb4e455),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd30fa2),
	.w1(32'h3c436fb6),
	.w2(32'h3c8d475c),
	.w3(32'hbbbe913e),
	.w4(32'h3bbab082),
	.w5(32'h3c6443a6),
	.w6(32'h3c890fd4),
	.w7(32'h3b317ee1),
	.w8(32'hbb49ad2f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59c1c4),
	.w1(32'hba8971ce),
	.w2(32'h3936e483),
	.w3(32'h3bca54b6),
	.w4(32'hbb115711),
	.w5(32'hbadd0e70),
	.w6(32'h3b100f98),
	.w7(32'hbb19a6e4),
	.w8(32'hbb8cc624),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06da84),
	.w1(32'h3c0987f3),
	.w2(32'hbacbb342),
	.w3(32'h39df5684),
	.w4(32'h3cac6a97),
	.w5(32'h39f7e8dd),
	.w6(32'h3bf0b5e1),
	.w7(32'h3b60fc50),
	.w8(32'h3be49efc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d1bc6),
	.w1(32'h3b13d99e),
	.w2(32'h3a65ca07),
	.w3(32'h3bc22d98),
	.w4(32'h3b8a32af),
	.w5(32'h3bd009e4),
	.w6(32'h3b1b54cc),
	.w7(32'h3c00ffba),
	.w8(32'h3c0cf5a3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8765c),
	.w1(32'hb984b725),
	.w2(32'hbc697df6),
	.w3(32'hbb51de9e),
	.w4(32'h3c1c98d5),
	.w5(32'hbb4ed03d),
	.w6(32'hbc01de2b),
	.w7(32'hbca43d6b),
	.w8(32'hbc86ef60),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f7692),
	.w1(32'h3b8670d8),
	.w2(32'hbca3df3e),
	.w3(32'hbc0834e5),
	.w4(32'h3ca51fde),
	.w5(32'h3ca0b99e),
	.w6(32'hbc140936),
	.w7(32'hbc8d36e3),
	.w8(32'hbc333973),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc979dee),
	.w1(32'h3b286685),
	.w2(32'h3b2ec70b),
	.w3(32'h3b816a55),
	.w4(32'hbac9fc09),
	.w5(32'hbac4f02e),
	.w6(32'h3b74a997),
	.w7(32'h3a79417e),
	.w8(32'hbb3534b4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ec1a4),
	.w1(32'h3c216944),
	.w2(32'h3c03ea96),
	.w3(32'h3b2d33f4),
	.w4(32'h3bc0fb19),
	.w5(32'h3ba767f8),
	.w6(32'h3c0288cc),
	.w7(32'h3bd5fc49),
	.w8(32'h3b4903c1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e9e46),
	.w1(32'h3a3b0fc9),
	.w2(32'hbb8bb805),
	.w3(32'h3a03a8fd),
	.w4(32'hb8cac185),
	.w5(32'hbb9811dc),
	.w6(32'hba63a006),
	.w7(32'h3b58529e),
	.w8(32'h3c24d561),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a153e),
	.w1(32'hba41c8c1),
	.w2(32'hbb50be57),
	.w3(32'hbb375bc9),
	.w4(32'h3b896b98),
	.w5(32'hbb3f1a95),
	.w6(32'h3b479752),
	.w7(32'hbbc7fce4),
	.w8(32'hbbb10158),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3944cf),
	.w1(32'hbae02739),
	.w2(32'h3b43fb2c),
	.w3(32'hbb80acaa),
	.w4(32'hbbddcfad),
	.w5(32'hbb9e8b54),
	.w6(32'h3b6c4ac5),
	.w7(32'h3c0080fc),
	.w8(32'h3b89350a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925037e),
	.w1(32'hbb1eb7d3),
	.w2(32'h3a9a160d),
	.w3(32'h3bf976fe),
	.w4(32'hb9f710f0),
	.w5(32'hbbae30c3),
	.w6(32'h3ba03f80),
	.w7(32'h3b5c001d),
	.w8(32'h3b122ee1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5d8f7),
	.w1(32'hbaad0a78),
	.w2(32'h395333c2),
	.w3(32'hba544a1d),
	.w4(32'hbbbe6e98),
	.w5(32'hbc20f315),
	.w6(32'hbb0f5e0d),
	.w7(32'h3b2f5f9a),
	.w8(32'h3bea253c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80c8e6),
	.w1(32'hbc065b6b),
	.w2(32'hbbee500a),
	.w3(32'h3b6a1c56),
	.w4(32'hbb6f766b),
	.w5(32'hbb685596),
	.w6(32'hbb21c9c9),
	.w7(32'h3b5cdd12),
	.w8(32'h3b36027d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4e7fe),
	.w1(32'h3c0c6d67),
	.w2(32'h3a110974),
	.w3(32'hbbf82e99),
	.w4(32'h3cb5725f),
	.w5(32'h3c8c78ea),
	.w6(32'hbc261a43),
	.w7(32'hbcb4e5b8),
	.w8(32'hbcdae1e9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc984e0c),
	.w1(32'h3aa176dc),
	.w2(32'hbc1b6e59),
	.w3(32'h3b918acd),
	.w4(32'h3ad94299),
	.w5(32'hbbba8719),
	.w6(32'h3b2a33c6),
	.w7(32'h39bcf6d6),
	.w8(32'hbb89dc49),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14501e),
	.w1(32'h3b05e6f5),
	.w2(32'h3ba95400),
	.w3(32'hbc33f330),
	.w4(32'hbbdfcd2b),
	.w5(32'hbc1a5205),
	.w6(32'hba8d5085),
	.w7(32'hbafb7d78),
	.w8(32'h3c822f21),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89855b),
	.w1(32'h3c0b5f95),
	.w2(32'h392db1ef),
	.w3(32'h3c01149d),
	.w4(32'h3bce9402),
	.w5(32'h3c962797),
	.w6(32'h3b300d3d),
	.w7(32'hbb8ade2c),
	.w8(32'hba404134),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc238d1e),
	.w1(32'hbcfde563),
	.w2(32'hbd01889c),
	.w3(32'h3c130450),
	.w4(32'hbbb10488),
	.w5(32'hbc97ad25),
	.w6(32'hbc3ca97c),
	.w7(32'h3be5c69c),
	.w8(32'h3ccced1f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56fb7b),
	.w1(32'h3b17376e),
	.w2(32'hbc247b6a),
	.w3(32'hbc8b3d55),
	.w4(32'hbb72392e),
	.w5(32'hbb898e26),
	.w6(32'h3b4894f4),
	.w7(32'hbaa24bdd),
	.w8(32'hbc02b16b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c8882),
	.w1(32'hbbe020b3),
	.w2(32'hbc821265),
	.w3(32'hba3273fb),
	.w4(32'hbbd19dee),
	.w5(32'hbc204562),
	.w6(32'hbad33263),
	.w7(32'hbb8c51cc),
	.w8(32'h3c19fed2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f69aa),
	.w1(32'hbb2dfa56),
	.w2(32'hbc251449),
	.w3(32'hbac3d78e),
	.w4(32'hb9cbedc4),
	.w5(32'hbaff9394),
	.w6(32'h3b7cab42),
	.w7(32'hb7c339ec),
	.w8(32'h3b9d07db),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4718b3),
	.w1(32'hbb4e2393),
	.w2(32'hbc7c2e44),
	.w3(32'hbab10759),
	.w4(32'h3c0e718b),
	.w5(32'h3b07b608),
	.w6(32'h3c249e87),
	.w7(32'hbb3e94ed),
	.w8(32'hbbb5e35f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b8d01),
	.w1(32'h3a32a531),
	.w2(32'h3c0c6391),
	.w3(32'h3c1f9650),
	.w4(32'hbbca6534),
	.w5(32'hbac3b1e4),
	.w6(32'h3c15f9f8),
	.w7(32'h3c67c139),
	.w8(32'h3c561373),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28b747),
	.w1(32'h3abf3b3f),
	.w2(32'h3b45ae43),
	.w3(32'h3ac21867),
	.w4(32'hbb1efdd3),
	.w5(32'h3a8145a3),
	.w6(32'hba928472),
	.w7(32'hbb7a041e),
	.w8(32'hbc05d616),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26122b),
	.w1(32'h3c423461),
	.w2(32'h3cc1de1b),
	.w3(32'hba1f9cba),
	.w4(32'h3c37de3e),
	.w5(32'h3c226d86),
	.w6(32'h3c3e1b46),
	.w7(32'h3c68416e),
	.w8(32'h3c0d3092),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932227),
	.w1(32'h3b88f9a6),
	.w2(32'h3baca95e),
	.w3(32'h3be0eb47),
	.w4(32'h3aecf356),
	.w5(32'h3a9f68cf),
	.w6(32'hbb9a5dae),
	.w7(32'h388a9b2f),
	.w8(32'h3a6eb9dc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb963c5),
	.w1(32'h3acad402),
	.w2(32'h3b98cfd7),
	.w3(32'h3bb9b1b4),
	.w4(32'h3b13a84e),
	.w5(32'h3babb563),
	.w6(32'h3ba70c85),
	.w7(32'h3bccd3db),
	.w8(32'h3b64641d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b855eaa),
	.w1(32'h3c4e18b7),
	.w2(32'hbb78e387),
	.w3(32'h3b3eafa6),
	.w4(32'h3c9b3a0f),
	.w5(32'h3c508f4b),
	.w6(32'hbb8f50a5),
	.w7(32'hbc6694e9),
	.w8(32'hbb6c5cde),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdd726),
	.w1(32'hbbd184db),
	.w2(32'h3b8b8453),
	.w3(32'h3c25e408),
	.w4(32'hbc304f1a),
	.w5(32'hbc2d94a0),
	.w6(32'h3b512cf0),
	.w7(32'h3c24ec06),
	.w8(32'h3c3b00cd),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ead1f),
	.w1(32'hbc7a1fd1),
	.w2(32'hbd048d24),
	.w3(32'hbb722e2a),
	.w4(32'hbbc804e6),
	.w5(32'hbc902591),
	.w6(32'hbc67da66),
	.w7(32'hbcac143b),
	.w8(32'hbc4e42ce),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb8378),
	.w1(32'hbba051f8),
	.w2(32'hbc215bc1),
	.w3(32'hbca56d2f),
	.w4(32'hbbed11dd),
	.w5(32'hbc665c1a),
	.w6(32'h39979fe4),
	.w7(32'hbc5baef9),
	.w8(32'h3a9f2dba),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b489704),
	.w1(32'h3b628794),
	.w2(32'h3a5a1c51),
	.w3(32'h3c3d6673),
	.w4(32'h3a158cde),
	.w5(32'hbb0bac7c),
	.w6(32'h3bbd54d0),
	.w7(32'h3b5a9b93),
	.w8(32'h3b596a61),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b8310),
	.w1(32'hbbc93ecd),
	.w2(32'hbbaf44a8),
	.w3(32'h3b01f6e7),
	.w4(32'h3b81b90d),
	.w5(32'hbaeb089e),
	.w6(32'hbaed4234),
	.w7(32'hbb2c0648),
	.w8(32'hbbfe8437),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d6549),
	.w1(32'hbc25c2a9),
	.w2(32'hbc9845dc),
	.w3(32'hbb7505d1),
	.w4(32'hbbc5fb91),
	.w5(32'hbc2207dd),
	.w6(32'hbb3e9511),
	.w7(32'hbb99daf8),
	.w8(32'hbb9cf506),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba637a2d),
	.w1(32'hbc30b05c),
	.w2(32'hbcc2fd2d),
	.w3(32'hbabcfd0b),
	.w4(32'hba77cb2c),
	.w5(32'hbc90ca16),
	.w6(32'hbb8d90c3),
	.w7(32'hbc0bdb73),
	.w8(32'hbbce8c9e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62c3e8),
	.w1(32'h3a1a400b),
	.w2(32'h3b0795aa),
	.w3(32'hbc0b7ab7),
	.w4(32'h3c0c225f),
	.w5(32'h3c4c8a20),
	.w6(32'hbc1b5e5a),
	.w7(32'hbc45bdc2),
	.w8(32'hbc51142b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41c990),
	.w1(32'hbae42d13),
	.w2(32'h3ab8dbe0),
	.w3(32'h3c52198c),
	.w4(32'h3a6f0457),
	.w5(32'hb9d212a5),
	.w6(32'hb67bc45c),
	.w7(32'hbaa07c08),
	.w8(32'hb7aecb37),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b731198),
	.w1(32'h3bf7d6f4),
	.w2(32'h39bb2c27),
	.w3(32'h39574a8f),
	.w4(32'h3ca5268e),
	.w5(32'h3caa2124),
	.w6(32'hba786641),
	.w7(32'hbc06184b),
	.w8(32'hbbc96416),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01fe1a),
	.w1(32'h3b3cd2a5),
	.w2(32'h3b53d94b),
	.w3(32'h3c707c41),
	.w4(32'h3b9c2c16),
	.w5(32'h3b5951b9),
	.w6(32'h3bad21f0),
	.w7(32'h3bfac6e8),
	.w8(32'h3b4c2229),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac794fe),
	.w1(32'hbb209fae),
	.w2(32'h3bd2aadc),
	.w3(32'hbae565c6),
	.w4(32'hbc2d891f),
	.w5(32'h3bba0ffc),
	.w6(32'hbb7dc8d5),
	.w7(32'hbbf65d07),
	.w8(32'h3a89cd47),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae42112),
	.w1(32'h3c75d81d),
	.w2(32'h3c903481),
	.w3(32'hbb2a84bf),
	.w4(32'hbc0e1e71),
	.w5(32'h3c212b89),
	.w6(32'h3c9d375c),
	.w7(32'h3ba247a1),
	.w8(32'h3afc71c2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd84d94),
	.w1(32'hbcbe13a5),
	.w2(32'hbd0dfed0),
	.w3(32'h3c382c42),
	.w4(32'hbc8ca4d2),
	.w5(32'hbcb79f6d),
	.w6(32'hbc4622a8),
	.w7(32'hbcc89021),
	.w8(32'hbcc72a82),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf319d3),
	.w1(32'hbcb87911),
	.w2(32'hbc0c776d),
	.w3(32'hbcda9030),
	.w4(32'hbc96ab4d),
	.w5(32'hbc32e249),
	.w6(32'hbc05f155),
	.w7(32'hbb72bb6b),
	.w8(32'h3b50a1b6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7712d5),
	.w1(32'h393bb7d2),
	.w2(32'hbabb5283),
	.w3(32'hbc4cce88),
	.w4(32'hbba90edf),
	.w5(32'hbc50faf8),
	.w6(32'h3bb25af1),
	.w7(32'h3b67a503),
	.w8(32'h3c207bf5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb16c41),
	.w1(32'hbaf8a6c6),
	.w2(32'hbb4603b9),
	.w3(32'hbb3399e8),
	.w4(32'h3b28ae51),
	.w5(32'h3b0a833e),
	.w6(32'hba8a780a),
	.w7(32'hbb2ed69c),
	.w8(32'hbb0e775b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e577b),
	.w1(32'h3c1cdd33),
	.w2(32'h3ace5c2b),
	.w3(32'hbad65a83),
	.w4(32'h3bb818c0),
	.w5(32'hba39590f),
	.w6(32'h3b489db6),
	.w7(32'h3ab9b9b8),
	.w8(32'h3a7af679),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af49841),
	.w1(32'hbb5d9e6f),
	.w2(32'h3b58d963),
	.w3(32'hbb82ef32),
	.w4(32'hbca601bb),
	.w5(32'hbcbc9b20),
	.w6(32'h3c35a995),
	.w7(32'h3c963a4f),
	.w8(32'h3b8f4056),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13c090),
	.w1(32'hbc025505),
	.w2(32'h3c127e26),
	.w3(32'hbc86fced),
	.w4(32'hbc9a0a77),
	.w5(32'hbc843181),
	.w6(32'h3a563108),
	.w7(32'h3be9532b),
	.w8(32'hbb165bd9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b8853),
	.w1(32'h3ac90a8f),
	.w2(32'h3b843f1c),
	.w3(32'h3ab8fd37),
	.w4(32'hbb5d9663),
	.w5(32'h3b271e71),
	.w6(32'h3ac6698c),
	.w7(32'h3c32fe64),
	.w8(32'h3c4ddd8e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9447ce),
	.w1(32'hba1f29cb),
	.w2(32'hba82a9aa),
	.w3(32'h3bc6e856),
	.w4(32'h3a043e3a),
	.w5(32'h3b07b320),
	.w6(32'hba34f3d7),
	.w7(32'hbb824cb1),
	.w8(32'h39880062),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd3c4),
	.w1(32'hbb8fcb95),
	.w2(32'hbbea0812),
	.w3(32'h3b87dda6),
	.w4(32'h3a3240a0),
	.w5(32'hba8cf6bf),
	.w6(32'hbb3dd6b5),
	.w7(32'h395dcfa1),
	.w8(32'h3b939be1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a672210),
	.w1(32'h3b369984),
	.w2(32'h3c19b8cd),
	.w3(32'hba7cfaed),
	.w4(32'hbabc4f2e),
	.w5(32'h3b378c75),
	.w6(32'h3bb059ae),
	.w7(32'h3b79fd60),
	.w8(32'h39f9cc0c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8e612),
	.w1(32'hbc60d79e),
	.w2(32'hbcca6c51),
	.w3(32'h3ba78bbe),
	.w4(32'hbbd20f4f),
	.w5(32'hbccc9f7f),
	.w6(32'hbb2475b2),
	.w7(32'hbc4d2f42),
	.w8(32'hbba53259),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf61682),
	.w1(32'h3b8b37f0),
	.w2(32'h3b6b978e),
	.w3(32'hbc71bd66),
	.w4(32'h3bceefc6),
	.w5(32'h3bff4f87),
	.w6(32'hbac478c2),
	.w7(32'hba3202bd),
	.w8(32'h39b78c9f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb044ec4),
	.w1(32'hbc517c80),
	.w2(32'hbcd26e36),
	.w3(32'h3b55c6b1),
	.w4(32'hbbb5a5cd),
	.w5(32'hbbb6621f),
	.w6(32'hbc22ddf9),
	.w7(32'hbcd21a3e),
	.w8(32'hbc47e4a7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1f513),
	.w1(32'hbb93fb5c),
	.w2(32'hbbd8b23d),
	.w3(32'hbbddea7e),
	.w4(32'h3b0644cf),
	.w5(32'hbc32af5b),
	.w6(32'hbbb42737),
	.w7(32'h3bbc65ed),
	.w8(32'h3bbd25de),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92d5b3),
	.w1(32'h3b94eb20),
	.w2(32'h398ff12f),
	.w3(32'hbb1a651c),
	.w4(32'h3a2f4092),
	.w5(32'h3c1a8216),
	.w6(32'hbbe08cb6),
	.w7(32'hbc5dad27),
	.w8(32'hbbee1e8b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af23a),
	.w1(32'h3c310b26),
	.w2(32'h3c191038),
	.w3(32'h3b64938d),
	.w4(32'h3bf27398),
	.w5(32'h3c14e584),
	.w6(32'hbbed87a9),
	.w7(32'hb9836a82),
	.w8(32'hbbb4ec27),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12df34),
	.w1(32'hbc1150d5),
	.w2(32'hbc2cfd39),
	.w3(32'hbc12087b),
	.w4(32'h3bc7eb1f),
	.w5(32'hbc0cb7fe),
	.w6(32'hbc4140e6),
	.w7(32'hbc2a34cf),
	.w8(32'hbba23245),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba294fb4),
	.w1(32'h3bfed4d0),
	.w2(32'h3bdb8fbd),
	.w3(32'hbbab9b3e),
	.w4(32'h3bbb57d9),
	.w5(32'hbad73767),
	.w6(32'h3bf9a639),
	.w7(32'h3b906ee2),
	.w8(32'h3accefff),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31b4c8),
	.w1(32'hbb920316),
	.w2(32'hbbd6edbf),
	.w3(32'hbc1a31a4),
	.w4(32'hb7bdd64a),
	.w5(32'hbb2c4629),
	.w6(32'h3b9b53c0),
	.w7(32'hba16fd04),
	.w8(32'h3c00c35a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b36ab),
	.w1(32'h3b48b564),
	.w2(32'hba1688d0),
	.w3(32'hbb519451),
	.w4(32'h3c464de7),
	.w5(32'h3be3afcb),
	.w6(32'hbb504e34),
	.w7(32'hbc032e3c),
	.w8(32'hbbf514de),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad73c9d),
	.w1(32'h3a451211),
	.w2(32'h3af80417),
	.w3(32'h3b088659),
	.w4(32'h3b9faca7),
	.w5(32'hba86f028),
	.w6(32'h3ad17bfa),
	.w7(32'h3b1eb623),
	.w8(32'h3b42dee7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ba49a),
	.w1(32'h3b21f6ec),
	.w2(32'h3b36835a),
	.w3(32'hbc026158),
	.w4(32'h3b3e48a7),
	.w5(32'h3a92ebd5),
	.w6(32'h3a701aac),
	.w7(32'hb9442a78),
	.w8(32'hbb113f8e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dfb19),
	.w1(32'h3ca0aa12),
	.w2(32'h3b2b3342),
	.w3(32'hbb44b4b8),
	.w4(32'h3c7f8809),
	.w5(32'h3c83c7fa),
	.w6(32'h3b6d42fe),
	.w7(32'hbcc4b3e6),
	.w8(32'hbcc58d97),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca29d1c),
	.w1(32'hbcc8c588),
	.w2(32'hbd1b9a35),
	.w3(32'h3bd63eef),
	.w4(32'hbc00c502),
	.w5(32'hbc86ffd8),
	.w6(32'hbc8cade3),
	.w7(32'hbcd8f0db),
	.w8(32'hbc82c0a7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf0916),
	.w1(32'h3c2886c3),
	.w2(32'h3c646521),
	.w3(32'hbc849c57),
	.w4(32'h3b74d8e3),
	.w5(32'h3a933074),
	.w6(32'h39780072),
	.w7(32'h3b140708),
	.w8(32'hba78a8bd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf0fef),
	.w1(32'hbc32be54),
	.w2(32'hbc0ceafa),
	.w3(32'hb93686d2),
	.w4(32'hbc525f98),
	.w5(32'hbbcaecf5),
	.w6(32'hba8da518),
	.w7(32'hbc850ee5),
	.w8(32'hbc3890c2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0fd6d),
	.w1(32'h3abdb55f),
	.w2(32'hbc859bdc),
	.w3(32'h3aa9530c),
	.w4(32'hba51b7c8),
	.w5(32'h3a373417),
	.w6(32'hbb24b135),
	.w7(32'hbbbf36e2),
	.w8(32'h3a0788ac),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75427c),
	.w1(32'hbc1cde29),
	.w2(32'hbc42d94b),
	.w3(32'hb83fa3ee),
	.w4(32'hbbc651fd),
	.w5(32'hbb337375),
	.w6(32'hbba3e8ed),
	.w7(32'hbb6427fc),
	.w8(32'h3a01eadf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24d6bd),
	.w1(32'h3ccf5354),
	.w2(32'h3ce373a3),
	.w3(32'hbbd95938),
	.w4(32'h3c8c7e66),
	.w5(32'h3cc3e3b6),
	.w6(32'h3c88c959),
	.w7(32'h3b105dae),
	.w8(32'h3bc13df6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0614af),
	.w1(32'h3c9ae38c),
	.w2(32'h3ba65df2),
	.w3(32'h3cc94fbc),
	.w4(32'h3c21bc75),
	.w5(32'h3c52954b),
	.w6(32'h3c033f01),
	.w7(32'h3b9309ee),
	.w8(32'hbbc133e1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a3aa4),
	.w1(32'h3c48b33e),
	.w2(32'h3bdee065),
	.w3(32'h3a660662),
	.w4(32'h3b9bdc17),
	.w5(32'h3bc4b0df),
	.w6(32'hb757eaaf),
	.w7(32'hbc02622b),
	.w8(32'hbbf34341),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb79925),
	.w1(32'hbc169f12),
	.w2(32'hbab40d84),
	.w3(32'hbb47fcce),
	.w4(32'h3a707fab),
	.w5(32'h3a7c9c74),
	.w6(32'h3b51d6d1),
	.w7(32'h3c64b029),
	.w8(32'h3c0cab16),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c257f1f),
	.w1(32'h3bd56dc7),
	.w2(32'hbb26ddf0),
	.w3(32'h3b9f5f1e),
	.w4(32'h3c0f4f60),
	.w5(32'h3aff3607),
	.w6(32'h3b726606),
	.w7(32'hbb55c0a2),
	.w8(32'hbb9caf1d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b8b20),
	.w1(32'hbacd0a57),
	.w2(32'hbb0e826f),
	.w3(32'hbc1b5c0f),
	.w4(32'hbc01d53c),
	.w5(32'hbbb4a232),
	.w6(32'h3a8df375),
	.w7(32'hbc2be84a),
	.w8(32'hbc1c3b59),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b737f59),
	.w1(32'hb9ca670a),
	.w2(32'hbaf426ea),
	.w3(32'hbc4230c7),
	.w4(32'h3b64bd9b),
	.w5(32'h3b8177e7),
	.w6(32'hbb01d0c2),
	.w7(32'hbb8c215f),
	.w8(32'h3a4e0f7f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbded30c),
	.w1(32'hbb759f4d),
	.w2(32'hbc2eb3f1),
	.w3(32'h3a92c0e9),
	.w4(32'hbc10b3ae),
	.w5(32'hbad1c74c),
	.w6(32'h3bd4b60d),
	.w7(32'h3ae16a94),
	.w8(32'h3be6b8e1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0888fa),
	.w1(32'h3b0bc520),
	.w2(32'hb89be2b3),
	.w3(32'h3b27788a),
	.w4(32'h3acc36ed),
	.w5(32'h3a5f5cfc),
	.w6(32'h3a7d9aa4),
	.w7(32'hbab63b15),
	.w8(32'h3a011e99),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40f270),
	.w1(32'hbb557c7a),
	.w2(32'hbbc3f90f),
	.w3(32'h3adef7f7),
	.w4(32'h3a5a5b05),
	.w5(32'hbac31507),
	.w6(32'hbb7121ab),
	.w7(32'hbb4b7b54),
	.w8(32'hb93b2014),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe023f),
	.w1(32'h3bedc24d),
	.w2(32'h3c7aa968),
	.w3(32'hbb56d48f),
	.w4(32'hbc9ea151),
	.w5(32'hbbfa45b4),
	.w6(32'h3caf375d),
	.w7(32'h3bf9b314),
	.w8(32'h3bdd2007),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c0eb1),
	.w1(32'h3c10ba50),
	.w2(32'h3b19b29e),
	.w3(32'h3bde172c),
	.w4(32'h3bd3be71),
	.w5(32'hb9cdcc9c),
	.w6(32'h3c0de587),
	.w7(32'h3ba409ee),
	.w8(32'hbb5c0114),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf12d58),
	.w1(32'hbbb9de40),
	.w2(32'hbc320cef),
	.w3(32'hbbff23ad),
	.w4(32'h3c796373),
	.w5(32'hba0f10fa),
	.w6(32'h3b281824),
	.w7(32'h3ad9d9a2),
	.w8(32'h3b7cc9ec),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bd52a),
	.w1(32'h3b9a29cc),
	.w2(32'h3c237982),
	.w3(32'hbb662492),
	.w4(32'h3b5b8d95),
	.w5(32'h3c03979c),
	.w6(32'h3b2c45f9),
	.w7(32'h3c273475),
	.w8(32'hbb2cca4e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc121fa1),
	.w1(32'h3ba517a9),
	.w2(32'h3b590bb7),
	.w3(32'hbaa44331),
	.w4(32'h3c17f246),
	.w5(32'h3c2205dc),
	.w6(32'h3a30765f),
	.w7(32'h3ac413f2),
	.w8(32'hbbf26252),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe242f8),
	.w1(32'h3b1ecffb),
	.w2(32'h3b90b892),
	.w3(32'hb9a2c877),
	.w4(32'hbb5752d5),
	.w5(32'hbb85e9a8),
	.w6(32'h3c5a0fa9),
	.w7(32'h3cc0cdc3),
	.w8(32'h3c6f5085),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b825bb0),
	.w1(32'hb9b02b13),
	.w2(32'h3bbd66bb),
	.w3(32'hbb88c578),
	.w4(32'hbc34a090),
	.w5(32'h3b8cd9b7),
	.w6(32'hbb3db8c7),
	.w7(32'hbc3394c8),
	.w8(32'h3aec32ce),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e70fc),
	.w1(32'hbc34719e),
	.w2(32'hbcb1f7c8),
	.w3(32'h3c415fbb),
	.w4(32'hbc8d0bf5),
	.w5(32'hbc8e1a85),
	.w6(32'hbbbf8635),
	.w7(32'hbc43f906),
	.w8(32'hbb6c8934),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a0c7f),
	.w1(32'h3bc67dee),
	.w2(32'h38593e6f),
	.w3(32'hbc3971a6),
	.w4(32'hbb92a7bf),
	.w5(32'h3b363998),
	.w6(32'h3bc3a647),
	.w7(32'hbba68344),
	.w8(32'hba8ef917),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ed86d),
	.w1(32'hbc1c2a41),
	.w2(32'hbc4e9338),
	.w3(32'h3c134514),
	.w4(32'hbb3ce648),
	.w5(32'hbc8238e0),
	.w6(32'hbc2ded1e),
	.w7(32'hbbba3be4),
	.w8(32'h3b04137b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab337a0),
	.w1(32'h3bf80b4f),
	.w2(32'h3b5c05cf),
	.w3(32'hbc2ded64),
	.w4(32'h3b6074f7),
	.w5(32'hbb3a5999),
	.w6(32'h3a31d140),
	.w7(32'h3b07cc30),
	.w8(32'hbc0a0fde),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3041f5),
	.w1(32'h37988211),
	.w2(32'hba5714b4),
	.w3(32'hbb7142ee),
	.w4(32'h3aeaaab1),
	.w5(32'h3af4dc4c),
	.w6(32'h3b869555),
	.w7(32'h3bb21e7c),
	.w8(32'h3bd18c25),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b450d95),
	.w1(32'h3c587846),
	.w2(32'h3be9f7bc),
	.w3(32'h3ba7ab02),
	.w4(32'h3a271ac7),
	.w5(32'h3b55af1a),
	.w6(32'h3c0b2981),
	.w7(32'hbad9a28e),
	.w8(32'h3a46a496),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd665b),
	.w1(32'hbadf374d),
	.w2(32'h3c60433e),
	.w3(32'hbc4f0e39),
	.w4(32'hbcd90901),
	.w5(32'hbc5d5c51),
	.w6(32'h3c14c287),
	.w7(32'h3be6a754),
	.w8(32'hbba0dca9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dd0c1),
	.w1(32'h3c20da9a),
	.w2(32'h3cb9a4b0),
	.w3(32'h3ad35195),
	.w4(32'hb961eae0),
	.w5(32'h3c5160d5),
	.w6(32'h3bbc540d),
	.w7(32'h3c3500c6),
	.w8(32'h3b7779be),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c5469),
	.w1(32'h3a799371),
	.w2(32'hbad279a8),
	.w3(32'h3c14847b),
	.w4(32'h3b3e00bc),
	.w5(32'h3a948c1e),
	.w6(32'hb9a3c777),
	.w7(32'h3ae8ec15),
	.w8(32'h3b72937e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a829e0f),
	.w1(32'h3c225baa),
	.w2(32'h3c413a05),
	.w3(32'h39920a71),
	.w4(32'h3bc80af4),
	.w5(32'h3c220c26),
	.w6(32'h3b97732a),
	.w7(32'h3b7f14dd),
	.w8(32'hba1f7fdb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ef907),
	.w1(32'hbbb43597),
	.w2(32'hbc00860e),
	.w3(32'h3c2f973e),
	.w4(32'hbbdae19d),
	.w5(32'hbbec4d20),
	.w6(32'hbb9ab21c),
	.w7(32'hbb4b525f),
	.w8(32'h389379fe),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a6ce5),
	.w1(32'h3c2b28ca),
	.w2(32'h3c110148),
	.w3(32'hbba212ee),
	.w4(32'h3c2d8649),
	.w5(32'h3c240c36),
	.w6(32'h3bae2283),
	.w7(32'h3aeb2b29),
	.w8(32'h3c09ed99),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf576d),
	.w1(32'hbc91bf86),
	.w2(32'hbc9d7b5a),
	.w3(32'h3b102276),
	.w4(32'hbbaf6815),
	.w5(32'hbc5369e9),
	.w6(32'hbc89d757),
	.w7(32'hbc464ad1),
	.w8(32'hbbf5d4a9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc408766),
	.w1(32'h3be30c9c),
	.w2(32'hbbdd9fae),
	.w3(32'hbc77750e),
	.w4(32'h3c6aa7ee),
	.w5(32'h3c45a31b),
	.w6(32'hbbd50f2d),
	.w7(32'hbc9733f4),
	.w8(32'hbc204d10),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc831c4b),
	.w1(32'h3a1f8166),
	.w2(32'hbb094258),
	.w3(32'h3a79d813),
	.w4(32'h3b60d033),
	.w5(32'h39f67473),
	.w6(32'hb797ad29),
	.w7(32'h3b4dfcfb),
	.w8(32'h3b626696),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95d975),
	.w1(32'hbc030db7),
	.w2(32'h3bc1cd3e),
	.w3(32'hba73b55c),
	.w4(32'hbc82a921),
	.w5(32'hbc52cc95),
	.w6(32'h3b045a80),
	.w7(32'h3bc431e9),
	.w8(32'h3bf23e68),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b3650),
	.w1(32'hb9421d01),
	.w2(32'hbb00b6c1),
	.w3(32'h3b633e85),
	.w4(32'h3baa510a),
	.w5(32'hbb3a3e97),
	.w6(32'h3ac29b47),
	.w7(32'h3b0bd33d),
	.w8(32'h3bb6f933),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7183c),
	.w1(32'hbc425ec6),
	.w2(32'hbcf61adb),
	.w3(32'h3bb4db2a),
	.w4(32'hbb007655),
	.w5(32'hbc3a51ba),
	.w6(32'hbc34e1ee),
	.w7(32'hbca4c151),
	.w8(32'hbc94c83a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca14cbb),
	.w1(32'h3abdf334),
	.w2(32'h3a986840),
	.w3(32'hbbca815f),
	.w4(32'h3c23cc01),
	.w5(32'h3ba18c0d),
	.w6(32'hbb3238e2),
	.w7(32'hbbdf056e),
	.w8(32'h3b86175e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f634cc),
	.w1(32'hbcb96391),
	.w2(32'hbd02427c),
	.w3(32'h3b5cb577),
	.w4(32'hbc418d70),
	.w5(32'hbc9b0985),
	.w6(32'hbc8ca79d),
	.w7(32'hbd036385),
	.w8(32'hbc8fdd1c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7df47),
	.w1(32'hbc2324a9),
	.w2(32'hbc82e59f),
	.w3(32'hbcab2951),
	.w4(32'hbba83f6f),
	.w5(32'hbbccfcd5),
	.w6(32'hbb104b7e),
	.w7(32'hbb5b8c0d),
	.w8(32'hbad8bd15),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5aea67),
	.w1(32'h3a2f0fc0),
	.w2(32'hba30e23d),
	.w3(32'hbb8be1da),
	.w4(32'h3b426295),
	.w5(32'h39935c55),
	.w6(32'hbaf97013),
	.w7(32'hbb0e466a),
	.w8(32'h3aa45aa7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dcf461),
	.w1(32'hb984eeee),
	.w2(32'h3bab0796),
	.w3(32'hb9333c83),
	.w4(32'h3b8424ea),
	.w5(32'h3c10c5c0),
	.w6(32'hb8256b6a),
	.w7(32'h3b4a7d92),
	.w8(32'h3b95e71f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba295d2),
	.w1(32'h3b9a3ee9),
	.w2(32'h3ce63d40),
	.w3(32'h3c300441),
	.w4(32'hbc5626cf),
	.w5(32'hbc6a6c60),
	.w6(32'h3cda51f4),
	.w7(32'h3c34adce),
	.w8(32'h39432c6e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccfc30a),
	.w1(32'hbc4a3237),
	.w2(32'hbc692bfc),
	.w3(32'h3bdd13ee),
	.w4(32'hbb0a1b20),
	.w5(32'hbc40bbb5),
	.w6(32'h3b4a3cfd),
	.w7(32'hbc86282b),
	.w8(32'hbc817c07),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560a49),
	.w1(32'hbb671c82),
	.w2(32'hbb1bb5da),
	.w3(32'hbbfed26a),
	.w4(32'hba503206),
	.w5(32'hb994a409),
	.w6(32'hbb2270e9),
	.w7(32'hbb12d7a9),
	.w8(32'h3acbf782),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98f234),
	.w1(32'h3929615e),
	.w2(32'h3b10393a),
	.w3(32'h3b308927),
	.w4(32'h3b3cc73c),
	.w5(32'h3b050587),
	.w6(32'h3beab4fd),
	.w7(32'h3c287a29),
	.w8(32'h3c13d3fd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule