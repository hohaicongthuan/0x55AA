module layer_10_featuremap_191(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380d6abe),
	.w1(32'hb53d66ee),
	.w2(32'h3724f008),
	.w3(32'h383987a0),
	.w4(32'h36ed0924),
	.w5(32'h3706e090),
	.w6(32'h38109665),
	.w7(32'h37e1e969),
	.w8(32'h37c251c2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac26306),
	.w1(32'hbac507ea),
	.w2(32'hbb2ecf2f),
	.w3(32'hba710269),
	.w4(32'hb990177d),
	.w5(32'hbb39bd6f),
	.w6(32'hbaaa18c6),
	.w7(32'hbaf43a1f),
	.w8(32'hbbbdd216),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371ce8d6),
	.w1(32'h37135b3f),
	.w2(32'h37841c92),
	.w3(32'h3707e9f5),
	.w4(32'h32a6581b),
	.w5(32'h371f2756),
	.w6(32'h377142ad),
	.w7(32'h36efa5c8),
	.w8(32'h379b4ce1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6268e7),
	.w1(32'h3a12a62d),
	.w2(32'h3a29b043),
	.w3(32'hb9261b03),
	.w4(32'hb9fc2a76),
	.w5(32'hba28b771),
	.w6(32'hb9bb4f52),
	.w7(32'hb950070b),
	.w8(32'hba00a7f2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39933284),
	.w1(32'h389e880e),
	.w2(32'hb98210a0),
	.w3(32'h39c9deef),
	.w4(32'h3999dad0),
	.w5(32'hb813ea77),
	.w6(32'h39c3471f),
	.w7(32'h39d05d10),
	.w8(32'h39495711),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3767e01a),
	.w1(32'h36fed02b),
	.w2(32'h3834e0cf),
	.w3(32'h37ebd69e),
	.w4(32'h3784f75a),
	.w5(32'h382ec949),
	.w6(32'h381a8bcf),
	.w7(32'h37339b94),
	.w8(32'h381675c6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a87fe),
	.w1(32'hbb9df820),
	.w2(32'hbb2d5c06),
	.w3(32'hbaefc743),
	.w4(32'hbbc77bc9),
	.w5(32'hbb814d5f),
	.w6(32'hb98214ec),
	.w7(32'hbb05826f),
	.w8(32'hba47555a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc811a66),
	.w1(32'hbc003c70),
	.w2(32'hbbadf20a),
	.w3(32'hbca2f530),
	.w4(32'hbc1fdfea),
	.w5(32'h36e0bad0),
	.w6(32'hbc83ecbf),
	.w7(32'hbba62689),
	.w8(32'h3ae11b4e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9fdee),
	.w1(32'hb9714d99),
	.w2(32'hba0b8e4f),
	.w3(32'hb8a117ac),
	.w4(32'hba294093),
	.w5(32'hba30b57b),
	.w6(32'hb834eef1),
	.w7(32'hba0fdb7a),
	.w8(32'hba7a9ea0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce49d2),
	.w1(32'hbb43218d),
	.w2(32'hbbd79fb7),
	.w3(32'hbb8e404e),
	.w4(32'hba9f0604),
	.w5(32'hbb20bb58),
	.w6(32'hbba11cd7),
	.w7(32'h3a88660c),
	.w8(32'hb93e718f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc78da),
	.w1(32'hb8a8d275),
	.w2(32'hba26241e),
	.w3(32'h38d6b040),
	.w4(32'h397b9b6e),
	.w5(32'hb9b8e462),
	.w6(32'hb81264dd),
	.w7(32'h392daf64),
	.w8(32'hb9a748da),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba529a35),
	.w1(32'h398f0483),
	.w2(32'hba421034),
	.w3(32'hb828325e),
	.w4(32'h3ab21610),
	.w5(32'hbad9c86b),
	.w6(32'h3a69b447),
	.w7(32'h3b4cfe63),
	.w8(32'h3b68c4e9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca4948),
	.w1(32'hbb299ac7),
	.w2(32'hbba37bc4),
	.w3(32'hbbcd9856),
	.w4(32'hbb1c230c),
	.w5(32'hbb462836),
	.w6(32'hbb592639),
	.w7(32'hb97730a6),
	.w8(32'h39d91e0d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09b8d1),
	.w1(32'hbb29a90f),
	.w2(32'hbb75ac25),
	.w3(32'hbaaa5bbf),
	.w4(32'hb94ad3b0),
	.w5(32'hb769e05a),
	.w6(32'hba78d871),
	.w7(32'hba676b97),
	.w8(32'hba49b27a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a111c63),
	.w1(32'h3a29801d),
	.w2(32'hba802ac0),
	.w3(32'h3a932040),
	.w4(32'h3ac4c560),
	.w5(32'hb9b221bc),
	.w6(32'h39689b5e),
	.w7(32'hba13fa7e),
	.w8(32'hbb5ab630),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda54e4),
	.w1(32'hbb30c9f7),
	.w2(32'hbb10c56f),
	.w3(32'hbbcb0e4b),
	.w4(32'h3ab0a48e),
	.w5(32'h3af405cf),
	.w6(32'hbbe863f5),
	.w7(32'h3adb1d13),
	.w8(32'h3a30d867),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927029f),
	.w1(32'hb84b7de0),
	.w2(32'hb8f5bfa7),
	.w3(32'hb91a9272),
	.w4(32'h392197a5),
	.w5(32'hb7277e23),
	.w6(32'hb9263213),
	.w7(32'h3922f4b5),
	.w8(32'h3822db93),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c7bd0),
	.w1(32'hbbdfc36e),
	.w2(32'hbc015186),
	.w3(32'hbc11981a),
	.w4(32'h394f29ea),
	.w5(32'hba653dda),
	.w6(32'hbc009200),
	.w7(32'h3b8948c5),
	.w8(32'h3bccf20b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7752d),
	.w1(32'hbb1deb9b),
	.w2(32'hbb40c524),
	.w3(32'hbb9e336c),
	.w4(32'hba3355a4),
	.w5(32'hba192496),
	.w6(32'hbb5a7424),
	.w7(32'h3ad43226),
	.w8(32'h3ada0c28),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c5c478),
	.w1(32'h3864f9fa),
	.w2(32'h390429ec),
	.w3(32'h386c15f3),
	.w4(32'h3945a920),
	.w5(32'h3955d280),
	.w6(32'hb7c8d3b9),
	.w7(32'h385371d8),
	.w8(32'hb856b20b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a8fbaa),
	.w1(32'hb88de62c),
	.w2(32'hb7396285),
	.w3(32'hb8ddd4c6),
	.w4(32'hb903fc21),
	.w5(32'hb8c3c667),
	.w6(32'hb824d698),
	.w7(32'hb689c93b),
	.w8(32'h3911307d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b86c5),
	.w1(32'h3a793361),
	.w2(32'hba608e8c),
	.w3(32'h3b420e46),
	.w4(32'h3a8c1df5),
	.w5(32'hbac08011),
	.w6(32'h3ad8784b),
	.w7(32'h399dbfa4),
	.w8(32'hbb099355),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a8d2c),
	.w1(32'hbb93bb40),
	.w2(32'hbb88dbab),
	.w3(32'hbbe0a404),
	.w4(32'hbb022c70),
	.w5(32'hbb7875a8),
	.w6(32'hbc2562fc),
	.w7(32'h3bc73cd1),
	.w8(32'h387a3e85),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb048201),
	.w1(32'hb9f119f6),
	.w2(32'hbba2a17c),
	.w3(32'h3a56939a),
	.w4(32'h3b061df6),
	.w5(32'hbaffbb4a),
	.w6(32'hba864eff),
	.w7(32'h3a35fe63),
	.w8(32'hbb80b5b3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21cc3d),
	.w1(32'h3b2657ba),
	.w2(32'hbb812d23),
	.w3(32'hb8b62184),
	.w4(32'h3abad29c),
	.w5(32'hbb9ad048),
	.w6(32'hbaf3d7c7),
	.w7(32'hbb204174),
	.w8(32'hbc32b9ad),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03037c),
	.w1(32'hb9bb7581),
	.w2(32'hb97976a1),
	.w3(32'h399ff361),
	.w4(32'hba052d69),
	.w5(32'hb9d5c409),
	.w6(32'h3978c02f),
	.w7(32'hb936dc74),
	.w8(32'hb9a8323d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e8cea),
	.w1(32'h391fd1c5),
	.w2(32'h397878e0),
	.w3(32'h38d183ea),
	.w4(32'h38e29dd4),
	.w5(32'h3944cc4b),
	.w6(32'h3925aaaa),
	.w7(32'h39273e3f),
	.w8(32'h3956ff93),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c185bec),
	.w1(32'hbbd598ed),
	.w2(32'hbbe18b9b),
	.w3(32'h3aa3038c),
	.w4(32'hbbe566c3),
	.w5(32'hbb90148b),
	.w6(32'h3c1a37ea),
	.w7(32'h3b6d209d),
	.w8(32'h3b1dc0d5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99531c),
	.w1(32'h3a900190),
	.w2(32'hba06a5c5),
	.w3(32'h3ae794df),
	.w4(32'h3ad4d998),
	.w5(32'hba4a3344),
	.w6(32'h395f5fce),
	.w7(32'h3aaed813),
	.w8(32'hb9d24ab5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cc99a),
	.w1(32'h3a2b6ded),
	.w2(32'hbb3274a7),
	.w3(32'h3b675080),
	.w4(32'hbb543d85),
	.w5(32'hbc02695f),
	.w6(32'h3ba34151),
	.w7(32'hbb027124),
	.w8(32'hbc319e7d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387419b8),
	.w1(32'h384b2d15),
	.w2(32'h38567cd5),
	.w3(32'h38353c77),
	.w4(32'h386d19df),
	.w5(32'h386a6199),
	.w6(32'h3860e02e),
	.w7(32'h38785ec0),
	.w8(32'h387df3f7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb740b381),
	.w1(32'h382e630a),
	.w2(32'h37fcc87e),
	.w3(32'h37a8874a),
	.w4(32'h3860e3aa),
	.w5(32'h385e47a6),
	.w6(32'h374069a0),
	.w7(32'h3869062e),
	.w8(32'h37de677b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb023aa7),
	.w1(32'hba2e3ca3),
	.w2(32'hbaffdcda),
	.w3(32'h39a6111f),
	.w4(32'h3af1a1a7),
	.w5(32'h39cd3662),
	.w6(32'hb9ccdca5),
	.w7(32'h3aa9b18c),
	.w8(32'h39816451),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba427b52),
	.w1(32'hba3b2fdd),
	.w2(32'hbb095aeb),
	.w3(32'hba4dd580),
	.w4(32'hb9738e01),
	.w5(32'hbadb0adf),
	.w6(32'hba974d09),
	.w7(32'hba97c23e),
	.w8(32'hbb3fd731),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a50a4),
	.w1(32'hb8165e2d),
	.w2(32'h39c759f7),
	.w3(32'hb8982a56),
	.w4(32'h39546fa6),
	.w5(32'h39e63d8a),
	.w6(32'hb9d332d9),
	.w7(32'h3a0cfbcc),
	.w8(32'h3a547063),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ef3da),
	.w1(32'hbb7723f1),
	.w2(32'hbafb9729),
	.w3(32'hbb108cac),
	.w4(32'hbb7f1aec),
	.w5(32'hbaa6ef3e),
	.w6(32'hbad2e16b),
	.w7(32'hb9f766f6),
	.w8(32'h3b0a5a98),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66e49b),
	.w1(32'hbbbe8b45),
	.w2(32'hbbf3db6e),
	.w3(32'hbaf0ccf0),
	.w4(32'hba5b2714),
	.w5(32'h3b2885cd),
	.w6(32'h3b78854f),
	.w7(32'h3bb83973),
	.w8(32'hbb58bb15),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38e3d8),
	.w1(32'h3a37ca83),
	.w2(32'hbc0cb9cc),
	.w3(32'h3c11ea44),
	.w4(32'h3b0a13dd),
	.w5(32'hbc1fb1e5),
	.w6(32'h3b2ae40b),
	.w7(32'hbbe23d56),
	.w8(32'hbca32913),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca595d9),
	.w1(32'h3bdcefc0),
	.w2(32'hbbdd29d1),
	.w3(32'h3c48513d),
	.w4(32'h3a6a7485),
	.w5(32'hbc8b01bc),
	.w6(32'h3bf7e3d2),
	.w7(32'hbb654542),
	.w8(32'hbcb14828),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb819f265),
	.w1(32'h38510c01),
	.w2(32'hba1dd450),
	.w3(32'hb99461ae),
	.w4(32'hba0ef762),
	.w5(32'hba8a6b8c),
	.w6(32'hba5046e4),
	.w7(32'hbaf8f15c),
	.w8(32'hbb50e1e4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361727ce),
	.w1(32'hb8869d92),
	.w2(32'h38e30836),
	.w3(32'hb7c65176),
	.w4(32'hb8c9a5a9),
	.w5(32'h3841d069),
	.w6(32'hb70c00f8),
	.w7(32'hb7e550ac),
	.w8(32'h391e8381),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fa4f62),
	.w1(32'h3892c9f5),
	.w2(32'h3919d108),
	.w3(32'h38ff235c),
	.w4(32'h3901861d),
	.w5(32'h39526a8b),
	.w6(32'h399cccfe),
	.w7(32'h39744cf9),
	.w8(32'h3972c113),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a2ee9),
	.w1(32'hb96a4a45),
	.w2(32'hba98f9e3),
	.w3(32'h39dc65c6),
	.w4(32'h3a966344),
	.w5(32'hba8f2a05),
	.w6(32'h3a317725),
	.w7(32'h3aad948f),
	.w8(32'hba6ac18d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a18dc),
	.w1(32'hbb74cee6),
	.w2(32'hbbc73189),
	.w3(32'hbc287e07),
	.w4(32'h3a679a22),
	.w5(32'hbb0b0634),
	.w6(32'hbbdcb581),
	.w7(32'h3b8c54a2),
	.w8(32'h3b8a74b7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bb15e),
	.w1(32'h3a68ca2c),
	.w2(32'hbb72bf4b),
	.w3(32'h3adfe0ca),
	.w4(32'h3b4bb706),
	.w5(32'hbb0af1dc),
	.w6(32'h3abb2428),
	.w7(32'h3ad1840c),
	.w8(32'hbbb2fa34),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b7edb),
	.w1(32'hbaac38b1),
	.w2(32'hbb84461d),
	.w3(32'hba3b7c8c),
	.w4(32'h3aa4be4d),
	.w5(32'h39d7d2a7),
	.w6(32'hbb0e48de),
	.w7(32'h3ad6e7ce),
	.w8(32'hbb14933d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee25a1),
	.w1(32'hb889351f),
	.w2(32'hbb7f6ff8),
	.w3(32'h398d57d8),
	.w4(32'h3b20000a),
	.w5(32'hba970393),
	.w6(32'hb9c5fe04),
	.w7(32'h3ac8601e),
	.w8(32'hbae8d434),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eae6f),
	.w1(32'hbbb680cf),
	.w2(32'hbc09da8c),
	.w3(32'hbc17c184),
	.w4(32'hbb47714c),
	.w5(32'hbb738ba2),
	.w6(32'hbbfb866d),
	.w7(32'h3b3e4ac2),
	.w8(32'h3bb24d7d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f12cc4),
	.w1(32'hb8d15c7b),
	.w2(32'hb8daf450),
	.w3(32'hb8180495),
	.w4(32'hb90ce7b4),
	.w5(32'hb8abf065),
	.w6(32'hb7b126e1),
	.w7(32'hb911147c),
	.w8(32'hb89bfcc8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94689a9),
	.w1(32'hb9af0464),
	.w2(32'hb96d64b2),
	.w3(32'hba81264a),
	.w4(32'hba537afe),
	.w5(32'hba1b51a8),
	.w6(32'hba8ce411),
	.w7(32'hba6bb145),
	.w8(32'hba6b1bab),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905f21a),
	.w1(32'h38223ba2),
	.w2(32'hb8703bee),
	.w3(32'h3922fa50),
	.w4(32'hb5f1713c),
	.w5(32'hb903f9ec),
	.w6(32'h38cbf791),
	.w7(32'hb9129a7d),
	.w8(32'hb913449d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43a481),
	.w1(32'hbb47bbc5),
	.w2(32'hbaf49050),
	.w3(32'hbb649a4d),
	.w4(32'hbae05fe2),
	.w5(32'hbb039fa0),
	.w6(32'hbb3fa207),
	.w7(32'h3a8bfa98),
	.w8(32'hba9104a8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3c788),
	.w1(32'hba2f1196),
	.w2(32'hba169f62),
	.w3(32'hba2b512c),
	.w4(32'h396df38b),
	.w5(32'h39a91a48),
	.w6(32'hba4345b3),
	.w7(32'h3a080795),
	.w8(32'h3a35e421),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49368a),
	.w1(32'hbb90fca5),
	.w2(32'hbbe9f8f9),
	.w3(32'hbbec4217),
	.w4(32'h3a992d36),
	.w5(32'hba92a7b6),
	.w6(32'hbb8a32f5),
	.w7(32'h3b995afa),
	.w8(32'h3b9c6063),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f9fbc),
	.w1(32'hb932bf52),
	.w2(32'hba82b7b3),
	.w3(32'hbae9c642),
	.w4(32'h3a2080b5),
	.w5(32'h383232fb),
	.w6(32'h397ebc43),
	.w7(32'h3aeb670e),
	.w8(32'h3a5c9bc2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366e33be),
	.w1(32'hb8ccd5c1),
	.w2(32'hb8a10fe4),
	.w3(32'h38030287),
	.w4(32'h38892bf2),
	.w5(32'hb85ed53c),
	.w6(32'h38f15f32),
	.w7(32'hb7f1c585),
	.w8(32'hb96c20b9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37decc3e),
	.w1(32'h3742e4b9),
	.w2(32'h37fc7efc),
	.w3(32'h36d1bf0d),
	.w4(32'hb657e794),
	.w5(32'h3691fdfd),
	.w6(32'h37e8c6d3),
	.w7(32'h36d168c6),
	.w8(32'hb70ea623),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63e452),
	.w1(32'h39903c35),
	.w2(32'hb9d6a594),
	.w3(32'h392f35f3),
	.w4(32'hb9cb0136),
	.w5(32'hba57de21),
	.w6(32'h39a97fb7),
	.w7(32'hb9a4947a),
	.w8(32'hba7268d2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdbcdd),
	.w1(32'h3a910295),
	.w2(32'h39926b29),
	.w3(32'h3ac2d11a),
	.w4(32'h3a9729e6),
	.w5(32'h38d8c011),
	.w6(32'h3a25f2af),
	.w7(32'h3a03b4f2),
	.w8(32'hb9c34e64),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398177ab),
	.w1(32'hb8ee1273),
	.w2(32'h3899459f),
	.w3(32'h391f3336),
	.w4(32'h38e609f6),
	.w5(32'hb8b93c8c),
	.w6(32'h39e1b8f2),
	.w7(32'h39a75a2d),
	.w8(32'h380ad2a9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdaabf),
	.w1(32'hbab5b9f2),
	.w2(32'hbb1482d6),
	.w3(32'hbb9b45a3),
	.w4(32'hb9467d00),
	.w5(32'hba218202),
	.w6(32'hbb3ffb26),
	.w7(32'h3aaa26a8),
	.w8(32'h3ab24001),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c9104),
	.w1(32'hbac3927b),
	.w2(32'hba974bfd),
	.w3(32'hbb848562),
	.w4(32'h3a1d089e),
	.w5(32'hb9a9e8ad),
	.w6(32'hbad5800f),
	.w7(32'h3bc7c98f),
	.w8(32'h3b80e4fb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366b2956),
	.w1(32'h372054be),
	.w2(32'h38d314f3),
	.w3(32'hb79b3ddf),
	.w4(32'hb5c64b37),
	.w5(32'h3894e91d),
	.w6(32'h37c2db6e),
	.w7(32'h37ef8134),
	.w8(32'h38bb17f4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382797ff),
	.w1(32'h37ca7ba3),
	.w2(32'h38936b4b),
	.w3(32'h37033dfe),
	.w4(32'h3602b774),
	.w5(32'h3833f77d),
	.w6(32'h382f5e66),
	.w7(32'h37822a2d),
	.w8(32'h3849c6bb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d9e110),
	.w1(32'h38185232),
	.w2(32'h3757738d),
	.w3(32'h37ba667a),
	.w4(32'h38844157),
	.w5(32'h384140b9),
	.w6(32'h381b2ce0),
	.w7(32'h389948c0),
	.w8(32'h3852e4e0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe4894),
	.w1(32'h3893957b),
	.w2(32'h3913814f),
	.w3(32'h38c03c4b),
	.w4(32'h384c0528),
	.w5(32'h390bd83f),
	.w6(32'h38c272a4),
	.w7(32'h38810600),
	.w8(32'h391a2864),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc102daa),
	.w1(32'h398315f0),
	.w2(32'hbb5f4cb8),
	.w3(32'hbbee756b),
	.w4(32'h3b50de2a),
	.w5(32'h3b21b6a8),
	.w6(32'hbbf4391a),
	.w7(32'h3bdfab56),
	.w8(32'h3c46c169),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc4105),
	.w1(32'h3777b10a),
	.w2(32'hbb37de3e),
	.w3(32'hbadde2b8),
	.w4(32'h3a7e4de7),
	.w5(32'h39aedc3e),
	.w6(32'hbbcdc5b3),
	.w7(32'h3a7eff25),
	.w8(32'hba6dfe61),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba30c4f),
	.w1(32'h379e0e77),
	.w2(32'hbbd18525),
	.w3(32'hbb6e8521),
	.w4(32'h3b81a0da),
	.w5(32'hbb1b63ac),
	.w6(32'hbb81be6f),
	.w7(32'h3bd764cb),
	.w8(32'h3a966cee),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02cd54),
	.w1(32'h3b642d72),
	.w2(32'hbbc9fe31),
	.w3(32'h3b5264b2),
	.w4(32'h3ad6027e),
	.w5(32'hbc07abae),
	.w6(32'hbaba874d),
	.w7(32'hbb489a9d),
	.w8(32'hbc8f98b9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370033e8),
	.w1(32'hb81569f1),
	.w2(32'h38c14dcb),
	.w3(32'h3609c616),
	.w4(32'hb7d2f394),
	.w5(32'h38dc46ac),
	.w6(32'h382c1018),
	.w7(32'h37cbacad),
	.w8(32'h3909cf4c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a8d5ab),
	.w1(32'h37f0dc3b),
	.w2(32'h393bccd2),
	.w3(32'h37e87177),
	.w4(32'hb64094d5),
	.w5(32'h393c616c),
	.w6(32'h38dee25b),
	.w7(32'h389678b3),
	.w8(32'h396fdd35),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c759e5),
	.w1(32'hb84d183d),
	.w2(32'h3920f0f0),
	.w3(32'h384cbe1b),
	.w4(32'hb80304c9),
	.w5(32'h392dd348),
	.w6(32'h38e533dd),
	.w7(32'h387486de),
	.w8(32'h397e3cac),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bcd9c),
	.w1(32'hb982f5a8),
	.w2(32'hba260089),
	.w3(32'hbaddf151),
	.w4(32'h3a3d6f86),
	.w5(32'h399a8820),
	.w6(32'hba75a25d),
	.w7(32'h3a44cd3b),
	.w8(32'h3a79669a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e8e533),
	.w1(32'h378dd100),
	.w2(32'h38ffc311),
	.w3(32'h37ebf0ef),
	.w4(32'h378a1155),
	.w5(32'h38f960df),
	.w6(32'h38d94335),
	.w7(32'h38c720c3),
	.w8(32'h39449053),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeccee7),
	.w1(32'hbb4d754d),
	.w2(32'hbb115662),
	.w3(32'hbb9f3df0),
	.w4(32'hbb328d1d),
	.w5(32'hbaba7b50),
	.w6(32'hbb348546),
	.w7(32'hb9a332f7),
	.w8(32'h3b4e971b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7130fb),
	.w1(32'hbc024aea),
	.w2(32'hbbc2effb),
	.w3(32'hbc210441),
	.w4(32'hbb391a4a),
	.w5(32'hba8cd722),
	.w6(32'hbc04645f),
	.w7(32'hbb27fdef),
	.w8(32'h3b44dfe7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb275fe8),
	.w1(32'hbb39d7d4),
	.w2(32'hbb72eed5),
	.w3(32'hbb46784e),
	.w4(32'hbae7e46f),
	.w5(32'hbb823b26),
	.w6(32'hbb05ee65),
	.w7(32'hbb4504ea),
	.w8(32'hbbd5f137),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32da5b),
	.w1(32'hb9522d90),
	.w2(32'hbb23955e),
	.w3(32'hbae24c21),
	.w4(32'h3afbddaa),
	.w5(32'h393a8523),
	.w6(32'hbb1234cf),
	.w7(32'h3b0d2180),
	.w8(32'h3ad8cb6c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895fa2),
	.w1(32'hbb1cfa0a),
	.w2(32'hbac2398e),
	.w3(32'hbb3a961e),
	.w4(32'hbb35f8a7),
	.w5(32'h3933f724),
	.w6(32'hbb2aef5a),
	.w7(32'hba023dae),
	.w8(32'h3b7e9708),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65bb3c),
	.w1(32'hb97cb28d),
	.w2(32'hbb02fce9),
	.w3(32'hba2b904c),
	.w4(32'h3aec4aa8),
	.w5(32'hb86f9bf1),
	.w6(32'h39522882),
	.w7(32'h3ad15e48),
	.w8(32'h36b2a376),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb34241),
	.w1(32'hbb20faea),
	.w2(32'hbb36b424),
	.w3(32'hbb7b1719),
	.w4(32'hbaaf7cd0),
	.w5(32'hbaf745ae),
	.w6(32'hbb2d8bbe),
	.w7(32'h3a853c20),
	.w8(32'h3aafe9c9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69fc873),
	.w1(32'h3711a3b4),
	.w2(32'h378746ca),
	.w3(32'hb70cf19b),
	.w4(32'h36d5a1a4),
	.w5(32'h37bc09da),
	.w6(32'h37b29bbf),
	.w7(32'h379906fd),
	.w8(32'h38213f6f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81484cb),
	.w1(32'hb85ccfdd),
	.w2(32'hb846e587),
	.w3(32'hb6c27e80),
	.w4(32'hb722e5f3),
	.w5(32'hb6149211),
	.w6(32'hb846a1c1),
	.w7(32'hb7c16b42),
	.w8(32'hb7a06337),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38935cfb),
	.w1(32'h37af5423),
	.w2(32'h391e7ae7),
	.w3(32'h391f5f4c),
	.w4(32'h37be97a6),
	.w5(32'h392ebbea),
	.w6(32'h38dda8a7),
	.w7(32'h380f1d57),
	.w8(32'h38f3fa20),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8950cf),
	.w1(32'h39b3a6db),
	.w2(32'hb975ff41),
	.w3(32'h39be300c),
	.w4(32'hb998f410),
	.w5(32'hba990350),
	.w6(32'h39b2827a),
	.w7(32'hba263af1),
	.w8(32'hbaac2320),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38d322),
	.w1(32'h3ab40e0d),
	.w2(32'hbb31951c),
	.w3(32'hb9b465e0),
	.w4(32'h3aee8090),
	.w5(32'hbae88698),
	.w6(32'hbaca973a),
	.w7(32'hb901ea79),
	.w8(32'hbbb0cc68),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a07493),
	.w1(32'h3a5e1893),
	.w2(32'h39a0b545),
	.w3(32'h388bb83c),
	.w4(32'h39e99cdd),
	.w5(32'hb8c6f2d4),
	.w6(32'hb949c027),
	.w7(32'h39a8012a),
	.w8(32'hb9967762),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5837cb),
	.w1(32'hb9ad0c68),
	.w2(32'h3957a975),
	.w3(32'hbad27b47),
	.w4(32'hba3514a7),
	.w5(32'h3a80aa9d),
	.w6(32'hbaf19c6e),
	.w7(32'h39a50200),
	.w8(32'hba5aec5a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc258eb7),
	.w1(32'hbb90592b),
	.w2(32'hbbcff06c),
	.w3(32'hbbeba70a),
	.w4(32'hba769f4e),
	.w5(32'hbb1c16e0),
	.w6(32'hbbfbad97),
	.w7(32'h3a4df3ae),
	.w8(32'h3b1fbdd9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0df688),
	.w1(32'h3b19978f),
	.w2(32'hbb371027),
	.w3(32'h3b85ec96),
	.w4(32'hba0aa6f2),
	.w5(32'hbc1113e1),
	.w6(32'h3b701523),
	.w7(32'hbae6186a),
	.w8(32'hbc2048ac),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc035b35),
	.w1(32'hbba10ef6),
	.w2(32'hbb3814aa),
	.w3(32'hbb01be3f),
	.w4(32'hbaa5e53e),
	.w5(32'hb9f96305),
	.w6(32'hbb7a29dd),
	.w7(32'h3b86f955),
	.w8(32'h3b413dcc),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58e1da),
	.w1(32'hb9fae57d),
	.w2(32'hbb51996d),
	.w3(32'h3a3d1539),
	.w4(32'hbb29933f),
	.w5(32'hbbcbb3d9),
	.w6(32'hb9f044b9),
	.w7(32'hbb407b19),
	.w8(32'hbbc1f72e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b4118),
	.w1(32'h3a0f50b9),
	.w2(32'hbb07d899),
	.w3(32'hba9c7fc0),
	.w4(32'h3bbf1964),
	.w5(32'h3bb59821),
	.w6(32'hbb556b49),
	.w7(32'h3ba2ddf2),
	.w8(32'h3bcc1d06),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4de211),
	.w1(32'hb9ffbbd8),
	.w2(32'hbae52db3),
	.w3(32'hb9dd7146),
	.w4(32'h3a736e86),
	.w5(32'hb8d5611b),
	.w6(32'hba6a1bdc),
	.w7(32'h3a10ca18),
	.w8(32'hba98f934),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b587023),
	.w1(32'hba24eb26),
	.w2(32'hbb6411b1),
	.w3(32'h3a950482),
	.w4(32'hbabed743),
	.w5(32'hbbd6b0b6),
	.w6(32'h3a2b9c62),
	.w7(32'hbb83c08f),
	.w8(32'hbc2a5961),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9277736),
	.w1(32'hb8af110f),
	.w2(32'hb9bf4d9c),
	.w3(32'hb3f25a18),
	.w4(32'hb8d29436),
	.w5(32'hb9d06b28),
	.w6(32'h381476bd),
	.w7(32'hb8865d77),
	.w8(32'h3763fbd2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd13b96),
	.w1(32'hbb2df566),
	.w2(32'hbbbe9856),
	.w3(32'hbb44200c),
	.w4(32'h3b00965a),
	.w5(32'hb9f8eab3),
	.w6(32'hbb6c6ee3),
	.w7(32'h3b04339f),
	.w8(32'h3a1fec6b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb811184),
	.w1(32'hb98cef09),
	.w2(32'hbacf51b4),
	.w3(32'hbb35c528),
	.w4(32'hb99ad5b8),
	.w5(32'hbab31467),
	.w6(32'hbadd8ac2),
	.w7(32'h3b6367c5),
	.w8(32'h3b80a28c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85318c),
	.w1(32'hbc1e931a),
	.w2(32'hbbd4953c),
	.w3(32'hbc3d5dca),
	.w4(32'hbbaa58ec),
	.w5(32'h3a66ede0),
	.w6(32'hbc31e8e5),
	.w7(32'h3af22cb1),
	.w8(32'h3a5cb0a5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70aeeb),
	.w1(32'h3b646e6b),
	.w2(32'hbb7ccbb4),
	.w3(32'h3c2e7287),
	.w4(32'h3b4e3e3e),
	.w5(32'hbbbd8210),
	.w6(32'h3b72f53e),
	.w7(32'hbb289999),
	.w8(32'hbc4e95eb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81a5a3),
	.w1(32'h3910a2b9),
	.w2(32'hbb7fc693),
	.w3(32'hbae7945e),
	.w4(32'hbab1def9),
	.w5(32'hbb639bd5),
	.w6(32'hbb182e9b),
	.w7(32'hbabc44b0),
	.w8(32'hbbe71d30),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fd862),
	.w1(32'hbba40512),
	.w2(32'hbb0a1d24),
	.w3(32'hbb314762),
	.w4(32'hb951faa4),
	.w5(32'h3b2460d2),
	.w6(32'h39d07466),
	.w7(32'h3c038c5c),
	.w8(32'h3c156bae),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba8be1),
	.w1(32'h388259a5),
	.w2(32'hb7649f55),
	.w3(32'h3a1bfc31),
	.w4(32'h3947520a),
	.w5(32'hb66f8790),
	.w6(32'h39573f4f),
	.w7(32'hb88e0f23),
	.w8(32'h3806176b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad3762),
	.w1(32'hbc1e8b86),
	.w2(32'hbc768b3a),
	.w3(32'hbc1b1ab9),
	.w4(32'hbb18b793),
	.w5(32'hbb25d655),
	.w6(32'hbc0c5dea),
	.w7(32'hb9b27d4b),
	.w8(32'hbbe715d4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66a9af),
	.w1(32'hbaeea10e),
	.w2(32'hbb6c2a10),
	.w3(32'hbaea7986),
	.w4(32'hbb53764e),
	.w5(32'hbb8fd549),
	.w6(32'hbb1c9994),
	.w7(32'hbb1bceba),
	.w8(32'hbb680627),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e47571),
	.w1(32'hb884561d),
	.w2(32'hb985ad88),
	.w3(32'h3a019bd5),
	.w4(32'h37f45169),
	.w5(32'hb919e75c),
	.w6(32'h39fbe087),
	.w7(32'h34d82f8a),
	.w8(32'hb97b0805),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c6d3f),
	.w1(32'hbae2da13),
	.w2(32'hbac6a708),
	.w3(32'hbad43205),
	.w4(32'hbaa75d9b),
	.w5(32'hba221084),
	.w6(32'hbacec746),
	.w7(32'h39264a48),
	.w8(32'hba0aa699),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ddd01),
	.w1(32'hbb63310a),
	.w2(32'hbb99d1b9),
	.w3(32'hbb7b9057),
	.w4(32'hbb3a4cf3),
	.w5(32'hbb4db1e9),
	.w6(32'hbb6c9e76),
	.w7(32'hbadb1450),
	.w8(32'hbb031c87),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a147870),
	.w1(32'hba2056c4),
	.w2(32'hbb624b3e),
	.w3(32'hba30df4b),
	.w4(32'hba7cb80c),
	.w5(32'hbb728a44),
	.w6(32'hba4454b5),
	.w7(32'hbaf1d9e9),
	.w8(32'hbbc001df),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f4439),
	.w1(32'hba04e0c9),
	.w2(32'hbbbbd59e),
	.w3(32'h3ae968d0),
	.w4(32'h37cf6c60),
	.w5(32'hbbfdc6f0),
	.w6(32'h3b4d9837),
	.w7(32'hba96b05c),
	.w8(32'hbc270c91),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09904d),
	.w1(32'h3a4b6b23),
	.w2(32'hb809f1e9),
	.w3(32'h3a1a25e1),
	.w4(32'h3ad2b39c),
	.w5(32'hba30d81c),
	.w6(32'h3a15ce19),
	.w7(32'hb96a4805),
	.w8(32'hbb7f842c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b563ae1),
	.w1(32'h3b243bc5),
	.w2(32'h3a0d0f7f),
	.w3(32'h3a25a8ff),
	.w4(32'h3a56c9aa),
	.w5(32'h3b234a8c),
	.w6(32'hbb519478),
	.w7(32'h3aacdeea),
	.w8(32'h3b3f1853),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c51bd),
	.w1(32'hbb2db5f4),
	.w2(32'hbb5ca3c3),
	.w3(32'hbb43d9f3),
	.w4(32'h3abb7952),
	.w5(32'h3b276a9b),
	.w6(32'hbba5ab67),
	.w7(32'h3b1abd8e),
	.w8(32'h3b24481d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9525f5d),
	.w1(32'hb9897fb3),
	.w2(32'hbae1dba0),
	.w3(32'hb9aa2bd0),
	.w4(32'hb90ee412),
	.w5(32'hbad6f4ec),
	.w6(32'hba38cd4f),
	.w7(32'hb97cdfb9),
	.w8(32'hbb0c7282),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92aa24e),
	.w1(32'hb8f866e1),
	.w2(32'hb8093f10),
	.w3(32'hb8c8879a),
	.w4(32'hb8694b6d),
	.w5(32'h360174fe),
	.w6(32'hb88d3842),
	.w7(32'hb89bed8a),
	.w8(32'hb7531c01),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f5d8f),
	.w1(32'hb94d65e0),
	.w2(32'hb96d499e),
	.w3(32'hba11c783),
	.w4(32'h37d82269),
	.w5(32'h397f8406),
	.w6(32'hba5006af),
	.w7(32'hb996e3f5),
	.w8(32'hb9e48b60),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e980d),
	.w1(32'h3949d8c5),
	.w2(32'h3922b779),
	.w3(32'hb88f43bb),
	.w4(32'h38c733e8),
	.w5(32'h38b77941),
	.w6(32'h37b8a15c),
	.w7(32'h38a32ba7),
	.w8(32'h38c9fcde),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915a856),
	.w1(32'h3995bb10),
	.w2(32'h37a8da27),
	.w3(32'h3980b416),
	.w4(32'h3939ba18),
	.w5(32'h38bebeae),
	.w6(32'h38de1e8b),
	.w7(32'h394deadf),
	.w8(32'h38eeb739),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d5f330),
	.w1(32'h3a8d5e1d),
	.w2(32'hbae90aea),
	.w3(32'h39758cc3),
	.w4(32'h3ad590e4),
	.w5(32'hba0c449a),
	.w6(32'hb943d1a8),
	.w7(32'h3ae43532),
	.w8(32'hbaa6af96),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a5594),
	.w1(32'h38e5d612),
	.w2(32'hba44d791),
	.w3(32'h3a81bf45),
	.w4(32'h3a19392a),
	.w5(32'hba0c0e02),
	.w6(32'h3a59a7a7),
	.w7(32'h3a18880e),
	.w8(32'hb9d4977e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb823924),
	.w1(32'hbaf82e45),
	.w2(32'hbb058d5d),
	.w3(32'hbb508c01),
	.w4(32'hbb3742b2),
	.w5(32'hb9c5f64c),
	.w6(32'hbb1c4cb6),
	.w7(32'hb8da540b),
	.w8(32'h3b272bd8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63dc1f),
	.w1(32'hba2204aa),
	.w2(32'hbaad5a4b),
	.w3(32'h3a8d64f5),
	.w4(32'hbac26853),
	.w5(32'hbb9ac4ff),
	.w6(32'h3acf3ed2),
	.w7(32'hbb9308ff),
	.w8(32'hbc2ad82e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886e624),
	.w1(32'h381ea156),
	.w2(32'h386af24d),
	.w3(32'h38adee25),
	.w4(32'h38a8fbff),
	.w5(32'h3906c6ff),
	.w6(32'h39286649),
	.w7(32'h38eac7c6),
	.w8(32'h388916af),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986dc6f),
	.w1(32'h39239987),
	.w2(32'hb8a49254),
	.w3(32'h39cc5591),
	.w4(32'h397d105e),
	.w5(32'h38763e99),
	.w6(32'h39402b84),
	.w7(32'h38c3b127),
	.w8(32'hb8d10ba8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380cc7b9),
	.w1(32'h3871e01a),
	.w2(32'h38479926),
	.w3(32'h382a2abb),
	.w4(32'h38974eeb),
	.w5(32'h385665ff),
	.w6(32'h384ea2f0),
	.w7(32'h38953d1b),
	.w8(32'h386353ee),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11ec37),
	.w1(32'hb8a18c7d),
	.w2(32'hb8b01eed),
	.w3(32'h393b5bdd),
	.w4(32'hba19a00b),
	.w5(32'hb9f72df4),
	.w6(32'hb95c5d88),
	.w7(32'hba5a7afe),
	.w8(32'hba8490e7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93a324),
	.w1(32'hbc02cbbb),
	.w2(32'hbb066b8b),
	.w3(32'hbbbe222b),
	.w4(32'hbc1d601b),
	.w5(32'h39ffa5e0),
	.w6(32'hbb9fc89c),
	.w7(32'hbb7d397e),
	.w8(32'h3afdff82),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6c3b1),
	.w1(32'hbb0a3444),
	.w2(32'hbb72f747),
	.w3(32'hbb69f97b),
	.w4(32'h3a564c6e),
	.w5(32'h398918b8),
	.w6(32'hbb52f373),
	.w7(32'h3b497275),
	.w8(32'h3b2fa3d4),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa97d0b),
	.w1(32'hba02739d),
	.w2(32'hba05fdf6),
	.w3(32'hb992e6cc),
	.w4(32'hb8c80c07),
	.w5(32'hb8d9ad63),
	.w6(32'hb986eba6),
	.w7(32'h3a067fe9),
	.w8(32'h3a531c20),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa437f),
	.w1(32'hba36c6dd),
	.w2(32'hbac49d95),
	.w3(32'hbaf5dec5),
	.w4(32'hb9879f62),
	.w5(32'h378cd9e9),
	.w6(32'hbb09e3cb),
	.w7(32'h3976ba8b),
	.w8(32'hb9a9fc92),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39693287),
	.w1(32'hb74c9c02),
	.w2(32'hba858d81),
	.w3(32'hb7991350),
	.w4(32'h3947b571),
	.w5(32'hba61f4ad),
	.w6(32'h39c28429),
	.w7(32'h3973910c),
	.w8(32'hbac77db7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27f6ba),
	.w1(32'hb9ed7102),
	.w2(32'hbabc3988),
	.w3(32'hbace19bf),
	.w4(32'h3ab08893),
	.w5(32'h3a86b6b0),
	.w6(32'hbaa537b1),
	.w7(32'h3af5e926),
	.w8(32'h3af8fe24),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb902d90),
	.w1(32'hbae1a659),
	.w2(32'hbb85df1f),
	.w3(32'hbb56ed99),
	.w4(32'h3a2484c9),
	.w5(32'hba42df0a),
	.w6(32'hba826843),
	.w7(32'h3a1e3d39),
	.w8(32'hbb076ccd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24b5f9),
	.w1(32'hbbb201cd),
	.w2(32'hbba82c72),
	.w3(32'hbbe752fd),
	.w4(32'hbb0618f4),
	.w5(32'hba40ea08),
	.w6(32'hbbb7ece4),
	.w7(32'h3b3ec6bc),
	.w8(32'h3ba9afa3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae524a0),
	.w1(32'h392f2694),
	.w2(32'hb954a0a2),
	.w3(32'h3a5d2f88),
	.w4(32'h39a0feb7),
	.w5(32'hbac6f096),
	.w6(32'h3a5c2f2e),
	.w7(32'hbafc2582),
	.w8(32'hbbb5c78a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a1662),
	.w1(32'hbac2b433),
	.w2(32'hba9ef115),
	.w3(32'hbacf1a68),
	.w4(32'h3aa61cdb),
	.w5(32'h3ad13216),
	.w6(32'hbb204e83),
	.w7(32'h3ac0113b),
	.w8(32'h39b6aa36),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd68c4),
	.w1(32'hbb663cca),
	.w2(32'hbb3193f8),
	.w3(32'hbb7dc9ff),
	.w4(32'hba51aee8),
	.w5(32'hba01265a),
	.w6(32'hbad63a5c),
	.w7(32'h3b69bc35),
	.w8(32'h3b91bfd5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0bc5d),
	.w1(32'h3a07c1bc),
	.w2(32'hba905cb4),
	.w3(32'hba3928f8),
	.w4(32'h39eeb9e6),
	.w5(32'h3983c672),
	.w6(32'hbb121fde),
	.w7(32'h3a142b3c),
	.w8(32'hbaa26bd6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25feb8),
	.w1(32'hbac6d62f),
	.w2(32'hbb0fd851),
	.w3(32'hba83f3d9),
	.w4(32'hb9f8c319),
	.w5(32'hb923c907),
	.w6(32'hbae2d840),
	.w7(32'h3a2fb31b),
	.w8(32'h3ac2b7ab),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d95d6),
	.w1(32'hb9a21b40),
	.w2(32'hba586aac),
	.w3(32'hb9b63891),
	.w4(32'hb86525cd),
	.w5(32'hba22ad03),
	.w6(32'hb9f2c165),
	.w7(32'hb92ffcb1),
	.w8(32'hba76bd94),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68b1ce),
	.w1(32'h39f744ff),
	.w2(32'hb9c68ce2),
	.w3(32'h3bbbef04),
	.w4(32'hbba6f9b4),
	.w5(32'hbc1dbc0e),
	.w6(32'h3b8a0e16),
	.w7(32'hbc0ca508),
	.w8(32'hbc7ec808),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa74b11),
	.w1(32'h39a2f63b),
	.w2(32'hba0074a8),
	.w3(32'hbadc12d9),
	.w4(32'h3a97e494),
	.w5(32'h3989df4e),
	.w6(32'hbadac64f),
	.w7(32'h3a565cc3),
	.w8(32'hba2939c1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916a736),
	.w1(32'hb8db3eb4),
	.w2(32'hb81ff4d4),
	.w3(32'hb971ce9f),
	.w4(32'hb943d246),
	.w5(32'h376c3e0e),
	.w6(32'hb980519b),
	.w7(32'hb8f8f637),
	.w8(32'h38957d2b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e4039),
	.w1(32'hb86e3372),
	.w2(32'h37f99c8a),
	.w3(32'h390d5e79),
	.w4(32'hb82577cf),
	.w5(32'h3786593b),
	.w6(32'h3963c181),
	.w7(32'hb83cfeaa),
	.w8(32'hb81a7ec2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6c18d),
	.w1(32'hba29e072),
	.w2(32'hba98b34a),
	.w3(32'hbaa80a78),
	.w4(32'hba0ea067),
	.w5(32'hb914c939),
	.w6(32'hba92e3d9),
	.w7(32'hb7185bf2),
	.w8(32'hb93b41c8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b19b0),
	.w1(32'hba828326),
	.w2(32'hbb39fc3c),
	.w3(32'h38f953ff),
	.w4(32'h3a47b9c4),
	.w5(32'hbb2fb25f),
	.w6(32'hb940e33c),
	.w7(32'hbaa4ca64),
	.w8(32'hbbf22a17),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912f59),
	.w1(32'hba278e0e),
	.w2(32'hbb30f4cd),
	.w3(32'hbbc97b5b),
	.w4(32'hbb2e3167),
	.w5(32'hbb2bd23d),
	.w6(32'hbb992cb8),
	.w7(32'hbafe634c),
	.w8(32'hbb3e28ba),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377ebeaa),
	.w1(32'hb6edd005),
	.w2(32'hb695cb93),
	.w3(32'h360cd7c6),
	.w4(32'h372c2b0c),
	.w5(32'h37f6246c),
	.w6(32'hb7d8bcca),
	.w7(32'hb5f0c8ca),
	.w8(32'h384e30f7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95ab75),
	.w1(32'hbadfed34),
	.w2(32'hbb887ee1),
	.w3(32'hbb359f32),
	.w4(32'hba008fd4),
	.w5(32'hbacd42c6),
	.w6(32'hbb5e0086),
	.w7(32'hba3f6c24),
	.w8(32'hb91e2a74),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb5224),
	.w1(32'hbaf6b6c1),
	.w2(32'hbb0223d2),
	.w3(32'hbaf96f90),
	.w4(32'hbaf41623),
	.w5(32'hbace9013),
	.w6(32'hbb275c43),
	.w7(32'hbafb3615),
	.w8(32'hbb39b097),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15a858),
	.w1(32'hbb93533b),
	.w2(32'hbb68455a),
	.w3(32'hbb701900),
	.w4(32'hbb430c66),
	.w5(32'hba2f45cb),
	.w6(32'hbb40170b),
	.w7(32'h3a9c679e),
	.w8(32'h3ba1ec0e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b4270),
	.w1(32'hbb32f86b),
	.w2(32'hbbddb20e),
	.w3(32'h3ab33190),
	.w4(32'h3a86662e),
	.w5(32'hbbcec544),
	.w6(32'h3bb647a6),
	.w7(32'h3a66b64c),
	.w8(32'hbbbb18f7),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf41f3),
	.w1(32'h39862fba),
	.w2(32'hba810042),
	.w3(32'h39665a26),
	.w4(32'h3960e36e),
	.w5(32'hbae777b5),
	.w6(32'h38abd990),
	.w7(32'h38c0f3ac),
	.w8(32'hbb0b77cf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a087225),
	.w1(32'h39b4809a),
	.w2(32'h39b6839e),
	.w3(32'h39849ea6),
	.w4(32'h392d746d),
	.w5(32'hb8d207af),
	.w6(32'h387350ce),
	.w7(32'hb8d9a887),
	.w8(32'hba06c91a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8699a0),
	.w1(32'h3b2e0dc7),
	.w2(32'h3990d8e0),
	.w3(32'h3b9badbd),
	.w4(32'h3b5fc3ad),
	.w5(32'h3a43fe40),
	.w6(32'h3b4d53ff),
	.w7(32'h3b4155d7),
	.w8(32'hb9d6fce8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0feca8),
	.w1(32'h3ae26f03),
	.w2(32'hbb17ce19),
	.w3(32'h3b0ec9ee),
	.w4(32'h3b293113),
	.w5(32'hbaf6a448),
	.w6(32'h3904d6ae),
	.w7(32'h3a9e061b),
	.w8(32'hbb81cca0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b8435),
	.w1(32'h3af6f634),
	.w2(32'hba42c19d),
	.w3(32'h3b110517),
	.w4(32'h3a879e00),
	.w5(32'hbb04a33d),
	.w6(32'h3a661bcd),
	.w7(32'h3989dfd9),
	.w8(32'hbb599da8),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fe891),
	.w1(32'hba84af96),
	.w2(32'hba0154c3),
	.w3(32'hbaa3d72e),
	.w4(32'hba1f7b73),
	.w5(32'hb924ea2f),
	.w6(32'hba7d474d),
	.w7(32'h3a026780),
	.w8(32'h3a8ce7e3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f29d92),
	.w1(32'hb91193f7),
	.w2(32'hb9243ad1),
	.w3(32'h3893a7bf),
	.w4(32'hb89df81a),
	.w5(32'hb813397e),
	.w6(32'hb7d35712),
	.w7(32'h3915b0c9),
	.w8(32'hb8bf2de5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bcfd1),
	.w1(32'hbb43d157),
	.w2(32'hbb3a01c9),
	.w3(32'hbac9de5b),
	.w4(32'h3906afa6),
	.w5(32'h3a7d8e41),
	.w6(32'hbb119678),
	.w7(32'h3a59d207),
	.w8(32'h3aec4271),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10c88a),
	.w1(32'hba705ef7),
	.w2(32'hba6ad7f7),
	.w3(32'hba0e8459),
	.w4(32'hba4e2bf9),
	.w5(32'hbaa14566),
	.w6(32'h3a3208a1),
	.w7(32'h393b1d07),
	.w8(32'hb8daa59d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b349329),
	.w1(32'h3a93d2d7),
	.w2(32'hba07789f),
	.w3(32'h3a74fc54),
	.w4(32'h39513e73),
	.w5(32'hb99fb29f),
	.w6(32'h39eaf3ef),
	.w7(32'h39ae36b1),
	.w8(32'hbac3fea4),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980b3e3),
	.w1(32'h38e74492),
	.w2(32'hb9777810),
	.w3(32'h399d5946),
	.w4(32'h397ede67),
	.w5(32'hb9055d15),
	.w6(32'h3974f967),
	.w7(32'h39737155),
	.w8(32'hb870cfac),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16a8bf),
	.w1(32'hba31439c),
	.w2(32'hbb331703),
	.w3(32'hbade8ff0),
	.w4(32'hbb597c36),
	.w5(32'hbb9a13f2),
	.w6(32'hbb037ec8),
	.w7(32'hbb58502e),
	.w8(32'hbbb3961a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38810dc7),
	.w1(32'h35a7a157),
	.w2(32'h37a8c6d3),
	.w3(32'h38ec1a04),
	.w4(32'h380c5b99),
	.w5(32'h381bac50),
	.w6(32'h391e0bf8),
	.w7(32'h38a5ae90),
	.w8(32'h386e6067),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97dfa19),
	.w1(32'hb90c7cd4),
	.w2(32'hb9a3c15e),
	.w3(32'hb8b44aed),
	.w4(32'hb721134c),
	.w5(32'hb94c7771),
	.w6(32'hb762c214),
	.w7(32'h37997ce8),
	.w8(32'hb8f5fd76),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53e335),
	.w1(32'h3a37109b),
	.w2(32'hbadf28cb),
	.w3(32'h3b3cc031),
	.w4(32'h3a965f50),
	.w5(32'hbb04173e),
	.w6(32'h3b291527),
	.w7(32'hb87b4497),
	.w8(32'hbb7a4d7f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac1e8d),
	.w1(32'hbb8cb1ef),
	.w2(32'hbb99510f),
	.w3(32'hbb757a77),
	.w4(32'hbb3f2c01),
	.w5(32'hbb372f02),
	.w6(32'hbbb2a285),
	.w7(32'hb9a98ab9),
	.w8(32'hb9eabdb6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa77e0),
	.w1(32'h3a9bd37e),
	.w2(32'hb9d40f5c),
	.w3(32'h3a64008a),
	.w4(32'h3a4be193),
	.w5(32'hba68f629),
	.w6(32'hb94ec547),
	.w7(32'h39d38440),
	.w8(32'hba565b0d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1629c),
	.w1(32'hb9a9e221),
	.w2(32'hbaf0f533),
	.w3(32'hba0cdb2c),
	.w4(32'hba693c1f),
	.w5(32'hbb26fd26),
	.w6(32'hb8eeaee0),
	.w7(32'hbae7f627),
	.w8(32'hbbb24f73),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a738373),
	.w1(32'h3a1ad713),
	.w2(32'hba7856fb),
	.w3(32'hb9d4527f),
	.w4(32'hb983fd03),
	.w5(32'hba9fed6c),
	.w6(32'h3a91a645),
	.w7(32'h3aaa588a),
	.w8(32'h3a6acaec),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcb6d3),
	.w1(32'h39e85cd5),
	.w2(32'hbb7a25a3),
	.w3(32'hbbba6ead),
	.w4(32'h3b67dead),
	.w5(32'hbb1e6505),
	.w6(32'hbb3a448c),
	.w7(32'h3bde52f8),
	.w8(32'h3b1fad9b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a9033),
	.w1(32'h38aeec06),
	.w2(32'hbba2257e),
	.w3(32'hba6cb6f4),
	.w4(32'h3b2dc5c0),
	.w5(32'hb97b989d),
	.w6(32'hba6b07d9),
	.w7(32'h3a9f4b43),
	.w8(32'h39829891),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe444a9),
	.w1(32'hbb3ba88c),
	.w2(32'hbb7f1c11),
	.w3(32'hbb9e31fe),
	.w4(32'h39818425),
	.w5(32'hb9db04a3),
	.w6(32'hbb866699),
	.w7(32'h3b173933),
	.w8(32'h3af549cf),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398daa02),
	.w1(32'h388c8b13),
	.w2(32'hb7249773),
	.w3(32'h39604164),
	.w4(32'h3932c382),
	.w5(32'h38f89adf),
	.w6(32'h398f767e),
	.w7(32'h390c18b1),
	.w8(32'h3892293e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae79118),
	.w1(32'hb997239b),
	.w2(32'hba71bc6f),
	.w3(32'hba7f0479),
	.w4(32'h3aaf5b82),
	.w5(32'h3ac82d62),
	.w6(32'hb91d6af6),
	.w7(32'h3b361e09),
	.w8(32'h3b657c93),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b42fc0),
	.w1(32'h3745b161),
	.w2(32'h38c25808),
	.w3(32'hb6a8a535),
	.w4(32'h33cf9dad),
	.w5(32'h38b7afe4),
	.w6(32'h382251fd),
	.w7(32'h38113a88),
	.w8(32'h390de272),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b973e),
	.w1(32'h3a162acd),
	.w2(32'h398bd377),
	.w3(32'hba0b78b2),
	.w4(32'h3a1de0b6),
	.w5(32'h388d5db8),
	.w6(32'hba9a2364),
	.w7(32'hb963de43),
	.w8(32'hb9612582),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8596c52),
	.w1(32'hb8053150),
	.w2(32'h398a874f),
	.w3(32'hba453b3c),
	.w4(32'hb6975a5f),
	.w5(32'hb9ca0632),
	.w6(32'h38c5694e),
	.w7(32'hb9b7c8a8),
	.w8(32'hba308031),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56c828),
	.w1(32'h398e10e6),
	.w2(32'hbab1f40d),
	.w3(32'hbb79da49),
	.w4(32'h3adc7f6f),
	.w5(32'h3a69770d),
	.w6(32'hbba3cb44),
	.w7(32'h3ae6957f),
	.w8(32'h3a4d80a9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710b4ff),
	.w1(32'hb6466dab),
	.w2(32'h37ea6f6f),
	.w3(32'hb6bc8873),
	.w4(32'hb77c6fcc),
	.w5(32'h37b42b63),
	.w6(32'hb49dcaa0),
	.w7(32'h36ee5fb8),
	.w8(32'h3806cdd9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ff644),
	.w1(32'hb742ffdf),
	.w2(32'h37e81153),
	.w3(32'hb82f9ab8),
	.w4(32'h37a11251),
	.w5(32'h37922d3c),
	.w6(32'h36d1111d),
	.w7(32'h375818ce),
	.w8(32'h3791f3b6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eca2c),
	.w1(32'hba06a7c3),
	.w2(32'hba98a10e),
	.w3(32'h3a1223bc),
	.w4(32'h3978b994),
	.w5(32'h3a54c6a4),
	.w6(32'h3a8fbd45),
	.w7(32'h398b91ca),
	.w8(32'h39823de7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89573b),
	.w1(32'hb907c897),
	.w2(32'hbb319361),
	.w3(32'hbada8c3f),
	.w4(32'h3b0d17da),
	.w5(32'hb9b8a9a6),
	.w6(32'hb9b1d7ef),
	.w7(32'h3b2cfb7d),
	.w8(32'h3a586a8b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf55a2c),
	.w1(32'hbb8e36b8),
	.w2(32'hbb3ffc63),
	.w3(32'hbbb42177),
	.w4(32'hbb917b63),
	.w5(32'h3a91dbd6),
	.w6(32'hba999918),
	.w7(32'hba87e8c2),
	.w8(32'hbb5e5c42),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc4ee4),
	.w1(32'h393f690c),
	.w2(32'hb9b6899b),
	.w3(32'h3999e457),
	.w4(32'h3888cf0e),
	.w5(32'hb984d482),
	.w6(32'hb966d813),
	.w7(32'hb9661737),
	.w8(32'hb9612343),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42fc08),
	.w1(32'hbabcc39e),
	.w2(32'hbb9573aa),
	.w3(32'hbc2da447),
	.w4(32'h3acf2638),
	.w5(32'h3a9085a2),
	.w6(32'hbb84b8f9),
	.w7(32'h3bd942e8),
	.w8(32'h3bea0786),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c0105),
	.w1(32'h37ae4110),
	.w2(32'hbbe8d740),
	.w3(32'h3ad3ecb3),
	.w4(32'h3b9b2a15),
	.w5(32'hbaae6674),
	.w6(32'h3b9c579b),
	.w7(32'h3bd26d40),
	.w8(32'hbaddda7f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac82f2a),
	.w1(32'hbab75bec),
	.w2(32'hba852361),
	.w3(32'hb9efe51f),
	.w4(32'hbaedddd5),
	.w5(32'hba8e3248),
	.w6(32'hb9c52c6d),
	.w7(32'hba91640f),
	.w8(32'h39d09668),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f14e7c),
	.w1(32'hb7b2d8cd),
	.w2(32'h36fd5c9e),
	.w3(32'hb839c9ae),
	.w4(32'hb84db57a),
	.w5(32'h37e7de53),
	.w6(32'hb8e13a98),
	.w7(32'h364a2e51),
	.w8(32'h382441be),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8232a57),
	.w1(32'h3643726c),
	.w2(32'hb8594324),
	.w3(32'hb81513df),
	.w4(32'h3775f83f),
	.w5(32'hb847382f),
	.w6(32'hb79f9c3d),
	.w7(32'hb7c87925),
	.w8(32'hb88ea4f3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cf644a),
	.w1(32'h3739acee),
	.w2(32'h3864b6b5),
	.w3(32'h3725cb5c),
	.w4(32'h35e3b5d6),
	.w5(32'h384d6485),
	.w6(32'h37edf1a1),
	.w7(32'h379eab8e),
	.w8(32'h38779a62),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba866c83),
	.w1(32'hbb223527),
	.w2(32'hbae3e2d6),
	.w3(32'hba3b61f1),
	.w4(32'hbb71118b),
	.w5(32'hbaf93803),
	.w6(32'hba82f3ca),
	.w7(32'hbad4b910),
	.w8(32'hb9acee41),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15fac0),
	.w1(32'hba5d9a0d),
	.w2(32'hbaf7ca77),
	.w3(32'hbaa4875c),
	.w4(32'h39bbc913),
	.w5(32'hba892ca9),
	.w6(32'hba2c7046),
	.w7(32'h3a9144e5),
	.w8(32'hbb046b00),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826437),
	.w1(32'hbb2202f0),
	.w2(32'hbb92a689),
	.w3(32'hbb66f68a),
	.w4(32'hbacd81ee),
	.w5(32'hbb72719b),
	.w6(32'hbac694e5),
	.w7(32'hbb1dda12),
	.w8(32'hbbed516d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f27f7),
	.w1(32'h3a802efc),
	.w2(32'h3796e0f8),
	.w3(32'hb973b7a7),
	.w4(32'hb8e3b775),
	.w5(32'hba1a7b59),
	.w6(32'h37e47b2e),
	.w7(32'hb9129f77),
	.w8(32'hba81a9f6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb951763),
	.w1(32'hbb8cb3ce),
	.w2(32'hbbc1e7ae),
	.w3(32'hbb2dde00),
	.w4(32'hba7da9c9),
	.w5(32'hbb43f96a),
	.w6(32'hbb6dcf48),
	.w7(32'h389bcf67),
	.w8(32'hbaf81550),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ad71a),
	.w1(32'hbab8a599),
	.w2(32'hbb01942b),
	.w3(32'hbb020a59),
	.w4(32'hbb0cbb9d),
	.w5(32'hbabc47ed),
	.w6(32'hbaf4b23d),
	.w7(32'hba562738),
	.w8(32'hb9784103),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38055c74),
	.w1(32'h37a6623f),
	.w2(32'h38bc1473),
	.w3(32'h36f00a04),
	.w4(32'h35e76bca),
	.w5(32'h389f03ff),
	.w6(32'h383825b2),
	.w7(32'h37f6c04c),
	.w8(32'h38ca9db9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4724e6),
	.w1(32'hbb073ffa),
	.w2(32'hbb20064c),
	.w3(32'hbac66db3),
	.w4(32'h38380065),
	.w5(32'h3a15a0eb),
	.w6(32'hbb08ceb8),
	.w7(32'h3a59c094),
	.w8(32'h3ad259b9),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ad77b),
	.w1(32'h383c4dff),
	.w2(32'h395791d2),
	.w3(32'h38158a07),
	.w4(32'h37958f46),
	.w5(32'h3947fce3),
	.w6(32'h39075e19),
	.w7(32'h38a98cc2),
	.w8(32'h396e18c9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c24dd),
	.w1(32'hbaf41880),
	.w2(32'hbb68ca95),
	.w3(32'hbabc9d08),
	.w4(32'hb9bc9923),
	.w5(32'hbb03dc64),
	.w6(32'hbb031c90),
	.w7(32'hb9911f3f),
	.w8(32'hbb0de29d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c13042),
	.w1(32'h3af611e9),
	.w2(32'hbb7ffd0a),
	.w3(32'h39c64c3b),
	.w4(32'h3b2c9da4),
	.w5(32'hbb6af1d7),
	.w6(32'hba62e11b),
	.w7(32'h3a6b6bd0),
	.w8(32'hbbd915d3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e4ba6),
	.w1(32'h3a22c7d2),
	.w2(32'hbb3b03ad),
	.w3(32'h3ae63f08),
	.w4(32'h3adaced4),
	.w5(32'hbb15ed69),
	.w6(32'h3a307bc3),
	.w7(32'h3965bd18),
	.w8(32'hbb97afcd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96055f),
	.w1(32'h3a8e06df),
	.w2(32'hb98241ed),
	.w3(32'h3aaa97dd),
	.w4(32'h3a8da1e7),
	.w5(32'hb9bc6204),
	.w6(32'h3a287046),
	.w7(32'h3a0df2ab),
	.w8(32'hba20038a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33edcc),
	.w1(32'hba9f2dba),
	.w2(32'hbba1be7a),
	.w3(32'h3a8f346a),
	.w4(32'h3ac22b80),
	.w5(32'hbb4f95cd),
	.w6(32'h3af8316f),
	.w7(32'hb9dbada8),
	.w8(32'hbbff0923),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75f6d2),
	.w1(32'hbaf9c369),
	.w2(32'hbb0b0cc0),
	.w3(32'hbb495268),
	.w4(32'hb95eb730),
	.w5(32'h39aa8ce2),
	.w6(32'hbb75cbd3),
	.w7(32'h3a0883ba),
	.w8(32'h3b0fe4cd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf3dc7),
	.w1(32'hbaade4e2),
	.w2(32'hbb57dd07),
	.w3(32'hbc12fa5c),
	.w4(32'hbb3ab60e),
	.w5(32'hbb427a6d),
	.w6(32'hbbc0325d),
	.w7(32'hbb3fd6d6),
	.w8(32'hbb84566f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d6375d),
	.w1(32'h3746eabc),
	.w2(32'h38b485ff),
	.w3(32'hb6d344b5),
	.w4(32'hb8003421),
	.w5(32'h3821bf7b),
	.w6(32'h38056f72),
	.w7(32'hb6c6818f),
	.w8(32'h387b3082),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39864607),
	.w1(32'h38db2e26),
	.w2(32'h3761a52f),
	.w3(32'hb904612a),
	.w4(32'hb9828b41),
	.w5(32'hba011550),
	.w6(32'hb8633d8c),
	.w7(32'hb7af6851),
	.w8(32'hb8dcf9e3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f1b54),
	.w1(32'hbb5ac8e5),
	.w2(32'hbbb2f0b6),
	.w3(32'hbafd77c6),
	.w4(32'hba09ecee),
	.w5(32'hb801d596),
	.w6(32'hbb316090),
	.w7(32'h3a1a95f2),
	.w8(32'hba6c00ab),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d195c),
	.w1(32'hbb030954),
	.w2(32'hbb904023),
	.w3(32'hbb026a24),
	.w4(32'hb9c96b58),
	.w5(32'hbae293ef),
	.w6(32'hbbb17a43),
	.w7(32'h393427e2),
	.w8(32'hbab316fe),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf0b09),
	.w1(32'h39deb6c3),
	.w2(32'hbb4bc458),
	.w3(32'hb9416939),
	.w4(32'h3ad9827a),
	.w5(32'hb9458840),
	.w6(32'hba84e202),
	.w7(32'h3ab96930),
	.w8(32'hbae23c75),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb322c54),
	.w1(32'hbac012d0),
	.w2(32'h3b06cd8f),
	.w3(32'hbb9e1ea1),
	.w4(32'hbba8c4fe),
	.w5(32'hba8b52b2),
	.w6(32'hba9542aa),
	.w7(32'h3b277d6f),
	.w8(32'h3c051b3b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bd57d),
	.w1(32'hb9966a00),
	.w2(32'hb9315c4f),
	.w3(32'hba472eff),
	.w4(32'hb9a7cc4a),
	.w5(32'h3a140837),
	.w6(32'hba89b536),
	.w7(32'hb9990c9f),
	.w8(32'h3a4709d0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1cfe4),
	.w1(32'hba8ae28e),
	.w2(32'hba0d0c84),
	.w3(32'hba6b8555),
	.w4(32'hb9811ec2),
	.w5(32'h3aa9b630),
	.w6(32'hba3100ee),
	.w7(32'h399ad5b6),
	.w8(32'h3a8220ab),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9313a7),
	.w1(32'hbbc8987a),
	.w2(32'hbb96e646),
	.w3(32'hbb97e201),
	.w4(32'hbbe6756f),
	.w5(32'hbbe27bb4),
	.w6(32'hbb798f4c),
	.w7(32'hbb20f602),
	.w8(32'hbb587d24),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc335632),
	.w1(32'hbb8ffeeb),
	.w2(32'hbbcac821),
	.w3(32'hbc0f0ac6),
	.w4(32'hbab1db86),
	.w5(32'hba4349ce),
	.w6(32'hbbcdf1df),
	.w7(32'h3b109528),
	.w8(32'h3b6e22a4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27fb31),
	.w1(32'hbbaedd65),
	.w2(32'hbb2489e8),
	.w3(32'hbbbcf68e),
	.w4(32'hbb4f0a3c),
	.w5(32'hba5c2d8c),
	.w6(32'hbbc7888c),
	.w7(32'h3a9ff062),
	.w8(32'h3ac0a518),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea28e6),
	.w1(32'h3b5e758a),
	.w2(32'h39629462),
	.w3(32'h3b2b3e8e),
	.w4(32'h39f84b93),
	.w5(32'hbb4e7ddd),
	.w6(32'h3a9218cb),
	.w7(32'hbad5fb62),
	.w8(32'hbbcb8de0),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a842b4a),
	.w1(32'hb9adc985),
	.w2(32'hbb8d3c58),
	.w3(32'h3ad0876a),
	.w4(32'h3ade31a8),
	.w5(32'hbb78ea7a),
	.w6(32'h3b057a2e),
	.w7(32'hba875534),
	.w8(32'hbbe9f308),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a578ca),
	.w1(32'h37ce62f5),
	.w2(32'h385069c1),
	.w3(32'h3745a4dc),
	.w4(32'h37a7ba98),
	.w5(32'h38298536),
	.w6(32'h380e6f5d),
	.w7(32'h38027978),
	.w8(32'h3830aad4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382771eb),
	.w1(32'h379139c6),
	.w2(32'h385509f3),
	.w3(32'h37d4187f),
	.w4(32'h375e99d1),
	.w5(32'h3860f1df),
	.w6(32'h381b4c04),
	.w7(32'h37e4ca39),
	.w8(32'h38899ff5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d93fdc),
	.w1(32'h39a2698a),
	.w2(32'h3a45f592),
	.w3(32'h39fb2fcc),
	.w4(32'h39b8e245),
	.w5(32'h3a93ca99),
	.w6(32'h3a079b01),
	.w7(32'h3a17b1e2),
	.w8(32'h3a51b7cc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37894544),
	.w1(32'hb6777f40),
	.w2(32'h3883e376),
	.w3(32'hb53dd2ff),
	.w4(32'hb76aa87c),
	.w5(32'h38534c32),
	.w6(32'h380abd6c),
	.w7(32'h37539d04),
	.w8(32'h389a667d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5484ab),
	.w1(32'hbaf5c465),
	.w2(32'hbb1220d5),
	.w3(32'hba7b586f),
	.w4(32'hbb3d1fe1),
	.w5(32'hbb37d72d),
	.w6(32'hba9a1998),
	.w7(32'hbabc4621),
	.w8(32'hba9cf12f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4eb0a),
	.w1(32'hbb106cef),
	.w2(32'hbb08bc50),
	.w3(32'hb7911a55),
	.w4(32'hba5e698a),
	.w5(32'h3abf7faf),
	.w6(32'hbb328ea0),
	.w7(32'hb98787a8),
	.w8(32'h3ab5078c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983b998),
	.w1(32'h391364f2),
	.w2(32'hba935e00),
	.w3(32'hb93a15c5),
	.w4(32'h39ccc3b7),
	.w5(32'hba481b85),
	.w6(32'h395bee07),
	.w7(32'h376ba29c),
	.w8(32'hbadda79d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38038de9),
	.w1(32'h37fb99ec),
	.w2(32'h383e6ecc),
	.w3(32'h38063bf6),
	.w4(32'h3857c4f0),
	.w5(32'h38a11744),
	.w6(32'h381a407f),
	.w7(32'h3848260c),
	.w8(32'h38820121),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73e95c),
	.w1(32'hbc0b6eaa),
	.w2(32'hbbc6ff49),
	.w3(32'hbc0d0f18),
	.w4(32'hbb722cf9),
	.w5(32'hb9f47c89),
	.w6(32'hbc010915),
	.w7(32'h3b27002e),
	.w8(32'h3bd11894),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb968418),
	.w1(32'hbae96ae1),
	.w2(32'hbaa40964),
	.w3(32'hbb2356ff),
	.w4(32'h39e5f7e4),
	.w5(32'h3a838bbe),
	.w6(32'hbb2ddd81),
	.w7(32'h3a1b4449),
	.w8(32'h3aebef5a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383c9b1c),
	.w1(32'hb9990e4a),
	.w2(32'hb94981a1),
	.w3(32'hb8bd761e),
	.w4(32'hba1519ac),
	.w5(32'hb99ff71b),
	.w6(32'hb8baee5b),
	.w7(32'hb9f78599),
	.w8(32'hba0a921c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eb7dc),
	.w1(32'hbb2cec64),
	.w2(32'hbb051d3f),
	.w3(32'hbb3020d4),
	.w4(32'hbab1e42c),
	.w5(32'hb97f936f),
	.w6(32'hbb2c3657),
	.w7(32'h39ef27e0),
	.w8(32'h3b2f10c1),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390fc284),
	.w1(32'h38b5c186),
	.w2(32'h388a483e),
	.w3(32'h38cbf2c2),
	.w4(32'h3888cf44),
	.w5(32'h388ac6e4),
	.w6(32'h386e9a0d),
	.w7(32'hb7baefb6),
	.w8(32'h37c15c9b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951e619),
	.w1(32'hb9d71f9f),
	.w2(32'hb9e12977),
	.w3(32'hb905d4c2),
	.w4(32'hb94f815b),
	.w5(32'hb9097fc2),
	.w6(32'hb9e946e6),
	.w7(32'hb99b86ad),
	.w8(32'hb949cac4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36da36c7),
	.w1(32'h37fd594d),
	.w2(32'h38483861),
	.w3(32'h3818d77f),
	.w4(32'h385be8ac),
	.w5(32'h385ca6a9),
	.w6(32'h386d2055),
	.w7(32'h38308df2),
	.w8(32'h3852543d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a04eb6),
	.w1(32'h3854f769),
	.w2(32'h385434c6),
	.w3(32'h3804ac11),
	.w4(32'h37aa70a1),
	.w5(32'h38903ba2),
	.w6(32'h3871440c),
	.w7(32'h3868fb11),
	.w8(32'h390f4d98),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b446967),
	.w1(32'h3ab8ce84),
	.w2(32'hb9abd508),
	.w3(32'h3a3f2214),
	.w4(32'h38c3605a),
	.w5(32'hbade26d6),
	.w6(32'hb914c585),
	.w7(32'hba75f983),
	.w8(32'hbb2c84c6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8df0e1),
	.w1(32'hb8209757),
	.w2(32'hbb337406),
	.w3(32'hbb52778b),
	.w4(32'h3b150ee8),
	.w5(32'h3a1765df),
	.w6(32'hbb8093e4),
	.w7(32'h3ba26aac),
	.w8(32'h3b8c7354),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad597c),
	.w1(32'hbb1784df),
	.w2(32'hbb550d67),
	.w3(32'hbb023e0d),
	.w4(32'h3aa77287),
	.w5(32'h3a56bd03),
	.w6(32'hba9e3705),
	.w7(32'h3b430b80),
	.w8(32'h3b75b080),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcee5d8),
	.w1(32'hbb890bed),
	.w2(32'hbb79775e),
	.w3(32'hbbac4888),
	.w4(32'hbb04a629),
	.w5(32'hba4f5ed0),
	.w6(32'hbb7b16b8),
	.w7(32'h3ab9fe7e),
	.w8(32'h3b3ee28f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397160cd),
	.w1(32'h38c72cc7),
	.w2(32'h364cff45),
	.w3(32'h3958f55f),
	.w4(32'h392f8b3c),
	.w5(32'h3874b0e9),
	.w6(32'h392feade),
	.w7(32'h39028917),
	.w8(32'h38129557),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf2930),
	.w1(32'hb90e2e7d),
	.w2(32'h383ec2c5),
	.w3(32'hb90d5919),
	.w4(32'h394bf0b7),
	.w5(32'h3a65f650),
	.w6(32'hb94a6784),
	.w7(32'hb766db46),
	.w8(32'h39d5405d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb706197b),
	.w1(32'hb73b1b5c),
	.w2(32'h37ff4d0a),
	.w3(32'hb7b55b66),
	.w4(32'hb756e2b0),
	.w5(32'h37d7cee9),
	.w6(32'h372c4438),
	.w7(32'hb62f712c),
	.w8(32'h38248f24),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3869fe9d),
	.w1(32'h37d88583),
	.w2(32'h3838beb6),
	.w3(32'h3868ae40),
	.w4(32'h37ca3745),
	.w5(32'h38358da7),
	.w6(32'h3860e435),
	.w7(32'h3742e6bc),
	.w8(32'h3819f4a7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb82b2),
	.w1(32'hbad8cd42),
	.w2(32'hbb34a1a8),
	.w3(32'hbb10faa9),
	.w4(32'h3b75378e),
	.w5(32'h3b0514d9),
	.w6(32'hbaa851d8),
	.w7(32'h3b9063b7),
	.w8(32'h3b7d1786),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb787c1db),
	.w1(32'hb86c45de),
	.w2(32'hb863d619),
	.w3(32'hb7a18d24),
	.w4(32'hb870c632),
	.w5(32'hb8608ec7),
	.w6(32'hb7f92f15),
	.w7(32'hb847234e),
	.w8(32'hb7fd8d8f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cb60c),
	.w1(32'h3aa9aa56),
	.w2(32'hba6c3f61),
	.w3(32'h3a58cc10),
	.w4(32'h3a6d5d8f),
	.w5(32'hba990324),
	.w6(32'h396949a4),
	.w7(32'h3a28792e),
	.w8(32'hbaade12e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5b7e7),
	.w1(32'hba88c75b),
	.w2(32'hbb21604f),
	.w3(32'hbadd9475),
	.w4(32'hba1ec7db),
	.w5(32'hba52ab43),
	.w6(32'hbaa25e2b),
	.w7(32'h3a678866),
	.w8(32'h395cefb0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e4b9b0),
	.w1(32'h3702eb0b),
	.w2(32'h37a5a9e1),
	.w3(32'h37d4a798),
	.w4(32'h368fb341),
	.w5(32'h37e61a53),
	.w6(32'h35c15aee),
	.w7(32'hb6d3b6ab),
	.w8(32'h37c48834),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae184b4),
	.w1(32'hba1b7de8),
	.w2(32'hba7628a7),
	.w3(32'hbac97777),
	.w4(32'hb87324fb),
	.w5(32'hb9805e63),
	.w6(32'hb93bc326),
	.w7(32'h39bd0c4a),
	.w8(32'hb8c0ca78),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939ab27),
	.w1(32'hb972c966),
	.w2(32'hb9c90a4f),
	.w3(32'hb89797e4),
	.w4(32'hb8c781b5),
	.w5(32'hb936b4aa),
	.w6(32'hb9851c3c),
	.w7(32'hb87e2a4f),
	.w8(32'hb7052c43),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3275f),
	.w1(32'hba8d9d42),
	.w2(32'hbb8ae2f1),
	.w3(32'hbb95bb18),
	.w4(32'h3b9f20c7),
	.w5(32'h3b35f7da),
	.w6(32'hbb49cb45),
	.w7(32'h3c14d6cf),
	.w8(32'h3c1d6084),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371d062c),
	.w1(32'hbb08f912),
	.w2(32'hbb458965),
	.w3(32'hb8473aff),
	.w4(32'hbb0faf13),
	.w5(32'hbb498b0a),
	.w6(32'hbab20851),
	.w7(32'hbb3368ff),
	.w8(32'hb8ae8056),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5df25a),
	.w1(32'h3b1fc762),
	.w2(32'hbae3506c),
	.w3(32'hb9f03199),
	.w4(32'hbb26aad7),
	.w5(32'hbafd1c76),
	.w6(32'hbb9c5ce8),
	.w7(32'hbaf77fa7),
	.w8(32'hbb03ea08),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule