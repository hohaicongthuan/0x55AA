module layer_10_featuremap_140(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71278c),
	.w1(32'h39c77596),
	.w2(32'hb9ff6876),
	.w3(32'h3b4c80db),
	.w4(32'h3b6e20f0),
	.w5(32'h3b5349c1),
	.w6(32'hba417370),
	.w7(32'hbb117c5e),
	.w8(32'hbb909a64),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98795f),
	.w1(32'h39387877),
	.w2(32'hb8ea66f5),
	.w3(32'hba759fd8),
	.w4(32'h3a637f0a),
	.w5(32'h3978758e),
	.w6(32'h3a54f192),
	.w7(32'h37fa8658),
	.w8(32'hb8e77d0d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39406d57),
	.w1(32'h38ad9acf),
	.w2(32'h3a858e6b),
	.w3(32'h384f0d2d),
	.w4(32'h39f7f0b4),
	.w5(32'h3ab13276),
	.w6(32'hb9e5d097),
	.w7(32'h39acf1bf),
	.w8(32'h3a84f96a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad98463),
	.w1(32'h3b3547ee),
	.w2(32'h3b25fcb8),
	.w3(32'h3b02d640),
	.w4(32'h3a86382f),
	.w5(32'h3a3508a9),
	.w6(32'h3a83890f),
	.w7(32'h3b14df3f),
	.w8(32'h3aaf6ced),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b098c4c),
	.w1(32'hbaa89eb7),
	.w2(32'hbb60d599),
	.w3(32'hb9816296),
	.w4(32'hbb5ed33b),
	.w5(32'hbb39cf46),
	.w6(32'hbaadd40f),
	.w7(32'hbac2e4bb),
	.w8(32'hba8b1d34),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01fbf5),
	.w1(32'h3b5a9c15),
	.w2(32'h3b7bb4ba),
	.w3(32'hbb2ae17a),
	.w4(32'h3b1e6243),
	.w5(32'h3b46dcd4),
	.w6(32'h3b0f789e),
	.w7(32'h3b38a0e1),
	.w8(32'h3b1b7be6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80720e),
	.w1(32'h3b12676c),
	.w2(32'h3a180d1b),
	.w3(32'h3b56c372),
	.w4(32'h3b1341c5),
	.w5(32'h3a03d832),
	.w6(32'h3b2b6ad5),
	.w7(32'h3ae5331e),
	.w8(32'h3a6b8767),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af2fad),
	.w1(32'h3b1f8c61),
	.w2(32'h3b2088e8),
	.w3(32'h38fc10a5),
	.w4(32'h3aaa05ec),
	.w5(32'h3b00fe69),
	.w6(32'h3afa1b9a),
	.w7(32'h3b0972d8),
	.w8(32'h3af185c7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a4100),
	.w1(32'h3affb32b),
	.w2(32'h3abeeda1),
	.w3(32'h3b19403c),
	.w4(32'h39e9d01e),
	.w5(32'h39e70ec9),
	.w6(32'h3a7ea9b0),
	.w7(32'h3a56be6a),
	.w8(32'h3a282bd0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5f60d),
	.w1(32'hbae6145e),
	.w2(32'hbb690987),
	.w3(32'h3a75e8eb),
	.w4(32'hba2f250a),
	.w5(32'hbb48c19f),
	.w6(32'h3902d41d),
	.w7(32'hbb0b5a9b),
	.w8(32'hbb178cc3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a94ee),
	.w1(32'h3a5e48e5),
	.w2(32'h39816a38),
	.w3(32'hbb5cd696),
	.w4(32'hbaa3b0ff),
	.w5(32'hba90f865),
	.w6(32'h3a43b6f7),
	.w7(32'h3abe274e),
	.w8(32'h38ce8093),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981d8b1),
	.w1(32'h3b15f5de),
	.w2(32'hb99f1a4e),
	.w3(32'hb9fc4c92),
	.w4(32'hba9300ca),
	.w5(32'hbaff118c),
	.w6(32'h3b98ef4a),
	.w7(32'h3b7d74d0),
	.w8(32'h3ad89ad9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4ed60),
	.w1(32'hbabdd45c),
	.w2(32'hb947fc54),
	.w3(32'hbb1c9daf),
	.w4(32'hba1fe2a0),
	.w5(32'h3913c785),
	.w6(32'hbb17d27c),
	.w7(32'hbacb56c3),
	.w8(32'hbab1617a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94bbf1e),
	.w1(32'h3adb1cf2),
	.w2(32'hb917e848),
	.w3(32'hb8b8c97b),
	.w4(32'h3a3d3fc9),
	.w5(32'hb9b5296d),
	.w6(32'h3b1466fc),
	.w7(32'h3ad4a153),
	.w8(32'h3a4d63c4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba447093),
	.w1(32'hb97d161d),
	.w2(32'hbb12722d),
	.w3(32'h3834eb81),
	.w4(32'hbb2df189),
	.w5(32'hbb2fd8a5),
	.w6(32'h3b3b273c),
	.w7(32'h3af4f61b),
	.w8(32'h3a7aecab),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a3b53),
	.w1(32'h3b162bfc),
	.w2(32'h3b34ac23),
	.w3(32'hbb30da52),
	.w4(32'h3a098f45),
	.w5(32'h3a8f598d),
	.w6(32'h3adfa906),
	.w7(32'h3ac2b424),
	.w8(32'h3ab95763),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcece6),
	.w1(32'h3a18df1e),
	.w2(32'hba220b3e),
	.w3(32'h3a2559ab),
	.w4(32'h3aa71e58),
	.w5(32'hbaae7b37),
	.w6(32'h39c5df29),
	.w7(32'hb90f2d8c),
	.w8(32'hba3164ea),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa6444),
	.w1(32'h3b3b9bf2),
	.w2(32'h3b1bbeff),
	.w3(32'hbaa34c26),
	.w4(32'h3b3f6d8c),
	.w5(32'h3ada7064),
	.w6(32'h3b55caa3),
	.w7(32'h3b1ce69b),
	.w8(32'h3acdbff8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae824ef),
	.w1(32'h38129c92),
	.w2(32'h3a01f109),
	.w3(32'h3a762dff),
	.w4(32'h39d14cb3),
	.w5(32'h3a48bcce),
	.w6(32'h3999720f),
	.w7(32'h39f3eaf9),
	.w8(32'h3a27e070),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73b4d2),
	.w1(32'h3b38b68c),
	.w2(32'h3ac9390d),
	.w3(32'h3a5c8777),
	.w4(32'h3ab165a2),
	.w5(32'h3a6b981e),
	.w6(32'h3b04e437),
	.w7(32'h3af78e1c),
	.w8(32'h3aa5c51b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a3285),
	.w1(32'hba6ccf69),
	.w2(32'hbb2692a7),
	.w3(32'h39083fa8),
	.w4(32'hbb6c21e0),
	.w5(32'hbb946a24),
	.w6(32'hba163550),
	.w7(32'hbac42fca),
	.w8(32'hbb3fe468),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a7f58),
	.w1(32'h38db2e87),
	.w2(32'hbb7fc189),
	.w3(32'hbba2c4b6),
	.w4(32'h3acf786e),
	.w5(32'hbb42cfb7),
	.w6(32'hbb55d49c),
	.w7(32'hbb87a667),
	.w8(32'hbb85766a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88566),
	.w1(32'hba1db652),
	.w2(32'hbb005c6d),
	.w3(32'hbb7150d0),
	.w4(32'h38f70f07),
	.w5(32'hbb0aa1c3),
	.w6(32'hb9c61965),
	.w7(32'hbae84a90),
	.w8(32'hb9f637e2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15db78),
	.w1(32'h3b38a819),
	.w2(32'h3b2e428e),
	.w3(32'hba19c679),
	.w4(32'h3ae72350),
	.w5(32'h3b06bdc7),
	.w6(32'h3b1a6d46),
	.w7(32'h3b24622c),
	.w8(32'h3aeffb40),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a8291),
	.w1(32'hbb314607),
	.w2(32'hbb307e68),
	.w3(32'h3b0780bd),
	.w4(32'hbb297705),
	.w5(32'hbb336cbb),
	.w6(32'hbb4b53e0),
	.w7(32'hbb33f087),
	.w8(32'hbb20f335),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ec5dc),
	.w1(32'h3ae2bd8a),
	.w2(32'h3af61813),
	.w3(32'hbb34359a),
	.w4(32'hba1af10d),
	.w5(32'hbaf8a68a),
	.w6(32'h3b27e31c),
	.w7(32'h3b955471),
	.w8(32'h3b7c8163),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce01e7),
	.w1(32'h3b1afb26),
	.w2(32'h3b007958),
	.w3(32'hbac5ede2),
	.w4(32'h3a0cc402),
	.w5(32'h3a3952b2),
	.w6(32'h3b05926a),
	.w7(32'h3b22373a),
	.w8(32'h3acc32ad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a887326),
	.w1(32'hb8db59d5),
	.w2(32'h3a34cf3b),
	.w3(32'h3a230294),
	.w4(32'hba79a0b3),
	.w5(32'h38c05e7b),
	.w6(32'hba2dac11),
	.w7(32'h3a189b9d),
	.w8(32'hb98d0856),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66a2451),
	.w1(32'hbbb5361b),
	.w2(32'hbbbda605),
	.w3(32'hba086817),
	.w4(32'hbb94dba2),
	.w5(32'hbb960896),
	.w6(32'hbbc42989),
	.w7(32'hbbc72024),
	.w8(32'hbb4dbc4b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb189486),
	.w1(32'h384c3577),
	.w2(32'hb98a7f1d),
	.w3(32'hba7d287c),
	.w4(32'h3998a65d),
	.w5(32'hb9e60673),
	.w6(32'h3a070a56),
	.w7(32'hb8ed32f2),
	.w8(32'hba4d6c76),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba887131),
	.w1(32'h398272b7),
	.w2(32'hb9a39e8d),
	.w3(32'hba564043),
	.w4(32'hba753b1d),
	.w5(32'hbac4a4b9),
	.w6(32'hb8e55717),
	.w7(32'hba10f46e),
	.w8(32'hba6042f2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f80d9),
	.w1(32'h3ab7aab0),
	.w2(32'h3b1df121),
	.w3(32'hbae08ab0),
	.w4(32'h39c00a1b),
	.w5(32'h3a8baba6),
	.w6(32'h3a2d90fd),
	.w7(32'h3ab022c6),
	.w8(32'h3ab393ad),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae766cd),
	.w1(32'h3a36a5b7),
	.w2(32'hbb542e53),
	.w3(32'h3a8a1da9),
	.w4(32'hba6e076a),
	.w5(32'hbb4a0f5e),
	.w6(32'h39b9c0c2),
	.w7(32'hbb2b3ecb),
	.w8(32'hbae22a39),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28b5c1),
	.w1(32'hb9fb5850),
	.w2(32'hba028964),
	.w3(32'hbb29d46e),
	.w4(32'hbadcdfa7),
	.w5(32'h3a1f98ff),
	.w6(32'hba2d08ce),
	.w7(32'hbabbe714),
	.w8(32'hba71126c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba088c7a),
	.w1(32'hbabb0eea),
	.w2(32'hba6b7c02),
	.w3(32'hb93e9f98),
	.w4(32'hba579a5c),
	.w5(32'hba7ee4b3),
	.w6(32'hba0a58d9),
	.w7(32'hba8c413a),
	.w8(32'hbab0100c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3e4e6),
	.w1(32'h3b1f2a7a),
	.w2(32'h3b37b232),
	.w3(32'hbadc3734),
	.w4(32'h38c5d409),
	.w5(32'h3a589ee0),
	.w6(32'h3ad4c362),
	.w7(32'h3b35a43f),
	.w8(32'h3b2279d6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b304761),
	.w1(32'h3a0b68ab),
	.w2(32'hba0b9c60),
	.w3(32'h3b091ad8),
	.w4(32'h3ad1560d),
	.w5(32'hb9186aba),
	.w6(32'h3a5a0d0d),
	.w7(32'hb981260f),
	.w8(32'hba59bddf),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9d05d),
	.w1(32'h3a8ede1e),
	.w2(32'hba2b439a),
	.w3(32'h3991cbac),
	.w4(32'h3aaca6fe),
	.w5(32'hb9efe83b),
	.w6(32'h3ac542b4),
	.w7(32'h3a50b896),
	.w8(32'hb702cde8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a8e1a3),
	.w1(32'h3b5d53b5),
	.w2(32'h3b3eb2af),
	.w3(32'hb9896de4),
	.w4(32'h3b0254d4),
	.w5(32'h3afc69a4),
	.w6(32'h3b1086d3),
	.w7(32'h3b466811),
	.w8(32'h3afbddba),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e19d9),
	.w1(32'h39fb0314),
	.w2(32'h3956367e),
	.w3(32'h3b1d82d1),
	.w4(32'h3a66b79d),
	.w5(32'h3a3cae32),
	.w6(32'h3a7c3843),
	.w7(32'h3a30cc8f),
	.w8(32'h39d0ee42),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10658b),
	.w1(32'hbaf44e26),
	.w2(32'hbb1cd6f4),
	.w3(32'h3a4dc113),
	.w4(32'hb9923684),
	.w5(32'hbac8628c),
	.w6(32'hbab421c7),
	.w7(32'hbb169e7d),
	.w8(32'hbaf5bc28),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1baf9a),
	.w1(32'h39f4d837),
	.w2(32'h3a3e28ad),
	.w3(32'hbaafb38f),
	.w4(32'hb93b03bf),
	.w5(32'h39cc316c),
	.w6(32'hb889b1d8),
	.w7(32'h39813b7d),
	.w8(32'h38408339),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ebc5b),
	.w1(32'hba2bdf69),
	.w2(32'h39065649),
	.w3(32'h393870e5),
	.w4(32'hb9b4df9c),
	.w5(32'hba326c02),
	.w6(32'hbaad006e),
	.w7(32'hb96667cd),
	.w8(32'hba3d0206),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e731f),
	.w1(32'hbad58cca),
	.w2(32'hbba9515e),
	.w3(32'hba12ea8a),
	.w4(32'hb8acebcc),
	.w5(32'hbb80fdfe),
	.w6(32'h3a8c8097),
	.w7(32'hbb337917),
	.w8(32'hbb46ca18),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb939b7b),
	.w1(32'h3b4c9d58),
	.w2(32'h3a4e67b1),
	.w3(32'hbb5c5356),
	.w4(32'h3b44073d),
	.w5(32'hb88bdd44),
	.w6(32'h3b758936),
	.w7(32'h3aeea622),
	.w8(32'h3aa418ac),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5a0d5),
	.w1(32'h3a76f172),
	.w2(32'hb95d4ef0),
	.w3(32'h393362cc),
	.w4(32'h3856dbb5),
	.w5(32'hba979c8f),
	.w6(32'h3a89709f),
	.w7(32'h3a351581),
	.w8(32'hb99e5d53),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9276ed),
	.w1(32'h3a5515e1),
	.w2(32'hbb31be7c),
	.w3(32'hbae409b4),
	.w4(32'hba0bfa2e),
	.w5(32'hbb01040b),
	.w6(32'h3aab8114),
	.w7(32'hba7ccc3d),
	.w8(32'hba3fa49f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae74d5f),
	.w1(32'hbac34b74),
	.w2(32'hbb0b1e7a),
	.w3(32'hbb34e41c),
	.w4(32'hba999d8d),
	.w5(32'hbaccca16),
	.w6(32'hbabc9e3d),
	.w7(32'hbb03e9b2),
	.w8(32'hbb2e3bc8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2201ec),
	.w1(32'h3ac232e6),
	.w2(32'h3af28d72),
	.w3(32'hbb1b929c),
	.w4(32'h3a56bf7c),
	.w5(32'h3a8ca262),
	.w6(32'h3a5e00fd),
	.w7(32'h3acd399f),
	.w8(32'h3ac52921),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5cfb8),
	.w1(32'h3ae2b086),
	.w2(32'h3abef8af),
	.w3(32'h3a729060),
	.w4(32'h3a4d0449),
	.w5(32'h3a829ea6),
	.w6(32'h3ad58514),
	.w7(32'h3ab88d86),
	.w8(32'h3a97e78d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e34f8),
	.w1(32'h3b20586b),
	.w2(32'h3a7d75fa),
	.w3(32'h3a904033),
	.w4(32'h3b14608b),
	.w5(32'h3a666f3e),
	.w6(32'h3b2b805f),
	.w7(32'h3aeb0347),
	.w8(32'h3af10a9e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a402b83),
	.w1(32'h3b805ac8),
	.w2(32'h3b9a6684),
	.w3(32'h3a2d5979),
	.w4(32'h3a2b1ce1),
	.w5(32'hb8a4b429),
	.w6(32'h3ba2ef89),
	.w7(32'h3b70b2ce),
	.w8(32'h395503e3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51ac20),
	.w1(32'h3b879540),
	.w2(32'h3ba41622),
	.w3(32'hbbf1bde7),
	.w4(32'h3b329f28),
	.w5(32'h3b6cb3f8),
	.w6(32'h3b3e58ce),
	.w7(32'h3b5f8a87),
	.w8(32'h3b288ba3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71e48d),
	.w1(32'hbac8a929),
	.w2(32'hbb4c5fe4),
	.w3(32'h3b487f4c),
	.w4(32'hbb056db2),
	.w5(32'hbb1499b6),
	.w6(32'hba6dbc20),
	.w7(32'hbb11676c),
	.w8(32'hbb043dfb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb186ee5),
	.w1(32'hbb03f380),
	.w2(32'hbae2a01a),
	.w3(32'hbafa8b4d),
	.w4(32'hbad0dbb0),
	.w5(32'hbafec0a6),
	.w6(32'hbafc3667),
	.w7(32'hbb113237),
	.w8(32'hbb312739),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb310604),
	.w1(32'hbb8fe86c),
	.w2(32'hbb5ce963),
	.w3(32'hbb3459e0),
	.w4(32'hbb22cf8f),
	.w5(32'hbb0a33ca),
	.w6(32'hbb931682),
	.w7(32'hbb752152),
	.w8(32'hbad7cbc1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4583a1),
	.w1(32'hb9b87d15),
	.w2(32'hb945fdad),
	.w3(32'hb9cde5d4),
	.w4(32'h38b5c9a6),
	.w5(32'hb81702cc),
	.w6(32'h3953a90e),
	.w7(32'h38c0731b),
	.w8(32'h38580aa7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f0709),
	.w1(32'hbb866dc6),
	.w2(32'hbb22e179),
	.w3(32'h37b6ea3f),
	.w4(32'hbbb6f2ec),
	.w5(32'hbb43ce94),
	.w6(32'hbb6ba589),
	.w7(32'hbabe2261),
	.w8(32'hbae7e5df),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801f4e),
	.w1(32'h39e6e219),
	.w2(32'h39af6123),
	.w3(32'hbb9137ed),
	.w4(32'h3a92f939),
	.w5(32'h3a31301b),
	.w6(32'h3a76192d),
	.w7(32'h3a0f7098),
	.w8(32'h3966a130),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39153143),
	.w1(32'h3b59008b),
	.w2(32'h3b57178c),
	.w3(32'h39e7c714),
	.w4(32'h3b136e9c),
	.w5(32'h3b2785d7),
	.w6(32'h3b21abe3),
	.w7(32'h3b3f39ed),
	.w8(32'h3b0a7a8c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a46a6),
	.w1(32'hb8f9a237),
	.w2(32'h398a8509),
	.w3(32'h3b2df6dd),
	.w4(32'h3a1f0d2e),
	.w5(32'h3a49b84d),
	.w6(32'h3a10c80b),
	.w7(32'h39f27ecc),
	.w8(32'h3a40e858),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a712e0f),
	.w1(32'h3ae94915),
	.w2(32'h39bff8b9),
	.w3(32'h3a6ed291),
	.w4(32'h3b0d6741),
	.w5(32'h3a7683d4),
	.w6(32'hb907ced0),
	.w7(32'hba260db6),
	.w8(32'hba4fc6d6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c738e2),
	.w1(32'h3a54d653),
	.w2(32'hbb4ccce0),
	.w3(32'h3a009506),
	.w4(32'h3a91c3f2),
	.w5(32'hbab4fb13),
	.w6(32'h39a415ea),
	.w7(32'hbb48364d),
	.w8(32'hba8eb117),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef7401),
	.w1(32'hbabe35c5),
	.w2(32'hbb5ebcdb),
	.w3(32'hba831c19),
	.w4(32'hb9cb3223),
	.w5(32'hbb25f6c9),
	.w6(32'h398438fe),
	.w7(32'hbae5ea8d),
	.w8(32'hbae3c9f4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c4280),
	.w1(32'h370d3791),
	.w2(32'hb9985d08),
	.w3(32'hbb2ee8cb),
	.w4(32'h3a1eb2a4),
	.w5(32'hb8e9f468),
	.w6(32'h3891c0c5),
	.w7(32'hb9bf9d2b),
	.w8(32'h39a1bb58),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e952c9),
	.w1(32'hbb4172c5),
	.w2(32'hbae3389b),
	.w3(32'h39878d32),
	.w4(32'hbb377c51),
	.w5(32'hba7925bc),
	.w6(32'hbb8a6c40),
	.w7(32'hbb19a6ee),
	.w8(32'hba9b04f8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf10eaa),
	.w1(32'h39c5439d),
	.w2(32'h3a77736b),
	.w3(32'hbb143de5),
	.w4(32'h3a367c4c),
	.w5(32'h3a6c2333),
	.w6(32'h39200663),
	.w7(32'h3a44dcbc),
	.w8(32'h39c50b69),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2534d0),
	.w1(32'hbb04f4b2),
	.w2(32'hbb5d898b),
	.w3(32'h3a1a197b),
	.w4(32'hba01ac23),
	.w5(32'hbb33915f),
	.w6(32'hba8c9604),
	.w7(32'hbb30c2c0),
	.w8(32'hbaf5b824),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bb1bd),
	.w1(32'h3b370d8e),
	.w2(32'h3b3e341d),
	.w3(32'hbb08b96c),
	.w4(32'h3a0ac6e0),
	.w5(32'h3a508f34),
	.w6(32'h3b094982),
	.w7(32'h3b1265c8),
	.w8(32'h39ddb64a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a684e8c),
	.w1(32'h3b1d6536),
	.w2(32'h3ac65e05),
	.w3(32'h3a7b6eea),
	.w4(32'h3b0037b1),
	.w5(32'h3aefadb6),
	.w6(32'h3b1b6321),
	.w7(32'h3b37d54f),
	.w8(32'h3aa0c84e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb808137f),
	.w1(32'h3a4241ea),
	.w2(32'h3a804a3c),
	.w3(32'h386e1d85),
	.w4(32'h3a8bcf6f),
	.w5(32'h3a44b9f1),
	.w6(32'h3abba606),
	.w7(32'h3a879a66),
	.w8(32'h3a1d1ff6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1665a),
	.w1(32'h3b13de00),
	.w2(32'h3b6617fc),
	.w3(32'h391a5011),
	.w4(32'h3a98ca4a),
	.w5(32'h3b1fdf20),
	.w6(32'h3af9f872),
	.w7(32'h3b38f12e),
	.w8(32'h3b177880),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09a08a),
	.w1(32'h3b4bfff6),
	.w2(32'h3b58e13a),
	.w3(32'h3b19ebed),
	.w4(32'h3af3ff29),
	.w5(32'h3b14b2f1),
	.w6(32'h3b1ec34e),
	.w7(32'h3b3dd4d8),
	.w8(32'h3b0ee543),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24ff83),
	.w1(32'h3b3853a9),
	.w2(32'h3b5c9af7),
	.w3(32'h3b150830),
	.w4(32'h39be352a),
	.w5(32'h3a79dcf1),
	.w6(32'h3b38a4d8),
	.w7(32'h3b5fdbcf),
	.w8(32'h3b0fa1d0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1897b4),
	.w1(32'hb8908c90),
	.w2(32'h39865f28),
	.w3(32'h3aa7e902),
	.w4(32'h3927574d),
	.w5(32'h37cbb341),
	.w6(32'hb8953738),
	.w7(32'hb9e258ad),
	.w8(32'hb847fe77),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8891236),
	.w1(32'h3b0f14ad),
	.w2(32'hba81e9f3),
	.w3(32'hb9e78dfb),
	.w4(32'h38fd1297),
	.w5(32'hbb08ef81),
	.w6(32'h3b98df79),
	.w7(32'h3b2d969b),
	.w8(32'h3b29a1b3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01e227),
	.w1(32'h3b3367eb),
	.w2(32'h3ae89060),
	.w3(32'hbb3d974b),
	.w4(32'h3ad83ad7),
	.w5(32'h3ab88107),
	.w6(32'h3b047906),
	.w7(32'h3aec8da5),
	.w8(32'h3ac6506c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae15fb9),
	.w1(32'h39d12f8f),
	.w2(32'h3ad80b05),
	.w3(32'h3b0b39eb),
	.w4(32'h3aa830b7),
	.w5(32'h3b15fdc4),
	.w6(32'h3a453f63),
	.w7(32'h3a999df5),
	.w8(32'h3b1f0199),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d3e2e),
	.w1(32'h3ad4c166),
	.w2(32'h3b188f8d),
	.w3(32'h3b3ffa1f),
	.w4(32'h3a46c73f),
	.w5(32'hba45b936),
	.w6(32'h3a738322),
	.w7(32'h3ad37919),
	.w8(32'h3a7abc67),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392395ac),
	.w1(32'hba7e3a43),
	.w2(32'hbacf989e),
	.w3(32'hba2e64e9),
	.w4(32'hbb48074d),
	.w5(32'hbb54ba96),
	.w6(32'hba805264),
	.w7(32'hbab6ced7),
	.w8(32'hbace99ec),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24a9a5),
	.w1(32'hbb088d15),
	.w2(32'hbb4ec454),
	.w3(32'hbb58a8b7),
	.w4(32'hb9c55242),
	.w5(32'hbaf03b41),
	.w6(32'hbaa60142),
	.w7(32'hbb3784de),
	.w8(32'hbab65889),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc07b8),
	.w1(32'hba6712d5),
	.w2(32'hba13d39a),
	.w3(32'hba8398b0),
	.w4(32'hb9b0a4af),
	.w5(32'hb8322172),
	.w6(32'hba400fa4),
	.w7(32'hba76441a),
	.w8(32'hba97341d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3752a4),
	.w1(32'hbb09e61e),
	.w2(32'hbae5d67f),
	.w3(32'hb99447dd),
	.w4(32'hbaec71b2),
	.w5(32'hbb0433ea),
	.w6(32'hbb0e2765),
	.w7(32'hbafe13e8),
	.w8(32'hbad84f1a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe7429),
	.w1(32'h3a4aafd4),
	.w2(32'h39668424),
	.w3(32'hbb020faa),
	.w4(32'h3a9f84e1),
	.w5(32'h3a2a1f58),
	.w6(32'h3a9c4426),
	.w7(32'h39ee4686),
	.w8(32'h3a088b61),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb75fd),
	.w1(32'hba7f6ae8),
	.w2(32'hb7622c94),
	.w3(32'h39cf0745),
	.w4(32'hbab6aef7),
	.w5(32'hb982b918),
	.w6(32'hba106566),
	.w7(32'hba7a6fbf),
	.w8(32'hbadb9629),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcaae3),
	.w1(32'h3abe1e8e),
	.w2(32'h3ada001f),
	.w3(32'hb9f0d7bf),
	.w4(32'h3aeb6524),
	.w5(32'h3aef14ac),
	.w6(32'h3a9addb0),
	.w7(32'h3ab42da7),
	.w8(32'h3ac8fde1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc8b86),
	.w1(32'hbab345da),
	.w2(32'hba1cc87e),
	.w3(32'h3ada8e5d),
	.w4(32'hbaa712ad),
	.w5(32'hba1ed533),
	.w6(32'h3993f0a7),
	.w7(32'h39a4df27),
	.w8(32'h3aa88dea),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396af497),
	.w1(32'h38257834),
	.w2(32'hba24b93a),
	.w3(32'h3a3cb800),
	.w4(32'hbaccc913),
	.w5(32'hbb022668),
	.w6(32'hb98904d8),
	.w7(32'hba5533cc),
	.w8(32'hbaddedf8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02c200),
	.w1(32'hbb7d0f6d),
	.w2(32'hbb72f505),
	.w3(32'hbb1c9ef5),
	.w4(32'hbb5691fb),
	.w5(32'hbb6cd2fd),
	.w6(32'hbb6a8e5e),
	.w7(32'hbb829c22),
	.w8(32'hbb85b4a1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8877fc),
	.w1(32'hb950c188),
	.w2(32'hb9d089f0),
	.w3(32'hbb87042d),
	.w4(32'hbb14ffec),
	.w5(32'hbb20b165),
	.w6(32'hba63e76e),
	.w7(32'hba5a769d),
	.w8(32'hba9c5a30),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade9e93),
	.w1(32'h3a80d457),
	.w2(32'h3a560c1b),
	.w3(32'hbb48e701),
	.w4(32'h38ca2245),
	.w5(32'hb9ff20e7),
	.w6(32'h3a0699cd),
	.w7(32'h39cff5ef),
	.w8(32'hba3e3adc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389237d6),
	.w1(32'h3aca4b4b),
	.w2(32'hb9c558fb),
	.w3(32'hb9f8352f),
	.w4(32'h3b0172d5),
	.w5(32'hb9665a9a),
	.w6(32'h3b2a7425),
	.w7(32'h3a8a7758),
	.w8(32'h39fae7fe),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942fefa),
	.w1(32'hbb0ce6ed),
	.w2(32'hbab391fd),
	.w3(32'hb9a0ca19),
	.w4(32'hba92a88a),
	.w5(32'hba57ef7a),
	.w6(32'hbaae6153),
	.w7(32'hbabb31b2),
	.w8(32'hbacb2816),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f9826),
	.w1(32'hbb944de6),
	.w2(32'hbbcb88b9),
	.w3(32'hba7a273c),
	.w4(32'hbb1845d6),
	.w5(32'hbb934a34),
	.w6(32'hbb6b2f95),
	.w7(32'hbbb5f3b8),
	.w8(32'hbb0b7ec1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1edb4e),
	.w1(32'hb98d67ca),
	.w2(32'h3a873cbd),
	.w3(32'hbaa2a4f8),
	.w4(32'h39027c74),
	.w5(32'h3a981706),
	.w6(32'hba36a5a3),
	.w7(32'h3807d99a),
	.w8(32'h3a24025b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac02000),
	.w1(32'h3ac6b127),
	.w2(32'h3a90af8e),
	.w3(32'h3ac19cf3),
	.w4(32'h3b5cb1e2),
	.w5(32'h3b4a7bc3),
	.w6(32'hba5645ca),
	.w7(32'hb9f8375a),
	.w8(32'hba079d29),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab49563),
	.w1(32'h38f910b5),
	.w2(32'h37d0820f),
	.w3(32'h3b41e23c),
	.w4(32'h38f28109),
	.w5(32'hba8d8196),
	.w6(32'hb9fed8a4),
	.w7(32'hba4ac216),
	.w8(32'hbae9662b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade4776),
	.w1(32'hba85b13f),
	.w2(32'hb9760da3),
	.w3(32'hbb2e2a56),
	.w4(32'hbac702e7),
	.w5(32'h39ac42a9),
	.w6(32'hbab676c4),
	.w7(32'hba349adf),
	.w8(32'h392b4edd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba361d5a),
	.w1(32'hba8f1e3f),
	.w2(32'hba00c328),
	.w3(32'hba0820cc),
	.w4(32'hba12f321),
	.w5(32'hb990c7cc),
	.w6(32'hba9e202b),
	.w7(32'hba44070a),
	.w8(32'hba8462cc),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7b10f),
	.w1(32'hbafc73df),
	.w2(32'hba59cc24),
	.w3(32'hb8c806f7),
	.w4(32'hba9ad8e8),
	.w5(32'hba3f9e80),
	.w6(32'hbb1a3443),
	.w7(32'hbb0eeb8a),
	.w8(32'hbae56748),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b34cab),
	.w1(32'hbaf6242c),
	.w2(32'hbb192c92),
	.w3(32'hb8f9e189),
	.w4(32'hbb7a2a40),
	.w5(32'hbb724d62),
	.w6(32'hbb10d477),
	.w7(32'hbae30725),
	.w8(32'hbb400d23),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95c709),
	.w1(32'hba841cff),
	.w2(32'hba9b8f67),
	.w3(32'hbb9ded98),
	.w4(32'hb9f993db),
	.w5(32'hbadeb915),
	.w6(32'hbb9413a9),
	.w7(32'hbb132f1b),
	.w8(32'hbab9db55),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c04d2),
	.w1(32'h3b84e9bd),
	.w2(32'h3b190962),
	.w3(32'hbb22928d),
	.w4(32'h3b17adc0),
	.w5(32'h3b01f750),
	.w6(32'h3b4b31eb),
	.w7(32'h3b32ba52),
	.w8(32'h3b0c650a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1267cd),
	.w1(32'h3b1d774b),
	.w2(32'h3b5ab006),
	.w3(32'h3b403659),
	.w4(32'h3a8392c7),
	.w5(32'h3ae8d738),
	.w6(32'h3b048511),
	.w7(32'h3b2b06fe),
	.w8(32'h3b1d074c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b191ee1),
	.w1(32'h3b0b763e),
	.w2(32'h3aad464d),
	.w3(32'h3b0a6d8c),
	.w4(32'h3aa6464c),
	.w5(32'h3a8d9151),
	.w6(32'h3ae6d55a),
	.w7(32'h3ab93841),
	.w8(32'h3aa03d12),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1a9c4),
	.w1(32'h3ac94098),
	.w2(32'h3a18a403),
	.w3(32'h3ac45075),
	.w4(32'hb94cdb7f),
	.w5(32'hb9a19405),
	.w6(32'h3ab8a7e1),
	.w7(32'h3aa2c807),
	.w8(32'h39f7683e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a627f),
	.w1(32'h39bd43a5),
	.w2(32'h3a1500e3),
	.w3(32'hb9afb13d),
	.w4(32'h3a62fb78),
	.w5(32'h3a76aa3f),
	.w6(32'h37b9b540),
	.w7(32'hb7e9832f),
	.w8(32'h39e3aaea),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae7955),
	.w1(32'h3a38109c),
	.w2(32'hb9a7da6c),
	.w3(32'h3aa46cbf),
	.w4(32'hba63fed8),
	.w5(32'hbb085232),
	.w6(32'h39decc5d),
	.w7(32'hb9c2b4f7),
	.w8(32'hbb09634a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf633fa),
	.w1(32'h3b0c42b9),
	.w2(32'h3a9da43a),
	.w3(32'hbb381eba),
	.w4(32'h3aadede8),
	.w5(32'h3a8fe22d),
	.w6(32'h3ad8ddbe),
	.w7(32'h3ab4c7c7),
	.w8(32'h3a960f27),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa39481),
	.w1(32'h3b7cc036),
	.w2(32'h3b162992),
	.w3(32'h3ad88327),
	.w4(32'h3b87079e),
	.w5(32'h3afdb26c),
	.w6(32'h3b9c9758),
	.w7(32'h3b1f54ff),
	.w8(32'h3b32d63b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e7095),
	.w1(32'h3b816110),
	.w2(32'h3b746e8c),
	.w3(32'h3b24fb52),
	.w4(32'h3affcac4),
	.w5(32'h3b041e99),
	.w6(32'h3b754040),
	.w7(32'h3b6db134),
	.w8(32'h3b38e789),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b257faf),
	.w1(32'h3a0ecd41),
	.w2(32'hbad2d0bc),
	.w3(32'h3a922abd),
	.w4(32'h3ac38fa0),
	.w5(32'hbac3030b),
	.w6(32'h39563d1a),
	.w7(32'hbb2dab4e),
	.w8(32'hbb2b3ef2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c120d),
	.w1(32'h3b42ef2a),
	.w2(32'h3b3f4377),
	.w3(32'hbb582c99),
	.w4(32'h3a942b88),
	.w5(32'h3a97ce3a),
	.w6(32'h3b287f9e),
	.w7(32'h3b319552),
	.w8(32'h3b02000d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b108bd2),
	.w1(32'h394123e6),
	.w2(32'h3a93e3bb),
	.w3(32'h3a89ed92),
	.w4(32'h3a1e1505),
	.w5(32'h3a403698),
	.w6(32'h3a485901),
	.w7(32'h3a3d8263),
	.w8(32'h3a6d97b6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4716c),
	.w1(32'h3adbfdd8),
	.w2(32'h3a11c75c),
	.w3(32'h3ad046bf),
	.w4(32'h3ae8e330),
	.w5(32'h39bbac84),
	.w6(32'h3acb34c3),
	.w7(32'h3a1b9ae3),
	.w8(32'h3a466c60),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e598b),
	.w1(32'h3b4b5b14),
	.w2(32'h3b03778a),
	.w3(32'h39f98284),
	.w4(32'h3af088fa),
	.w5(32'h3add6bf6),
	.w6(32'h3b1e957b),
	.w7(32'h3b12061f),
	.w8(32'h3b017248),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8ed6f),
	.w1(32'h3b2d5377),
	.w2(32'h3b4e71fa),
	.w3(32'h3b0f651d),
	.w4(32'h3ad699be),
	.w5(32'h3b1e4adc),
	.w6(32'h3b06bc4e),
	.w7(32'h3b31a2e4),
	.w8(32'h3b1541db),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a11ed),
	.w1(32'h3b3b9bc6),
	.w2(32'h3b56dbc8),
	.w3(32'h3b2ad492),
	.w4(32'h3ada6377),
	.w5(32'h3b21f6ee),
	.w6(32'h3b094c8e),
	.w7(32'h3b300570),
	.w8(32'h3b15f902),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f8004),
	.w1(32'h3a7bfac2),
	.w2(32'hbad18af8),
	.w3(32'h3b399577),
	.w4(32'h3b54f08a),
	.w5(32'hb9137aa8),
	.w6(32'hbb71b38c),
	.w7(32'hbb790155),
	.w8(32'hbb85c8a1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab911d5),
	.w1(32'hba91c529),
	.w2(32'hbaf0e429),
	.w3(32'hba444da6),
	.w4(32'hba369cea),
	.w5(32'hbac8c960),
	.w6(32'hba93d154),
	.w7(32'hbaaaaec7),
	.w8(32'hba42bdf6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97d7ee),
	.w1(32'h3b8b6b65),
	.w2(32'h3bc1fb53),
	.w3(32'hbaa54546),
	.w4(32'h3af03ed1),
	.w5(32'h3b4bc848),
	.w6(32'h3b6b4159),
	.w7(32'h3bb221ad),
	.w8(32'h3b9e0740),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b072),
	.w1(32'h3b97df55),
	.w2(32'h3bb478a1),
	.w3(32'h3b6d4730),
	.w4(32'h3b4641f0),
	.w5(32'h3b84e004),
	.w6(32'h3b66e67a),
	.w7(32'h3b977bb4),
	.w8(32'h3b1890dc),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31a999),
	.w1(32'h3b4ac2b4),
	.w2(32'h3b402406),
	.w3(32'h3af3d3f2),
	.w4(32'h3b074cc0),
	.w5(32'h3b176abb),
	.w6(32'h3b18661e),
	.w7(32'h3b2d1b8b),
	.w8(32'h3b00eba2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ec789),
	.w1(32'h3abe2103),
	.w2(32'hbb193915),
	.w3(32'h3b271ae9),
	.w4(32'h3b92bf5e),
	.w5(32'h386d23ac),
	.w6(32'hbb4b9296),
	.w7(32'hbb46e724),
	.w8(32'hbb87b97e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb887b4f),
	.w1(32'h3b6492fc),
	.w2(32'h3b9f6afe),
	.w3(32'hbb15179a),
	.w4(32'h3b48077a),
	.w5(32'h3b8912ed),
	.w6(32'h3b0b4e92),
	.w7(32'h3b4038f5),
	.w8(32'h3b2b1336),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e03f5),
	.w1(32'h3aa44869),
	.w2(32'h3a4442ec),
	.w3(32'h3b943492),
	.w4(32'hbaa0b1ae),
	.w5(32'hbad46fc9),
	.w6(32'h3a9b4898),
	.w7(32'h3a3612a1),
	.w8(32'hb9c38e88),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1071d6),
	.w1(32'h379316da),
	.w2(32'hb7855da7),
	.w3(32'hbaeb4c52),
	.w4(32'h37a930f8),
	.w5(32'hb6085631),
	.w6(32'h384da537),
	.w7(32'h35a33a64),
	.w8(32'hb81e9fd6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d25bcf),
	.w1(32'hb75bf290),
	.w2(32'hb9028af0),
	.w3(32'hb8a4669d),
	.w4(32'h380af038),
	.w5(32'hb8b443b1),
	.w6(32'h384b0f84),
	.w7(32'hb792fd3d),
	.w8(32'hb80e9df6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388877f3),
	.w1(32'h38f9e255),
	.w2(32'h39018f06),
	.w3(32'h39245600),
	.w4(32'h393132df),
	.w5(32'h3914a326),
	.w6(32'h39271601),
	.w7(32'h386aab51),
	.w8(32'h37cbeeb4),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371adffb),
	.w1(32'hb6849d7c),
	.w2(32'hb6f74b10),
	.w3(32'hb612494a),
	.w4(32'hb5f80223),
	.w5(32'hb714eb2e),
	.w6(32'hb69b54b6),
	.w7(32'hb74285ec),
	.w8(32'hb7711c61),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aed298),
	.w1(32'h37b7c6a4),
	.w2(32'hb60aeff2),
	.w3(32'h381b14e0),
	.w4(32'h366d32ef),
	.w5(32'hb8677c5e),
	.w6(32'hb8c391b0),
	.w7(32'hb888ebaf),
	.w8(32'hb86f0abf),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb743cd95),
	.w1(32'h36e16594),
	.w2(32'hb648876e),
	.w3(32'h3720bc1f),
	.w4(32'h377e99cf),
	.w5(32'h35d91399),
	.w6(32'hb6b1a9a4),
	.w7(32'hb716858f),
	.w8(32'hb7cc560c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb715eb90),
	.w1(32'hb8670b6d),
	.w2(32'hb882a76f),
	.w3(32'h372b3376),
	.w4(32'hb770f9d6),
	.w5(32'hb819eef9),
	.w6(32'hb7b922ef),
	.w7(32'hb7e1be59),
	.w8(32'hb7da5038),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7adf79d),
	.w1(32'h37b20e52),
	.w2(32'hb5abfb4a),
	.w3(32'hb7b7e26b),
	.w4(32'hb732de1f),
	.w5(32'h35d0da78),
	.w6(32'hb83d7309),
	.w7(32'h37aa548e),
	.w8(32'hb7c8e9a2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75c9d0a),
	.w1(32'hb90648ed),
	.w2(32'hb8edbfb7),
	.w3(32'h38f84541),
	.w4(32'hb85cd920),
	.w5(32'hb7146ed9),
	.w6(32'h384fe4dd),
	.w7(32'hb943f2b9),
	.w8(32'hb9558cf8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384b0096),
	.w1(32'hb6a59069),
	.w2(32'hb82cd814),
	.w3(32'h387d5a7c),
	.w4(32'h378a7a6c),
	.w5(32'hb8159c52),
	.w6(32'h38b316ad),
	.w7(32'hb67332d0),
	.w8(32'hb894dc38),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360c5bda),
	.w1(32'hb893cb80),
	.w2(32'h379cdf13),
	.w3(32'h38735187),
	.w4(32'hb801f443),
	.w5(32'h3813d380),
	.w6(32'h38b225c4),
	.w7(32'hb8b9becf),
	.w8(32'h36d11f41),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85a1eae),
	.w1(32'hb7644e05),
	.w2(32'hb8dc8a02),
	.w3(32'h38d8e1ed),
	.w4(32'h38778ca8),
	.w5(32'hb88e5e6b),
	.w6(32'h36bde39c),
	.w7(32'hb6b7d55e),
	.w8(32'hb906eb1f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385c4bc2),
	.w1(32'h385fe840),
	.w2(32'hb94c2ffb),
	.w3(32'h382047ed),
	.w4(32'h3820b9bb),
	.w5(32'hb94f5d04),
	.w6(32'h38242836),
	.w7(32'hb7f34ee2),
	.w8(32'hb996ffc9),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb793522c),
	.w1(32'hb90cc6ac),
	.w2(32'h35609af3),
	.w3(32'h39001b93),
	.w4(32'hb83f3ce2),
	.w5(32'h3713796e),
	.w6(32'h385726ed),
	.w7(32'hb8b6b9b3),
	.w8(32'hb88ed601),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377f4a73),
	.w1(32'hb7bc0476),
	.w2(32'hb85fd2f1),
	.w3(32'h3813e0a7),
	.w4(32'hb77f067b),
	.w5(32'hb82dd14b),
	.w6(32'h375a01a0),
	.w7(32'hb82790e4),
	.w8(32'hb887d247),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38efb13c),
	.w1(32'h384b2b6e),
	.w2(32'h37956e15),
	.w3(32'h392c7b19),
	.w4(32'h39049488),
	.w5(32'hb5435501),
	.w6(32'h39959e46),
	.w7(32'h38e273b0),
	.w8(32'h37578424),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5487ccc),
	.w1(32'h368ad149),
	.w2(32'h383a59dd),
	.w3(32'h387739aa),
	.w4(32'h3734493f),
	.w5(32'h37a8e26a),
	.w6(32'h380b66b5),
	.w7(32'h378f419c),
	.w8(32'h3806bd16),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c766bc),
	.w1(32'hb5fad2c6),
	.w2(32'hb58ed8fb),
	.w3(32'h374c8239),
	.w4(32'h35b48c0b),
	.w5(32'h31078ab5),
	.w6(32'h37221d66),
	.w7(32'hb5c51b6d),
	.w8(32'hb6bf9d0d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4ec503f),
	.w1(32'hb6759eb6),
	.w2(32'hb704d6a6),
	.w3(32'h36102740),
	.w4(32'hb572a36e),
	.w5(32'hb6fb6f22),
	.w6(32'hb427158f),
	.w7(32'h354de5b8),
	.w8(32'hb5939358),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb744fba9),
	.w1(32'h378cd3dd),
	.w2(32'h36edb777),
	.w3(32'h365eac96),
	.w4(32'h3709ff5f),
	.w5(32'hb71d10c2),
	.w6(32'hb784c64d),
	.w7(32'hb7ccfcaa),
	.w8(32'hb799efaf),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9a01a),
	.w1(32'hb795fbbc),
	.w2(32'h3818d883),
	.w3(32'hb5a75e72),
	.w4(32'hb824d56f),
	.w5(32'h38910e22),
	.w6(32'hb55f4459),
	.w7(32'hb6eedca2),
	.w8(32'h37c75b1e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390dd1bd),
	.w1(32'h3905eb1b),
	.w2(32'h37eb27fd),
	.w3(32'h39668edb),
	.w4(32'h39086b7f),
	.w5(32'h3871ae49),
	.w6(32'h3852d5cf),
	.w7(32'hb8247703),
	.w8(32'hb8f43e80),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5195102),
	.w1(32'hb49a6ae6),
	.w2(32'hb5eaecee),
	.w3(32'hb5c1415b),
	.w4(32'hb609aba3),
	.w5(32'hb3f9713e),
	.w6(32'hb6b74364),
	.w7(32'hb70de3e8),
	.w8(32'hb6db23a4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ae72c8),
	.w1(32'hb8cd588a),
	.w2(32'h37a1dbfa),
	.w3(32'h3918fbfd),
	.w4(32'hb8938ea8),
	.w5(32'h385a4a53),
	.w6(32'h38d7e1cb),
	.w7(32'hb8b4948d),
	.w8(32'hb8fdc668),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3711a895),
	.w1(32'hb91bec60),
	.w2(32'h39116851),
	.w3(32'hb908ddec),
	.w4(32'hb98ea42a),
	.w5(32'h38f5afbf),
	.w6(32'hb7646539),
	.w7(32'hb9692be2),
	.w8(32'h3905693b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389de845),
	.w1(32'h37682bf6),
	.w2(32'hb93413ea),
	.w3(32'h3904b2a0),
	.w4(32'h380b782c),
	.w5(32'hb877c3f7),
	.w6(32'h3971634d),
	.w7(32'h36bedb9d),
	.w8(32'hb94392c8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37207a46),
	.w1(32'hb7fe090f),
	.w2(32'h34052b86),
	.w3(32'h3925da1a),
	.w4(32'h37e1488d),
	.w5(32'hb7f80583),
	.w6(32'h39386394),
	.w7(32'h383425fe),
	.w8(32'hb7b4541d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38045faa),
	.w1(32'hb8269231),
	.w2(32'h37112096),
	.w3(32'hb8aaec1a),
	.w4(32'hb896a138),
	.w5(32'hb6331334),
	.w6(32'hb94924dd),
	.w7(32'hb932b70a),
	.w8(32'hb8ead22b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807b6a1),
	.w1(32'h3972b2e7),
	.w2(32'h390c0486),
	.w3(32'hb989030e),
	.w4(32'h373e567f),
	.w5(32'hb8f14e72),
	.w6(32'hb9cb8cba),
	.w7(32'hb92b3d9a),
	.w8(32'hb9228ff2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0a2e3),
	.w1(32'h382b16ae),
	.w2(32'hb9017f0d),
	.w3(32'h39bc456e),
	.w4(32'h378a1f86),
	.w5(32'hb97bf16e),
	.w6(32'h39c664e6),
	.w7(32'hb8b3a667),
	.w8(32'hb9b1ce1f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365a5123),
	.w1(32'h38c9cf44),
	.w2(32'h3835e419),
	.w3(32'hb8c65b16),
	.w4(32'hb8f810ee),
	.w5(32'hb81f3cce),
	.w6(32'hb9078938),
	.w7(32'hb95e6af2),
	.w8(32'hb87748d7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386bcb8a),
	.w1(32'h38869d11),
	.w2(32'h37c54222),
	.w3(32'h38932030),
	.w4(32'h38ac6a13),
	.w5(32'h37e64e70),
	.w6(32'h388b3dac),
	.w7(32'h38c53369),
	.w8(32'h37ab7d7c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ab1635),
	.w1(32'hb79d39a0),
	.w2(32'hb809eb9a),
	.w3(32'hb7a308b3),
	.w4(32'hb6bb8d60),
	.w5(32'hb74ce587),
	.w6(32'hb721bce3),
	.w7(32'hb72c6b5c),
	.w8(32'hb80ea613),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb686dbf0),
	.w1(32'hb5cb6dd2),
	.w2(32'h36974889),
	.w3(32'hb6a5392d),
	.w4(32'hb6664002),
	.w5(32'h36a248ce),
	.w6(32'hb55f55d3),
	.w7(32'hb6831059),
	.w8(32'h35dfaf54),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359309c1),
	.w1(32'h37c63fb4),
	.w2(32'h3863580a),
	.w3(32'h38b082d3),
	.w4(32'h37edb0f0),
	.w5(32'h38d0d44f),
	.w6(32'hb7195032),
	.w7(32'hb60f9882),
	.w8(32'hb7b51bf0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c7d251),
	.w1(32'hb78de643),
	.w2(32'hb69623fb),
	.w3(32'h37ac202f),
	.w4(32'hb6a80f1c),
	.w5(32'hb762a112),
	.w6(32'h373fd16a),
	.w7(32'h36bfda64),
	.w8(32'hb77a870b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38afadd3),
	.w1(32'h378db7e5),
	.w2(32'h37dda93c),
	.w3(32'h39299a9e),
	.w4(32'h38a757f0),
	.w5(32'h3686b5d4),
	.w6(32'h392f5cae),
	.w7(32'h388248d0),
	.w8(32'hb6a02b8d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac1fd9),
	.w1(32'h38610189),
	.w2(32'hb8ca944f),
	.w3(32'h391b663d),
	.w4(32'h38048926),
	.w5(32'hb898ba74),
	.w6(32'h3956b001),
	.w7(32'h38937af7),
	.w8(32'hb8ccc18b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83fab08),
	.w1(32'h38d051e4),
	.w2(32'h37925a1d),
	.w3(32'hb84f2d50),
	.w4(32'h38951554),
	.w5(32'hb70dd52e),
	.w6(32'hb92eaffa),
	.w7(32'hb808e31e),
	.w8(32'hb8bdae94),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f78c3),
	.w1(32'hb838a335),
	.w2(32'hb8606e27),
	.w3(32'hb898392c),
	.w4(32'hb83b316a),
	.w5(32'hb8339bc5),
	.w6(32'hb8c70c35),
	.w7(32'hb89cce89),
	.w8(32'hb887a1e7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e1812b),
	.w1(32'h3842b070),
	.w2(32'hb7b596de),
	.w3(32'hb80f83dc),
	.w4(32'h381c8856),
	.w5(32'h36fe3c6f),
	.w6(32'h36120f66),
	.w7(32'h38690086),
	.w8(32'h379098e8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970b7a9),
	.w1(32'h38e502ae),
	.w2(32'hb73e86c6),
	.w3(32'h39ddde94),
	.w4(32'h395d1b4c),
	.w5(32'h3871e623),
	.w6(32'h397dcc82),
	.w7(32'h38d97b1b),
	.w8(32'hb81e3bb8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38559657),
	.w1(32'hb61f3a5d),
	.w2(32'hb7fea3f7),
	.w3(32'h3983cb22),
	.w4(32'hb9050543),
	.w5(32'hb85d8cac),
	.w6(32'h3942fb40),
	.w7(32'hb987d6db),
	.w8(32'hb926de66),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82a35bb),
	.w1(32'h33d65ecf),
	.w2(32'hb935951c),
	.w3(32'hb8e80875),
	.w4(32'hb82fba17),
	.w5(32'hb90d9d43),
	.w6(32'hb8a90c4e),
	.w7(32'hb7b89086),
	.w8(32'hb9111bda),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9492176),
	.w1(32'hb98b19c0),
	.w2(32'hb8d8300c),
	.w3(32'hb981a624),
	.w4(32'hb9a23732),
	.w5(32'hb893164e),
	.w6(32'hb92a5b62),
	.w7(32'hb9c483cc),
	.w8(32'hb8df3d2b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7351e4c),
	.w1(32'h37a87117),
	.w2(32'hb6afa701),
	.w3(32'hb5b3f2c4),
	.w4(32'h371a9c28),
	.w5(32'hb7bfd57f),
	.w6(32'hb732648f),
	.w7(32'h371f4fb9),
	.w8(32'hb7ab9f72),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd2acc),
	.w1(32'h38c98ad2),
	.w2(32'hb994e745),
	.w3(32'h3a152408),
	.w4(32'h39a87326),
	.w5(32'hb9b374c6),
	.w6(32'h3a08a9e5),
	.w7(32'h390cef99),
	.w8(32'hb9e95985),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38024226),
	.w1(32'hb783a8e8),
	.w2(32'hb98dcfdc),
	.w3(32'h381a98e8),
	.w4(32'hb7a7e7f1),
	.w5(32'hb97851e2),
	.w6(32'hb750a13d),
	.w7(32'hb85fc9e0),
	.w8(32'hb97388fc),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b9cbc),
	.w1(32'hb906e200),
	.w2(32'h38bf248c),
	.w3(32'h390b38d1),
	.w4(32'hb9a145c4),
	.w5(32'hb89f26b6),
	.w6(32'hb7ca7fad),
	.w7(32'hb9dd5343),
	.w8(32'hb9920b54),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3897f103),
	.w1(32'hb8892794),
	.w2(32'hb8ba249b),
	.w3(32'h38c0c071),
	.w4(32'hb6366158),
	.w5(32'hb8c3c194),
	.w6(32'h39241861),
	.w7(32'hb7c3c6df),
	.w8(32'hb9121a02),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e4bfc7),
	.w1(32'hb6d154ee),
	.w2(32'hb72201fb),
	.w3(32'h3934dac9),
	.w4(32'h37d4a609),
	.w5(32'h38584ffd),
	.w6(32'h39189dad),
	.w7(32'hb776f9ca),
	.w8(32'hb88fbddf),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73530d4),
	.w1(32'hb2d93cca),
	.w2(32'h35047cc5),
	.w3(32'hb724e3d4),
	.w4(32'h36073c74),
	.w5(32'h36ff8aa0),
	.w6(32'hb5b7744b),
	.w7(32'h35cccc4b),
	.w8(32'h36f6743e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371e0163),
	.w1(32'h378fabcb),
	.w2(32'hb849dd0a),
	.w3(32'h3717b798),
	.w4(32'hb5d6a38c),
	.w5(32'hb8a603cd),
	.w6(32'h3800a9f8),
	.w7(32'h376d5c6d),
	.w8(32'hb893e967),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363ec8bb),
	.w1(32'h37fb9479),
	.w2(32'h358b4175),
	.w3(32'hb6893517),
	.w4(32'h383b49dc),
	.w5(32'h37599d4b),
	.w6(32'h37d51712),
	.w7(32'h38193426),
	.w8(32'h36e03f11),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389eea21),
	.w1(32'hb7123581),
	.w2(32'hb89fd5b1),
	.w3(32'h38bf3c70),
	.w4(32'h3806b0d7),
	.w5(32'hb8816544),
	.w6(32'h383ea244),
	.w7(32'hb82564fd),
	.w8(32'hb8f5ca08),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a649b9),
	.w1(32'hb716157d),
	.w2(32'hb6f23eff),
	.w3(32'h35d4ce69),
	.w4(32'hb716317f),
	.w5(32'hb6cc07c7),
	.w6(32'hb75d0f50),
	.w7(32'hb74fa0b2),
	.w8(32'hb70cc5c5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74cd190),
	.w1(32'h371777e1),
	.w2(32'h373a9892),
	.w3(32'hb681d9b9),
	.w4(32'hb6464163),
	.w5(32'hb71af7ea),
	.w6(32'h36d5294e),
	.w7(32'hb70a757a),
	.w8(32'h37183037),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6706ff0),
	.w1(32'h36b5df3d),
	.w2(32'hb79fb93c),
	.w3(32'hb797a636),
	.w4(32'hb60da1f0),
	.w5(32'hb70f251c),
	.w6(32'hb740ed5d),
	.w7(32'hb6752cb8),
	.w8(32'hb7d8b5c5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7da90ba),
	.w1(32'hb80e127d),
	.w2(32'hb941aeb5),
	.w3(32'hb6569c30),
	.w4(32'hb883a29f),
	.w5(32'hb93ab49d),
	.w6(32'hb86185c1),
	.w7(32'hb8c19d28),
	.w8(32'hb95c3422),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ca307c),
	.w1(32'h37cef048),
	.w2(32'hb8702c2a),
	.w3(32'hb53b9598),
	.w4(32'h3836c1d1),
	.w5(32'hb85e9939),
	.w6(32'hb3be5a6e),
	.w7(32'h36d2f751),
	.w8(32'hb84d26a2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a24957),
	.w1(32'hb82683a7),
	.w2(32'hb8de6538),
	.w3(32'hb7c0e70a),
	.w4(32'hb54f7354),
	.w5(32'hb8ae121b),
	.w6(32'h3678da59),
	.w7(32'h379cd31a),
	.w8(32'hb8d6d41f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79c4144),
	.w1(32'hb9a54d9d),
	.w2(32'h38816c3d),
	.w3(32'h38e102a0),
	.w4(32'hb9094365),
	.w5(32'h37390343),
	.w6(32'hb9056d33),
	.w7(32'hba00633f),
	.w8(32'hb9e53099),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398fb455),
	.w1(32'h393e70a0),
	.w2(32'hb65175cf),
	.w3(32'h3989f130),
	.w4(32'h38733da9),
	.w5(32'hb8b1371b),
	.w6(32'h39167dca),
	.w7(32'hb76557be),
	.w8(32'hb90e21c7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360c7405),
	.w1(32'hb8730496),
	.w2(32'hb8f299f2),
	.w3(32'h376bb08d),
	.w4(32'hb8114aa8),
	.w5(32'hb8f09a6d),
	.w6(32'h378cc983),
	.w7(32'hb83d1861),
	.w8(32'hb902fd1f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bcb471),
	.w1(32'h369adc53),
	.w2(32'hb68add20),
	.w3(32'h3669f053),
	.w4(32'hb6fc72e5),
	.w5(32'hb723099f),
	.w6(32'hb3a8c0ab),
	.w7(32'hb71d93b5),
	.w8(32'hb7b6f741),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dce856),
	.w1(32'h389fe96d),
	.w2(32'h3758a267),
	.w3(32'h378c7ef7),
	.w4(32'h379d0a38),
	.w5(32'h3685b5de),
	.w6(32'hb649a0df),
	.w7(32'h36ab7ba6),
	.w8(32'h376c8c48),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3588a1fe),
	.w1(32'h3649f755),
	.w2(32'h36274393),
	.w3(32'hb6e49f96),
	.w4(32'h3669b482),
	.w5(32'h36a440d7),
	.w6(32'hb6ea4626),
	.w7(32'hb6939889),
	.w8(32'h3682b7b4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373cbcc1),
	.w1(32'hb73f16b4),
	.w2(32'h358e9737),
	.w3(32'h38468399),
	.w4(32'hb6a8beea),
	.w5(32'h3610a10d),
	.w6(32'h380bffc9),
	.w7(32'h364d8e1b),
	.w8(32'h3802f9e7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36311a41),
	.w1(32'h37d9b5c5),
	.w2(32'hb79fc493),
	.w3(32'hb823af28),
	.w4(32'h382ad43d),
	.w5(32'hb887b1de),
	.w6(32'hb8434acf),
	.w7(32'hb8d11cd9),
	.w8(32'hb899edcd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c1d4f),
	.w1(32'h393bb852),
	.w2(32'hb725821a),
	.w3(32'h39860f2e),
	.w4(32'h3981053d),
	.w5(32'h38072789),
	.w6(32'h39322610),
	.w7(32'h38e7e247),
	.w8(32'hb8e09c40),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d17f31),
	.w1(32'h3826dffe),
	.w2(32'hb82e131b),
	.w3(32'hb7ddb48b),
	.w4(32'h3832d22d),
	.w5(32'hb8af93c1),
	.w6(32'h3797ef19),
	.w7(32'hb5878d1a),
	.w8(32'hb8c87393),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eca3c8),
	.w1(32'hb908dbfe),
	.w2(32'hb9a6b811),
	.w3(32'h3970e14b),
	.w4(32'hb7914b12),
	.w5(32'hb986a939),
	.w6(32'h396937e5),
	.w7(32'h3796b197),
	.w8(32'hb98c0120),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3837ebb5),
	.w1(32'h37e35406),
	.w2(32'hb847d99c),
	.w3(32'h387209c1),
	.w4(32'h37c0f1ef),
	.w5(32'hb86fde5b),
	.w6(32'h38664e1c),
	.w7(32'h379f1501),
	.w8(32'hb86aaa54),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37022ad7),
	.w1(32'h3524c448),
	.w2(32'h36c8a63e),
	.w3(32'h3722e7ed),
	.w4(32'h369bde65),
	.w5(32'h373c80e4),
	.w6(32'h36d64eb8),
	.w7(32'h365b9b2c),
	.w8(32'h370d028a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c14799),
	.w1(32'hb787d4d8),
	.w2(32'hb79026b7),
	.w3(32'hb78b2041),
	.w4(32'hb78c0665),
	.w5(32'hb77c8f39),
	.w6(32'hb7f393c5),
	.w7(32'hb8304aef),
	.w8(32'hb8172b04),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb722243f),
	.w1(32'hb58b7941),
	.w2(32'h37a96ae2),
	.w3(32'hb6dafef8),
	.w4(32'hb43741c8),
	.w5(32'h37b425b2),
	.w6(32'hb6ed5566),
	.w7(32'h32b6a97e),
	.w8(32'h379b7d7b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c934f7),
	.w1(32'hb7c0a20d),
	.w2(32'hb9244829),
	.w3(32'h390fdaad),
	.w4(32'h384d4843),
	.w5(32'hb8ee9de5),
	.w6(32'h38a82fe9),
	.w7(32'h385e79fe),
	.w8(32'hb8f013df),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3877c8c9),
	.w1(32'h3944f338),
	.w2(32'h38bcf429),
	.w3(32'hb231a5a0),
	.w4(32'h39373bc7),
	.w5(32'h3843acb4),
	.w6(32'h378992c1),
	.w7(32'h391e2db1),
	.w8(32'h37c8fe9a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68a456f),
	.w1(32'hb83b2d86),
	.w2(32'hb9808dc6),
	.w3(32'h37917339),
	.w4(32'hb7be196c),
	.w5(32'hb97ca4aa),
	.w6(32'h37f75683),
	.w7(32'hb7f137f6),
	.w8(32'hb97f0f74),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3757c099),
	.w1(32'h381a65cd),
	.w2(32'hb928e838),
	.w3(32'h38079e8e),
	.w4(32'h38558bf3),
	.w5(32'hb90a9b1e),
	.w6(32'h379bfd9e),
	.w7(32'h3842e4e1),
	.w8(32'hb913a22e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b562e7),
	.w1(32'hb8bb2d21),
	.w2(32'hb8bfaaa4),
	.w3(32'h388ccd94),
	.w4(32'hb8df80b8),
	.w5(32'hb8db1171),
	.w6(32'hb6fbed91),
	.w7(32'hb903264d),
	.w8(32'hb91f9846),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5ac8e),
	.w1(32'hb8f44f93),
	.w2(32'hb809f0df),
	.w3(32'h391186cf),
	.w4(32'hb87e016d),
	.w5(32'h35ec75b2),
	.w6(32'h392e8456),
	.w7(32'hb8395807),
	.w8(32'hb80115c1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39162937),
	.w1(32'h386e1286),
	.w2(32'hb864c963),
	.w3(32'h399ac42b),
	.w4(32'h390024fc),
	.w5(32'hb728fe64),
	.w6(32'h397d7cc1),
	.w7(32'h3833568c),
	.w8(32'hb9523246),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73f6288),
	.w1(32'hb66b4a67),
	.w2(32'h36223d39),
	.w3(32'hb76321b3),
	.w4(32'h36700ac4),
	.w5(32'h371654a5),
	.w6(32'hb4773db6),
	.w7(32'hb5f74791),
	.w8(32'h376b2bf7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c3c6bc),
	.w1(32'h3610726a),
	.w2(32'h36a887d6),
	.w3(32'h36946795),
	.w4(32'h368258c0),
	.w5(32'h36a3d4c9),
	.w6(32'h368a1050),
	.w7(32'h3679c817),
	.w8(32'hb5aa2017),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a1891),
	.w1(32'h3754b260),
	.w2(32'hb98badf1),
	.w3(32'h383a2022),
	.w4(32'hb7287140),
	.w5(32'hb980be8b),
	.w6(32'hb712ad60),
	.w7(32'hb895f066),
	.w8(32'hb991ec7f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bc52e9),
	.w1(32'hb8125656),
	.w2(32'hb893e556),
	.w3(32'h38ce0f47),
	.w4(32'hb82c4607),
	.w5(32'hb85aeb04),
	.w6(32'h37478703),
	.w7(32'hb93b8d40),
	.w8(32'hb930e996),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d90571),
	.w1(32'h37912810),
	.w2(32'hb7e8feda),
	.w3(32'h39820d2b),
	.w4(32'h388d8baa),
	.w5(32'h389b4695),
	.w6(32'h39591a45),
	.w7(32'h381ad052),
	.w8(32'h37fd38f8),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84baff2),
	.w1(32'hb84dc34f),
	.w2(32'hb812e079),
	.w3(32'h37c2b195),
	.w4(32'h371368cc),
	.w5(32'h3680334b),
	.w6(32'hb7f943e8),
	.w7(32'hb8450838),
	.w8(32'hb8716d0a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361b8a73),
	.w1(32'hb674edc3),
	.w2(32'h36b953e7),
	.w3(32'hb622002b),
	.w4(32'hb6f10fc4),
	.w5(32'h36a4c209),
	.w6(32'hb6b279ce),
	.w7(32'hb6f264b7),
	.w8(32'h36534326),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384e446b),
	.w1(32'h37fbdbd3),
	.w2(32'h37712962),
	.w3(32'h381df7f1),
	.w4(32'h3810ee06),
	.w5(32'h3743412d),
	.w6(32'h383f2c85),
	.w7(32'h37cc7974),
	.w8(32'h37bcb655),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82f2f67),
	.w1(32'h383a0e83),
	.w2(32'hb8c1b3b3),
	.w3(32'hb7a764a6),
	.w4(32'h385ba003),
	.w5(32'hb7ae0b5c),
	.w6(32'hb739b763),
	.w7(32'h38665c63),
	.w8(32'hb7657795),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36505c35),
	.w1(32'h38a177f2),
	.w2(32'h37d16ccc),
	.w3(32'hb6add952),
	.w4(32'h38d5673a),
	.w5(32'h38a9fc4f),
	.w6(32'hb86c5f1c),
	.w7(32'h3739e3a9),
	.w8(32'hb8d0ac54),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c48870),
	.w1(32'hb82a9337),
	.w2(32'hb866aeae),
	.w3(32'h37f4823d),
	.w4(32'h3887b6a0),
	.w5(32'h380da39b),
	.w6(32'hb731a869),
	.w7(32'hb8241858),
	.w8(32'hb89dc70c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383cf95e),
	.w1(32'h38925d70),
	.w2(32'hb8936cb0),
	.w3(32'h37c5b945),
	.w4(32'h3858c229),
	.w5(32'hb8c92a91),
	.w6(32'h35d59695),
	.w7(32'h37a4f8fe),
	.w8(32'hb9017b72),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37906ca6),
	.w1(32'hb805844f),
	.w2(32'hb8592183),
	.w3(32'h386c5242),
	.w4(32'hb82039b3),
	.w5(32'hb847cebf),
	.w6(32'h3703c1e9),
	.w7(32'hb80ef3ab),
	.w8(32'hb8b18d6c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb703c677),
	.w1(32'hb63ac9e6),
	.w2(32'hb63a6b3e),
	.w3(32'hb746ef4a),
	.w4(32'h36c06d21),
	.w5(32'h369b52e1),
	.w6(32'hb3f25e97),
	.w7(32'h35fc6e1a),
	.w8(32'h36c2a7a5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34fe9be0),
	.w1(32'hb6e52969),
	.w2(32'h3680811e),
	.w3(32'h366cca26),
	.w4(32'hb77ba53c),
	.w5(32'hb7564987),
	.w6(32'hb721d0bf),
	.w7(32'hb34a2504),
	.w8(32'h36cd3178),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f7fc5c),
	.w1(32'hb6b4bd1c),
	.w2(32'hb74c3e1c),
	.w3(32'hb799ddba),
	.w4(32'hb72ad520),
	.w5(32'hb79c0e1b),
	.w6(32'hb6fcb566),
	.w7(32'hb7009b28),
	.w8(32'hb7637034),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7899bc0),
	.w1(32'hb710c1ad),
	.w2(32'h372351d4),
	.w3(32'hb79cf73e),
	.w4(32'h34236115),
	.w5(32'h370ab751),
	.w6(32'hb6eef26d),
	.w7(32'h364c13f7),
	.w8(32'h36a7969d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381396c0),
	.w1(32'h37b27556),
	.w2(32'hb8645fc8),
	.w3(32'h380d60e7),
	.w4(32'h37a96e8f),
	.w5(32'hb8518a6e),
	.w6(32'h38166ec6),
	.w7(32'h36f50109),
	.w8(32'hb85fe9c3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3875a040),
	.w1(32'hb9356f65),
	.w2(32'h38aea5d2),
	.w3(32'h39815b5d),
	.w4(32'hb70c6d39),
	.w5(32'h38ab1e86),
	.w6(32'h39851759),
	.w7(32'h382b3390),
	.w8(32'h386bfd60),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78897d2),
	.w1(32'hb8552b5b),
	.w2(32'h37893002),
	.w3(32'h38733292),
	.w4(32'h37bc5d88),
	.w5(32'h380771ef),
	.w6(32'h3883a53b),
	.w7(32'h37982191),
	.w8(32'h37d2b8a4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3743e906),
	.w1(32'hb6b919e8),
	.w2(32'hb50b07aa),
	.w3(32'h371ace75),
	.w4(32'hb706830c),
	.w5(32'hb78a4cd9),
	.w6(32'hb788bc96),
	.w7(32'hb7754f65),
	.w8(32'hb6c140e2),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3851c826),
	.w1(32'hb77be870),
	.w2(32'hb925edf3),
	.w3(32'h38972114),
	.w4(32'h38216950),
	.w5(32'hb8b42831),
	.w6(32'h379352bd),
	.w7(32'hb880abad),
	.w8(32'hb97c43e8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a80202),
	.w1(32'hb834ca72),
	.w2(32'hb70c8383),
	.w3(32'hb789b3cb),
	.w4(32'hb80577c7),
	.w5(32'h37519adb),
	.w6(32'hb843d0bf),
	.w7(32'hb88aaffe),
	.w8(32'hb8f114f7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a4f0dd),
	.w1(32'hb695f6f6),
	.w2(32'hb5bd7b98),
	.w3(32'hb6a7de97),
	.w4(32'hb6841fe3),
	.w5(32'h35e80dab),
	.w6(32'hb432fd09),
	.w7(32'hb5d415c8),
	.w8(32'h35c15069),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389196ac),
	.w1(32'h37d521f0),
	.w2(32'hb8e2785e),
	.w3(32'h38df58a1),
	.w4(32'h388b85db),
	.w5(32'hb8acc95c),
	.w6(32'h3881149f),
	.w7(32'hb6d3a2d9),
	.w8(32'hb92d2a1f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3785180c),
	.w1(32'hb65f42af),
	.w2(32'hb60db20e),
	.w3(32'h369dad0d),
	.w4(32'h36358b57),
	.w5(32'hb6e9f3fa),
	.w6(32'h3601366d),
	.w7(32'hb5898a33),
	.w8(32'hb64d3799),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380926db),
	.w1(32'hb7d420e9),
	.w2(32'h37beb355),
	.w3(32'h36f78180),
	.w4(32'hb88f1a22),
	.w5(32'hb70975f9),
	.w6(32'hb7c2f0dc),
	.w7(32'hb8c67ca8),
	.w8(32'hb52d3b83),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dc469f),
	.w1(32'h3616d934),
	.w2(32'h36a57f4a),
	.w3(32'hb69c44f8),
	.w4(32'h3611ed9e),
	.w5(32'h36e81fa6),
	.w6(32'h3601f7ae),
	.w7(32'h3681a5ce),
	.w8(32'h369c3dd2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5321dd6),
	.w1(32'hb7318846),
	.w2(32'hb77e02aa),
	.w3(32'hb6673fea),
	.w4(32'hb7389823),
	.w5(32'hb7446ccf),
	.w6(32'hb76e9512),
	.w7(32'hb76aaac4),
	.w8(32'hb6c9ae9b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3843c619),
	.w1(32'h382c8909),
	.w2(32'hb7303acd),
	.w3(32'h36df6942),
	.w4(32'h37719f84),
	.w5(32'hb735d0c3),
	.w6(32'h3809e34f),
	.w7(32'h376ed477),
	.w8(32'hb80f9e87),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3887e093),
	.w1(32'hb88e8b3f),
	.w2(32'hb61005a0),
	.w3(32'h398cccd4),
	.w4(32'h384b9055),
	.w5(32'h3878ca67),
	.w6(32'h39762435),
	.w7(32'hb77517fe),
	.w8(32'hb872f9e2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76b1282),
	.w1(32'h380dc011),
	.w2(32'h3846a330),
	.w3(32'h37fa4119),
	.w4(32'hb7fd8344),
	.w5(32'hb7741cdf),
	.w6(32'hb7d0c6b1),
	.w7(32'hb8cb8e7a),
	.w8(32'hb8e0bc0f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909c67f),
	.w1(32'hb8ae4868),
	.w2(32'hb87c0cf6),
	.w3(32'h393e62ff),
	.w4(32'hb87e0638),
	.w5(32'h38096ce0),
	.w6(32'h390cfd77),
	.w7(32'hb8aacd9c),
	.w8(32'hb91be8d6),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3852525c),
	.w1(32'h382d4d24),
	.w2(32'hb829c2ef),
	.w3(32'h3859e322),
	.w4(32'h384e0658),
	.w5(32'hb826e5b3),
	.w6(32'h387db3eb),
	.w7(32'h386b7bdc),
	.w8(32'hb81dc46f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368926a7),
	.w1(32'hb683c3b2),
	.w2(32'hb6fbb8c1),
	.w3(32'h36f28c04),
	.w4(32'hb688947e),
	.w5(32'hb66e8d7f),
	.w6(32'h35167f3a),
	.w7(32'hb67580b6),
	.w8(32'hb68abf08),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3738211a),
	.w1(32'h372ea994),
	.w2(32'hb5b94802),
	.w3(32'h36d2bd6e),
	.w4(32'h36b5b2ac),
	.w5(32'h371c2e00),
	.w6(32'h339303d0),
	.w7(32'h36ad3447),
	.w8(32'h370f1e22),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3626daf3),
	.w1(32'h36e248e3),
	.w2(32'hb56f8d2d),
	.w3(32'hb5ae40db),
	.w4(32'hb46b0d51),
	.w5(32'hb52bec30),
	.w6(32'h3607bd41),
	.w7(32'hb4533e5f),
	.w8(32'hb6a7f6de),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8570309),
	.w1(32'hb83c9746),
	.w2(32'hb72bb89f),
	.w3(32'hb6b570a4),
	.w4(32'hb8185054),
	.w5(32'hb82026ff),
	.w6(32'hb81c7740),
	.w7(32'hb89dd76a),
	.w8(32'hb8f76e7d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38205a8e),
	.w1(32'hb74e560b),
	.w2(32'hb53a6724),
	.w3(32'h3858ca4d),
	.w4(32'hb7d8f692),
	.w5(32'hb62f9a89),
	.w6(32'h37d12eba),
	.w7(32'hb8481f22),
	.w8(32'hb7d96d39),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b2f3c),
	.w1(32'h399cbc58),
	.w2(32'hb918defe),
	.w3(32'h3975a161),
	.w4(32'h39a0784e),
	.w5(32'hb885fd26),
	.w6(32'h391f0008),
	.w7(32'h39571553),
	.w8(32'hb8e1590e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ad2335),
	.w1(32'h37c4c014),
	.w2(32'hb86f2e96),
	.w3(32'h3801e63a),
	.w4(32'h38325c4a),
	.w5(32'hb82a856d),
	.w6(32'h3875ae14),
	.w7(32'h38a1746b),
	.w8(32'hb7d5cb36),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c82ee1),
	.w1(32'h36184ae5),
	.w2(32'hb745077f),
	.w3(32'h37dec2fb),
	.w4(32'hb7946ead),
	.w5(32'hb80904d2),
	.w6(32'h380b5e81),
	.w7(32'hb75c1682),
	.w8(32'hb8339df0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3731041c),
	.w1(32'hb796ba85),
	.w2(32'h36c7ed92),
	.w3(32'h3857cd86),
	.w4(32'h3744d0d5),
	.w5(32'hb6904e88),
	.w6(32'h377abbca),
	.w7(32'hb7ce56e0),
	.w8(32'hb83be061),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3780c357),
	.w1(32'hb5ca0c3e),
	.w2(32'hb7d9836c),
	.w3(32'hb76d5d95),
	.w4(32'hb75767b2),
	.w5(32'hb7b10daf),
	.w6(32'h35ae4987),
	.w7(32'hb6d2df3b),
	.w8(32'hb784bfb9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f1b0fc),
	.w1(32'h3727dd78),
	.w2(32'hb90fcee8),
	.w3(32'h38ddb58a),
	.w4(32'h38be55a8),
	.w5(32'hb8fab678),
	.w6(32'h37e16c23),
	.w7(32'hb7bd5a1e),
	.w8(32'hb9299b68),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f33d20),
	.w1(32'h390de879),
	.w2(32'hba07bd74),
	.w3(32'hb7503116),
	.w4(32'h3828fe1f),
	.w5(32'hb9e17db0),
	.w6(32'hb81be293),
	.w7(32'hba5151be),
	.w8(32'hba1b5f2f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b22f3),
	.w1(32'hbb26888f),
	.w2(32'hbb6a5833),
	.w3(32'hba04bce1),
	.w4(32'hbb3f56f5),
	.w5(32'hbb4e0fa3),
	.w6(32'hbb3c1809),
	.w7(32'hbb53a73c),
	.w8(32'hbb568937),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule