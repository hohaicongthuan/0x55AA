module layer_10_featuremap_375(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f0736),
	.w1(32'hbc0bd2a1),
	.w2(32'h3bc48bae),
	.w3(32'hbb01fd61),
	.w4(32'hbb21c9d1),
	.w5(32'h3ca41ca7),
	.w6(32'hbb0a89f6),
	.w7(32'hbbead33a),
	.w8(32'h3b214225),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa3f5d),
	.w1(32'hbbd4163b),
	.w2(32'hbc2bb5a2),
	.w3(32'hbc7d0cef),
	.w4(32'h3a025b69),
	.w5(32'h3b743584),
	.w6(32'hbc9a3894),
	.w7(32'h3b25a219),
	.w8(32'h3ab3a035),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fddcd),
	.w1(32'h3c19be24),
	.w2(32'h3c8b1eee),
	.w3(32'hb995516c),
	.w4(32'hbbfce471),
	.w5(32'hbb1a15f8),
	.w6(32'hbba71bcc),
	.w7(32'hbb7925c7),
	.w8(32'hbc36b839),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9984b7),
	.w1(32'h3c5de079),
	.w2(32'h3b948d81),
	.w3(32'hbb77610c),
	.w4(32'hbcc0f16f),
	.w5(32'hbad8bb38),
	.w6(32'hbc4cfbbc),
	.w7(32'hbbe549ce),
	.w8(32'h3b7b2991),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35267f),
	.w1(32'h3c2efe89),
	.w2(32'hbbb25081),
	.w3(32'hbcbfa542),
	.w4(32'hbb8e551b),
	.w5(32'h36eddc48),
	.w6(32'h3c756264),
	.w7(32'hba183a37),
	.w8(32'hbd14876f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbb714),
	.w1(32'h3b43a297),
	.w2(32'h3b8c3d84),
	.w3(32'hbb21099e),
	.w4(32'hbaafea74),
	.w5(32'h3c19b1ff),
	.w6(32'hbbdc6284),
	.w7(32'hbb42e4ec),
	.w8(32'hbbdc8d2d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd52164),
	.w1(32'h3b9e28c2),
	.w2(32'hba4dcaeb),
	.w3(32'h3b6d1812),
	.w4(32'h3be3f5a7),
	.w5(32'hbc53605f),
	.w6(32'hbc854a63),
	.w7(32'hbb598e93),
	.w8(32'hbcb2c025),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc654aa9),
	.w1(32'hbbe8822f),
	.w2(32'hbc40a94a),
	.w3(32'hbc5f5f35),
	.w4(32'hbcf44753),
	.w5(32'hbc46bd97),
	.w6(32'hbc7e712a),
	.w7(32'hbb72a271),
	.w8(32'hbc00aaf2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1e6e8),
	.w1(32'hbb310e16),
	.w2(32'hbc9032c1),
	.w3(32'h3b99ed6d),
	.w4(32'h3c46fe2a),
	.w5(32'hbb9df7eb),
	.w6(32'hbc380212),
	.w7(32'h3beba876),
	.w8(32'hbb3b70cf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f4b77),
	.w1(32'hbb58cd6a),
	.w2(32'hbd0f1c23),
	.w3(32'hbc0a0e2c),
	.w4(32'h3be6dcb8),
	.w5(32'hbb967626),
	.w6(32'hbcb4b521),
	.w7(32'h3c9cc674),
	.w8(32'hbc1d515f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc359f21),
	.w1(32'h3a8a553c),
	.w2(32'hbbab3a5f),
	.w3(32'h3c0cb034),
	.w4(32'hbb9d41d5),
	.w5(32'h3b068b94),
	.w6(32'h3b99679a),
	.w7(32'hba86b20d),
	.w8(32'h3a8f57e9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a0ba5),
	.w1(32'h3bc385db),
	.w2(32'hbb071df2),
	.w3(32'h3701b58e),
	.w4(32'h3c93b88b),
	.w5(32'hbbcb3e1d),
	.w6(32'hbbcb66c0),
	.w7(32'h3a6b6566),
	.w8(32'hbc925253),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28d05b),
	.w1(32'h3c63b7f9),
	.w2(32'hbc946897),
	.w3(32'hbbbd33d0),
	.w4(32'hbb6d456a),
	.w5(32'h39e1541f),
	.w6(32'h3c47e92f),
	.w7(32'h3c17b96e),
	.w8(32'hbca44531),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a390960),
	.w1(32'h3c0af4a9),
	.w2(32'h3b73d677),
	.w3(32'hbb4336d9),
	.w4(32'hbaefa19b),
	.w5(32'hbc1e7740),
	.w6(32'h3ca5e9fb),
	.w7(32'hbbdeefca),
	.w8(32'hba8edcda),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f2bbd),
	.w1(32'h3baa7295),
	.w2(32'hbc0b9530),
	.w3(32'h3c5e727e),
	.w4(32'h3bf90105),
	.w5(32'h3962a4ce),
	.w6(32'hbc925874),
	.w7(32'h3c47008d),
	.w8(32'hbb2a0e60),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc749669),
	.w1(32'h3b00b05e),
	.w2(32'hbc894eaa),
	.w3(32'hbc1452e4),
	.w4(32'h3b048691),
	.w5(32'hbc5db758),
	.w6(32'hbbc6a37f),
	.w7(32'hbae18bc4),
	.w8(32'hbc90740b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf969b5),
	.w1(32'hbb958547),
	.w2(32'h3b244ec5),
	.w3(32'h3b04f17a),
	.w4(32'h39c3ae6e),
	.w5(32'hb9564e2d),
	.w6(32'hbaa9acc2),
	.w7(32'hbbafe8b1),
	.w8(32'hb8b6afc2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf87e7),
	.w1(32'hbca6f6b5),
	.w2(32'hbcdddd1c),
	.w3(32'hbcefac79),
	.w4(32'hbb464bc1),
	.w5(32'hbc597cb5),
	.w6(32'hbc9ba449),
	.w7(32'hbd22ca75),
	.w8(32'hbc70bee1),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10bdce),
	.w1(32'hbcc80b5e),
	.w2(32'h3b494ab4),
	.w3(32'hbc4b101f),
	.w4(32'hbbfbbd6f),
	.w5(32'h3c2827ce),
	.w6(32'hbbec055a),
	.w7(32'h3afdab70),
	.w8(32'hbbb60067),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bdc8d),
	.w1(32'hbb5c4221),
	.w2(32'hbad56763),
	.w3(32'hbc443668),
	.w4(32'h3cf2da30),
	.w5(32'hb9ded411),
	.w6(32'hbab8998c),
	.w7(32'h3a822a22),
	.w8(32'h3c60c88b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfeaeee),
	.w1(32'h3b322ac7),
	.w2(32'h3cdfd27e),
	.w3(32'hbb680afa),
	.w4(32'h3b991ca4),
	.w5(32'hbb080d4b),
	.w6(32'hbc6cd7e1),
	.w7(32'hba09dcac),
	.w8(32'h3c393435),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf4adc),
	.w1(32'hbb9e4899),
	.w2(32'hbc27d907),
	.w3(32'h39af5367),
	.w4(32'h3bb46868),
	.w5(32'hbaad6cac),
	.w6(32'hbce17cfa),
	.w7(32'h3bcd74ac),
	.w8(32'h3c15d6b4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1db918),
	.w1(32'hbae3c5c4),
	.w2(32'hbd2335ab),
	.w3(32'hbce5b23d),
	.w4(32'h3b883e0a),
	.w5(32'hbc7d7f88),
	.w6(32'hbcb8c9ca),
	.w7(32'hba9d3c83),
	.w8(32'hbcc4909b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda3c1b),
	.w1(32'h3ac2a28b),
	.w2(32'hbce7b693),
	.w3(32'hbbe952ce),
	.w4(32'h3b104c7d),
	.w5(32'hbaa9a423),
	.w6(32'hbc01b964),
	.w7(32'h395eeb7e),
	.w8(32'hbc45fe44),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce80b1b),
	.w1(32'h3c013a56),
	.w2(32'hbc025468),
	.w3(32'hbc7ab130),
	.w4(32'h3c1176d3),
	.w5(32'h3a281874),
	.w6(32'hbc9b5406),
	.w7(32'h3c9a6805),
	.w8(32'hbcab6785),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5836ac),
	.w1(32'hbb1689f8),
	.w2(32'h3c0e4696),
	.w3(32'hbc737622),
	.w4(32'hbb0d6836),
	.w5(32'hbb090fd9),
	.w6(32'h3b85b786),
	.w7(32'hbb027410),
	.w8(32'hbc880301),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8441d9a),
	.w1(32'h3bf6063d),
	.w2(32'h3bf2c570),
	.w3(32'h3bf1ccb7),
	.w4(32'hb9abb393),
	.w5(32'h3b51d3d6),
	.w6(32'h3b5df558),
	.w7(32'h3c3eb2d2),
	.w8(32'h3bacc934),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0e2e3),
	.w1(32'hbb51035e),
	.w2(32'h3c8c1783),
	.w3(32'hbb8e04e7),
	.w4(32'h3c0000a7),
	.w5(32'h3cbad3a9),
	.w6(32'h3bcc927d),
	.w7(32'hbc054d63),
	.w8(32'hbb8a20bc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc230ad8),
	.w1(32'hbbf0fd7d),
	.w2(32'hbdaf69f0),
	.w3(32'hbc481645),
	.w4(32'hbc2f98a2),
	.w5(32'h3bc05d69),
	.w6(32'hba6b49c0),
	.w7(32'hbb1aa12e),
	.w8(32'h3b828b91),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b579782),
	.w1(32'h3b938cf8),
	.w2(32'h3b8d2ce8),
	.w3(32'hbc1a3d29),
	.w4(32'hbdb1486b),
	.w5(32'h3c1be0a8),
	.w6(32'hbc8c0989),
	.w7(32'h3c35cb23),
	.w8(32'h3b1f28f1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a8e8c),
	.w1(32'h3ba10b5c),
	.w2(32'h3bb02a03),
	.w3(32'h3c231ae4),
	.w4(32'hb8e66e8d),
	.w5(32'hb969d0a1),
	.w6(32'h3bd892c0),
	.w7(32'h3c49e0a3),
	.w8(32'h3cc26933),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c983f),
	.w1(32'hbb3eb6e8),
	.w2(32'h3b58b3b2),
	.w3(32'hb9e887ac),
	.w4(32'h3caa1f82),
	.w5(32'h3c204143),
	.w6(32'h3ba3328b),
	.w7(32'h3c15f6de),
	.w8(32'h3bb91bc2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec6b00),
	.w1(32'hbc385c88),
	.w2(32'h3c3ef5f5),
	.w3(32'h3c0851c2),
	.w4(32'h3bec8539),
	.w5(32'hbb923825),
	.w6(32'hbaffcfcd),
	.w7(32'hbaeceb31),
	.w8(32'hbbdb25f8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bf00b),
	.w1(32'hbc409afd),
	.w2(32'hbb4faa0c),
	.w3(32'h39e757c4),
	.w4(32'hbbb4237f),
	.w5(32'hbbda1f75),
	.w6(32'hbb9bf4b1),
	.w7(32'h3a92e9b9),
	.w8(32'hbc03f4bb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a032c),
	.w1(32'h3b7a680e),
	.w2(32'h385dd903),
	.w3(32'hbbe68315),
	.w4(32'hbcbd287d),
	.w5(32'h3beea720),
	.w6(32'h3bf9dddb),
	.w7(32'hbb99fff8),
	.w8(32'h3bedd431),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dd710),
	.w1(32'h3ccea37a),
	.w2(32'hbadbdf0e),
	.w3(32'h3bade1b0),
	.w4(32'hbc820fb6),
	.w5(32'hbc8e0e3c),
	.w6(32'h3d015d05),
	.w7(32'hbc0045c4),
	.w8(32'hbb7116c3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2b9c2),
	.w1(32'hbbc530e4),
	.w2(32'hbb358db2),
	.w3(32'hba733dcc),
	.w4(32'hbc9346be),
	.w5(32'h3cd2c8d8),
	.w6(32'h3b6c29c7),
	.w7(32'h3c4b116e),
	.w8(32'hbca8f13f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b3f04),
	.w1(32'hbb95862a),
	.w2(32'hbb43459f),
	.w3(32'hbd3fa470),
	.w4(32'h3c0cfe30),
	.w5(32'hbbc77717),
	.w6(32'hbcb64d63),
	.w7(32'h3c4f3851),
	.w8(32'h3b463f8e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd48ab02),
	.w1(32'h3ca2eb87),
	.w2(32'hbc8af36c),
	.w3(32'hbaabb11d),
	.w4(32'h3cc720e7),
	.w5(32'h380be22e),
	.w6(32'hbcac1d5d),
	.w7(32'h3bd8d98f),
	.w8(32'h3a876d2b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75e68c),
	.w1(32'h3be83500),
	.w2(32'hbc5b624c),
	.w3(32'hbbe265ec),
	.w4(32'hbd98e8a0),
	.w5(32'h3a4a18d1),
	.w6(32'hbcfa0bfa),
	.w7(32'hbae32ec7),
	.w8(32'hbb413bc9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba917a13),
	.w1(32'h3bd61c40),
	.w2(32'h3ac0c98b),
	.w3(32'hbab473f6),
	.w4(32'hbb95bddc),
	.w5(32'h3b0b8992),
	.w6(32'h3bb1d996),
	.w7(32'h3af4a073),
	.w8(32'hbb19683a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0baffc),
	.w1(32'hbc929096),
	.w2(32'hbbe0d001),
	.w3(32'hbb6ab157),
	.w4(32'h3db0a17e),
	.w5(32'h3baff640),
	.w6(32'hbbbacfaf),
	.w7(32'h39bc7fc9),
	.w8(32'h3bafd95d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc12555),
	.w1(32'hbaaf8512),
	.w2(32'hbb1dbd41),
	.w3(32'hbc53e58b),
	.w4(32'h3c5dfdf0),
	.w5(32'hbc110ade),
	.w6(32'hbc610747),
	.w7(32'h3bb8bca0),
	.w8(32'h39f96e6e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82b684),
	.w1(32'hbbfc9ab7),
	.w2(32'hbc610e20),
	.w3(32'hbc84ccb9),
	.w4(32'hba7a3d75),
	.w5(32'hbb05b61d),
	.w6(32'hbcc16942),
	.w7(32'h3c8484aa),
	.w8(32'hbc03b139),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf6be24),
	.w1(32'h3d89c4e6),
	.w2(32'hbc823109),
	.w3(32'hbc1d3add),
	.w4(32'h3c3589a3),
	.w5(32'h3c3e23f1),
	.w6(32'hbc0361bd),
	.w7(32'h3c83fc4b),
	.w8(32'hbad32d6b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccf49ad),
	.w1(32'h3c059aad),
	.w2(32'hbca44999),
	.w3(32'hbc3a6fd3),
	.w4(32'h3c8eb065),
	.w5(32'hbdc4a098),
	.w6(32'hbd6e09a3),
	.w7(32'h3cbde79d),
	.w8(32'hbc8dc0eb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd141401),
	.w1(32'h3c2905b1),
	.w2(32'hbc850af1),
	.w3(32'hbddf0dc6),
	.w4(32'h3c511478),
	.w5(32'hbd49f6ba),
	.w6(32'hbcbf7363),
	.w7(32'h3be2892d),
	.w8(32'hbbf3c25e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd45440),
	.w1(32'hbb8b00c5),
	.w2(32'hbcd79c69),
	.w3(32'hbb6c2623),
	.w4(32'hbd93406e),
	.w5(32'hbc2c1817),
	.w6(32'h3b9a959c),
	.w7(32'hbbcbce4b),
	.w8(32'h3be22d7e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca8b37),
	.w1(32'h3b11d8ec),
	.w2(32'h3bb7916b),
	.w3(32'h3b182431),
	.w4(32'h3b559a4d),
	.w5(32'hbb992005),
	.w6(32'hbb0d0bb8),
	.w7(32'h3c040ba8),
	.w8(32'h3c27e4b1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cf952),
	.w1(32'hbc542992),
	.w2(32'h3a6eff07),
	.w3(32'hba84d17a),
	.w4(32'h3c474b60),
	.w5(32'hbbff7244),
	.w6(32'h3c4e3ecc),
	.w7(32'hbc1d9c25),
	.w8(32'hbab44c99),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ed97c),
	.w1(32'h3b534a3c),
	.w2(32'h3ba0e523),
	.w3(32'hbb7889dd),
	.w4(32'h3b46d9f8),
	.w5(32'h3b107cb5),
	.w6(32'hbc00b517),
	.w7(32'hbc1e9b26),
	.w8(32'hbab2f40b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19663b),
	.w1(32'h3c0a704a),
	.w2(32'hbc782e6b),
	.w3(32'h3c5542ba),
	.w4(32'hbc4da7df),
	.w5(32'hbba83df2),
	.w6(32'hbd2c9ef5),
	.w7(32'h3abd849e),
	.w8(32'hbc74432d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842622),
	.w1(32'hbac7d3b2),
	.w2(32'hb9649256),
	.w3(32'hbb7583bf),
	.w4(32'hbb89bd88),
	.w5(32'h3bdbc849),
	.w6(32'hbb253645),
	.w7(32'hbbe45b72),
	.w8(32'h3c3bb57d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf03e8b),
	.w1(32'h3c8c2da1),
	.w2(32'hbc5d03cc),
	.w3(32'hbb9eb94a),
	.w4(32'hbb1f5e88),
	.w5(32'hbca1a761),
	.w6(32'hbbb22325),
	.w7(32'h3c52b010),
	.w8(32'hbcbb6f21),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5a1d3),
	.w1(32'h3bc33912),
	.w2(32'hbbab05aa),
	.w3(32'hbc7a620f),
	.w4(32'hbc665cfc),
	.w5(32'h3c60ad33),
	.w6(32'hbb32237e),
	.w7(32'h3bb35ca7),
	.w8(32'h39c62627),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbba2e),
	.w1(32'hb993b37d),
	.w2(32'hbbe5baaf),
	.w3(32'h38aee49b),
	.w4(32'hbc1f521c),
	.w5(32'h3b5ce3ef),
	.w6(32'h3bd0e3b7),
	.w7(32'h3bac6168),
	.w8(32'h3c2229b5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd145074),
	.w1(32'hba2830f7),
	.w2(32'hbbac90d5),
	.w3(32'h3bdaae19),
	.w4(32'h3b39b527),
	.w5(32'hbbf96f16),
	.w6(32'hbcc01c12),
	.w7(32'hba8e6483),
	.w8(32'hb94b5943),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c296176),
	.w1(32'h3a4007f9),
	.w2(32'hbb9fec76),
	.w3(32'h3caaceb0),
	.w4(32'h3bdc3413),
	.w5(32'h3b85903a),
	.w6(32'h3bd0be2d),
	.w7(32'hbb51c89f),
	.w8(32'hbc9b925b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f3271),
	.w1(32'hb99f81e9),
	.w2(32'h3a641e7e),
	.w3(32'h3c952da7),
	.w4(32'hbab3f708),
	.w5(32'hb9cba071),
	.w6(32'hbb28ef91),
	.w7(32'hbb14b045),
	.w8(32'h3b4cba35),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08ffb8),
	.w1(32'h3c959f89),
	.w2(32'h3c7616a9),
	.w3(32'hbbfeb5bb),
	.w4(32'h3ae8667d),
	.w5(32'h3a7649b6),
	.w6(32'hba17b4a6),
	.w7(32'hbb8a356a),
	.w8(32'hbb9c2b64),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4afc63),
	.w1(32'h3a8d8182),
	.w2(32'hbbc65e02),
	.w3(32'hbc6e19fa),
	.w4(32'hbbbc1528),
	.w5(32'hbb2e6b5b),
	.w6(32'hbd2385b9),
	.w7(32'hba5e22de),
	.w8(32'hba5207ab),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83f16a),
	.w1(32'hbc462708),
	.w2(32'hbb7cc607),
	.w3(32'hbca2ee9c),
	.w4(32'hbc093279),
	.w5(32'h3c9bbbd3),
	.w6(32'hbcae99ef),
	.w7(32'hbbf31907),
	.w8(32'hbb81a83e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6e35e),
	.w1(32'h3c2115b7),
	.w2(32'h3a20a137),
	.w3(32'h3ad2f215),
	.w4(32'hbad204ac),
	.w5(32'h3be8aa65),
	.w6(32'hbb492640),
	.w7(32'h39e2f4d7),
	.w8(32'hbb321106),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf4ded),
	.w1(32'hbd2644a1),
	.w2(32'h3cddce58),
	.w3(32'h3bb789f8),
	.w4(32'h3bc6c5cd),
	.w5(32'h3c1ff9e6),
	.w6(32'hbb95bdb8),
	.w7(32'hbb290b41),
	.w8(32'h3bf50f93),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49f8dc),
	.w1(32'hbc1d31e0),
	.w2(32'hbb6a65b2),
	.w3(32'h3bfc9d5c),
	.w4(32'h3bd0436a),
	.w5(32'hbc501ae7),
	.w6(32'hbbd3ebbf),
	.w7(32'hba4b5257),
	.w8(32'hbca4a798),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e22436),
	.w1(32'hb929cafc),
	.w2(32'hba000aa4),
	.w3(32'hb8e5e65e),
	.w4(32'hbb355e4b),
	.w5(32'hba36d5e7),
	.w6(32'h3c931dc8),
	.w7(32'hbc95f52f),
	.w8(32'hbaa1c6e3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b987eb),
	.w1(32'hbb6ffe19),
	.w2(32'hbc855dc8),
	.w3(32'hbcd661a1),
	.w4(32'hbd3615fe),
	.w5(32'hbbb56bfd),
	.w6(32'hbc02c948),
	.w7(32'h3bf2b30b),
	.w8(32'hbc91987f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce13cb7),
	.w1(32'hbbc3d8e5),
	.w2(32'hbcf65e24),
	.w3(32'hbc217dd2),
	.w4(32'h3b56cee9),
	.w5(32'hbc94478b),
	.w6(32'hbc69d8cb),
	.w7(32'h3c15b56c),
	.w8(32'hbc321e8c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72ac60),
	.w1(32'h3aeae963),
	.w2(32'hbbfef543),
	.w3(32'hbc866efd),
	.w4(32'h3b94796e),
	.w5(32'hbbf7b537),
	.w6(32'hbc8ec119),
	.w7(32'h3be24b7d),
	.w8(32'hbcbfae67),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01724e),
	.w1(32'h3c5a0574),
	.w2(32'hbc43f48f),
	.w3(32'hbc28f1eb),
	.w4(32'h3ca980ef),
	.w5(32'h3c76128f),
	.w6(32'hbcc7204c),
	.w7(32'h3d118faa),
	.w8(32'h3cb12dd3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabb446),
	.w1(32'hbc80fa8f),
	.w2(32'h3b8f35f0),
	.w3(32'hbc668baf),
	.w4(32'h3c3edbc5),
	.w5(32'h3b9be962),
	.w6(32'h3bfe1b87),
	.w7(32'h3c802bac),
	.w8(32'h3b823389),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3617a9),
	.w1(32'h3b92b319),
	.w2(32'h3b4ae402),
	.w3(32'hbb80553a),
	.w4(32'hbbb40753),
	.w5(32'h3bc2564c),
	.w6(32'hba827ca7),
	.w7(32'h3b09bb46),
	.w8(32'hbb88455b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e674e),
	.w1(32'h3bdd2fb0),
	.w2(32'h3bb4653f),
	.w3(32'hbb4bf41f),
	.w4(32'h3b5febbf),
	.w5(32'h3d31eff4),
	.w6(32'h3b9ce87a),
	.w7(32'h3bcc0527),
	.w8(32'h3bdd1fce),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8432e),
	.w1(32'h3a8d0afc),
	.w2(32'hbd0bfa36),
	.w3(32'hbbd45789),
	.w4(32'h3ba1c910),
	.w5(32'hbc00778e),
	.w6(32'h3c16d65a),
	.w7(32'hbc030f5b),
	.w8(32'h3a560e0c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cacf6),
	.w1(32'hbca8d8f3),
	.w2(32'h3bceca44),
	.w3(32'hbb8ed121),
	.w4(32'h3d12cbdf),
	.w5(32'hbb916bbb),
	.w6(32'hbd854559),
	.w7(32'hbbe7e6c9),
	.w8(32'h3ca1b8b6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96066d),
	.w1(32'hbc1281d9),
	.w2(32'hbae804f2),
	.w3(32'hbbeda34f),
	.w4(32'hbbc76d5f),
	.w5(32'hbbf0043e),
	.w6(32'h3c6b736d),
	.w7(32'hbb0e1d7b),
	.w8(32'h3bff468e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf0a30),
	.w1(32'hbcdb08be),
	.w2(32'hbc242c56),
	.w3(32'hbc2e479e),
	.w4(32'h3c1b3190),
	.w5(32'hbbb96476),
	.w6(32'hbc1b2999),
	.w7(32'hbb9cc5bb),
	.w8(32'hbbca128f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc84169),
	.w1(32'hbc00637e),
	.w2(32'hbc0944b1),
	.w3(32'h3ae485ab),
	.w4(32'h3c0f9a9e),
	.w5(32'hba80403c),
	.w6(32'h3b7c99f6),
	.w7(32'h3b84fad5),
	.w8(32'hbbf5fe46),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d78d7),
	.w1(32'hbb2c22cd),
	.w2(32'hbbe30fba),
	.w3(32'h3c978dfb),
	.w4(32'h3a3f7ef3),
	.w5(32'hb9b72d92),
	.w6(32'hbb855ad4),
	.w7(32'h3a481d59),
	.w8(32'h3bdcd89f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0f717),
	.w1(32'h3bc34eff),
	.w2(32'hbc3c12f8),
	.w3(32'hba770f51),
	.w4(32'h3ba92cb4),
	.w5(32'hbc50e12b),
	.w6(32'h3a1cbf96),
	.w7(32'h3d28b941),
	.w8(32'hbb62a731),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe970a1),
	.w1(32'h3c36c442),
	.w2(32'hbc08d19f),
	.w3(32'hbb98ed2f),
	.w4(32'hbc1e30e8),
	.w5(32'h3c548bbe),
	.w6(32'hbbf1bd21),
	.w7(32'h3c3a65cc),
	.w8(32'h3c0cbf22),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc5527),
	.w1(32'h3c38408f),
	.w2(32'hbb1a6720),
	.w3(32'hba0d68c2),
	.w4(32'hbc335373),
	.w5(32'hbc6881e9),
	.w6(32'hbc007255),
	.w7(32'h3b4a4906),
	.w8(32'hbb7bcef2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a306da7),
	.w1(32'h3b39af36),
	.w2(32'h3b95cdfd),
	.w3(32'h3b7e98e8),
	.w4(32'hbba450a6),
	.w5(32'hbb8c6057),
	.w6(32'hbb66c5ac),
	.w7(32'hbb7c0dd4),
	.w8(32'hbaf90cd4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd857af),
	.w1(32'h3b5d6dda),
	.w2(32'hbbe2f47a),
	.w3(32'h3bb0c822),
	.w4(32'hbb1108df),
	.w5(32'hbb68446c),
	.w6(32'h39b797cb),
	.w7(32'hbb22e19f),
	.w8(32'hbc3bd216),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb21493),
	.w1(32'h3b1a177d),
	.w2(32'hbce76a7d),
	.w3(32'hbb52259c),
	.w4(32'hbb8c2f9e),
	.w5(32'hbbefe219),
	.w6(32'hbc1ef2e2),
	.w7(32'h3973d6eb),
	.w8(32'hbb653698),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac696a2),
	.w1(32'h39a0f2b1),
	.w2(32'hbbb5592a),
	.w3(32'h3c10150d),
	.w4(32'hbb9b757d),
	.w5(32'hbbd014f5),
	.w6(32'hba6b86b0),
	.w7(32'h3c92bb5d),
	.w8(32'h3ade6fe4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc986500),
	.w1(32'h3aee1870),
	.w2(32'hbc188369),
	.w3(32'h3c22e319),
	.w4(32'h3bfab058),
	.w5(32'hbaf5dfbb),
	.w6(32'hbbe2fc69),
	.w7(32'hbc0a2ca0),
	.w8(32'hbb11cb85),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8795c7),
	.w1(32'h3b15a474),
	.w2(32'h39bb2e89),
	.w3(32'h3c20d69b),
	.w4(32'h38a1684a),
	.w5(32'h3cc4f1e3),
	.w6(32'hbc5a53d4),
	.w7(32'h39b1f862),
	.w8(32'hbadef46f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc603d9b),
	.w1(32'hbc721bf9),
	.w2(32'hbbe94e2f),
	.w3(32'hbc1d66d9),
	.w4(32'h3c354a8b),
	.w5(32'hbbfc455a),
	.w6(32'hbba9a1bd),
	.w7(32'h3bf2f647),
	.w8(32'h3b6e78ac),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8f61f),
	.w1(32'hbb8b5889),
	.w2(32'hbcbcf367),
	.w3(32'hbcad472a),
	.w4(32'hbd7dfd0f),
	.w5(32'hbc7801e6),
	.w6(32'hbca6ef99),
	.w7(32'h3a8c90f1),
	.w8(32'hbc31fefa),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe58c),
	.w1(32'h383d4709),
	.w2(32'h3ae5c71a),
	.w3(32'hbb2b4675),
	.w4(32'h3c0cd40c),
	.w5(32'h3bbe806b),
	.w6(32'hbd6cdeac),
	.w7(32'h3c4fb4c8),
	.w8(32'hbc1ea724),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a6253),
	.w1(32'hbb2e45fd),
	.w2(32'hbbf6304b),
	.w3(32'hbb08ba74),
	.w4(32'hbb51f12d),
	.w5(32'h3d27c036),
	.w6(32'hbc381c39),
	.w7(32'hbb40ce1d),
	.w8(32'hbc95fbfb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2cc2b),
	.w1(32'h3b526907),
	.w2(32'hbb948408),
	.w3(32'hbc391ffe),
	.w4(32'h3c5cb7d0),
	.w5(32'h387578e8),
	.w6(32'h3c2b8d04),
	.w7(32'h3c0bcb08),
	.w8(32'h3aaefb6b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e6e09),
	.w1(32'h3c6d1bee),
	.w2(32'hbb65cc10),
	.w3(32'hbca86db1),
	.w4(32'h3c4b612d),
	.w5(32'hbc5c3605),
	.w6(32'hbca2b78b),
	.w7(32'hbc09f8f6),
	.w8(32'hbc547073),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce5c15),
	.w1(32'hbcc28704),
	.w2(32'hbb618532),
	.w3(32'hbc7c2e30),
	.w4(32'h3c24ed4e),
	.w5(32'hbc72e8a9),
	.w6(32'hba7cf5f4),
	.w7(32'hbc143b00),
	.w8(32'hbc4da88a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48ebf2),
	.w1(32'hbb312584),
	.w2(32'h3baec337),
	.w3(32'hbbdc769f),
	.w4(32'h3cb7ed92),
	.w5(32'hbca9f06c),
	.w6(32'hbc5e9eeb),
	.w7(32'h3c527023),
	.w8(32'h3b43b85f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18f9c5),
	.w1(32'hbb12d340),
	.w2(32'hbb611a14),
	.w3(32'hbb80545c),
	.w4(32'hb97ad3dc),
	.w5(32'hbc237c8e),
	.w6(32'h39c3305d),
	.w7(32'hb87a4e99),
	.w8(32'hba93e9df),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c5185),
	.w1(32'hbbc1820d),
	.w2(32'hbc8e559c),
	.w3(32'hbb357917),
	.w4(32'h3c8161f8),
	.w5(32'hba2dd974),
	.w6(32'hbc546813),
	.w7(32'h3c5a4253),
	.w8(32'hbb875201),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bacac),
	.w1(32'h3c80401e),
	.w2(32'hbca0e1a2),
	.w3(32'hbc2ee7c6),
	.w4(32'h3892026b),
	.w5(32'h3c0a9476),
	.w6(32'hbc3c7907),
	.w7(32'h3bd0a4c5),
	.w8(32'hbb660151),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8468b9),
	.w1(32'hbc2da171),
	.w2(32'hbcc2717c),
	.w3(32'hbc1835be),
	.w4(32'h3a376918),
	.w5(32'hbc77eaa0),
	.w6(32'hbc2dee09),
	.w7(32'hbaf2e92e),
	.w8(32'hbc061ee6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8181e),
	.w1(32'hbbeec1dc),
	.w2(32'h3b32d922),
	.w3(32'hbcb084bb),
	.w4(32'h3c41c7e0),
	.w5(32'h39f0c8bb),
	.w6(32'hbcc37371),
	.w7(32'hba5363ec),
	.w8(32'hbc5b9c0e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cbde1),
	.w1(32'h3c2cb52b),
	.w2(32'h3b340270),
	.w3(32'hbc23fe4b),
	.w4(32'h3c9cefaf),
	.w5(32'h3900e5e8),
	.w6(32'h3b726106),
	.w7(32'h3c8fcb85),
	.w8(32'h3aa7d9b3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc714f9d),
	.w1(32'h3ab526c3),
	.w2(32'hbbab1e8e),
	.w3(32'hbcfd1cd9),
	.w4(32'h3bd04bac),
	.w5(32'hbca30a24),
	.w6(32'hbbba9e31),
	.w7(32'hbc810d54),
	.w8(32'hbd90d452),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1e96b),
	.w1(32'h3c9a64bb),
	.w2(32'h3c2e5ee7),
	.w3(32'h3b06f7de),
	.w4(32'h3c74d4a4),
	.w5(32'hbbb408f8),
	.w6(32'h3bd53e9f),
	.w7(32'hbbe28e00),
	.w8(32'hbbf8033f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca200d1),
	.w1(32'hbc360af4),
	.w2(32'hbc9f8ee0),
	.w3(32'hbbc3f94c),
	.w4(32'hbc60be65),
	.w5(32'h3d1509c7),
	.w6(32'h3c1e2c35),
	.w7(32'h36a7c260),
	.w8(32'h3be3478a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba985a99),
	.w1(32'hbb837ab5),
	.w2(32'hbb3bd55f),
	.w3(32'hbc08b858),
	.w4(32'hbbced91b),
	.w5(32'h3c014a49),
	.w6(32'hbc2a5bc2),
	.w7(32'hb942baf1),
	.w8(32'hbb9646b3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd87720),
	.w1(32'h3b09d06a),
	.w2(32'h3be1dbb9),
	.w3(32'hbba6f6b4),
	.w4(32'hbb08e7cf),
	.w5(32'hbba5d8a6),
	.w6(32'hba1644ac),
	.w7(32'hbbe8ac15),
	.w8(32'h3b399d20),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff4b2f),
	.w1(32'hb9d9d3cb),
	.w2(32'hbb46f379),
	.w3(32'h3ac1d0c8),
	.w4(32'hbb37f091),
	.w5(32'h3b6d4089),
	.w6(32'h3bd9cc08),
	.w7(32'h3a62b7a5),
	.w8(32'hbb7f21b1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c5ce1),
	.w1(32'hbb1c0606),
	.w2(32'hbc26f621),
	.w3(32'hbc60ff79),
	.w4(32'h3aaa4e3f),
	.w5(32'hbc470b26),
	.w6(32'hbcca7638),
	.w7(32'hbbd824ad),
	.w8(32'hbc23d9f0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc981665),
	.w1(32'h3c2a944e),
	.w2(32'h3c1e98d3),
	.w3(32'hbc4e50de),
	.w4(32'h3b86132d),
	.w5(32'hbc9774d1),
	.w6(32'hbc871860),
	.w7(32'h3c04cfbc),
	.w8(32'h3c39412a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7302b),
	.w1(32'hbcad6555),
	.w2(32'hbc4f156a),
	.w3(32'h3b8242ae),
	.w4(32'hbb9263ad),
	.w5(32'hbb512481),
	.w6(32'hbcb4805e),
	.w7(32'hbc214ac3),
	.w8(32'hbad7aae9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e699a),
	.w1(32'hbb02907f),
	.w2(32'hbc29d278),
	.w3(32'hbb62e3ff),
	.w4(32'h3bec2b53),
	.w5(32'hbb851614),
	.w6(32'hbbbb6e76),
	.w7(32'h3b32d11a),
	.w8(32'hb9b66b01),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fa6d1),
	.w1(32'h3b4198b2),
	.w2(32'h3c504f21),
	.w3(32'h39ffc3af),
	.w4(32'hbb26292b),
	.w5(32'hbbdc0426),
	.w6(32'hbaac0857),
	.w7(32'h3c2a55a8),
	.w8(32'hbc0059c9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd17d33c),
	.w1(32'h3bd308ce),
	.w2(32'hbc882b5c),
	.w3(32'hbafd4880),
	.w4(32'h3c07768d),
	.w5(32'h3b3139da),
	.w6(32'hbbdfca5a),
	.w7(32'hbd2e5fd6),
	.w8(32'hbb4b2e9d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a45dc),
	.w1(32'hbc8bd041),
	.w2(32'h3bb4ea0f),
	.w3(32'hbc0c9d54),
	.w4(32'h3a9e6c5d),
	.w5(32'hbbfa0630),
	.w6(32'hbc6abf25),
	.w7(32'h3cbe1bce),
	.w8(32'h3af3a116),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60d624),
	.w1(32'hbbfd2b43),
	.w2(32'h3c3149c4),
	.w3(32'h3c115a64),
	.w4(32'hbbec7c4d),
	.w5(32'hbbad3113),
	.w6(32'h3c7cdd04),
	.w7(32'hba3f3c0d),
	.w8(32'h3bc1debb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb902c12),
	.w1(32'hbcc09b18),
	.w2(32'hbca77488),
	.w3(32'h3bd0e7d3),
	.w4(32'hbb961dcc),
	.w5(32'hbb6d6fa3),
	.w6(32'h3b983a1f),
	.w7(32'h3b81e392),
	.w8(32'hbb994e06),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda0b98),
	.w1(32'h3b67c1b1),
	.w2(32'h3ab66b71),
	.w3(32'h3d16191f),
	.w4(32'hb970ff4f),
	.w5(32'hbc281aa8),
	.w6(32'hbcac6584),
	.w7(32'h3d2d505b),
	.w8(32'hbcdc4c6e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13870d),
	.w1(32'h3b89dbee),
	.w2(32'hbc45cd6d),
	.w3(32'h3cc8a06d),
	.w4(32'hbc0ac77b),
	.w5(32'hbc90bc04),
	.w6(32'h3bf40aaa),
	.w7(32'h3b25a1dd),
	.w8(32'h3c36dbdc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be837bb),
	.w1(32'hbb2ad610),
	.w2(32'h3b1dbc10),
	.w3(32'hbb927dae),
	.w4(32'h3c920ba1),
	.w5(32'hbbe743e1),
	.w6(32'hbc33747b),
	.w7(32'h3c61e7e4),
	.w8(32'hbc101dd6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36416b),
	.w1(32'h3bb87b15),
	.w2(32'h3b75eb53),
	.w3(32'h3b0fa4a3),
	.w4(32'hba618a00),
	.w5(32'hbc217ca9),
	.w6(32'hbc58c493),
	.w7(32'hbb4f25c1),
	.w8(32'hbd0dcb23),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb24d99),
	.w1(32'h3b92dab3),
	.w2(32'hbb6697d2),
	.w3(32'h3b9340a3),
	.w4(32'h3b966722),
	.w5(32'hbc3b1982),
	.w6(32'hbb0483cb),
	.w7(32'h3b5cddfe),
	.w8(32'h3aa8dda9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08d047),
	.w1(32'h3aca0f4a),
	.w2(32'hbb9c4557),
	.w3(32'hbbd9b46c),
	.w4(32'hbb63279a),
	.w5(32'hbbb50c38),
	.w6(32'hbad15936),
	.w7(32'hbb0775a0),
	.w8(32'h3c3ec3c6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9452bb),
	.w1(32'h3c34b054),
	.w2(32'h3b7b7317),
	.w3(32'hbab282dd),
	.w4(32'h3a99d416),
	.w5(32'hbb8186d9),
	.w6(32'h3cea22dc),
	.w7(32'hbc8fce71),
	.w8(32'h3aa97f84),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5d0e8),
	.w1(32'hbb21f082),
	.w2(32'hbb6cdecd),
	.w3(32'hbabb655b),
	.w4(32'hbb823dc3),
	.w5(32'hbba4f2c7),
	.w6(32'hbc8ebb68),
	.w7(32'hbbba2e9f),
	.w8(32'h3a04b811),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a8107),
	.w1(32'hb938f750),
	.w2(32'hbc5a8340),
	.w3(32'h3b4191e1),
	.w4(32'h3b063522),
	.w5(32'hbc44f2e8),
	.w6(32'hbc46a99e),
	.w7(32'h3bbe5978),
	.w8(32'h3c7e4312),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80b91b),
	.w1(32'h3bb915d7),
	.w2(32'hbcaf92c5),
	.w3(32'h3c908087),
	.w4(32'hbc5e71e7),
	.w5(32'h3bdd8e41),
	.w6(32'hbb93051e),
	.w7(32'hbbf7f7e3),
	.w8(32'hbc298d71),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c3946),
	.w1(32'hbb2ec47b),
	.w2(32'hbc963e4b),
	.w3(32'h3b2c9b6d),
	.w4(32'hbcd4da1d),
	.w5(32'hbc83dba2),
	.w6(32'hbb014744),
	.w7(32'hbc535ec8),
	.w8(32'hbc9e04a5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc99b93),
	.w1(32'hbb84b2ab),
	.w2(32'hbc7399f6),
	.w3(32'hbc41f600),
	.w4(32'h3c0de546),
	.w5(32'h3cdfbf68),
	.w6(32'h3b825f04),
	.w7(32'hbb8f0d54),
	.w8(32'h399c7b14),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf0c655),
	.w1(32'h3a988ba8),
	.w2(32'h3bea5ecf),
	.w3(32'hbb979e38),
	.w4(32'hb93bbc63),
	.w5(32'hbb872368),
	.w6(32'h3b1c498a),
	.w7(32'h392bd114),
	.w8(32'h3c12a41f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22a957),
	.w1(32'h3b0c9d50),
	.w2(32'hbb3e750b),
	.w3(32'hbc45c87d),
	.w4(32'hbbcba353),
	.w5(32'h3bd9d440),
	.w6(32'hbbc44326),
	.w7(32'h3a980c3b),
	.w8(32'hbc924517),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc278ea6),
	.w1(32'hbc3014d2),
	.w2(32'hbc10ce4f),
	.w3(32'hbb920f3e),
	.w4(32'hbb514537),
	.w5(32'hb924d477),
	.w6(32'hbc938d06),
	.w7(32'hbb04669d),
	.w8(32'hbb9d7596),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c87d9),
	.w1(32'h3b17ec9f),
	.w2(32'hbaab88a8),
	.w3(32'hbc98fa56),
	.w4(32'hbc9f2459),
	.w5(32'hbbff644f),
	.w6(32'hbb8c4946),
	.w7(32'hbba79449),
	.w8(32'hbc476a2b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc983d36),
	.w1(32'hbaeee27f),
	.w2(32'hbba88e7c),
	.w3(32'h3b959679),
	.w4(32'hba84a014),
	.w5(32'hbb406bbc),
	.w6(32'hbc385705),
	.w7(32'h3c1ac645),
	.w8(32'hbca72922),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca005b2),
	.w1(32'hbc69e5fc),
	.w2(32'hbca0c92a),
	.w3(32'hbc04daab),
	.w4(32'h3c161e81),
	.w5(32'hbc440555),
	.w6(32'hba5a2900),
	.w7(32'hbbd9fca7),
	.w8(32'hbc2e5629),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a6c05),
	.w1(32'h3b0a5675),
	.w2(32'h3bc03b18),
	.w3(32'hbc99edac),
	.w4(32'h3ab11a2b),
	.w5(32'h3b99d542),
	.w6(32'hbb8bfead),
	.w7(32'h3c38f2d5),
	.w8(32'h39801389),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dde4e),
	.w1(32'hbc354727),
	.w2(32'h3afd6777),
	.w3(32'hbc011b94),
	.w4(32'h3ba136cd),
	.w5(32'hba0b66f7),
	.w6(32'hbaadf4e6),
	.w7(32'hbb56396d),
	.w8(32'hbbb50c50),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca083d0),
	.w1(32'h3b849e3a),
	.w2(32'h3b3b93fb),
	.w3(32'hbbfe7938),
	.w4(32'h3b01281c),
	.w5(32'hbc490b1e),
	.w6(32'hbc80975c),
	.w7(32'hbb07d27e),
	.w8(32'hbabeaa3a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3df0),
	.w1(32'hbb1b9bb4),
	.w2(32'h39a6769e),
	.w3(32'hbb39e9eb),
	.w4(32'h3c666994),
	.w5(32'h3b5a6c62),
	.w6(32'hbcb75d67),
	.w7(32'h3b7636c8),
	.w8(32'hbc4ac69f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23aea4),
	.w1(32'hbbdedb63),
	.w2(32'hbca75756),
	.w3(32'hbad7f71f),
	.w4(32'h3c64e560),
	.w5(32'hbc675bcd),
	.w6(32'hbc11ac9c),
	.w7(32'hbb8525db),
	.w8(32'h3c6524a7),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cc3bc),
	.w1(32'h3c57a827),
	.w2(32'hbb2b0d05),
	.w3(32'hbc1c2bb2),
	.w4(32'h3bc7b7fd),
	.w5(32'hbb163fd6),
	.w6(32'h3c1d3aef),
	.w7(32'hbaef244d),
	.w8(32'hba162e04),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc550252),
	.w1(32'h3c9a59eb),
	.w2(32'hbc23eb2f),
	.w3(32'hbcafa9c8),
	.w4(32'h3cd9bbd4),
	.w5(32'hbbcb529a),
	.w6(32'hbb97dfc4),
	.w7(32'h3cafe600),
	.w8(32'hbb28087d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3b5ef),
	.w1(32'hbbb2c3b4),
	.w2(32'h3ba91eff),
	.w3(32'hbc58f838),
	.w4(32'hbcdf526d),
	.w5(32'hbacaa8e8),
	.w6(32'hbbfaa0bf),
	.w7(32'h3b8f1586),
	.w8(32'h3a8b7d96),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c21dc),
	.w1(32'hbc07c648),
	.w2(32'h3a284f19),
	.w3(32'h3bf2e8b1),
	.w4(32'hb99b356e),
	.w5(32'h3a0f1076),
	.w6(32'h3c412aab),
	.w7(32'hbb08243a),
	.w8(32'hbb0b0970),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74bc4b),
	.w1(32'h3c592705),
	.w2(32'hbae665d5),
	.w3(32'h3a512e9d),
	.w4(32'hbc37f256),
	.w5(32'h3bb5c278),
	.w6(32'h3b6a7cad),
	.w7(32'hbbcdaf90),
	.w8(32'hbb61a014),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fe588),
	.w1(32'hbc16aff4),
	.w2(32'h3b908a8d),
	.w3(32'hbb99c9e8),
	.w4(32'h3c19273b),
	.w5(32'h3c1bffe1),
	.w6(32'hbc51b114),
	.w7(32'hbbd1eb8b),
	.w8(32'h3b0359c3),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc196ab),
	.w1(32'hbc1bf1b5),
	.w2(32'h3b24c833),
	.w3(32'hbc82229f),
	.w4(32'h3c233a66),
	.w5(32'hb999fe58),
	.w6(32'hbc3bdb83),
	.w7(32'hbc1c0e3c),
	.w8(32'hbbc6a464),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fd4fd),
	.w1(32'hb9e8b24d),
	.w2(32'hbc7a5f1e),
	.w3(32'h3c6924ea),
	.w4(32'h3b12ddec),
	.w5(32'hbc428830),
	.w6(32'hbb4a24a2),
	.w7(32'h3c82e67d),
	.w8(32'hbbdbcb22),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef49cb),
	.w1(32'h3ca8eaf0),
	.w2(32'hbc00beaa),
	.w3(32'h3b92234f),
	.w4(32'hbb97cbab),
	.w5(32'h3b6e0b02),
	.w6(32'hbb7baba6),
	.w7(32'h3b6a91bf),
	.w8(32'hbb8d8932),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0183d1),
	.w1(32'h3ba03550),
	.w2(32'h3b92a718),
	.w3(32'hbbabee34),
	.w4(32'h3b4717fa),
	.w5(32'hbbe641bc),
	.w6(32'hbba9129d),
	.w7(32'h3b864877),
	.w8(32'hbba1b274),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d494f),
	.w1(32'hb79b4582),
	.w2(32'hbc228e37),
	.w3(32'hbbaae2e9),
	.w4(32'h3ca65275),
	.w5(32'h3b4758ea),
	.w6(32'hbb62e051),
	.w7(32'hbbe79431),
	.w8(32'hbcf41d4f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a1e66),
	.w1(32'h3c1bdf3f),
	.w2(32'hbc37aa3b),
	.w3(32'hbc0dafc7),
	.w4(32'h3a1ac973),
	.w5(32'h3a54ec35),
	.w6(32'h3abc496a),
	.w7(32'h3ab35493),
	.w8(32'hbd10015a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc38a),
	.w1(32'h3c1ea8f9),
	.w2(32'hbc7c5a37),
	.w3(32'hbb9a515a),
	.w4(32'h3cb5f49b),
	.w5(32'hb9cee2bf),
	.w6(32'hbba340e4),
	.w7(32'h3cbf60b9),
	.w8(32'h3b662ac1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0d7fa),
	.w1(32'hbb8a4852),
	.w2(32'h3b5bc5ef),
	.w3(32'h3d039ce9),
	.w4(32'h3afc2238),
	.w5(32'hbb17825c),
	.w6(32'hbc47f681),
	.w7(32'hba30bd2a),
	.w8(32'h3c78eab4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b486290),
	.w1(32'hb9c02a9b),
	.w2(32'h3bb881f5),
	.w3(32'hbbbbd98e),
	.w4(32'h3c102fe1),
	.w5(32'hbb52e3a9),
	.w6(32'h3ccb508c),
	.w7(32'h3b9b1432),
	.w8(32'hbb811820),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf24750),
	.w1(32'h3c2bdbfc),
	.w2(32'hbab81698),
	.w3(32'hbb736584),
	.w4(32'hbcdca472),
	.w5(32'h3c6a601d),
	.w6(32'hbcd3da1e),
	.w7(32'h3cb93735),
	.w8(32'h3adac734),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5c636),
	.w1(32'h3b57a638),
	.w2(32'hbc69b7d0),
	.w3(32'hbc60648a),
	.w4(32'h3b017c88),
	.w5(32'hbbb4d400),
	.w6(32'hbc207694),
	.w7(32'h3b134b8b),
	.w8(32'hbb2a6d9f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fefbae),
	.w1(32'hbb8b05a3),
	.w2(32'hba5d3da0),
	.w3(32'hbbaf81c3),
	.w4(32'h3a135f56),
	.w5(32'hbc17da19),
	.w6(32'hba7eb699),
	.w7(32'h3bd914d9),
	.w8(32'hbb2bc250),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74086b),
	.w1(32'h3b8bbc93),
	.w2(32'hbb41e04d),
	.w3(32'hbc7dff16),
	.w4(32'hbb095acd),
	.w5(32'hbbafd98a),
	.w6(32'hb9189dc5),
	.w7(32'h3bc149c2),
	.w8(32'h3b4e7753),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fabf2),
	.w1(32'h3b21bd40),
	.w2(32'h3c66415a),
	.w3(32'hb98b5115),
	.w4(32'h3935373a),
	.w5(32'h3ca34614),
	.w6(32'h3bf2059c),
	.w7(32'h3b884bf3),
	.w8(32'hbb942f02),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19291f),
	.w1(32'hbba723f6),
	.w2(32'hbc1d01e3),
	.w3(32'hb9f59b4a),
	.w4(32'h3c0f0aac),
	.w5(32'hbc011f1b),
	.w6(32'hba7707f1),
	.w7(32'hbc56dfa7),
	.w8(32'h3c25103a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b3947),
	.w1(32'hbb9ac29d),
	.w2(32'hbcbc2ee1),
	.w3(32'h3c17ee2c),
	.w4(32'hbbe5b801),
	.w5(32'h3b4d9349),
	.w6(32'hbc6ee768),
	.w7(32'h3b7f2bf6),
	.w8(32'h3bfbeeaa),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9800fa6),
	.w1(32'h3c318be4),
	.w2(32'h3ab55b42),
	.w3(32'hbca2f61a),
	.w4(32'hba7d9d0e),
	.w5(32'h3a0c776a),
	.w6(32'hbc2c36e9),
	.w7(32'hbbb9cbda),
	.w8(32'hbccf22e7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9375d6),
	.w1(32'h3bbc22a6),
	.w2(32'hbb0737e5),
	.w3(32'hbbbbebcf),
	.w4(32'hbb9121e0),
	.w5(32'h3a9b47c1),
	.w6(32'h3b293786),
	.w7(32'h3b7add79),
	.w8(32'hbc30b442),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850aef),
	.w1(32'hba9bbf65),
	.w2(32'hbb2f6106),
	.w3(32'hbb72efd3),
	.w4(32'hba84b161),
	.w5(32'hbbe9d9dc),
	.w6(32'h3a5f85ac),
	.w7(32'hba0017d4),
	.w8(32'hbc8bf6a4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4910c),
	.w1(32'h3b29ee95),
	.w2(32'hbb39bccb),
	.w3(32'hbc33e161),
	.w4(32'hb7a99b8f),
	.w5(32'h3bfd7dcb),
	.w6(32'hbb050687),
	.w7(32'hbb77a793),
	.w8(32'h3bb76c6a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe4def),
	.w1(32'h3b3e2f61),
	.w2(32'hbc222bf9),
	.w3(32'hbbff7a3c),
	.w4(32'h3b60e44e),
	.w5(32'h39ecf69d),
	.w6(32'h3a58f504),
	.w7(32'h3aeb677e),
	.w8(32'h3b28f6b8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcf2ee),
	.w1(32'h3b1c74c5),
	.w2(32'hbc24f519),
	.w3(32'h3c0ee081),
	.w4(32'h3c208ecc),
	.w5(32'hba06a631),
	.w6(32'hbb00796a),
	.w7(32'hbbd8941a),
	.w8(32'h3c3591cb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca241f7),
	.w1(32'h3c16d208),
	.w2(32'hbc630f5e),
	.w3(32'hbbfd60cf),
	.w4(32'h3b950afc),
	.w5(32'hbc92d1b7),
	.w6(32'hbc327b0b),
	.w7(32'h3bd6ac97),
	.w8(32'hbb9924a2),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac64e54),
	.w1(32'hbb49e39a),
	.w2(32'hbb9ddc9c),
	.w3(32'hbba1fbf6),
	.w4(32'hba5abb89),
	.w5(32'hbad1e130),
	.w6(32'h3aa991fb),
	.w7(32'hbc8138e3),
	.w8(32'hbb585b75),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c9f0a),
	.w1(32'hbbe26ec7),
	.w2(32'hbc055821),
	.w3(32'hbb78d143),
	.w4(32'hbbbc84c5),
	.w5(32'hbadddc56),
	.w6(32'h3b2f5336),
	.w7(32'h3c0e836e),
	.w8(32'hba142877),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbceaf25),
	.w1(32'hbb5af952),
	.w2(32'h3a3e822a),
	.w3(32'h3b9b3e94),
	.w4(32'h3b8e64d8),
	.w5(32'h39810934),
	.w6(32'hba232d76),
	.w7(32'h3c072535),
	.w8(32'h3b8a83d7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8ca2d),
	.w1(32'hbc25bea5),
	.w2(32'hbcda5bbf),
	.w3(32'hbbf9795a),
	.w4(32'h3c4af85b),
	.w5(32'hbc82dcbe),
	.w6(32'hbcbc19a1),
	.w7(32'h3ba16c19),
	.w8(32'hbc843635),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62aa64),
	.w1(32'hba984ff9),
	.w2(32'hbca45b4f),
	.w3(32'hbbc25e1e),
	.w4(32'h3a27af30),
	.w5(32'hbc70ff8d),
	.w6(32'hbb01b29d),
	.w7(32'h3c30828d),
	.w8(32'hbbab888d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3d125),
	.w1(32'hbc2e749b),
	.w2(32'hbbf4116c),
	.w3(32'hbc8eb431),
	.w4(32'h3c9454d3),
	.w5(32'hbca8fb36),
	.w6(32'hbbc6fbc9),
	.w7(32'h3af90e83),
	.w8(32'hbc3d5a7c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5946e4),
	.w1(32'hbaa6d73a),
	.w2(32'h3a46ed84),
	.w3(32'hb9e69b26),
	.w4(32'hbaecb136),
	.w5(32'h3bbf666f),
	.w6(32'h3c6c8907),
	.w7(32'hbbbe6852),
	.w8(32'hbc05ae0d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc31eb8),
	.w1(32'h3b1c95c2),
	.w2(32'hbb588aa2),
	.w3(32'hbad2f096),
	.w4(32'hbc8e8484),
	.w5(32'hbc1ca99a),
	.w6(32'hbb0343d0),
	.w7(32'h3c02373c),
	.w8(32'h3b8ce048),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba223f04),
	.w1(32'hbc6700e8),
	.w2(32'hb977c758),
	.w3(32'hbbebc7c1),
	.w4(32'h3bfdb326),
	.w5(32'h3c0703fe),
	.w6(32'hbb17f8d1),
	.w7(32'hbc3b9f20),
	.w8(32'hbc027b6d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf08815),
	.w1(32'h3b96ca44),
	.w2(32'h3a3bd6ef),
	.w3(32'hbb7a488f),
	.w4(32'h3a7a5694),
	.w5(32'h3ba013de),
	.w6(32'hbaf34c30),
	.w7(32'hbb28b835),
	.w8(32'hbbba8edc),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5082e),
	.w1(32'hbbbed377),
	.w2(32'hbc5d1db0),
	.w3(32'hbc85d9eb),
	.w4(32'h3cab3dcb),
	.w5(32'h3cf992f7),
	.w6(32'hbad1ddb7),
	.w7(32'hbb80fbeb),
	.w8(32'h3c6f869e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc571a30),
	.w1(32'hbaef9e0d),
	.w2(32'hbc3ba6d5),
	.w3(32'hbc53022d),
	.w4(32'h3b886c71),
	.w5(32'h3c29fdc6),
	.w6(32'hba4dc45d),
	.w7(32'h3c0574cf),
	.w8(32'h3b12627e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038330),
	.w1(32'h3c3fd6ad),
	.w2(32'h3bf2a14c),
	.w3(32'h3bb94bd2),
	.w4(32'h3b991932),
	.w5(32'h3b3e5754),
	.w6(32'h3bfd57d1),
	.w7(32'h3bb080a2),
	.w8(32'h3bf0e607),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc391054),
	.w1(32'hbb190c8f),
	.w2(32'h3c3cbca2),
	.w3(32'hbbb15376),
	.w4(32'hba5bef94),
	.w5(32'hbb6ed2db),
	.w6(32'h3934bcfd),
	.w7(32'hbc6960fc),
	.w8(32'h3bbd5e1b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14bb8d),
	.w1(32'hbc1688c9),
	.w2(32'hbbd0a83e),
	.w3(32'hba846a37),
	.w4(32'hbc0c88c0),
	.w5(32'hbb82f5c9),
	.w6(32'hbb904880),
	.w7(32'h3af5e60b),
	.w8(32'hbceaa043),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e2ca1),
	.w1(32'h3c174a3d),
	.w2(32'hbc93cbfb),
	.w3(32'hbc96ee7c),
	.w4(32'hbb8c372e),
	.w5(32'hbc97748f),
	.w6(32'hbc8cc00e),
	.w7(32'h3c95eb4f),
	.w8(32'hbacf27af),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd8223),
	.w1(32'h3b17c39c),
	.w2(32'h39e21969),
	.w3(32'hba69d14e),
	.w4(32'h3a2f1015),
	.w5(32'hbc532ec7),
	.w6(32'h3c01b10a),
	.w7(32'h3b85b791),
	.w8(32'hbc2eb291),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b281c63),
	.w1(32'h3aafcfa3),
	.w2(32'hbb280e45),
	.w3(32'hbb7f2e37),
	.w4(32'h3b1c0754),
	.w5(32'h3c05b70d),
	.w6(32'h39dd2c74),
	.w7(32'h3c1a4547),
	.w8(32'hbb1c1d8a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93632e),
	.w1(32'hb927330e),
	.w2(32'hbc4cc10e),
	.w3(32'hbc473096),
	.w4(32'h3bac4365),
	.w5(32'hbbc48144),
	.w6(32'hbbdd3f82),
	.w7(32'hbb208054),
	.w8(32'hbc29f6ec),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc75ae),
	.w1(32'hbbec38fa),
	.w2(32'hbbe27e84),
	.w3(32'hbca1dc6f),
	.w4(32'h3c0da4e2),
	.w5(32'h3d28b98c),
	.w6(32'hbc7bd65f),
	.w7(32'h3c93666e),
	.w8(32'h3a8ed31f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be435c1),
	.w1(32'hbbc45fe0),
	.w2(32'hb9f22cf9),
	.w3(32'hbbc49f4e),
	.w4(32'hbbc0e06c),
	.w5(32'hbb0001d6),
	.w6(32'h3d3ca19e),
	.w7(32'h37cef9d3),
	.w8(32'h3cb34b3c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b087b0a),
	.w1(32'hbaab3485),
	.w2(32'hbbab740f),
	.w3(32'hbc64154b),
	.w4(32'h3bda362e),
	.w5(32'hbad92729),
	.w6(32'hbc000ba4),
	.w7(32'hbc487b4e),
	.w8(32'hbb81189e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb499cfe),
	.w1(32'hbb92e17d),
	.w2(32'h3cd05087),
	.w3(32'hbc3c1388),
	.w4(32'h3c2709a3),
	.w5(32'hbb245568),
	.w6(32'hbb365b93),
	.w7(32'hbc45ebfb),
	.w8(32'hbbe7310b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd5d92),
	.w1(32'hbac17ac9),
	.w2(32'hbb5549eb),
	.w3(32'h3b15a08e),
	.w4(32'hbbfaa466),
	.w5(32'h3b933a3b),
	.w6(32'h3af282a9),
	.w7(32'hbbc3fb7f),
	.w8(32'h398d8a81),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f9543),
	.w1(32'hbc55a32b),
	.w2(32'hbc8f2d79),
	.w3(32'h3b03c133),
	.w4(32'hbc100d89),
	.w5(32'hbba0da31),
	.w6(32'hbb964814),
	.w7(32'h3c5e4f40),
	.w8(32'hbc449625),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7880e9),
	.w1(32'hbb32b8f3),
	.w2(32'hbc77c91e),
	.w3(32'hbbeddec9),
	.w4(32'hbbd04ccd),
	.w5(32'hbba6a2cf),
	.w6(32'hbcb333fc),
	.w7(32'h3c617df2),
	.w8(32'h3ba24e51),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90bc12),
	.w1(32'hbc02123c),
	.w2(32'hbc12782e),
	.w3(32'h3a89b44c),
	.w4(32'hbb0f4330),
	.w5(32'h3b567411),
	.w6(32'hbc31ac24),
	.w7(32'h3b8062db),
	.w8(32'h3a0fd58d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc825908),
	.w1(32'hbc9f6853),
	.w2(32'hbc0f85a3),
	.w3(32'hbbc3ea3c),
	.w4(32'hbb669435),
	.w5(32'h3bf68f41),
	.w6(32'hbc0403b4),
	.w7(32'h3c032817),
	.w8(32'h3bbc5d43),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb004da),
	.w1(32'hbbaad250),
	.w2(32'hbb795ff5),
	.w3(32'hbbe2cb77),
	.w4(32'h3a14fc7c),
	.w5(32'hbc24832a),
	.w6(32'hbc13f0dd),
	.w7(32'hbb9a9115),
	.w8(32'hbc27df40),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc046eb4),
	.w1(32'hbaebafa6),
	.w2(32'hbbcc5d7f),
	.w3(32'hbb5b550c),
	.w4(32'h3c49fc2f),
	.w5(32'hbb795346),
	.w6(32'hbbbe821e),
	.w7(32'h3b54fc87),
	.w8(32'h3bf58a42),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7d227),
	.w1(32'h3bc6ac33),
	.w2(32'hbc07b469),
	.w3(32'hba1ec39a),
	.w4(32'hbb800604),
	.w5(32'h3bfde7dc),
	.w6(32'h3bc61889),
	.w7(32'hbb659651),
	.w8(32'h3bd90a41),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac2616),
	.w1(32'hb9c61101),
	.w2(32'hbcc944e6),
	.w3(32'hbc5f7ee2),
	.w4(32'h3bec12dc),
	.w5(32'hbce94d8e),
	.w6(32'hba433fcf),
	.w7(32'hbbcabadd),
	.w8(32'hba8fbef2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba91871),
	.w1(32'h3d2fc744),
	.w2(32'hbb90ebe8),
	.w3(32'h3c3c664c),
	.w4(32'h394378b5),
	.w5(32'h3d03f097),
	.w6(32'h3c1d9fce),
	.w7(32'h3b960ad8),
	.w8(32'h3c9536ab),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbd5a0),
	.w1(32'hbb3fdbc4),
	.w2(32'hbbfb5841),
	.w3(32'h3bf749b1),
	.w4(32'h3b2455bd),
	.w5(32'hbb5aac12),
	.w6(32'hbd58e4f4),
	.w7(32'hbca716ce),
	.w8(32'h3b68b2bc),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc127bc2),
	.w1(32'hba8761b6),
	.w2(32'hbba9e257),
	.w3(32'hbb8caf08),
	.w4(32'h3c1f302c),
	.w5(32'hbb204394),
	.w6(32'hbc9ade0d),
	.w7(32'hbc377ec2),
	.w8(32'hbbb5983e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1dd90d),
	.w1(32'hbb4cf5e6),
	.w2(32'h3ab322ab),
	.w3(32'hbc235656),
	.w4(32'hbb2bf432),
	.w5(32'hbc2530b2),
	.w6(32'hbc673ab1),
	.w7(32'h3be0a28a),
	.w8(32'h3b2b2b43),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89b10b),
	.w1(32'h3ab90040),
	.w2(32'hbb4f0bb2),
	.w3(32'hbc38bb7c),
	.w4(32'hbbafb794),
	.w5(32'h3bd4fbd2),
	.w6(32'hbbbfcc1f),
	.w7(32'h3ba96322),
	.w8(32'h3bd7c257),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01f890),
	.w1(32'hbcf4beb1),
	.w2(32'hbb857b74),
	.w3(32'hbbc4c29e),
	.w4(32'h3c063049),
	.w5(32'hbb69c693),
	.w6(32'hbc816bf0),
	.w7(32'h3c4b25a6),
	.w8(32'hbb33c034),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce12237),
	.w1(32'h3bb01a63),
	.w2(32'hb94a6703),
	.w3(32'hbc2b1934),
	.w4(32'h3af02a9f),
	.w5(32'h3c1412c4),
	.w6(32'hbc0647c4),
	.w7(32'hbb3099e2),
	.w8(32'h3b27a1c6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98864a),
	.w1(32'h3adbe1fb),
	.w2(32'hbc232154),
	.w3(32'hbd0c0ae5),
	.w4(32'h3c2b0b60),
	.w5(32'h3b958c28),
	.w6(32'hbc875e01),
	.w7(32'h3bdea85f),
	.w8(32'hbc05ac82),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ca7f5),
	.w1(32'h3c79bf1e),
	.w2(32'h3bdc6b63),
	.w3(32'h3c642efa),
	.w4(32'hbc24bcde),
	.w5(32'h3a137bec),
	.w6(32'hbc4027c8),
	.w7(32'hbc466c7a),
	.w8(32'hbc40c1a7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b655eb6),
	.w1(32'hbb805a79),
	.w2(32'h39a96123),
	.w3(32'h3b81f9b8),
	.w4(32'hbbf6ba50),
	.w5(32'hbd547e0d),
	.w6(32'h3bdf4455),
	.w7(32'hbd5f9387),
	.w8(32'h39563e88),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37f60e),
	.w1(32'h3b8753a9),
	.w2(32'hbbb91ffb),
	.w3(32'hbd1c2f64),
	.w4(32'hbb1839a6),
	.w5(32'hbbf74b57),
	.w6(32'hbc879f05),
	.w7(32'h3b709c92),
	.w8(32'hbc09dc0b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b72ce),
	.w1(32'h3c54e3c5),
	.w2(32'hbc8d3472),
	.w3(32'hbbf05582),
	.w4(32'hbcf218c1),
	.w5(32'hbba9735a),
	.w6(32'hbc21ff75),
	.w7(32'h3d2989c4),
	.w8(32'hbc2c2019),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac73d2),
	.w1(32'hbb19e380),
	.w2(32'hbc6a3748),
	.w3(32'hbc872de0),
	.w4(32'hbba58a66),
	.w5(32'h3a9f5c39),
	.w6(32'hbc68a125),
	.w7(32'h3c0d5b26),
	.w8(32'h3c03b882),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d378c),
	.w1(32'h3b66ef8a),
	.w2(32'hbafd02a4),
	.w3(32'hbc0a7818),
	.w4(32'hbc10b5fa),
	.w5(32'hbbf66d57),
	.w6(32'hba978988),
	.w7(32'hba914112),
	.w8(32'hbac94063),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b817ba5),
	.w1(32'hb799cccc),
	.w2(32'h3b19da55),
	.w3(32'h3b4741df),
	.w4(32'hb598f214),
	.w5(32'h3c894c6f),
	.w6(32'hbbd965e5),
	.w7(32'h38d4753a),
	.w8(32'hba765555),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5897),
	.w1(32'h3c57034f),
	.w2(32'h3b191705),
	.w3(32'hbb986524),
	.w4(32'hba0ec0a0),
	.w5(32'hbb53bc5d),
	.w6(32'h3b15f50a),
	.w7(32'h3a900c23),
	.w8(32'h3b3660c7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba4d5d),
	.w1(32'hbbf4e0c1),
	.w2(32'hbc6a9a6b),
	.w3(32'h3c56f13e),
	.w4(32'h3b824c73),
	.w5(32'hbc5e6350),
	.w6(32'hbb591819),
	.w7(32'hbba499b6),
	.w8(32'h3b4dccf9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194e38),
	.w1(32'h3b28b159),
	.w2(32'hbcaaaf7a),
	.w3(32'h3bd4f511),
	.w4(32'hbc76948d),
	.w5(32'hbb9c3a80),
	.w6(32'hbbe45c59),
	.w7(32'hbb57cc6f),
	.w8(32'hbbbb44e0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af471b9),
	.w1(32'hbc1d4746),
	.w2(32'hbc0f6d11),
	.w3(32'hbad7d512),
	.w4(32'hbc30b566),
	.w5(32'hbc70e562),
	.w6(32'hbb97e623),
	.w7(32'hbbce1e1b),
	.w8(32'hbba652de),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5026e),
	.w1(32'hbc2d619c),
	.w2(32'h3ad7e9c2),
	.w3(32'hbb698943),
	.w4(32'hbbcdcab8),
	.w5(32'h3a3dd86d),
	.w6(32'hbaa7e9b8),
	.w7(32'h3bc092fb),
	.w8(32'hbc4168d0),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09c5e4),
	.w1(32'h3b382cb7),
	.w2(32'hbbc2d1c4),
	.w3(32'hbc7738e2),
	.w4(32'h3c1836d7),
	.w5(32'h3ca012b5),
	.w6(32'hbb644ec8),
	.w7(32'h3b9b496e),
	.w8(32'hba8bd626),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb72b76),
	.w1(32'hbb37dfa6),
	.w2(32'hbc019652),
	.w3(32'h3b52aced),
	.w4(32'h3b9ff50a),
	.w5(32'hba622538),
	.w6(32'hb8c00f58),
	.w7(32'h3c944335),
	.w8(32'hbbcff9ff),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b707ddd),
	.w1(32'h3bd90371),
	.w2(32'hbc01c3e9),
	.w3(32'h3af868f1),
	.w4(32'hbc3f6911),
	.w5(32'h3c0b47d0),
	.w6(32'hb99670ac),
	.w7(32'h3c4abb08),
	.w8(32'h3a1e04f1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb1d58),
	.w1(32'hbb4c5733),
	.w2(32'h3b3f6dc5),
	.w3(32'h3cbc61d2),
	.w4(32'hbbc8c627),
	.w5(32'h3b1434dd),
	.w6(32'hbcf4fa68),
	.w7(32'h3c252661),
	.w8(32'hbb1d241c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd072ce),
	.w1(32'hbbfa5f23),
	.w2(32'hbac2cf94),
	.w3(32'hbaf1e251),
	.w4(32'h3c0ab179),
	.w5(32'h3bf686f8),
	.w6(32'hbc284a64),
	.w7(32'hbbbccdad),
	.w8(32'h3b328571),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0059f),
	.w1(32'hbbdf470a),
	.w2(32'hbad40adf),
	.w3(32'hbb4826bb),
	.w4(32'h3c0bf9b5),
	.w5(32'hbca5e6b9),
	.w6(32'h3c2238a6),
	.w7(32'hbb70fe0d),
	.w8(32'h3d13ed26),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4155eb),
	.w1(32'hbba37469),
	.w2(32'hbc8f24e3),
	.w3(32'hbc503556),
	.w4(32'hbb9f4090),
	.w5(32'h3d33f92f),
	.w6(32'hba9420d7),
	.w7(32'h3b143bdf),
	.w8(32'hbc1ffbef),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc887bbb),
	.w1(32'hbba2cb8c),
	.w2(32'h3ac1307d),
	.w3(32'hbbe0356d),
	.w4(32'hbb4a952a),
	.w5(32'h3b3fb01e),
	.w6(32'hbbfd6360),
	.w7(32'hbc80e03d),
	.w8(32'hbc9e3890),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08714f),
	.w1(32'h39904849),
	.w2(32'h3aa37c4f),
	.w3(32'hbbbca1d6),
	.w4(32'hbc2d06e4),
	.w5(32'hbbf64542),
	.w6(32'hbbc738cf),
	.w7(32'h3ab04480),
	.w8(32'h3aa0fb8c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01eb1d),
	.w1(32'hba70248e),
	.w2(32'hbc8e2f62),
	.w3(32'hb9470500),
	.w4(32'h398fef5b),
	.w5(32'hbc9035f4),
	.w6(32'hbc56a67e),
	.w7(32'h3c51147a),
	.w8(32'h3bf6e56a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bba79),
	.w1(32'hbc04b03b),
	.w2(32'hba0e4616),
	.w3(32'hbbb7f4bc),
	.w4(32'h3b9d9fae),
	.w5(32'hbc96c6f3),
	.w6(32'hbbd7807f),
	.w7(32'hbb62e1c2),
	.w8(32'hbb3351b0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7209b),
	.w1(32'h3a930273),
	.w2(32'hbb56b0bb),
	.w3(32'h3b16e1d3),
	.w4(32'hbc2a3f5d),
	.w5(32'hbc40512f),
	.w6(32'h3b59c6c3),
	.w7(32'hbb4f12a8),
	.w8(32'hbb8008d4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadadcf5),
	.w1(32'hbbaa7842),
	.w2(32'hbd19e9df),
	.w3(32'hbba50abd),
	.w4(32'hbba31b7a),
	.w5(32'hbba77554),
	.w6(32'h3bb092ac),
	.w7(32'hbae449b3),
	.w8(32'hbbb736b5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5124c2),
	.w1(32'h3d064f2f),
	.w2(32'h3bd43627),
	.w3(32'h3b7454df),
	.w4(32'h3c248095),
	.w5(32'hbc5df5f5),
	.w6(32'hbb6c189d),
	.w7(32'hbbc361d7),
	.w8(32'h3b8cc861),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bada708),
	.w1(32'hbb933182),
	.w2(32'hbafc5901),
	.w3(32'h395e1dd9),
	.w4(32'hbbb47be4),
	.w5(32'h3b0d83fc),
	.w6(32'h3c22a82b),
	.w7(32'hbc5d0b74),
	.w8(32'h3ce05ca2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b0d58),
	.w1(32'hbbbd1fd3),
	.w2(32'h3bd11ddb),
	.w3(32'hbc049e99),
	.w4(32'h3a2a41cc),
	.w5(32'h3cd46b00),
	.w6(32'h3cfc276d),
	.w7(32'h3c6bc595),
	.w8(32'hba274c81),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe1b55),
	.w1(32'hba93ca44),
	.w2(32'h3bf8b7e9),
	.w3(32'h3c16d046),
	.w4(32'hbb87cc52),
	.w5(32'h3c3e6dc4),
	.w6(32'h3b86f6b3),
	.w7(32'hbbf90a86),
	.w8(32'hb657f98f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b1a3c),
	.w1(32'h3bb57fc8),
	.w2(32'h3a0482d5),
	.w3(32'h3b325975),
	.w4(32'hbac687c3),
	.w5(32'h3a3e6a68),
	.w6(32'hbbe29d18),
	.w7(32'h3c08daa8),
	.w8(32'hbbeeddd4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca7679),
	.w1(32'h3b0ed3e9),
	.w2(32'hbca13892),
	.w3(32'hbbf40641),
	.w4(32'h3ab4d660),
	.w5(32'hbc8a9d54),
	.w6(32'hbb5e1b33),
	.w7(32'hbc4911c7),
	.w8(32'hbc3f0d92),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17efa1),
	.w1(32'h3cb38fe4),
	.w2(32'hbbc62216),
	.w3(32'hbc2c1944),
	.w4(32'hbb14e81d),
	.w5(32'h3d1e0ad0),
	.w6(32'hbc1f32d7),
	.w7(32'hbab48936),
	.w8(32'hbc024f42),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc855499),
	.w1(32'hbb82bce1),
	.w2(32'hbc6e1e92),
	.w3(32'h3bf717ed),
	.w4(32'hbaa1602d),
	.w5(32'hbbb9782a),
	.w6(32'hbc712dc3),
	.w7(32'hbc5ea95b),
	.w8(32'hbc39e559),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a651206),
	.w1(32'hbae75caa),
	.w2(32'hbb733284),
	.w3(32'hbb07d5fe),
	.w4(32'hbb38859d),
	.w5(32'hbc0bed68),
	.w6(32'h3b02b427),
	.w7(32'hbb8f31be),
	.w8(32'hbade7275),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd36b25),
	.w1(32'hbacd513c),
	.w2(32'hbc5e87c9),
	.w3(32'h3bdcf4b9),
	.w4(32'hbcf0299b),
	.w5(32'h3bc0d6af),
	.w6(32'hbb662001),
	.w7(32'hbb505def),
	.w8(32'h3cbfa2ea),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360e07eb),
	.w1(32'hbbbc41ef),
	.w2(32'h3ba5137b),
	.w3(32'h39ab0528),
	.w4(32'h35a539e6),
	.w5(32'hba9ea3cc),
	.w6(32'hbbbc1f0d),
	.w7(32'hbb38ed45),
	.w8(32'hbd79348b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc015cab),
	.w1(32'h3b6adf02),
	.w2(32'hbaf763e5),
	.w3(32'hbc8b7569),
	.w4(32'hbc5128e8),
	.w5(32'h3ba4010e),
	.w6(32'hbb292f4c),
	.w7(32'hbb607147),
	.w8(32'h3c82bdd9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98f570),
	.w1(32'h3a845eca),
	.w2(32'hbb8d53d7),
	.w3(32'hbb1153f6),
	.w4(32'hba9c3908),
	.w5(32'h3b9b0496),
	.w6(32'hbc1d0194),
	.w7(32'h3a4e1948),
	.w8(32'hbc14ec67),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21598d),
	.w1(32'hbba69c2d),
	.w2(32'hbaa7831d),
	.w3(32'h3b3c8244),
	.w4(32'hbc868a9d),
	.w5(32'hbb0eadaa),
	.w6(32'hbaed45f9),
	.w7(32'h39984782),
	.w8(32'hbb0f5368),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a9e88),
	.w1(32'h3b852185),
	.w2(32'h3920c626),
	.w3(32'hbbe026d5),
	.w4(32'h3bb31107),
	.w5(32'hbc3c36eb),
	.w6(32'hbcc36113),
	.w7(32'h3b6939fb),
	.w8(32'hbc0340c0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9494cf),
	.w1(32'hbc13f02b),
	.w2(32'hbbd5725e),
	.w3(32'hbb9968b4),
	.w4(32'h3bb2952a),
	.w5(32'h3a23da79),
	.w6(32'h3accbcfb),
	.w7(32'h3b6a35f4),
	.w8(32'hb916dc70),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a277541),
	.w1(32'hbcb65396),
	.w2(32'h3bec1e88),
	.w3(32'hbb949881),
	.w4(32'hbb06835e),
	.w5(32'hbbc92cf6),
	.w6(32'h3ce49239),
	.w7(32'hbc1fa4f1),
	.w8(32'h3c58f2d8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e5c9e),
	.w1(32'h3a5dd722),
	.w2(32'hbc37c959),
	.w3(32'hbbe8cb6a),
	.w4(32'hbaa65394),
	.w5(32'hbb093ebb),
	.w6(32'hbb136f5f),
	.w7(32'hbb75ce6b),
	.w8(32'hbc6f28bb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f6a22),
	.w1(32'hbb945a88),
	.w2(32'h3b34c0e0),
	.w3(32'hbb733bb2),
	.w4(32'hbd0a7aa3),
	.w5(32'hbb2f33f6),
	.w6(32'hbbd42add),
	.w7(32'hbb48f0d2),
	.w8(32'h3a9fc155),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ea8db),
	.w1(32'hbc53a302),
	.w2(32'hbc48dae8),
	.w3(32'hbc6af344),
	.w4(32'hbc13f6f5),
	.w5(32'hbb82f527),
	.w6(32'hbc0fb871),
	.w7(32'hbbbceda4),
	.w8(32'h3a94a35c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb384257),
	.w1(32'h3b050022),
	.w2(32'hbc59e4c7),
	.w3(32'hbb4a3508),
	.w4(32'hba81ab4f),
	.w5(32'h3a47428f),
	.w6(32'h3c9e7bcb),
	.w7(32'hbba0b6f1),
	.w8(32'hbcb07940),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39437784),
	.w1(32'h3d0b51d3),
	.w2(32'h3c25909a),
	.w3(32'hbb921707),
	.w4(32'h3b50d074),
	.w5(32'h3be0b448),
	.w6(32'hbd302c65),
	.w7(32'h3b91c796),
	.w8(32'h3ac5dc12),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule