module layer_10_featuremap_342(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb889269),
	.w1(32'hbc09d5c7),
	.w2(32'hbba8ba67),
	.w3(32'hbaa983d2),
	.w4(32'hbb8623cd),
	.w5(32'h3b170afd),
	.w6(32'hbbc3ab6f),
	.w7(32'hbaf2d6a5),
	.w8(32'h3b970a68),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d9122),
	.w1(32'h3c010679),
	.w2(32'h3bb5d073),
	.w3(32'h3bcf2920),
	.w4(32'hbb621970),
	.w5(32'h3b5de8f1),
	.w6(32'h3c4e8529),
	.w7(32'h38034bb3),
	.w8(32'h3b2abd01),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c546b37),
	.w1(32'h3c4d6bf6),
	.w2(32'h3b696309),
	.w3(32'h3b22fcc7),
	.w4(32'h3b9d7083),
	.w5(32'hbb02867c),
	.w6(32'h3b8ee253),
	.w7(32'h3ca7901e),
	.w8(32'hbb82c784),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb627ae7),
	.w1(32'hba758586),
	.w2(32'h3992c4cb),
	.w3(32'hbacbff42),
	.w4(32'hbbd6b99a),
	.w5(32'h3a9cd763),
	.w6(32'h3c4be660),
	.w7(32'hbabbf186),
	.w8(32'hbc013d11),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a509),
	.w1(32'h3a259d9d),
	.w2(32'h3b93b842),
	.w3(32'hbb2232bd),
	.w4(32'h3be02cbd),
	.w5(32'hb98c0bea),
	.w6(32'h3c1b94b0),
	.w7(32'h3acc8045),
	.w8(32'hb9ac3bff),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d954f),
	.w1(32'hbb2c08c6),
	.w2(32'hbaa536c5),
	.w3(32'h3ac644c5),
	.w4(32'h3a8c2f94),
	.w5(32'hbb215f78),
	.w6(32'h3c8b6b7d),
	.w7(32'h3c08a3f1),
	.w8(32'h3a0f5ac7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e88ed),
	.w1(32'hbb0958c1),
	.w2(32'hbb85f044),
	.w3(32'h3a84fd88),
	.w4(32'hbbd2930a),
	.w5(32'hbbffb7f4),
	.w6(32'h3c66b0f7),
	.w7(32'h3afc5cc3),
	.w8(32'hbb837429),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc563104),
	.w1(32'hbc537f56),
	.w2(32'hbc1348ec),
	.w3(32'hbb885e08),
	.w4(32'hbbd5b60d),
	.w5(32'hbbacd96d),
	.w6(32'hba2608a4),
	.w7(32'hbb00c8f2),
	.w8(32'hbc054839),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f4434),
	.w1(32'hbba31c34),
	.w2(32'hbb08700b),
	.w3(32'hbb7c7bdb),
	.w4(32'hbba1bf60),
	.w5(32'hb92bbf5d),
	.w6(32'hbb487843),
	.w7(32'hbaaf2f92),
	.w8(32'hba8441cc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc446858),
	.w1(32'hbbe318df),
	.w2(32'hbb8a6d2b),
	.w3(32'hbaf09829),
	.w4(32'hbb1c177c),
	.w5(32'hbaad7df9),
	.w6(32'h3c3a6a10),
	.w7(32'h3b793148),
	.w8(32'hb902401c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba936c),
	.w1(32'hba3bf546),
	.w2(32'hbb480eca),
	.w3(32'h3b53c76a),
	.w4(32'hba943431),
	.w5(32'h3b06c156),
	.w6(32'h3d03d715),
	.w7(32'h3b695a05),
	.w8(32'h3b95f2ec),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066064),
	.w1(32'h3c1b28f1),
	.w2(32'hbb015662),
	.w3(32'h3b77e96e),
	.w4(32'h3c0ac203),
	.w5(32'hbad93205),
	.w6(32'hbc271c4b),
	.w7(32'h3c5ed95f),
	.w8(32'hbb9f0bf4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ed99e),
	.w1(32'hbc24d0e9),
	.w2(32'h3b0d0b03),
	.w3(32'hbc40f7c0),
	.w4(32'hbc3c320b),
	.w5(32'hbb3f7c3d),
	.w6(32'hbbf3f57a),
	.w7(32'hbb8b00b4),
	.w8(32'hbc344cb4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b9f23),
	.w1(32'h3b580bdb),
	.w2(32'h3aa3d7d3),
	.w3(32'h3b89c766),
	.w4(32'hbbc9a793),
	.w5(32'h39528251),
	.w6(32'h3c3b807b),
	.w7(32'h3b32412c),
	.w8(32'h3baa82b5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8834a6),
	.w1(32'hbb125b60),
	.w2(32'hbb387ab2),
	.w3(32'h3be40928),
	.w4(32'hbb2e145c),
	.w5(32'hbbe9874f),
	.w6(32'h3c8e97dc),
	.w7(32'h3c2ba3bf),
	.w8(32'hbc105394),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02c5a2),
	.w1(32'hbb77aad3),
	.w2(32'hbb68979b),
	.w3(32'hbb6a2814),
	.w4(32'hbac6c5ea),
	.w5(32'hbb763e41),
	.w6(32'h3bf05b95),
	.w7(32'hbb249953),
	.w8(32'hbbdc71d9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a8afb),
	.w1(32'hbbfcaca2),
	.w2(32'hbbcda199),
	.w3(32'h3a8ffb81),
	.w4(32'hbaf09073),
	.w5(32'hbb6856dd),
	.w6(32'h3b42b67e),
	.w7(32'h3a4395ee),
	.w8(32'hba6f1982),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e401c),
	.w1(32'hbbe3012d),
	.w2(32'hbc0356c8),
	.w3(32'hbbbddc0d),
	.w4(32'hbc38c2ba),
	.w5(32'hbc0a49bd),
	.w6(32'hbbe364b8),
	.w7(32'hbbf35dbf),
	.w8(32'h3c5c40f3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99bd57),
	.w1(32'hbc05c2bc),
	.w2(32'h3a71e4bc),
	.w3(32'h3b89780e),
	.w4(32'hba0ad43d),
	.w5(32'h3a13a871),
	.w6(32'h3c34d8c7),
	.w7(32'h3c59f0d9),
	.w8(32'hbab0c081),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad80795),
	.w1(32'h3bbce122),
	.w2(32'h3b654526),
	.w3(32'h3b510ba7),
	.w4(32'h3b063618),
	.w5(32'hbb2cc896),
	.w6(32'h3b4ac7b8),
	.w7(32'h3b86f266),
	.w8(32'hbba525b8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a8f61),
	.w1(32'hbab6f1e4),
	.w2(32'hbab52870),
	.w3(32'hba0ce0f5),
	.w4(32'hbbd4f01e),
	.w5(32'h3b0ff324),
	.w6(32'h3ba46c6b),
	.w7(32'hbb0a6cf9),
	.w8(32'hbb181f67),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10e825),
	.w1(32'hbba1e3e7),
	.w2(32'h3aacf795),
	.w3(32'hbc1883ff),
	.w4(32'hbbd45a51),
	.w5(32'h3acca236),
	.w6(32'hbb8c0e58),
	.w7(32'hbaa8cb23),
	.w8(32'h3c0c4d28),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b651730),
	.w1(32'h3b05ebff),
	.w2(32'h3b9dbc3b),
	.w3(32'h3a84637d),
	.w4(32'h3c02bc21),
	.w5(32'hbbe2bf96),
	.w6(32'hbace324c),
	.w7(32'h3c18379c),
	.w8(32'hbb89ce2a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba18550),
	.w1(32'hbb1c450d),
	.w2(32'hbb8a8b86),
	.w3(32'h3bcc431d),
	.w4(32'hbc23fcb7),
	.w5(32'hbc17644d),
	.w6(32'h3c9be770),
	.w7(32'hbc1b070e),
	.w8(32'hbada886e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe27d4e),
	.w1(32'h38f4ac77),
	.w2(32'h3aeffc60),
	.w3(32'hbbbfdb33),
	.w4(32'hbb585d5e),
	.w5(32'h3be55663),
	.w6(32'hbbece033),
	.w7(32'hbb0a0831),
	.w8(32'h3c05b3bc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb122fa3),
	.w1(32'h3a00f888),
	.w2(32'h3b6d8d4c),
	.w3(32'h3c43bb77),
	.w4(32'h3aa061a8),
	.w5(32'h3b0f83a5),
	.w6(32'h3c873cb3),
	.w7(32'h3c0c5aaf),
	.w8(32'h3ad75ad7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8753a5),
	.w1(32'hbb9c95b4),
	.w2(32'hbb4e433f),
	.w3(32'hb98b40f5),
	.w4(32'hba88106f),
	.w5(32'hbb98ad9e),
	.w6(32'h3c01d2bd),
	.w7(32'h3bb200f0),
	.w8(32'hbc1c0611),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17927f),
	.w1(32'hbc428e23),
	.w2(32'hbbdb50dd),
	.w3(32'hbc07d835),
	.w4(32'hbbab782a),
	.w5(32'h3b3910ee),
	.w6(32'hbc5e034a),
	.w7(32'hbb716a2b),
	.w8(32'h39c9e71f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb370d01),
	.w1(32'hbb9464c2),
	.w2(32'hbae0cbe6),
	.w3(32'h3acaeed6),
	.w4(32'hbc0829d2),
	.w5(32'hbb258003),
	.w6(32'h3bb4ad24),
	.w7(32'hbb359fd0),
	.w8(32'hbc1290d4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda23e0),
	.w1(32'hbb3e174f),
	.w2(32'hbbb5e204),
	.w3(32'hbb706639),
	.w4(32'hbbb781eb),
	.w5(32'hbc580b07),
	.w6(32'hbbbc0dfa),
	.w7(32'hbb8684d9),
	.w8(32'hbbb2952f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b940dc6),
	.w1(32'hb82a1400),
	.w2(32'hba98ccb1),
	.w3(32'h3ac7af13),
	.w4(32'hbb0b1e4e),
	.w5(32'hb778d087),
	.w6(32'hbc1566a8),
	.w7(32'hbbbf9722),
	.w8(32'h3c00ffd2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8adfa),
	.w1(32'h3c4d937d),
	.w2(32'h3bc9e478),
	.w3(32'hbb56210e),
	.w4(32'h3a501aef),
	.w5(32'hbb60d114),
	.w6(32'hbc39994b),
	.w7(32'hbbcabe88),
	.w8(32'h3ca9a2e0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc43172),
	.w1(32'hbbe43893),
	.w2(32'h3ba8b629),
	.w3(32'h3cbcdbe2),
	.w4(32'h3c30ce28),
	.w5(32'hbaffca41),
	.w6(32'hbc464321),
	.w7(32'h3a842831),
	.w8(32'h3b8647ff),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb774aef),
	.w1(32'h3bbce6fa),
	.w2(32'hb9bd0426),
	.w3(32'h3bcf9aaa),
	.w4(32'hbb8fdc6d),
	.w5(32'h3aea9309),
	.w6(32'h3ae77432),
	.w7(32'h3b66f0bb),
	.w8(32'h3b741280),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7bb54),
	.w1(32'hbaf01c2d),
	.w2(32'hb9816008),
	.w3(32'h3a982143),
	.w4(32'h3bb88d07),
	.w5(32'h3bd0c1df),
	.w6(32'h3aa4d7e3),
	.w7(32'h3b9e46d3),
	.w8(32'h3a3f6629),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd10347),
	.w1(32'hbb61f740),
	.w2(32'hbbae493b),
	.w3(32'h3b394c0d),
	.w4(32'hb9d23828),
	.w5(32'h3c16c1b0),
	.w6(32'h399670e1),
	.w7(32'h3a62f860),
	.w8(32'h39b44694),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83862a),
	.w1(32'h3be7d200),
	.w2(32'h3b7e00b2),
	.w3(32'h3c847b2b),
	.w4(32'h3be56613),
	.w5(32'hb8952c55),
	.w6(32'hbcb35152),
	.w7(32'hbbad8f6c),
	.w8(32'h3aa4b8d0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb983220),
	.w1(32'hbb0fe4cb),
	.w2(32'h3b0b3783),
	.w3(32'hbbb2e083),
	.w4(32'h3a567708),
	.w5(32'h3b5ca303),
	.w6(32'h3cb51de9),
	.w7(32'h3c6a5287),
	.w8(32'hbabb7d2b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdfb4b),
	.w1(32'hbb92efe1),
	.w2(32'h3b72e5c3),
	.w3(32'hbbbeab4b),
	.w4(32'hbbbfc221),
	.w5(32'h3c04b3b7),
	.w6(32'h3aeb3ce7),
	.w7(32'h3a9ab81d),
	.w8(32'h3ac0550b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7b701),
	.w1(32'hbbe7706f),
	.w2(32'h3b6e116f),
	.w3(32'hbbfd1d38),
	.w4(32'h3a023914),
	.w5(32'hbb28d715),
	.w6(32'hbbb4d3e7),
	.w7(32'h3acc814c),
	.w8(32'hbb2bb576),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadff1de),
	.w1(32'hbc1eed87),
	.w2(32'hbb6b3a52),
	.w3(32'hbc0fc331),
	.w4(32'hbc045cab),
	.w5(32'h3bc08342),
	.w6(32'hbc61e886),
	.w7(32'hbb67b0a6),
	.w8(32'h3b6ee368),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993826),
	.w1(32'h3b542e12),
	.w2(32'h3b670ba5),
	.w3(32'h3bfae8ad),
	.w4(32'h3a8a23dd),
	.w5(32'hbc1527d8),
	.w6(32'h3c85ad1e),
	.w7(32'h3c409e93),
	.w8(32'hbbbf7293),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4363c7),
	.w1(32'hbbc8ce85),
	.w2(32'hbbaaa6f6),
	.w3(32'hbc116847),
	.w4(32'hbc0e6346),
	.w5(32'hbba79b7a),
	.w6(32'h3c121b12),
	.w7(32'h3b559274),
	.w8(32'hbba6e8f3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc361103),
	.w1(32'hbc9ece70),
	.w2(32'hbc314940),
	.w3(32'h3baecc36),
	.w4(32'hbbd2a843),
	.w5(32'hbb331283),
	.w6(32'h3d283d89),
	.w7(32'hbb9f822b),
	.w8(32'h3b9fcd18),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393aa7bd),
	.w1(32'hbb4d10da),
	.w2(32'hbb20979c),
	.w3(32'h3bdb07a8),
	.w4(32'h3b9c7eb2),
	.w5(32'hbb75ab5a),
	.w6(32'h3c01b89b),
	.w7(32'h3bc4d62c),
	.w8(32'hbb921884),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08f205),
	.w1(32'hbc0872fd),
	.w2(32'hbc33cd23),
	.w3(32'hbbe96a0b),
	.w4(32'hbc2e1cb5),
	.w5(32'hbbbccb28),
	.w6(32'hbbb6873b),
	.w7(32'hbc0ec69b),
	.w8(32'h3a8886ef),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be2c93),
	.w1(32'h3a1f2ba4),
	.w2(32'hbbb1d21a),
	.w3(32'h3b1c2207),
	.w4(32'hbb1cb155),
	.w5(32'h3ba756d2),
	.w6(32'h3b49852a),
	.w7(32'hba8de339),
	.w8(32'h3b8afc37),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f0b9b),
	.w1(32'h3a5276d6),
	.w2(32'h3ba0dfd0),
	.w3(32'hbbb8f37f),
	.w4(32'hbaab43f2),
	.w5(32'h3a707c7d),
	.w6(32'hbc2770d6),
	.w7(32'hbb9266d3),
	.w8(32'h3b860f28),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e69ccc),
	.w1(32'h3adb865a),
	.w2(32'hbb100a07),
	.w3(32'hbaaba9ef),
	.w4(32'hbbfe483e),
	.w5(32'h3badff95),
	.w6(32'h3ba85508),
	.w7(32'hbb8865e1),
	.w8(32'h3ab0f9a5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b560450),
	.w1(32'hbb2fee68),
	.w2(32'h3a94c016),
	.w3(32'hbb780662),
	.w4(32'hbb3dbf87),
	.w5(32'h3a7f8948),
	.w6(32'hbab5523b),
	.w7(32'h3aba099b),
	.w8(32'hbb86e4bf),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac811c1),
	.w1(32'h3b0c7362),
	.w2(32'h3a591318),
	.w3(32'hbb86cfd0),
	.w4(32'h3a702d20),
	.w5(32'hbb87eb35),
	.w6(32'h3b09f034),
	.w7(32'hbbd3922c),
	.w8(32'h3bf1d79c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c77b7),
	.w1(32'hbbf2d9f3),
	.w2(32'hbb69c334),
	.w3(32'hbb9bc6de),
	.w4(32'hbbec86e2),
	.w5(32'h3b06c668),
	.w6(32'h3c78c061),
	.w7(32'h3c1e90d8),
	.w8(32'hbb2948d0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b916153),
	.w1(32'h3ba6732a),
	.w2(32'h3b459aa2),
	.w3(32'h3bca4c95),
	.w4(32'h3b6d4879),
	.w5(32'h3b8f54fe),
	.w6(32'h3c93f7f6),
	.w7(32'h3b8ba84d),
	.w8(32'h3c84c110),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840920),
	.w1(32'hba37a506),
	.w2(32'h3a541a9b),
	.w3(32'hbbf51a02),
	.w4(32'h3b8629b0),
	.w5(32'hbc01e735),
	.w6(32'hbc1a55fb),
	.w7(32'h3c79982b),
	.w8(32'hba2ed8de),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ea5cc),
	.w1(32'h3c088e66),
	.w2(32'hbb005251),
	.w3(32'hbad4cfbf),
	.w4(32'h3aec75cc),
	.w5(32'h3bdc0b25),
	.w6(32'hbb796b83),
	.w7(32'hbaf99481),
	.w8(32'h3bbc1b9d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d90b6),
	.w1(32'h3c1a81b4),
	.w2(32'h3b874d3d),
	.w3(32'h3b548a9e),
	.w4(32'hb7361a78),
	.w5(32'hbb786f30),
	.w6(32'h3c92e031),
	.w7(32'hba217394),
	.w8(32'hba544d50),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f3da1),
	.w1(32'hbb89900b),
	.w2(32'hbb9518b8),
	.w3(32'hbbc7f8c6),
	.w4(32'hbb78130f),
	.w5(32'h3aa190fb),
	.w6(32'hbc1375e7),
	.w7(32'hbb6878a1),
	.w8(32'hbc06b541),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d65fc9),
	.w1(32'h3b8f0ed0),
	.w2(32'hbb624a3d),
	.w3(32'hb9b90b5f),
	.w4(32'h3ab04fbe),
	.w5(32'hb8979796),
	.w6(32'h3bc80616),
	.w7(32'h3b833dce),
	.w8(32'hbadba70f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba359847),
	.w1(32'hbb86ff74),
	.w2(32'hbaac7d4c),
	.w3(32'hbb5aeabf),
	.w4(32'hbba5bb0c),
	.w5(32'h3b412eba),
	.w6(32'hbb9e4a55),
	.w7(32'h3ab7292d),
	.w8(32'hb986b930),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f50ab8),
	.w1(32'hbbf212c7),
	.w2(32'h3aedd70f),
	.w3(32'hbc04eb3f),
	.w4(32'hbbc3103b),
	.w5(32'hba10af5d),
	.w6(32'hb99ea4d0),
	.w7(32'h3af8f803),
	.w8(32'hb9ba403b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4a8c8),
	.w1(32'hbbc74bcd),
	.w2(32'h39872d4b),
	.w3(32'hbb3fc7be),
	.w4(32'hbb9cae76),
	.w5(32'h3b27a812),
	.w6(32'h3ae15a97),
	.w7(32'h39599693),
	.w8(32'h3b2d82fd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9ccae),
	.w1(32'hbbc585d0),
	.w2(32'hbb998e7c),
	.w3(32'h3ae905f0),
	.w4(32'hbc011dca),
	.w5(32'hbb1991dc),
	.w6(32'h3c8c4b66),
	.w7(32'hba2883a2),
	.w8(32'h3a88f80b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7dbdeb),
	.w1(32'hbb9f0cc6),
	.w2(32'hbba068fd),
	.w3(32'hbb984130),
	.w4(32'h3bc77f1d),
	.w5(32'hbabfd8cc),
	.w6(32'hbb9de479),
	.w7(32'hbb16107d),
	.w8(32'h3b13fb1a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae01690),
	.w1(32'h38f8f808),
	.w2(32'hbb6ac399),
	.w3(32'hba80b138),
	.w4(32'h3bb2b488),
	.w5(32'h396c9440),
	.w6(32'h39fd297a),
	.w7(32'h3bdc80b9),
	.w8(32'hbb6ece9c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fd64c),
	.w1(32'h3c111a6c),
	.w2(32'hbaa4230d),
	.w3(32'h3a71066c),
	.w4(32'h3b7103b4),
	.w5(32'h3bedd010),
	.w6(32'h3b36ef9d),
	.w7(32'h3b99c47c),
	.w8(32'h3be3b02c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959958b),
	.w1(32'hbb992402),
	.w2(32'hb9d85e6a),
	.w3(32'h394aed0d),
	.w4(32'hb9e3a8fe),
	.w5(32'h3b651b92),
	.w6(32'h3bbe619e),
	.w7(32'h3acb969b),
	.w8(32'h3ab31155),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfa15e),
	.w1(32'hbb6f8aa8),
	.w2(32'hbb8ae34e),
	.w3(32'h3b6b7b5c),
	.w4(32'h3b31a02f),
	.w5(32'h3af44fd9),
	.w6(32'h3c2337d6),
	.w7(32'h3c0b0584),
	.w8(32'h3b2aaf9b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5793a),
	.w1(32'h39e1ba39),
	.w2(32'hbb22fc93),
	.w3(32'h3b952939),
	.w4(32'hba7a9d3d),
	.w5(32'hbb2b0cc3),
	.w6(32'h3c96620e),
	.w7(32'h3b14d2eb),
	.w8(32'h3c4c9d63),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58ffee),
	.w1(32'h3bf7c292),
	.w2(32'h3b9d7772),
	.w3(32'h3bafc07c),
	.w4(32'h3ba7764a),
	.w5(32'h3a7a69f0),
	.w6(32'h3b8ea8c5),
	.w7(32'h3c884672),
	.w8(32'h3c558208),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab87ab8),
	.w1(32'hbb53fd9e),
	.w2(32'hbafb6da2),
	.w3(32'h3b94bdaf),
	.w4(32'hb9aedd95),
	.w5(32'h3bbf9875),
	.w6(32'h397f24c4),
	.w7(32'h3bb6216b),
	.w8(32'h3bbd289c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b451c03),
	.w1(32'h3c0be184),
	.w2(32'h3c0f6828),
	.w3(32'h3c2c80b5),
	.w4(32'h3bb495fb),
	.w5(32'h3aa0da71),
	.w6(32'h39a1131e),
	.w7(32'h3c2d02e8),
	.w8(32'hbb0b7243),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a8b82),
	.w1(32'h3bd4d6e9),
	.w2(32'hbbaad432),
	.w3(32'h39e96a8d),
	.w4(32'h3b1759a7),
	.w5(32'hbac884dd),
	.w6(32'h3c1cc484),
	.w7(32'h3ade9aae),
	.w8(32'hba590504),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98637e),
	.w1(32'hbb9f3f13),
	.w2(32'hbbd36b1a),
	.w3(32'hbb8fe7c2),
	.w4(32'hbbb3bfcb),
	.w5(32'hbad8bfcd),
	.w6(32'h3c15e659),
	.w7(32'h3bc5dbfc),
	.w8(32'hbb67afb0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f6140),
	.w1(32'hbaa47486),
	.w2(32'h3b80b11d),
	.w3(32'h3bf70cbc),
	.w4(32'hb9325ee9),
	.w5(32'h3af1f172),
	.w6(32'hbb964600),
	.w7(32'h3c053880),
	.w8(32'hba0363f1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bac8b0),
	.w1(32'hbb07f235),
	.w2(32'hbbca6abb),
	.w3(32'h3b5f8e7f),
	.w4(32'hbb00151e),
	.w5(32'hbb825e96),
	.w6(32'h3c35a36b),
	.w7(32'h3b9cfbc5),
	.w8(32'hbb043807),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff3379),
	.w1(32'hba96d025),
	.w2(32'hba92639b),
	.w3(32'hbbd891bf),
	.w4(32'hbbc64b20),
	.w5(32'h3a99dfa5),
	.w6(32'hbb84769c),
	.w7(32'hbb765fed),
	.w8(32'h3b1aa217),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb180f),
	.w1(32'hbb41ba4f),
	.w2(32'h3a863949),
	.w3(32'hbb826705),
	.w4(32'hbb5b37a6),
	.w5(32'hba4e2b4b),
	.w6(32'h3b140503),
	.w7(32'hb96b70bb),
	.w8(32'hbb2f635f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc340991),
	.w1(32'hbc073743),
	.w2(32'hbbb9c2be),
	.w3(32'h3b077904),
	.w4(32'h3aa275b8),
	.w5(32'h39a43919),
	.w6(32'h3be87860),
	.w7(32'hbb25977b),
	.w8(32'h3ad4e13d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16eeca),
	.w1(32'h38a097ee),
	.w2(32'hbaea65aa),
	.w3(32'h3aece0cc),
	.w4(32'h3b2422e7),
	.w5(32'hbb93dfd0),
	.w6(32'h3bf4f9a6),
	.w7(32'h3bc1109e),
	.w8(32'hbb4b3b04),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf61ac),
	.w1(32'hbc2bb2b1),
	.w2(32'hbc0ee8f1),
	.w3(32'hbbe176f9),
	.w4(32'hbbfb787c),
	.w5(32'h3b659995),
	.w6(32'h3becee32),
	.w7(32'h39a78138),
	.w8(32'h3b80bac7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1672d1),
	.w1(32'h3c023d29),
	.w2(32'h3c57f4ef),
	.w3(32'hbaae1576),
	.w4(32'h3b069266),
	.w5(32'hbbcd7d4e),
	.w6(32'h3b5c3e7c),
	.w7(32'h3c01b538),
	.w8(32'hba64d12f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc431d75),
	.w1(32'hbbffe83e),
	.w2(32'hbb9cbb83),
	.w3(32'hbba7a90d),
	.w4(32'hbb719e98),
	.w5(32'hbacc1e79),
	.w6(32'hbc0a0af2),
	.w7(32'hbac9022a),
	.w8(32'h3aa1335b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa60a02),
	.w1(32'hba9830be),
	.w2(32'hb8f6c168),
	.w3(32'h3b0101f4),
	.w4(32'h3acb1f2e),
	.w5(32'h3ba2f5d5),
	.w6(32'h3c1bea36),
	.w7(32'hbb0f859d),
	.w8(32'h3bb98daf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc222a8),
	.w1(32'h3a88a615),
	.w2(32'hbb560c02),
	.w3(32'h3bdef74e),
	.w4(32'h3c25b05a),
	.w5(32'hbb659b56),
	.w6(32'h3c7265ef),
	.w7(32'hbada3a09),
	.w8(32'h3b872996),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9f923),
	.w1(32'hbb8d4e83),
	.w2(32'h3a432d56),
	.w3(32'h3a7c6fe0),
	.w4(32'h3b4f6b6a),
	.w5(32'hbb76569a),
	.w6(32'hbbd2934c),
	.w7(32'hbb65a24c),
	.w8(32'h3b2fdc17),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab25e9d),
	.w1(32'hbba76fe8),
	.w2(32'hbb07f9de),
	.w3(32'hbb1d53b9),
	.w4(32'hbbb8cd00),
	.w5(32'h3bc1fd71),
	.w6(32'h3cc6b20c),
	.w7(32'h3bbdc036),
	.w8(32'h3bc87f8e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baca8e4),
	.w1(32'h3befbd32),
	.w2(32'hba1a451c),
	.w3(32'h3bf6abd1),
	.w4(32'h3c21d5e6),
	.w5(32'h3b80224e),
	.w6(32'h3b10042a),
	.w7(32'h3cc46cbe),
	.w8(32'h3ba2d2cd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959ba5e),
	.w1(32'hbb26e40d),
	.w2(32'h3b01fdbb),
	.w3(32'h3b5f9622),
	.w4(32'h3bec6d2e),
	.w5(32'hbb855794),
	.w6(32'h3b0d8f83),
	.w7(32'h3b1d072d),
	.w8(32'hbbe450ce),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14bd91),
	.w1(32'hbc3c44f7),
	.w2(32'hbc0278d3),
	.w3(32'hbb7848d8),
	.w4(32'hbc0d8d82),
	.w5(32'hbadaed74),
	.w6(32'h3b9b16d2),
	.w7(32'hbb01e43b),
	.w8(32'hbc005308),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3239d1),
	.w1(32'h3a343674),
	.w2(32'hbc237ba1),
	.w3(32'hbb8304cb),
	.w4(32'hbc1b7ac8),
	.w5(32'h3978e456),
	.w6(32'hbbdc333a),
	.w7(32'hbc66ccad),
	.w8(32'h3b19753a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd35c01),
	.w1(32'h3b9ef20b),
	.w2(32'hb79dc350),
	.w3(32'hbaeb96b7),
	.w4(32'h3b037da7),
	.w5(32'h3b65e379),
	.w6(32'h3ac97685),
	.w7(32'hba21b0df),
	.w8(32'h3bbf4a47),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76b615),
	.w1(32'h3bb9f7e6),
	.w2(32'hb825da2d),
	.w3(32'h3c5fd426),
	.w4(32'hbb3aa963),
	.w5(32'h3c3d024e),
	.w6(32'h3cbfbbdb),
	.w7(32'hbbfa8e62),
	.w8(32'h3be16a26),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39171890),
	.w1(32'h3c63a123),
	.w2(32'h3ae1490a),
	.w3(32'h3b827605),
	.w4(32'h38fc8d0c),
	.w5(32'hbaceea01),
	.w6(32'h3af2cfa9),
	.w7(32'hbb97be78),
	.w8(32'h3b12b625),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba992fa0),
	.w1(32'h3c3a29d3),
	.w2(32'hbb1b3ba5),
	.w3(32'h3c56a709),
	.w4(32'h3b4b8a46),
	.w5(32'hbaa1d76e),
	.w6(32'h3cb5fbf7),
	.w7(32'h3c70cb2b),
	.w8(32'h3b84abab),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5edb8),
	.w1(32'hba98eac5),
	.w2(32'hba42db5d),
	.w3(32'h3baa5eff),
	.w4(32'hbacdc70b),
	.w5(32'hbb4c97d8),
	.w6(32'h3c3e3c59),
	.w7(32'h3bd17d2b),
	.w8(32'h3c50d929),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1cf76),
	.w1(32'hb9b3bdc1),
	.w2(32'hba62c981),
	.w3(32'h3c3c8a67),
	.w4(32'h3c0e8122),
	.w5(32'h3abd6a41),
	.w6(32'h3cc074d5),
	.w7(32'h3c800c17),
	.w8(32'hbac2f24c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf714a),
	.w1(32'hba8e8687),
	.w2(32'h3ac75b75),
	.w3(32'h3a000978),
	.w4(32'h3c059a99),
	.w5(32'h3aa3c8bf),
	.w6(32'h3a1b4467),
	.w7(32'hbbacd6d7),
	.w8(32'h3c878b3d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0330ab),
	.w1(32'h3b144766),
	.w2(32'h3c22cf94),
	.w3(32'h3c836ff7),
	.w4(32'h3a9880bf),
	.w5(32'h3a6f8913),
	.w6(32'hbb3679d5),
	.w7(32'h3b0a0692),
	.w8(32'h3b38cd5c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7399c3),
	.w1(32'h3b77f35c),
	.w2(32'h3b806923),
	.w3(32'h3b4d8dff),
	.w4(32'h3b854e73),
	.w5(32'h3b37b5ac),
	.w6(32'h3b6d322a),
	.w7(32'h3bb5f112),
	.w8(32'h3ad24a09),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5827),
	.w1(32'hbb4dc1f6),
	.w2(32'hbb5d87ba),
	.w3(32'hbbcee1ee),
	.w4(32'hbba4acc4),
	.w5(32'hbad5bfde),
	.w6(32'hbba03389),
	.w7(32'hbb86e2b3),
	.w8(32'hbb42fc91),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b673f30),
	.w1(32'h3c0947f3),
	.w2(32'h3ab4c38d),
	.w3(32'h3bf1e60f),
	.w4(32'h3bc2cc5f),
	.w5(32'hbc03d373),
	.w6(32'h3b925982),
	.w7(32'h3bbc6775),
	.w8(32'hbb90334b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c71a0),
	.w1(32'hbb8ac65c),
	.w2(32'hbb074915),
	.w3(32'hbb83d268),
	.w4(32'hbb20892f),
	.w5(32'hbb9d84f3),
	.w6(32'hbb5f9cf6),
	.w7(32'hbab77568),
	.w8(32'hbb874553),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2066bb),
	.w1(32'hb98cd8e7),
	.w2(32'hbba7d513),
	.w3(32'h384d95cf),
	.w4(32'hbad96030),
	.w5(32'hbb90c7fd),
	.w6(32'hbaeab017),
	.w7(32'hbabd59c0),
	.w8(32'hbb6e301b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf6637),
	.w1(32'hbbc0d5fb),
	.w2(32'hbb7e60dc),
	.w3(32'hbbb2fbbe),
	.w4(32'hbba73c86),
	.w5(32'hbb4daf37),
	.w6(32'hbbd1ff09),
	.w7(32'hbb86fc72),
	.w8(32'hbb37419c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc205fad),
	.w1(32'hbb8d425e),
	.w2(32'hbbb2f54c),
	.w3(32'hbbc5cc4b),
	.w4(32'hbb80f491),
	.w5(32'hba4c8f79),
	.w6(32'hbc1ec7df),
	.w7(32'hbbe349cc),
	.w8(32'hb9e5da0a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa080a),
	.w1(32'hbb405be6),
	.w2(32'hbb6e8a2f),
	.w3(32'hbbbc00f5),
	.w4(32'hbb0f5829),
	.w5(32'h3bf5b079),
	.w6(32'hbb1afd0f),
	.w7(32'hbb14cae2),
	.w8(32'h3b80fa61),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf7d8f),
	.w1(32'hb9dea697),
	.w2(32'h39962c19),
	.w3(32'h3aae6179),
	.w4(32'hba62d65f),
	.w5(32'hbab4f433),
	.w6(32'hbaa2fd0d),
	.w7(32'hbb21f9b0),
	.w8(32'h3a93688d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923bd8a),
	.w1(32'h3ae85bf4),
	.w2(32'hb87521af),
	.w3(32'hbabc93f3),
	.w4(32'hbb267d06),
	.w5(32'hb9b8b997),
	.w6(32'h3ae595ac),
	.w7(32'h368bbe76),
	.w8(32'hb708a28e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc182439),
	.w1(32'hbb929a85),
	.w2(32'hba5a02ba),
	.w3(32'hbacdf185),
	.w4(32'hbb062e78),
	.w5(32'hbb57d5c1),
	.w6(32'hba592c08),
	.w7(32'hb9d2b245),
	.w8(32'hbb6634e9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc043996),
	.w1(32'hbb0c7239),
	.w2(32'h3a49063f),
	.w3(32'hbb47565d),
	.w4(32'hbb7297a4),
	.w5(32'hbb090fab),
	.w6(32'h3a88b6a0),
	.w7(32'h3a5da44e),
	.w8(32'hb8f7d230),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c2a09),
	.w1(32'hbab6c8b7),
	.w2(32'hba86a9f9),
	.w3(32'hbb4de81d),
	.w4(32'hbb5bbdff),
	.w5(32'hbaec4fb0),
	.w6(32'hbb3d073a),
	.w7(32'hbb3cba8b),
	.w8(32'hbaf0ec72),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e6553),
	.w1(32'h39c4140d),
	.w2(32'hbb323179),
	.w3(32'hbae02600),
	.w4(32'hbb463894),
	.w5(32'h3a5b8e9c),
	.w6(32'hbad76e6e),
	.w7(32'hbb15be38),
	.w8(32'h3ae1133b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa36c69),
	.w1(32'h3995b2c8),
	.w2(32'h39f3ca55),
	.w3(32'hbb159771),
	.w4(32'hbb1238f8),
	.w5(32'h3ae3c8b7),
	.w6(32'hbb67b4e5),
	.w7(32'hbb57edbb),
	.w8(32'h39e667a3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25c0e6),
	.w1(32'hbb6df581),
	.w2(32'hbba7207f),
	.w3(32'h3b32f73e),
	.w4(32'hba26bc36),
	.w5(32'hbb7dfd2b),
	.w6(32'h3a07d011),
	.w7(32'hbb4097b7),
	.w8(32'hbb84babe),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88cbdc),
	.w1(32'hbb59a192),
	.w2(32'hbb333bf7),
	.w3(32'hba07c642),
	.w4(32'h3a816d24),
	.w5(32'hbb8c9238),
	.w6(32'hbab3b3d8),
	.w7(32'hbb6b4748),
	.w8(32'hbb2ca37c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa66343),
	.w1(32'hba5b9c61),
	.w2(32'hbb0a95ab),
	.w3(32'hba84bcc7),
	.w4(32'hbb0180c1),
	.w5(32'h3b8c1b64),
	.w6(32'hbb25b10e),
	.w7(32'hbaab0335),
	.w8(32'h3b56bb59),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33ce4c),
	.w1(32'h3b765280),
	.w2(32'h3b9320b3),
	.w3(32'h3ad986d2),
	.w4(32'h3b456c52),
	.w5(32'h3a341149),
	.w6(32'h3b301bab),
	.w7(32'h3b937664),
	.w8(32'h3b8d1dda),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ac4a),
	.w1(32'h3b147130),
	.w2(32'hbadd6436),
	.w3(32'hba2b1f09),
	.w4(32'hbaa87ad1),
	.w5(32'hbafef1ae),
	.w6(32'h3aecb51d),
	.w7(32'h39a7515d),
	.w8(32'hbb8f2efd),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb853c7f),
	.w1(32'hbb0a0752),
	.w2(32'hbae51689),
	.w3(32'hbb002b71),
	.w4(32'hbadff9ff),
	.w5(32'h3a3bfb71),
	.w6(32'hbb71af06),
	.w7(32'hbb17ace5),
	.w8(32'h39b9b2df),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcf3b9),
	.w1(32'hbbaa9a65),
	.w2(32'hbb95e417),
	.w3(32'h3a80787a),
	.w4(32'h3a351bb4),
	.w5(32'hb9f40186),
	.w6(32'hb9874fae),
	.w7(32'h39406f7b),
	.w8(32'h39a425a6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85407fa),
	.w1(32'hb93b4c0e),
	.w2(32'hb995f29b),
	.w3(32'h3b630ebf),
	.w4(32'h3ae2e43a),
	.w5(32'hbb97998b),
	.w6(32'h38edb0a9),
	.w7(32'h398bba20),
	.w8(32'hbba8bd6a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9729d1),
	.w1(32'hbbac9798),
	.w2(32'hbaaa922f),
	.w3(32'hbbac040e),
	.w4(32'hba635793),
	.w5(32'hbb945adc),
	.w6(32'hbbc25b70),
	.w7(32'hbab40b1c),
	.w8(32'hb9735f08),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d6f0a),
	.w1(32'h39370ff8),
	.w2(32'h3a9d4e0c),
	.w3(32'hbbd0d333),
	.w4(32'hbb5c82e6),
	.w5(32'hbb04e3b4),
	.w6(32'hbb828c72),
	.w7(32'hbb6f3ea0),
	.w8(32'hbbac95e9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb619e13),
	.w1(32'hbaa2bf5f),
	.w2(32'h3aa99af5),
	.w3(32'hba93291e),
	.w4(32'hb925a26b),
	.w5(32'hbbabb5a0),
	.w6(32'hba37c3c8),
	.w7(32'hbaaa8906),
	.w8(32'hbac1d73f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31d21f),
	.w1(32'hbaa7956f),
	.w2(32'hba910040),
	.w3(32'hbb14a232),
	.w4(32'hbb7e9136),
	.w5(32'h3a6051ee),
	.w6(32'hb9ac4389),
	.w7(32'h39a81180),
	.w8(32'h3bbb4f4b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b072e11),
	.w1(32'h3b71836e),
	.w2(32'h3a9bee32),
	.w3(32'h3a21b650),
	.w4(32'hba6f11a9),
	.w5(32'hbb7abfa7),
	.w6(32'h3b6c3963),
	.w7(32'h397ad1c6),
	.w8(32'hbacebaf6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add12c8),
	.w1(32'h3afdef29),
	.w2(32'h3ab25548),
	.w3(32'hbae72401),
	.w4(32'h3ab1b758),
	.w5(32'h3a1141d6),
	.w6(32'hbaa725b2),
	.w7(32'h3a0f4069),
	.w8(32'hbab525ff),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba21994),
	.w1(32'hbb76dec9),
	.w2(32'hbb80c81c),
	.w3(32'hbad6f135),
	.w4(32'h3902732b),
	.w5(32'hbbb62a38),
	.w6(32'hbaef2faa),
	.w7(32'hbb1aeb92),
	.w8(32'hbb53e427),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11b235),
	.w1(32'hbbe0f72b),
	.w2(32'hbb65aa89),
	.w3(32'hbb744a33),
	.w4(32'hbbba512e),
	.w5(32'hbb9a4152),
	.w6(32'hb9d36f46),
	.w7(32'hbafe89fc),
	.w8(32'hbb794ecd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb261d80),
	.w1(32'hbb4eb493),
	.w2(32'hbae2135b),
	.w3(32'hbb7c2e73),
	.w4(32'hbb49c5d7),
	.w5(32'hbba59988),
	.w6(32'hbbb40f30),
	.w7(32'hbba9cf4e),
	.w8(32'hb9db78e7),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c98c8),
	.w1(32'hbb2b75bb),
	.w2(32'hbb7722cb),
	.w3(32'h3a6be658),
	.w4(32'hbb331a52),
	.w5(32'hb9fdbb32),
	.w6(32'hbb5b69f3),
	.w7(32'hbb08cdd8),
	.w8(32'hb8b98ce3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb4bb0),
	.w1(32'hbaa8082d),
	.w2(32'hba90d5e0),
	.w3(32'hba8875f8),
	.w4(32'hb8c000d7),
	.w5(32'hbba030f2),
	.w6(32'hbac7662d),
	.w7(32'hb9a6ba85),
	.w8(32'hbb880fd1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7ceac),
	.w1(32'hbbb15c12),
	.w2(32'hbbee08ae),
	.w3(32'hbbbf7a87),
	.w4(32'hbb8a9a36),
	.w5(32'hbb8f5d58),
	.w6(32'hbbf08561),
	.w7(32'hbbd2ff1e),
	.w8(32'hbb498d05),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2a671),
	.w1(32'hb92ed8e6),
	.w2(32'hbabf1b90),
	.w3(32'hbb43c1e8),
	.w4(32'hbae237da),
	.w5(32'hbb1f4d53),
	.w6(32'hba973fa0),
	.w7(32'hba5d2d1f),
	.w8(32'hbaae34fa),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba411ae),
	.w1(32'hbb17417c),
	.w2(32'hb9f94bb2),
	.w3(32'hbb867ae8),
	.w4(32'h39897378),
	.w5(32'hbac0b56c),
	.w6(32'hbb98c77f),
	.w7(32'h3a8aa3bf),
	.w8(32'hb9cb9b23),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6718a9),
	.w1(32'hbb73ff9f),
	.w2(32'hbaf048f6),
	.w3(32'h3a161829),
	.w4(32'hbb1c4e99),
	.w5(32'hba29687e),
	.w6(32'hbaebfc8b),
	.w7(32'hba87b238),
	.w8(32'hba36349e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd0ab),
	.w1(32'hba98cb44),
	.w2(32'hb899a565),
	.w3(32'hbb1913c6),
	.w4(32'hbaa6cee0),
	.w5(32'hbb17ade8),
	.w6(32'hbb557d67),
	.w7(32'hba30efc5),
	.w8(32'hbb15e444),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b9386),
	.w1(32'hba3adbb9),
	.w2(32'hbad92aad),
	.w3(32'hbb463c29),
	.w4(32'hb9c09424),
	.w5(32'hbb9a110a),
	.w6(32'hbb4d11aa),
	.w7(32'h3a65bc77),
	.w8(32'hb9dd6b30),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f1475),
	.w1(32'hba83cbc3),
	.w2(32'hb9027bb5),
	.w3(32'hbb78998e),
	.w4(32'hba7b4fd4),
	.w5(32'h3bc696ab),
	.w6(32'hbaf7e086),
	.w7(32'h3a7f4271),
	.w8(32'h3b8e5e57),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03f6a0),
	.w1(32'hbbbac933),
	.w2(32'hbb7008bf),
	.w3(32'h3c0dc47d),
	.w4(32'h3acbed5d),
	.w5(32'hbb9fe5b9),
	.w6(32'hbabfc040),
	.w7(32'hbab2e9b9),
	.w8(32'hbbc60103),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb801e1),
	.w1(32'hbbc89247),
	.w2(32'hbbb36067),
	.w3(32'hbbb33582),
	.w4(32'hbb14d5d9),
	.w5(32'h3abb1d71),
	.w6(32'hbbc508c5),
	.w7(32'hbb88439d),
	.w8(32'h3b16ccd9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d21a1f),
	.w1(32'h3ae06a6c),
	.w2(32'hbadced23),
	.w3(32'hbaae0df8),
	.w4(32'hbb3d6cab),
	.w5(32'h3a2a48c4),
	.w6(32'hba9e33d3),
	.w7(32'hbb84d4c9),
	.w8(32'hb9a9ea08),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f0078),
	.w1(32'h3a173f32),
	.w2(32'h3a1ce540),
	.w3(32'h3a931f2e),
	.w4(32'h3a5bedad),
	.w5(32'h3bae9b0f),
	.w6(32'hba0c79b5),
	.w7(32'h3a06e6a1),
	.w8(32'h3bcb08cd),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc70aaf),
	.w1(32'h3b2ae895),
	.w2(32'hbae473bc),
	.w3(32'hb9b834c3),
	.w4(32'hbb5f14fd),
	.w5(32'hb94b192f),
	.w6(32'hba79c634),
	.w7(32'hbb5443e7),
	.w8(32'h3a6e195c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9166c00),
	.w1(32'hba870905),
	.w2(32'hbb1e0853),
	.w3(32'hba19414e),
	.w4(32'hbac3e120),
	.w5(32'hba5d6ecd),
	.w6(32'h3a475048),
	.w7(32'hbb3c93f5),
	.w8(32'hba825b5e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0485a2),
	.w1(32'hba5695e9),
	.w2(32'hba484fd0),
	.w3(32'hbb43f0e9),
	.w4(32'hba1d9f6b),
	.w5(32'hbb03016b),
	.w6(32'hba9ec730),
	.w7(32'hbac42a8b),
	.w8(32'hbaf71a07),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07a35a),
	.w1(32'hb957afec),
	.w2(32'hbb48cabc),
	.w3(32'hba50306a),
	.w4(32'hb91cb685),
	.w5(32'h3b87d0fe),
	.w6(32'hb937e4e2),
	.w7(32'hba5742ee),
	.w8(32'h3c0246c3),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe114f1),
	.w1(32'hbad3a631),
	.w2(32'hb9dba47b),
	.w3(32'hba8a3f1b),
	.w4(32'h39dc396d),
	.w5(32'h3b269b6c),
	.w6(32'hbb1ab275),
	.w7(32'hbb43813b),
	.w8(32'h3bacb7af),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05be34),
	.w1(32'h3b3597c9),
	.w2(32'hbb0e4c39),
	.w3(32'hbb1b3190),
	.w4(32'hbb958e42),
	.w5(32'h3b9974f9),
	.w6(32'hbab9d9b4),
	.w7(32'hbb849d4c),
	.w8(32'h3b82cc7e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a4ec6),
	.w1(32'h3a87b26a),
	.w2(32'h3aa23379),
	.w3(32'h3b44aab4),
	.w4(32'h3b17bfce),
	.w5(32'h3a78cdf8),
	.w6(32'h3b6c3ecb),
	.w7(32'h3b65c78b),
	.w8(32'h3aa2cba4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf4fe1),
	.w1(32'hbbd1f123),
	.w2(32'hbb8cd62b),
	.w3(32'hbb006bdd),
	.w4(32'hbb820cdc),
	.w5(32'h3b2a9717),
	.w6(32'hbb814ba4),
	.w7(32'hbb87bcbc),
	.w8(32'h3b0f5ea1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba652b74),
	.w1(32'hbb625e5b),
	.w2(32'hbb58f1e7),
	.w3(32'hbbe3073e),
	.w4(32'hbba05a14),
	.w5(32'hbae93af3),
	.w6(32'hbbfbdc85),
	.w7(32'hbb3a86e9),
	.w8(32'h38bcbaa9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79553f),
	.w1(32'hba6e1993),
	.w2(32'hbb3d74ed),
	.w3(32'h3acbe38a),
	.w4(32'h3acfd68e),
	.w5(32'hbbbd05fc),
	.w6(32'h3a8dc559),
	.w7(32'h3a639bb2),
	.w8(32'hbaa8e78c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22558b),
	.w1(32'h3afe2223),
	.w2(32'h3b1f8c19),
	.w3(32'hbaa9d2c9),
	.w4(32'h3a73b21a),
	.w5(32'hbab509b3),
	.w6(32'hba683702),
	.w7(32'h3a8d9c33),
	.w8(32'hb999886d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa75e52),
	.w1(32'hb8d4d8db),
	.w2(32'h3abd0764),
	.w3(32'hbb23bb09),
	.w4(32'hbab5206a),
	.w5(32'hbb0f73f9),
	.w6(32'hbb3b9650),
	.w7(32'hbafadcdd),
	.w8(32'hbb1afb99),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97f6d7),
	.w1(32'h3a81763f),
	.w2(32'h38aeed6e),
	.w3(32'h3a97b5af),
	.w4(32'hbb43759b),
	.w5(32'hbb04f754),
	.w6(32'h3b959a43),
	.w7(32'h3a5d8ede),
	.w8(32'h3b36b00b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4da0a6),
	.w1(32'h3b83b84f),
	.w2(32'hb8f168b6),
	.w3(32'hbaa2a115),
	.w4(32'h3aa7cefa),
	.w5(32'hbbd62af3),
	.w6(32'h3a74ee8f),
	.w7(32'h3ad8850d),
	.w8(32'hbb9e3d25),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3c8e1),
	.w1(32'hbb00ca7c),
	.w2(32'hba0610ee),
	.w3(32'hbb12faf9),
	.w4(32'h3888e4aa),
	.w5(32'h3b3f69bd),
	.w6(32'hbaec1b03),
	.w7(32'hb9fc384a),
	.w8(32'h3bb45e23),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba540928),
	.w1(32'h3b94c10d),
	.w2(32'h3ba2eebc),
	.w3(32'h3af676ad),
	.w4(32'h3b0775f0),
	.w5(32'h3b89f25a),
	.w6(32'h3bd8af0b),
	.w7(32'h3bbabc30),
	.w8(32'h3af42689),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba2048),
	.w1(32'hba5b441e),
	.w2(32'hbab78a23),
	.w3(32'h3c314910),
	.w4(32'h3c21c3ac),
	.w5(32'hbb8b93d7),
	.w6(32'h3b353d20),
	.w7(32'h3ae58266),
	.w8(32'hbbb3bb60),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b75c9),
	.w1(32'hbb4fd45f),
	.w2(32'hbb5e21a3),
	.w3(32'hbb759263),
	.w4(32'hb9fbb430),
	.w5(32'hb9e8428b),
	.w6(32'hbb65c6df),
	.w7(32'hba3a979f),
	.w8(32'hbae983bd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab881fa),
	.w1(32'hbb4f2df3),
	.w2(32'hbaeb053f),
	.w3(32'hbb5bd0f4),
	.w4(32'hbb079b51),
	.w5(32'hbb0e19a3),
	.w6(32'hba71bf1a),
	.w7(32'hba57529c),
	.w8(32'hba00683c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb835f1f4),
	.w1(32'hba93cd15),
	.w2(32'hbb8d07ec),
	.w3(32'hbadb2809),
	.w4(32'hbab0a3dc),
	.w5(32'h398de476),
	.w6(32'h3a1b7021),
	.w7(32'hbac39913),
	.w8(32'hbaa16ec8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99495c4),
	.w1(32'hbb66566c),
	.w2(32'hbb16b304),
	.w3(32'hbb0101f6),
	.w4(32'hbb3362bb),
	.w5(32'h3a5f19f9),
	.w6(32'hbb30eec5),
	.w7(32'hbb4a2fda),
	.w8(32'h3b9d8cb8),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14c607),
	.w1(32'h3b88384e),
	.w2(32'h3b97f243),
	.w3(32'hba80ff44),
	.w4(32'hb70da73c),
	.w5(32'hbb64a26d),
	.w6(32'h3b8b8db7),
	.w7(32'h38ee25bd),
	.w8(32'hba971a10),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7139ae),
	.w1(32'hbb6079a1),
	.w2(32'hbb3251ac),
	.w3(32'hbbb0e0ed),
	.w4(32'hbaecfd69),
	.w5(32'hba87b8e0),
	.w6(32'hbbb60937),
	.w7(32'hba1444a9),
	.w8(32'hbb50ab40),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fb96d),
	.w1(32'hbb1d95d0),
	.w2(32'hb9bc4748),
	.w3(32'hbaac4a1f),
	.w4(32'hbb06f693),
	.w5(32'hb9a2f95c),
	.w6(32'hba98fe84),
	.w7(32'hbb0e0d8d),
	.w8(32'h3b1893fa),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5b0a6),
	.w1(32'h3b8e490f),
	.w2(32'h3ad53a21),
	.w3(32'h3b5f7461),
	.w4(32'h3b84b9d9),
	.w5(32'h3b0045df),
	.w6(32'h3bba47d2),
	.w7(32'h3bc5750d),
	.w8(32'h39167c06),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f39d8),
	.w1(32'hbb436b1d),
	.w2(32'hbadb05a9),
	.w3(32'h398a57e0),
	.w4(32'hbb7fc657),
	.w5(32'hbbe520d3),
	.w6(32'h3aa898ed),
	.w7(32'h39d459be),
	.w8(32'hba744715),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb087dbd),
	.w1(32'hb96e3314),
	.w2(32'h3ae9ae9a),
	.w3(32'hba8541cf),
	.w4(32'h3aa0ee54),
	.w5(32'h3a38d1eb),
	.w6(32'hbb19772c),
	.w7(32'h3a6cdf3f),
	.w8(32'h3acd7a63),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf0c1d),
	.w1(32'hbb6e4ef5),
	.w2(32'hbb6a1f0a),
	.w3(32'hbb803e32),
	.w4(32'hbb467cf6),
	.w5(32'hbba45cdb),
	.w6(32'hbb4b30c5),
	.w7(32'hba367025),
	.w8(32'hbbb37acb),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96d6b3),
	.w1(32'hbb5dd982),
	.w2(32'hbb771dfa),
	.w3(32'hbbad0a56),
	.w4(32'hbba3c7ac),
	.w5(32'h3af35ecc),
	.w6(32'hbba3b53a),
	.w7(32'hbbabd45e),
	.w8(32'h3abec5b4),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb11fa),
	.w1(32'hbc06e215),
	.w2(32'hbb74b571),
	.w3(32'hbadf4d4b),
	.w4(32'hba8cce6f),
	.w5(32'hbb17acf1),
	.w6(32'hbb9a32d0),
	.w7(32'h3a0b75dd),
	.w8(32'h390af1eb),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adae026),
	.w1(32'h3baac0f4),
	.w2(32'h3b82bf50),
	.w3(32'hb9b270af),
	.w4(32'hb95915d0),
	.w5(32'h3abba4a8),
	.w6(32'h3bc03ce5),
	.w7(32'h3b824a5f),
	.w8(32'h3af63c44),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb62b71),
	.w1(32'hbbbadff7),
	.w2(32'hbb9c7452),
	.w3(32'hba9f11e4),
	.w4(32'hbbbce894),
	.w5(32'hb9d452ae),
	.w6(32'hbb28d4f2),
	.w7(32'hbb759275),
	.w8(32'h394ab69a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed59f2),
	.w1(32'h3ab6b28a),
	.w2(32'h3b1c59ce),
	.w3(32'h3a1bb531),
	.w4(32'h3ac93a9f),
	.w5(32'hbb616ec7),
	.w6(32'hb9ea2a60),
	.w7(32'hb99592b1),
	.w8(32'hbbaa2782),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86fde2),
	.w1(32'hbb67b2e7),
	.w2(32'hbbb4cea5),
	.w3(32'hba9c2a2f),
	.w4(32'hbb3ba0bf),
	.w5(32'h3ae75ce4),
	.w6(32'hbb3e8bd1),
	.w7(32'hbb2b373f),
	.w8(32'h3b3e0d13),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2c152),
	.w1(32'h3b636795),
	.w2(32'h3b512ff8),
	.w3(32'h3b76ff00),
	.w4(32'h3b956866),
	.w5(32'hba98b53e),
	.w6(32'h3b897781),
	.w7(32'h3b90a07c),
	.w8(32'hbb3a5e8a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47de98),
	.w1(32'hb8a3279c),
	.w2(32'hb9749828),
	.w3(32'h3996a0ba),
	.w4(32'hbb004364),
	.w5(32'hbadc6d0a),
	.w6(32'hbacde5f9),
	.w7(32'hb9d79518),
	.w8(32'hbb1c0843),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f795e),
	.w1(32'hbb07a128),
	.w2(32'hbb2549c5),
	.w3(32'hba424cb6),
	.w4(32'hba781037),
	.w5(32'hb9fcdc66),
	.w6(32'hbb21a15c),
	.w7(32'hbb26455c),
	.w8(32'hba406bd1),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc39572),
	.w1(32'hbb7b3248),
	.w2(32'hbacbf8c7),
	.w3(32'hbaf34d41),
	.w4(32'hbb5b3db2),
	.w5(32'hba797336),
	.w6(32'hbb66e8de),
	.w7(32'hbb057579),
	.w8(32'h3aa55073),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39925e79),
	.w1(32'h39534f15),
	.w2(32'h3a60e2c4),
	.w3(32'h3b807498),
	.w4(32'hb7b1ff20),
	.w5(32'h3a97401e),
	.w6(32'h3a666fe6),
	.w7(32'hbaf85808),
	.w8(32'h3b47ae20),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b540a99),
	.w1(32'h3b50fa63),
	.w2(32'hb8b3ff46),
	.w3(32'h3afcab7f),
	.w4(32'h3a3b20c6),
	.w5(32'hbb7974af),
	.w6(32'h3a69b19f),
	.w7(32'hba03a2f7),
	.w8(32'hbaf32b67),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5c65c),
	.w1(32'hb9d63eb7),
	.w2(32'hba94aeff),
	.w3(32'hbae0fb42),
	.w4(32'hbb28e844),
	.w5(32'h3b8d5c88),
	.w6(32'hb96fe9f2),
	.w7(32'hba74ee2b),
	.w8(32'h3b292962),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e65f5),
	.w1(32'h3b00f76c),
	.w2(32'hbaaa48bd),
	.w3(32'h3b1d5e10),
	.w4(32'hb9de8704),
	.w5(32'h3acbb576),
	.w6(32'h3a9012aa),
	.w7(32'hb9058fb6),
	.w8(32'h3bc2cc69),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc7cfa),
	.w1(32'h3b322cbe),
	.w2(32'h39f747f8),
	.w3(32'h3b26608b),
	.w4(32'hba853d7c),
	.w5(32'h3aba422c),
	.w6(32'h3a70560b),
	.w7(32'hbab6990a),
	.w8(32'h3ab5cf29),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a720c5),
	.w1(32'h3b0878b1),
	.w2(32'h3b598a58),
	.w3(32'h3b195e60),
	.w4(32'h3b7d0cca),
	.w5(32'hba4570d3),
	.w6(32'h3b1c2e35),
	.w7(32'h3b95120d),
	.w8(32'hbb5fef1e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d35c4),
	.w1(32'hbb9cab76),
	.w2(32'hb9dd72ae),
	.w3(32'hbc0bcfd3),
	.w4(32'h3a4cb77c),
	.w5(32'hb9eccf45),
	.w6(32'hbc18edd5),
	.w7(32'h3bce0ea9),
	.w8(32'h3ae1c93b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6827a),
	.w1(32'h3a1f6dbf),
	.w2(32'h3b32eda3),
	.w3(32'h3b4aafe4),
	.w4(32'h3aa0b6cc),
	.w5(32'hba55ba8b),
	.w6(32'h3b1ccc17),
	.w7(32'h3b1445df),
	.w8(32'hbad428a0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc8b15),
	.w1(32'h3b1aaccd),
	.w2(32'h3b12d015),
	.w3(32'h3a98070c),
	.w4(32'h3b0f1eae),
	.w5(32'hbb122ce3),
	.w6(32'hb9473af9),
	.w7(32'hbaa085bc),
	.w8(32'hba7c614e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e9b17),
	.w1(32'hbacad3eb),
	.w2(32'hbb13e011),
	.w3(32'hbacc8da0),
	.w4(32'hba63463f),
	.w5(32'hba7eec87),
	.w6(32'hba9aa10b),
	.w7(32'hbad39d11),
	.w8(32'hba34a75c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd7439),
	.w1(32'hba8e113d),
	.w2(32'hb9f40884),
	.w3(32'h3993d687),
	.w4(32'hba9a0d46),
	.w5(32'hbb297dd3),
	.w6(32'hb941d5e7),
	.w7(32'hba9fc16c),
	.w8(32'hba99017f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed665d),
	.w1(32'hba4252ef),
	.w2(32'hbb336dfc),
	.w3(32'hba28919d),
	.w4(32'hbac93520),
	.w5(32'hbb1d99d6),
	.w6(32'hb9e5c530),
	.w7(32'hba6d32e2),
	.w8(32'hba5a2d10),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b233a0a),
	.w1(32'h3acfa2d8),
	.w2(32'hb9897936),
	.w3(32'h39bea070),
	.w4(32'hb9604700),
	.w5(32'hbb00264f),
	.w6(32'hbb1e8f5d),
	.w7(32'hbb11b984),
	.w8(32'h3ad1ce56),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a288c2c),
	.w1(32'hbae9823e),
	.w2(32'hbb021030),
	.w3(32'h3a2e03de),
	.w4(32'hbb35e889),
	.w5(32'hbbc5c36c),
	.w6(32'hbb01f24e),
	.w7(32'hbb14c68b),
	.w8(32'hbb92447b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cda7a),
	.w1(32'hbbfda328),
	.w2(32'hbba4640a),
	.w3(32'hbbc34408),
	.w4(32'hbba707a4),
	.w5(32'hbba4bc53),
	.w6(32'hbc29c2c2),
	.w7(32'hbbeedae2),
	.w8(32'hbb90259e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25e90f),
	.w1(32'hba29d229),
	.w2(32'hbb51ddc3),
	.w3(32'hbaea2fdd),
	.w4(32'hbbb27bad),
	.w5(32'hbab7717e),
	.w6(32'hbb5f4b54),
	.w7(32'hbb832871),
	.w8(32'hbbb39e6a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d4417),
	.w1(32'hbc070cc5),
	.w2(32'hbbd1c50a),
	.w3(32'hbbfca0b5),
	.w4(32'hbb9e95c7),
	.w5(32'hb9f00cf5),
	.w6(32'hbbdfbcb3),
	.w7(32'hbb813310),
	.w8(32'h3b3d1612),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e392d),
	.w1(32'hbab09880),
	.w2(32'hba59b719),
	.w3(32'hbac75ce9),
	.w4(32'h38c738b0),
	.w5(32'h3b69f661),
	.w6(32'hba9488d3),
	.w7(32'h39c0ae7a),
	.w8(32'h3b7a917e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15668e),
	.w1(32'hbbb765f3),
	.w2(32'hbba48f72),
	.w3(32'hbb2976cc),
	.w4(32'hbbc927c7),
	.w5(32'h3b42e9ea),
	.w6(32'hbb462d10),
	.w7(32'hbb293d57),
	.w8(32'hbb18d804),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a3c8a),
	.w1(32'hbb4b2b69),
	.w2(32'hbaba25f8),
	.w3(32'h36aaf262),
	.w4(32'hbac2f7f7),
	.w5(32'hbb4cb16d),
	.w6(32'hbb1c22ca),
	.w7(32'hbb77ab2d),
	.w8(32'hbb825ff4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e825f),
	.w1(32'hbb89ab3b),
	.w2(32'hbb5a8e57),
	.w3(32'hbb4e1769),
	.w4(32'hbac12ea2),
	.w5(32'hbb1f143a),
	.w6(32'hbb5278ae),
	.w7(32'hbb03c366),
	.w8(32'h3a321f76),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ccd92),
	.w1(32'hbb82c46d),
	.w2(32'hbb311208),
	.w3(32'hbb1b6c5b),
	.w4(32'hbb5aa78d),
	.w5(32'hbb6a0bca),
	.w6(32'hbb1f2093),
	.w7(32'hbb066bf7),
	.w8(32'hbb5a95ec),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45d12a),
	.w1(32'hbb184808),
	.w2(32'hba4c59d1),
	.w3(32'hbb9a606e),
	.w4(32'hba2fa643),
	.w5(32'h394140d1),
	.w6(32'hbbb3c78a),
	.w7(32'hbaf525bf),
	.w8(32'h3a4c2ea3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67f691),
	.w1(32'hbb1627fb),
	.w2(32'hbb35a116),
	.w3(32'hbb20ba93),
	.w4(32'hbb2b616b),
	.w5(32'h3aae01d8),
	.w6(32'hbb278950),
	.w7(32'hbae5cd10),
	.w8(32'hb9d9c2f6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4368ad),
	.w1(32'hbb6e2a0d),
	.w2(32'hbb84a7a3),
	.w3(32'hbb58c6b4),
	.w4(32'hbb3b8e40),
	.w5(32'hbb2e7bf2),
	.w6(32'hbb8cc292),
	.w7(32'hbb7a27ac),
	.w8(32'hbb583e26),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75b942),
	.w1(32'hbb883c9f),
	.w2(32'hbb54de3e),
	.w3(32'hbb851b4f),
	.w4(32'hbb9bba3b),
	.w5(32'hbad08318),
	.w6(32'hbbc073ea),
	.w7(32'hbb3fdd8e),
	.w8(32'hb9df8efe),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c9adf),
	.w1(32'hba0b2a11),
	.w2(32'hb9de263f),
	.w3(32'hbb29b0e9),
	.w4(32'hbb71c98a),
	.w5(32'hbac89942),
	.w6(32'hba08eb22),
	.w7(32'hbada3872),
	.w8(32'hba9f9904),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57e856),
	.w1(32'hbc5aad50),
	.w2(32'hbc0a06bf),
	.w3(32'hbbd19b02),
	.w4(32'hbb990918),
	.w5(32'hbb2be441),
	.w6(32'hbc0c0785),
	.w7(32'hbb6bc748),
	.w8(32'hbbc1a5e6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2b1a0),
	.w1(32'hbaeb9fac),
	.w2(32'hbb2c7f1d),
	.w3(32'hba9d7ff1),
	.w4(32'hba73fae5),
	.w5(32'hbb01d318),
	.w6(32'h3a015d1f),
	.w7(32'h39893498),
	.w8(32'hbadae345),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4202e),
	.w1(32'hba4a778d),
	.w2(32'h3a213635),
	.w3(32'hbaeafb63),
	.w4(32'hbaa0ebf1),
	.w5(32'hbbeba7fa),
	.w6(32'hbb207daf),
	.w7(32'h39f10459),
	.w8(32'hbb8c1b5f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95cc9f),
	.w1(32'hbb914aed),
	.w2(32'hbb4392fc),
	.w3(32'hbbb7893f),
	.w4(32'hbb0acfd8),
	.w5(32'hbb0b7fd2),
	.w6(32'hbb9b5670),
	.w7(32'h396b9508),
	.w8(32'hb969e05b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb535959),
	.w1(32'hbb40fca6),
	.w2(32'hbb2a5c4e),
	.w3(32'hbad4a0cd),
	.w4(32'hbb816253),
	.w5(32'hbc059b5c),
	.w6(32'hbace1a6b),
	.w7(32'hba4ec10d),
	.w8(32'h3a70cd6c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c8327),
	.w1(32'h3a3f9d96),
	.w2(32'h3940e480),
	.w3(32'hbac53e87),
	.w4(32'hbb3476d6),
	.w5(32'h3b36bebd),
	.w6(32'h37c2e465),
	.w7(32'h399a76df),
	.w8(32'h3ba95bf2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c7873f),
	.w1(32'h3af2f9ca),
	.w2(32'h3a9716c8),
	.w3(32'h3bdac35b),
	.w4(32'hbaabbdc4),
	.w5(32'hba597524),
	.w6(32'h3b058e8a),
	.w7(32'hba9025b2),
	.w8(32'h3ade495a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a9c1e),
	.w1(32'hba007406),
	.w2(32'hba291f41),
	.w3(32'hba50bc1f),
	.w4(32'h39a89db2),
	.w5(32'h3a97ae66),
	.w6(32'h39ac7a68),
	.w7(32'hba09279f),
	.w8(32'h3aa320f6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac02c76),
	.w1(32'h3ae78199),
	.w2(32'h3a8b9cd5),
	.w3(32'h3a8b3991),
	.w4(32'h3a8b1c04),
	.w5(32'hbc1aeff4),
	.w6(32'h3a8101bd),
	.w7(32'h3a2c3555),
	.w8(32'hbbf0eaeb),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02fffc),
	.w1(32'hbb718c24),
	.w2(32'hbac34d57),
	.w3(32'hbbe8f12a),
	.w4(32'hbb028de8),
	.w5(32'hbb6b031d),
	.w6(32'hbbb17f30),
	.w7(32'hbaefb166),
	.w8(32'hbb606b71),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4787ec),
	.w1(32'hbc4cedb2),
	.w2(32'hbb91d909),
	.w3(32'hbc7ac0e8),
	.w4(32'hbba533d7),
	.w5(32'hbb77aa7c),
	.w6(32'hbc86f9ad),
	.w7(32'hbac0454e),
	.w8(32'hbb6d4d20),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f186d),
	.w1(32'hbb22dd0e),
	.w2(32'hbacf8650),
	.w3(32'hba9bc09e),
	.w4(32'h3b9c9e8d),
	.w5(32'hb910892f),
	.w6(32'hbba8cf1d),
	.w7(32'h39e8f261),
	.w8(32'h3a602cf8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb029948),
	.w1(32'hbb0cd41d),
	.w2(32'hbaa0a1e6),
	.w3(32'h3a033833),
	.w4(32'h394ea54f),
	.w5(32'hbb62bddf),
	.w6(32'hbb31ea5a),
	.w7(32'hbba56e67),
	.w8(32'hbb398d1c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb91fcd),
	.w1(32'hbadea3fb),
	.w2(32'hbb0f4b10),
	.w3(32'hba990c0b),
	.w4(32'hbb21bb31),
	.w5(32'hbb66938e),
	.w6(32'hb9e3594d),
	.w7(32'hba28f892),
	.w8(32'hbae544b3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2145b2),
	.w1(32'hbb81ca1e),
	.w2(32'hbad56dde),
	.w3(32'hbb22b2a4),
	.w4(32'hbb10a6d8),
	.w5(32'hba95552e),
	.w6(32'hbb7b0184),
	.w7(32'hba212342),
	.w8(32'hb9fb2355),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae480c4),
	.w1(32'hbbb42fb0),
	.w2(32'hbac724c1),
	.w3(32'h3b088187),
	.w4(32'h3b01c3e7),
	.w5(32'hbb370c1f),
	.w6(32'hbb3c7e95),
	.w7(32'hba3c1730),
	.w8(32'hbb8b4cf8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb360023),
	.w1(32'hba5619de),
	.w2(32'h3972329f),
	.w3(32'hba644fcf),
	.w4(32'h3a3817d2),
	.w5(32'h3a91aa54),
	.w6(32'hbb54945c),
	.w7(32'hba1028b5),
	.w8(32'hbabfce2d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84e7e1),
	.w1(32'hbb151d4a),
	.w2(32'hbb232b9f),
	.w3(32'hbb3d29f1),
	.w4(32'hbb723343),
	.w5(32'hba537fd4),
	.w6(32'hbb9c1314),
	.w7(32'hbb840a9d),
	.w8(32'hbaa542fb),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7f2d6),
	.w1(32'h3a2bcfcb),
	.w2(32'h3a3d066a),
	.w3(32'hbaa0f0f8),
	.w4(32'hba47a623),
	.w5(32'h3b0daa66),
	.w6(32'hbb120b0c),
	.w7(32'hba52cebb),
	.w8(32'h3a97f63b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a051dda),
	.w1(32'hba76d173),
	.w2(32'hbb4f8afd),
	.w3(32'h3b1425a2),
	.w4(32'h378d8aad),
	.w5(32'hbb37b054),
	.w6(32'h3ab05735),
	.w7(32'h3a69c4dd),
	.w8(32'hbb22ef92),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb527302),
	.w1(32'hbb51d14b),
	.w2(32'hbad150e1),
	.w3(32'hb9680cbf),
	.w4(32'hbaad6b72),
	.w5(32'hbb4eec0e),
	.w6(32'hba0488d4),
	.w7(32'hba07e448),
	.w8(32'hbb981701),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a62e34),
	.w1(32'hba97ce44),
	.w2(32'hbb7d3732),
	.w3(32'hbb25a421),
	.w4(32'hbb173d04),
	.w5(32'hbafe5eec),
	.w6(32'hb9aa65fe),
	.w7(32'h3a2ca0d4),
	.w8(32'hbb91fea2),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0a26d),
	.w1(32'hbb897c25),
	.w2(32'hbb5c7eab),
	.w3(32'hbb7297d8),
	.w4(32'h3a7db5ac),
	.w5(32'h3ace7c3f),
	.w6(32'hbb9ba5f5),
	.w7(32'h3a8be1dd),
	.w8(32'h3adbb817),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f398d),
	.w1(32'hb9b4be25),
	.w2(32'h38ec8c59),
	.w3(32'h3ad2b029),
	.w4(32'h3ab21d99),
	.w5(32'hbb934d5d),
	.w6(32'hb98ba5e0),
	.w7(32'h3a440091),
	.w8(32'hbbfe5360),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe28742),
	.w1(32'hbbd24725),
	.w2(32'hbbc18e30),
	.w3(32'hbb9e9dea),
	.w4(32'hbb5843e7),
	.w5(32'h3bc3e4b1),
	.w6(32'hbc0a6ef1),
	.w7(32'hbc13ebfc),
	.w8(32'h3bf09925),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7d31b),
	.w1(32'hba127a5e),
	.w2(32'hba88c0ec),
	.w3(32'h3abf97b3),
	.w4(32'h3a93eae3),
	.w5(32'hbb9492ba),
	.w6(32'h3b28a6c2),
	.w7(32'h3ab8748b),
	.w8(32'hbb83cebc),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb146b77),
	.w1(32'hba493650),
	.w2(32'h392507d0),
	.w3(32'h3af97d9b),
	.w4(32'hbae4965d),
	.w5(32'hb966b200),
	.w6(32'hba0735b4),
	.w7(32'h396fefdf),
	.w8(32'h38d572f0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a603afa),
	.w1(32'h3b03e363),
	.w2(32'h3a0f0b3c),
	.w3(32'hb73e18bd),
	.w4(32'hba5fe3b0),
	.w5(32'hba3e0342),
	.w6(32'h3b40d654),
	.w7(32'h3add4fa0),
	.w8(32'hbab91ab8),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9114a07),
	.w1(32'h3a6ec337),
	.w2(32'h3a2f2b6d),
	.w3(32'hb961c2e9),
	.w4(32'hb8ac5d2f),
	.w5(32'h3ae460f2),
	.w6(32'hbaf7e082),
	.w7(32'hba20c7fc),
	.w8(32'h3ba5b51e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe54c7),
	.w1(32'h3c35d33e),
	.w2(32'h3c24b50e),
	.w3(32'h3a9b814d),
	.w4(32'h3b581201),
	.w5(32'hb9d7baed),
	.w6(32'h3be735de),
	.w7(32'h3c35203f),
	.w8(32'h3b1b4f83),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d759f),
	.w1(32'h38f6dec3),
	.w2(32'hbaf193c2),
	.w3(32'h3b13ed33),
	.w4(32'h3b2c36cd),
	.w5(32'hbab8db1b),
	.w6(32'h3ab90f35),
	.w7(32'h3aef579d),
	.w8(32'hbb257100),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9741a4),
	.w1(32'hbb0a19fc),
	.w2(32'hbb3da8e1),
	.w3(32'hbb55d964),
	.w4(32'hbb9d5554),
	.w5(32'h3a103aa0),
	.w6(32'hba77054e),
	.w7(32'h3a81e7af),
	.w8(32'h3b7569f1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b973e9e),
	.w1(32'h3bd8263d),
	.w2(32'h3bbf6348),
	.w3(32'h3b87d572),
	.w4(32'h3b8b55c9),
	.w5(32'hba23bc08),
	.w6(32'h3b32cdad),
	.w7(32'h3b6203bb),
	.w8(32'hbbd358d9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadec923),
	.w1(32'hbaf661cb),
	.w2(32'hba7af895),
	.w3(32'h3ad98269),
	.w4(32'h3aa3acfd),
	.w5(32'h37348652),
	.w6(32'hbbe61bce),
	.w7(32'hbb2dd599),
	.w8(32'h3af09c0f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83e8ca),
	.w1(32'h3ac8d712),
	.w2(32'hbb3c0d8a),
	.w3(32'h39da572c),
	.w4(32'hbb2b75b0),
	.w5(32'hba308c88),
	.w6(32'hb81b08db),
	.w7(32'hbafb4689),
	.w8(32'hba80ec6a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3921e0),
	.w1(32'h3b6ca10b),
	.w2(32'h3aedd978),
	.w3(32'hba1053fb),
	.w4(32'hba9fe358),
	.w5(32'h3b18277c),
	.w6(32'h3aa0af12),
	.w7(32'h3b43c625),
	.w8(32'h3aeac05c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80c92d),
	.w1(32'h3aaff673),
	.w2(32'h3b567a1c),
	.w3(32'h3b1c1353),
	.w4(32'h3b1cfc3a),
	.w5(32'hbb2529f8),
	.w6(32'h3aea9c2a),
	.w7(32'h3ba6c1a7),
	.w8(32'hbbce6f3f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccd28e),
	.w1(32'hbbcbdb78),
	.w2(32'hbb2c6903),
	.w3(32'hbb1a1262),
	.w4(32'hbb718452),
	.w5(32'hbac7e293),
	.w6(32'hbb823e3a),
	.w7(32'hbb5d50e8),
	.w8(32'hbba516ad),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb275384),
	.w1(32'hbb4d3b28),
	.w2(32'hbb49c461),
	.w3(32'hbaab75e0),
	.w4(32'hbae96229),
	.w5(32'hbbdc476a),
	.w6(32'hbb9eb11a),
	.w7(32'hbb7d6e89),
	.w8(32'hbbb774d1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94e553),
	.w1(32'hbb68690a),
	.w2(32'hbb8adbb2),
	.w3(32'hbbb1ebb1),
	.w4(32'hbbbe26f4),
	.w5(32'hba956888),
	.w6(32'hbbc52144),
	.w7(32'hbbc1a243),
	.w8(32'hbb6628d6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38afea4f),
	.w1(32'h3ba1e794),
	.w2(32'h3b48c53b),
	.w3(32'hbaa49d5a),
	.w4(32'hbb0271e0),
	.w5(32'hba8faa3f),
	.w6(32'hbb243171),
	.w7(32'hba3190bf),
	.w8(32'h3aa42a6e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948479b),
	.w1(32'h3b34c0e8),
	.w2(32'hbab45462),
	.w3(32'hbaf6a625),
	.w4(32'h399b03cc),
	.w5(32'h3b644222),
	.w6(32'h395c9d59),
	.w7(32'hbb273712),
	.w8(32'h3ba1465e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380e2299),
	.w1(32'hbb64fc07),
	.w2(32'h393b7873),
	.w3(32'h3b8ef375),
	.w4(32'h3b147ba6),
	.w5(32'hbb115527),
	.w6(32'h3bab6cb9),
	.w7(32'h3a635784),
	.w8(32'h3b42fa44),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b19641),
	.w1(32'hba58a912),
	.w2(32'h39c19aa6),
	.w3(32'hbaeac15b),
	.w4(32'h3a1b0a4a),
	.w5(32'h3b52fd6b),
	.w6(32'hbb102e9b),
	.w7(32'h3b77fe81),
	.w8(32'h3a2e3650),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4f3c1),
	.w1(32'h3c1d9ca7),
	.w2(32'h3bc9db01),
	.w3(32'h3bc56cfd),
	.w4(32'h3b357cf7),
	.w5(32'hbb2392aa),
	.w6(32'hbb57a1d1),
	.w7(32'hbb2649f0),
	.w8(32'hbad13bf9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39119c3e),
	.w1(32'hb9059c45),
	.w2(32'hbb33485b),
	.w3(32'hba87b09f),
	.w4(32'hba9b56c8),
	.w5(32'h3a431628),
	.w6(32'hb941530b),
	.w7(32'hbb618ab5),
	.w8(32'h3b83702d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92f2ac),
	.w1(32'h3b062382),
	.w2(32'h3b694705),
	.w3(32'h3b1f9040),
	.w4(32'h3a7146ea),
	.w5(32'hbae80f53),
	.w6(32'h3c089f78),
	.w7(32'h3be6e9f5),
	.w8(32'hbad1680f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54b0ef),
	.w1(32'h38305b02),
	.w2(32'hbb1df0aa),
	.w3(32'hbaceacfb),
	.w4(32'hbb152665),
	.w5(32'h3c1e9473),
	.w6(32'hbb46c46e),
	.w7(32'hbb8e96f3),
	.w8(32'h3c1e13ae),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule