module layer_8_featuremap_235(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9be9cd),
	.w1(32'hbab852b0),
	.w2(32'hbc179b60),
	.w3(32'hb92307e1),
	.w4(32'hbb986db6),
	.w5(32'hbb52c516),
	.w6(32'hbb8256eb),
	.w7(32'hbc3baa96),
	.w8(32'hba14ff6b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb869ac1),
	.w1(32'hbcb9f0c2),
	.w2(32'hbd0443b5),
	.w3(32'hbb953bcb),
	.w4(32'h3c4f5d70),
	.w5(32'h3c24599f),
	.w6(32'hbb96858e),
	.w7(32'hbc890ecd),
	.w8(32'h3bc19de4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8949b9),
	.w1(32'h3b7344c2),
	.w2(32'h3b0ac80a),
	.w3(32'h3cf66641),
	.w4(32'h3a93e615),
	.w5(32'h3b5c493e),
	.w6(32'h3bd25e59),
	.w7(32'h3a5f84bf),
	.w8(32'h3bb7ace9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad981de),
	.w1(32'hbad528d0),
	.w2(32'hb9a8f852),
	.w3(32'h3c15beee),
	.w4(32'h3b7cfe4f),
	.w5(32'h3ae7c302),
	.w6(32'hbb7c0086),
	.w7(32'hbb037415),
	.w8(32'hba1a04b6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3df124),
	.w1(32'hbce172a6),
	.w2(32'hbda0bfe7),
	.w3(32'h3a2a38d3),
	.w4(32'h3c501de2),
	.w5(32'hbcef001e),
	.w6(32'h3c01e411),
	.w7(32'hbcea5020),
	.w8(32'h3b8cf4b3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1221cd),
	.w1(32'hbbcb65c3),
	.w2(32'hbb4d67c7),
	.w3(32'h3c20a949),
	.w4(32'hbc0f6e56),
	.w5(32'h3aa47611),
	.w6(32'hbc02cf7d),
	.w7(32'hbb42fc53),
	.w8(32'hbad4e887),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ea1cd),
	.w1(32'h3c3d73a5),
	.w2(32'h3c84b28c),
	.w3(32'h3b278edb),
	.w4(32'hbb82928b),
	.w5(32'hb82f14ba),
	.w6(32'hba961f79),
	.w7(32'h3ba811e9),
	.w8(32'hbc12c7b2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36c55f),
	.w1(32'hbb7698b3),
	.w2(32'hbaf92a3b),
	.w3(32'hbc47552a),
	.w4(32'hbb7df549),
	.w5(32'h3b22721b),
	.w6(32'hbbb9db21),
	.w7(32'hbbfaa4c2),
	.w8(32'hbb963053),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e6790),
	.w1(32'hbcfb7a0e),
	.w2(32'hbd8d5e31),
	.w3(32'h3a906ac4),
	.w4(32'h3be7cb7a),
	.w5(32'hbca1ff59),
	.w6(32'h3aab21bd),
	.w7(32'hbd06528a),
	.w8(32'hbb7dac64),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf9c7f8),
	.w1(32'hbbfec26d),
	.w2(32'hbbf88a9b),
	.w3(32'h3c862e90),
	.w4(32'hbc6a6530),
	.w5(32'hbb9e206e),
	.w6(32'hbb9687da),
	.w7(32'hbbfcdf20),
	.w8(32'hbb64b006),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba24234),
	.w1(32'hbb9c4dd8),
	.w2(32'hbbe182cb),
	.w3(32'hbb7cfd9d),
	.w4(32'hba40a7e2),
	.w5(32'hbaa6a199),
	.w6(32'hbbfe5596),
	.w7(32'hbc3a40ad),
	.w8(32'hbc5a11bb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896cfb),
	.w1(32'hbaa66071),
	.w2(32'h399f7fc4),
	.w3(32'hbbb11305),
	.w4(32'hbbe2a633),
	.w5(32'hbb8b1cd3),
	.w6(32'hb95770ba),
	.w7(32'hbb5f7f7e),
	.w8(32'hbbd3f746),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc009f18),
	.w1(32'hbc3ad105),
	.w2(32'hbbaaddf0),
	.w3(32'hbc0a7b70),
	.w4(32'hbc3db493),
	.w5(32'hbb8396d8),
	.w6(32'hbbdabea6),
	.w7(32'hbbbe8bd1),
	.w8(32'hba9cbe82),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb108cb9),
	.w1(32'h3a9a4b19),
	.w2(32'h3aea1b92),
	.w3(32'hbc1460bc),
	.w4(32'hb9d5829a),
	.w5(32'hba5a981d),
	.w6(32'h3a1510cd),
	.w7(32'hbb95b817),
	.w8(32'h3b622ffb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89d1bd),
	.w1(32'h3d2d3d4d),
	.w2(32'h3dc76548),
	.w3(32'h3b9392ba),
	.w4(32'h3b4ee2cc),
	.w5(32'h3d4506a2),
	.w6(32'h3c180d1f),
	.w7(32'h3d21a983),
	.w8(32'h3c45b3cb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d742c1b),
	.w1(32'hbb5ef5ee),
	.w2(32'hbb58f38d),
	.w3(32'h3c93cd16),
	.w4(32'hba8b50c9),
	.w5(32'h3a75d313),
	.w6(32'hbb088ab8),
	.w7(32'h3aa521d5),
	.w8(32'h39450c8c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88efb8),
	.w1(32'hba47b07d),
	.w2(32'h3b3b8846),
	.w3(32'hbc20283a),
	.w4(32'h3bb51a75),
	.w5(32'hbc1c6979),
	.w6(32'hbb202707),
	.w7(32'h38b77b37),
	.w8(32'hbb6d21ac),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8ff7),
	.w1(32'hbbb86c13),
	.w2(32'hbbc622f5),
	.w3(32'h3ab70e25),
	.w4(32'hbb8d0018),
	.w5(32'hba84b1cf),
	.w6(32'hba566b33),
	.w7(32'hbb1f3890),
	.w8(32'hbb390902),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997205f),
	.w1(32'hbb9fb632),
	.w2(32'hbadd49d6),
	.w3(32'hbb506a41),
	.w4(32'hbc2b0b86),
	.w5(32'hbb401541),
	.w6(32'hbbf7c588),
	.w7(32'hbc159f8e),
	.w8(32'h39ef5065),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad39e70),
	.w1(32'h3c89fb3d),
	.w2(32'h3d1012a1),
	.w3(32'hbacf3e09),
	.w4(32'hbc7c2084),
	.w5(32'hba9403d0),
	.w6(32'hbc10d4c9),
	.w7(32'h3c016434),
	.w8(32'hbc5b2727),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c229e6f),
	.w1(32'hba581528),
	.w2(32'h3b3a2850),
	.w3(32'hbca43e8a),
	.w4(32'hbbb0ff18),
	.w5(32'hbb8e050d),
	.w6(32'hbac07f1b),
	.w7(32'hbc03eb58),
	.w8(32'hbb8051b6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b8314),
	.w1(32'hbb81c3b5),
	.w2(32'h3aaa1eca),
	.w3(32'h3b7c37b6),
	.w4(32'hba6f180d),
	.w5(32'hba1df332),
	.w6(32'hbbedea45),
	.w7(32'h3b24c94c),
	.w8(32'hbb8e5a2a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397efd7e),
	.w1(32'hba3a351a),
	.w2(32'hbb1d2a63),
	.w3(32'h3b366ab4),
	.w4(32'hba8ae5ef),
	.w5(32'hbbbb440f),
	.w6(32'h39ae9fdc),
	.w7(32'hbab65c65),
	.w8(32'hbb81a871),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa140ef),
	.w1(32'hbbedb2a9),
	.w2(32'hba2a2a9b),
	.w3(32'hbbcde6df),
	.w4(32'hbbb8063e),
	.w5(32'hbbe7eb80),
	.w6(32'hbb0af546),
	.w7(32'h3b195c2a),
	.w8(32'h3a024105),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09419f),
	.w1(32'h39856d8e),
	.w2(32'hbb0239ff),
	.w3(32'hbbb95887),
	.w4(32'hbc046971),
	.w5(32'hbc186de5),
	.w6(32'h3aa1be52),
	.w7(32'h3b2311d4),
	.w8(32'h3a0721ad),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6efab),
	.w1(32'hbc3025f0),
	.w2(32'hbc2c39cf),
	.w3(32'hbc06f63f),
	.w4(32'hbc45735b),
	.w5(32'hbba078a8),
	.w6(32'hbc20adb2),
	.w7(32'hbc183bba),
	.w8(32'hbbc853da),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d519f),
	.w1(32'hbbd60f72),
	.w2(32'hbb48ff52),
	.w3(32'hbc3a298d),
	.w4(32'hba51e212),
	.w5(32'h3925bd0c),
	.w6(32'hbc11f8a8),
	.w7(32'hbbd9fd33),
	.w8(32'hbbfb3825),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb946070),
	.w1(32'hbb837c39),
	.w2(32'hbba61beb),
	.w3(32'hbb9635b7),
	.w4(32'h3c028171),
	.w5(32'h3b66f3e8),
	.w6(32'hbc4b4c41),
	.w7(32'hbc0b19bf),
	.w8(32'hbb852c85),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61023c),
	.w1(32'hbc1715ed),
	.w2(32'h3a3361b5),
	.w3(32'h39e46642),
	.w4(32'hbbc1fdae),
	.w5(32'h3bb354ca),
	.w6(32'hbb86c439),
	.w7(32'hbbd3b6c1),
	.w8(32'h3a988f20),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46d20a),
	.w1(32'hbb459547),
	.w2(32'h3bfb4dad),
	.w3(32'h3c805601),
	.w4(32'hbc06536c),
	.w5(32'h3bab986b),
	.w6(32'hba158dbc),
	.w7(32'hbb9944a7),
	.w8(32'hbb180a4f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e757d),
	.w1(32'h3aa48a5b),
	.w2(32'hbb406fc4),
	.w3(32'h3ba4d24e),
	.w4(32'h3c03e066),
	.w5(32'h3bf9dbf2),
	.w6(32'h3a931ed4),
	.w7(32'hbb8e407c),
	.w8(32'hbb53d3ae),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402c27),
	.w1(32'hbbd28061),
	.w2(32'hbb0627b2),
	.w3(32'h3be3afe2),
	.w4(32'hba61fd5b),
	.w5(32'h3b52c68a),
	.w6(32'hbc10319a),
	.w7(32'hbc176bbb),
	.w8(32'hbb62a95d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2fffc),
	.w1(32'h3a151a61),
	.w2(32'hbc151668),
	.w3(32'h3be06db2),
	.w4(32'hb820ef36),
	.w5(32'hbab960fb),
	.w6(32'hbacad36a),
	.w7(32'hbb92bc3a),
	.w8(32'hbb450c56),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb846a9c),
	.w1(32'hbb48e1c3),
	.w2(32'hbb20341c),
	.w3(32'hbb2e29b6),
	.w4(32'h3b466302),
	.w5(32'h3b15c2b9),
	.w6(32'hbb67b81f),
	.w7(32'h3b3f1be1),
	.w8(32'hbb754eef),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58fe70),
	.w1(32'h3b55f2a6),
	.w2(32'h3c4145fb),
	.w3(32'hbbdae741),
	.w4(32'h3b3902d5),
	.w5(32'h3b5268a1),
	.w6(32'hbb569917),
	.w7(32'hbb4a6aa9),
	.w8(32'hba40e749),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60eb25),
	.w1(32'h3b7f007b),
	.w2(32'hba46b852),
	.w3(32'hbaddf029),
	.w4(32'hbae0235f),
	.w5(32'hbb41ad8b),
	.w6(32'h3b8600f2),
	.w7(32'h38c7e802),
	.w8(32'hbab47734),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dc811),
	.w1(32'h3b065cd8),
	.w2(32'hbae7a4f5),
	.w3(32'hb9e37ea7),
	.w4(32'h3afaef71),
	.w5(32'hba1c7bba),
	.w6(32'hba227deb),
	.w7(32'hbb5873c1),
	.w8(32'hbb743845),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38959e3a),
	.w1(32'h3b7cacb5),
	.w2(32'h3d0a38a5),
	.w3(32'h3a94a23b),
	.w4(32'h3b43d3db),
	.w5(32'h3cd4dc27),
	.w6(32'h3b7aeaa3),
	.w7(32'h3c194de7),
	.w8(32'h3c33f23f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce78d59),
	.w1(32'h39ecd637),
	.w2(32'h3b260628),
	.w3(32'h3ca8497e),
	.w4(32'hba4eba72),
	.w5(32'hba33a1c5),
	.w6(32'hb9cb397a),
	.w7(32'hbb11a340),
	.w8(32'hbb86943b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd61b42),
	.w1(32'hbb4f5589),
	.w2(32'h39b96c5d),
	.w3(32'hbae6e39c),
	.w4(32'hbb843eed),
	.w5(32'hbb781786),
	.w6(32'hbb0b37ca),
	.w7(32'hbb55556c),
	.w8(32'hbb3f003f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038cda),
	.w1(32'hbb25d7c3),
	.w2(32'h3c0d07c9),
	.w3(32'hbc2d6594),
	.w4(32'hbb4e8e62),
	.w5(32'h3c128f26),
	.w6(32'hbbb78ad6),
	.w7(32'h3ab0ee1c),
	.w8(32'hbb938c41),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3815ecef),
	.w1(32'h3bae1cb0),
	.w2(32'h3b7a6dc6),
	.w3(32'hbacf8001),
	.w4(32'h3c0119be),
	.w5(32'h3bf77f32),
	.w6(32'hb903aabf),
	.w7(32'hba84544c),
	.w8(32'hbc40ec02),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d47ef),
	.w1(32'hbc02fcda),
	.w2(32'hbc40686f),
	.w3(32'hbc1469f6),
	.w4(32'hbb99dcf6),
	.w5(32'hbbbfdf11),
	.w6(32'hbb9c8ca7),
	.w7(32'hbc0eaec1),
	.w8(32'hbc134376),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e2591),
	.w1(32'hbb8a1ae8),
	.w2(32'hbbb3724f),
	.w3(32'hbbb67cde),
	.w4(32'hbb99f439),
	.w5(32'hbaa77cb1),
	.w6(32'hbb914fa6),
	.w7(32'hba3efcfd),
	.w8(32'hba5ada8d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08efd2),
	.w1(32'hbb7845ed),
	.w2(32'h3b51b6f4),
	.w3(32'hbbe8b0b8),
	.w4(32'hbc15fecf),
	.w5(32'h3a07f6f1),
	.w6(32'hbb16e627),
	.w7(32'hbad5bc48),
	.w8(32'h3b84771f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb3fdd),
	.w1(32'h3bb6d1bb),
	.w2(32'h3d86d62e),
	.w3(32'h3b707a9f),
	.w4(32'hbca1aa5e),
	.w5(32'h3d201758),
	.w6(32'hbd06573a),
	.w7(32'h3c5e3e07),
	.w8(32'hbcbd471c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3061c),
	.w1(32'hba94d99f),
	.w2(32'hb9f08bc3),
	.w3(32'hbb351604),
	.w4(32'hbb465f20),
	.w5(32'hbb17b7a2),
	.w6(32'h3ace556a),
	.w7(32'h3ac15948),
	.w8(32'hb965ed39),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04cb62),
	.w1(32'hbad83808),
	.w2(32'hbbaebc90),
	.w3(32'hbb5f5f88),
	.w4(32'hbbaedd4a),
	.w5(32'h3b7ae6e2),
	.w6(32'hbba7f1f0),
	.w7(32'hbbaefca0),
	.w8(32'hbb169174),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1c1e6),
	.w1(32'hbb7280c5),
	.w2(32'hba4f2c2a),
	.w3(32'hbb62b482),
	.w4(32'h3b9cc980),
	.w5(32'hb8bb27ee),
	.w6(32'hbb27f219),
	.w7(32'hbb9245ae),
	.w8(32'hbac9cb9b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987c6bc),
	.w1(32'hbb33be5c),
	.w2(32'hbad475f7),
	.w3(32'h3b5bd59e),
	.w4(32'h3a7f6dd4),
	.w5(32'h3681010a),
	.w6(32'hbaf42a53),
	.w7(32'hbb84de52),
	.w8(32'h3ab6444a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e75cc),
	.w1(32'hbb70a435),
	.w2(32'h3d3ab472),
	.w3(32'hbb477d28),
	.w4(32'hbb293d44),
	.w5(32'h3cce3dc2),
	.w6(32'hbbb6a6fd),
	.w7(32'h3c23190f),
	.w8(32'hba80fdcb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c333ffb),
	.w1(32'h3b92891b),
	.w2(32'h3a941e1f),
	.w3(32'h3af4e343),
	.w4(32'h3b0347d7),
	.w5(32'h3b910566),
	.w6(32'h3b28ad6b),
	.w7(32'hb8dada69),
	.w8(32'hbac9e8ff),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a800580),
	.w1(32'hbc7a8930),
	.w2(32'h3ce0cd68),
	.w3(32'h3a4fe3ec),
	.w4(32'h3ba0eb01),
	.w5(32'h3d4103c8),
	.w6(32'hbc707b23),
	.w7(32'hb925ee0a),
	.w8(32'h3bd012fa),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02b10d),
	.w1(32'hbb9bc46c),
	.w2(32'hbba9d544),
	.w3(32'h3d1c3287),
	.w4(32'hbc13e89d),
	.w5(32'hbb1b4be8),
	.w6(32'hbc17a9b0),
	.w7(32'hbbba5398),
	.w8(32'h3aa385bc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fd1e4),
	.w1(32'hbb696a48),
	.w2(32'hbb22ef0a),
	.w3(32'h3b506b7c),
	.w4(32'hbc032e30),
	.w5(32'h39b61d0e),
	.w6(32'h3aa16206),
	.w7(32'h387e7b56),
	.w8(32'hbaabf8cc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c7588),
	.w1(32'hbb697058),
	.w2(32'h3adc3ffe),
	.w3(32'hbb246ade),
	.w4(32'h3a40bbd9),
	.w5(32'hb732a323),
	.w6(32'hbb77a646),
	.w7(32'hbb24565a),
	.w8(32'hb794a8e1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d0e15),
	.w1(32'hbbba9a3b),
	.w2(32'hbc185768),
	.w3(32'hbb1255d0),
	.w4(32'hbb03fb94),
	.w5(32'hbc4e3f4b),
	.w6(32'hbae3f93a),
	.w7(32'hbbaa0b9a),
	.w8(32'hbb9ab8ba),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1afba2),
	.w1(32'h39fc3dbf),
	.w2(32'h3a56c458),
	.w3(32'hbbb5f98a),
	.w4(32'h3aed4217),
	.w5(32'h3bc6bc1d),
	.w6(32'hbb12c497),
	.w7(32'hbb2a78c5),
	.w8(32'hbbd501fd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5aa3b2),
	.w1(32'h3bee5aca),
	.w2(32'h3ca9fc0b),
	.w3(32'hba5651f4),
	.w4(32'h3bd02c17),
	.w5(32'h3cb2ec45),
	.w6(32'hbab354d6),
	.w7(32'h3bfe2fda),
	.w8(32'h3baf08c7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e59f9),
	.w1(32'hbaaf8384),
	.w2(32'h3a127975),
	.w3(32'h3c577a61),
	.w4(32'hbaaed8c3),
	.w5(32'hbaf45f41),
	.w6(32'hbbcdead8),
	.w7(32'hbac92255),
	.w8(32'h3a69892f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ae1d1),
	.w1(32'hbbf4adea),
	.w2(32'h3a81c9df),
	.w3(32'hbb0e88a0),
	.w4(32'hba9b4876),
	.w5(32'h3b40fb2f),
	.w6(32'h3b0682ee),
	.w7(32'hba540d97),
	.w8(32'hba564b9d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae16103),
	.w1(32'hb82a2127),
	.w2(32'h3c1651df),
	.w3(32'h3ae6edc7),
	.w4(32'h39ab3f7d),
	.w5(32'h3c22e090),
	.w6(32'hbb72f490),
	.w7(32'hb9ba0a2b),
	.w8(32'hbbe48d04),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c262d35),
	.w1(32'hbc6e5972),
	.w2(32'hbca8f42d),
	.w3(32'h3c3efb5c),
	.w4(32'hbc30710d),
	.w5(32'hbc96ef78),
	.w6(32'hbc880fa8),
	.w7(32'hbcde9190),
	.w8(32'hbcd45708),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f21b9),
	.w1(32'hbb9a8298),
	.w2(32'hbb3a61ee),
	.w3(32'hbc51709f),
	.w4(32'hbb2d7af9),
	.w5(32'hba6edca1),
	.w6(32'hb9ed335d),
	.w7(32'hba84f009),
	.w8(32'hbbd0420d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f56e6),
	.w1(32'h3cc31ae5),
	.w2(32'h3d8fefaf),
	.w3(32'hbba8d0bb),
	.w4(32'h3c50b835),
	.w5(32'h3d563264),
	.w6(32'h3b978528),
	.w7(32'h3cd71206),
	.w8(32'h3c75bd05),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d54d3c4),
	.w1(32'hbbb6d90b),
	.w2(32'hba1ea84b),
	.w3(32'h3d0527b0),
	.w4(32'hbba6aabb),
	.w5(32'hbbdd1f41),
	.w6(32'hbae374ac),
	.w7(32'hb9a8cc8b),
	.w8(32'hbbbe89e5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb073f1b),
	.w1(32'hb79bba6d),
	.w2(32'hbabd9152),
	.w3(32'hbb90ece0),
	.w4(32'hba6eed15),
	.w5(32'h3a8bbe5e),
	.w6(32'hbac56144),
	.w7(32'h3abe69c4),
	.w8(32'h3b933b5a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc2857),
	.w1(32'h3b35691a),
	.w2(32'hba173862),
	.w3(32'h3b5cfd0a),
	.w4(32'hbb0e2ec8),
	.w5(32'hbbd70c14),
	.w6(32'h3b2430ba),
	.w7(32'hb924150c),
	.w8(32'h3b58b6a8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5e348),
	.w1(32'hbacb8d0e),
	.w2(32'h3b047e00),
	.w3(32'h3aba0c80),
	.w4(32'hbbd10579),
	.w5(32'h3b214f82),
	.w6(32'hbb052fd6),
	.w7(32'hba73cfc6),
	.w8(32'hbb3c9e14),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43cb77),
	.w1(32'h3af0338d),
	.w2(32'h3b79c6a2),
	.w3(32'hba75ae0b),
	.w4(32'h3bf66200),
	.w5(32'h3ac41b42),
	.w6(32'h380ed816),
	.w7(32'hbb9fd9d8),
	.w8(32'hbb5692b9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e9721),
	.w1(32'hbba17b2c),
	.w2(32'h3a210008),
	.w3(32'h3aa6fdcc),
	.w4(32'hbc28ae5b),
	.w5(32'h3b1a94f0),
	.w6(32'hbb43dae7),
	.w7(32'h399a379b),
	.w8(32'h3b6f4d30),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c340a44),
	.w1(32'hb9c188c9),
	.w2(32'hbb63f47c),
	.w3(32'h3c31764a),
	.w4(32'hbbc2761b),
	.w5(32'hbb3b3379),
	.w6(32'hbb14ac90),
	.w7(32'hbaba5d65),
	.w8(32'hbb9c32c6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11c22a),
	.w1(32'h3aff2255),
	.w2(32'hba87cf94),
	.w3(32'h3b255986),
	.w4(32'hbbcb56b6),
	.w5(32'hbb636007),
	.w6(32'hbaddc0f4),
	.w7(32'hb8e42f71),
	.w8(32'hbbf94e9f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee2519),
	.w1(32'hbb818821),
	.w2(32'hb9007fa2),
	.w3(32'hbbd3d2ff),
	.w4(32'hbb91acde),
	.w5(32'hb9e3dc90),
	.w6(32'hbb7bae3d),
	.w7(32'h3a76d78d),
	.w8(32'hb970c8f8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab94c09),
	.w1(32'h3c1a3c8e),
	.w2(32'h3bf39f4c),
	.w3(32'hbb0e541f),
	.w4(32'h3bb9a2ff),
	.w5(32'h3b36c762),
	.w6(32'hbb9ea310),
	.w7(32'h3a7b196a),
	.w8(32'hba9a136f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb5049),
	.w1(32'hbba0d123),
	.w2(32'h3bbe98ac),
	.w3(32'hbb99bd7c),
	.w4(32'hbbce62cf),
	.w5(32'h3b184607),
	.w6(32'hbb30a051),
	.w7(32'h39570097),
	.w8(32'h3b304fef),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1faa0c),
	.w1(32'hbbc0179f),
	.w2(32'hbb81ed0a),
	.w3(32'h3a405306),
	.w4(32'hba8215a0),
	.w5(32'hbbc5802e),
	.w6(32'hba6d2c01),
	.w7(32'hbb392222),
	.w8(32'hbb2c266a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba10924),
	.w1(32'h3a8d89c6),
	.w2(32'hb9963959),
	.w3(32'hb9af3eff),
	.w4(32'h3aad28f9),
	.w5(32'hbb016d24),
	.w6(32'h3a9c1f74),
	.w7(32'hba2ca386),
	.w8(32'hbaad6396),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922acda),
	.w1(32'hbba37779),
	.w2(32'hbb184036),
	.w3(32'hbb21d4f8),
	.w4(32'hbb9e852a),
	.w5(32'h39b49ba4),
	.w6(32'hb9eb8027),
	.w7(32'h3b7f7c21),
	.w8(32'hbaac09e5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb021cee),
	.w1(32'hba977411),
	.w2(32'hbb6379a4),
	.w3(32'hbb1bf801),
	.w4(32'h3b1a0111),
	.w5(32'h3b562212),
	.w6(32'hbaf0ead9),
	.w7(32'hbbe7a672),
	.w8(32'h3ae1127c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddd5f1),
	.w1(32'hb90cde9b),
	.w2(32'h3b50f501),
	.w3(32'hbb59cc58),
	.w4(32'hb9b6acda),
	.w5(32'h3a16dfb5),
	.w6(32'h3a7bc1fe),
	.w7(32'h3b5d2f25),
	.w8(32'h3b47769f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b248056),
	.w1(32'hba3e6587),
	.w2(32'h3a1bebeb),
	.w3(32'h39e5b60c),
	.w4(32'h3ad5af9a),
	.w5(32'hba57e322),
	.w6(32'h398d4b44),
	.w7(32'hbb635603),
	.w8(32'hb8183a2e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d14353),
	.w1(32'h3a026ea0),
	.w2(32'hbabe6ab7),
	.w3(32'h3a5b469b),
	.w4(32'h3a48b758),
	.w5(32'hbab7ace2),
	.w6(32'hbae5e3b9),
	.w7(32'hbbbb70ba),
	.w8(32'h39e6a9ed),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6548ba),
	.w1(32'hbb46d844),
	.w2(32'hbb56648a),
	.w3(32'h3ad23cfb),
	.w4(32'hbb7a0b2d),
	.w5(32'hbb359e72),
	.w6(32'hbad2a7bf),
	.w7(32'h3a87f73c),
	.w8(32'hbb80d532),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72c4a5),
	.w1(32'h3b589faa),
	.w2(32'h3ad8b4d2),
	.w3(32'h3b7cc372),
	.w4(32'h3aa3d389),
	.w5(32'hb9f2eb6b),
	.w6(32'h3b8ad2c1),
	.w7(32'hbb23495f),
	.w8(32'hbb647512),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf30f4),
	.w1(32'h3b57a10e),
	.w2(32'h3c0307cc),
	.w3(32'h3a237e6d),
	.w4(32'h3b7a2e5c),
	.w5(32'h3c0c669f),
	.w6(32'hbb7f4a71),
	.w7(32'hbad8a2fd),
	.w8(32'h3a8601c0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bc37b),
	.w1(32'hbb193d67),
	.w2(32'hba917606),
	.w3(32'h3c00b814),
	.w4(32'hbb5f3b53),
	.w5(32'h3a926c5d),
	.w6(32'h3b2c0d79),
	.w7(32'h3b314e1b),
	.w8(32'hb90790cf),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb802a3e),
	.w1(32'hba94168a),
	.w2(32'h3ace652f),
	.w3(32'hbad0f9f7),
	.w4(32'hbbeab6e3),
	.w5(32'hbbec020d),
	.w6(32'h3b511c40),
	.w7(32'hb5785ece),
	.w8(32'h3af4ea9b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58dd72),
	.w1(32'h3ad49911),
	.w2(32'h3b9eba6a),
	.w3(32'hbbf9b510),
	.w4(32'hbbafdb53),
	.w5(32'hbbcb69f8),
	.w6(32'hb979d3c9),
	.w7(32'hbb04cd3e),
	.w8(32'h3847d935),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75a41a),
	.w1(32'h3b1cb06e),
	.w2(32'hbb4574f3),
	.w3(32'hbba7d4d1),
	.w4(32'h3b83f6c2),
	.w5(32'h3b669187),
	.w6(32'h3b21bca0),
	.w7(32'hbb2ab506),
	.w8(32'hb927a30a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fe54e),
	.w1(32'hbae5ffa7),
	.w2(32'hbb4f779f),
	.w3(32'hbb08a5c8),
	.w4(32'hba42f370),
	.w5(32'hbb440e4f),
	.w6(32'hbbc63305),
	.w7(32'hbb69b79f),
	.w8(32'hbb959a88),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf247cf),
	.w1(32'hbbe93ff0),
	.w2(32'hbada2629),
	.w3(32'hbb8b53aa),
	.w4(32'hbb357016),
	.w5(32'hbb13a104),
	.w6(32'hbaf68fae),
	.w7(32'hbb1d44a2),
	.w8(32'hbb0918e7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11ea6d),
	.w1(32'h3bd67607),
	.w2(32'hbb484f97),
	.w3(32'h39ae4b5f),
	.w4(32'h3c4343eb),
	.w5(32'h3bc863f6),
	.w6(32'h3c0d64f1),
	.w7(32'h3babad98),
	.w8(32'h3c0fcdc6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf0fe6),
	.w1(32'hbc4638e4),
	.w2(32'hbcc9ab0e),
	.w3(32'h3c32daff),
	.w4(32'h3bbf4564),
	.w5(32'hbb87d3b1),
	.w6(32'hbb32cb08),
	.w7(32'hbc42fd6e),
	.w8(32'hbb350612),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27e1bd),
	.w1(32'hbb9005fe),
	.w2(32'hbae855f3),
	.w3(32'h3bb83bb3),
	.w4(32'hba5cb7f7),
	.w5(32'hbb891848),
	.w6(32'hbbc2a86d),
	.w7(32'h3a9076c5),
	.w8(32'h3a010de7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37c511),
	.w1(32'h3a2d7d4e),
	.w2(32'hbb09f07b),
	.w3(32'h3b6aeeee),
	.w4(32'h3b137912),
	.w5(32'hbaaf39fa),
	.w6(32'hb79d9da6),
	.w7(32'hbb08ff1b),
	.w8(32'h3a72a904),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49a69e),
	.w1(32'h39b99c88),
	.w2(32'hbbcb2c7d),
	.w3(32'h3ad270ef),
	.w4(32'hba34fdea),
	.w5(32'h39ec6780),
	.w6(32'h3b7694cf),
	.w7(32'hb9a3fffa),
	.w8(32'hbb3b338f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6d742),
	.w1(32'h3a2a4725),
	.w2(32'h3baabdb6),
	.w3(32'h3b82e67f),
	.w4(32'hbb752c84),
	.w5(32'h3bac2dd8),
	.w6(32'hbb769417),
	.w7(32'h3ba6b5ce),
	.w8(32'h3ac320f5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb424e03),
	.w1(32'hbbb45346),
	.w2(32'hbbafb6b0),
	.w3(32'hbb29b30c),
	.w4(32'hbbca80d7),
	.w5(32'h39cd2d50),
	.w6(32'h39933032),
	.w7(32'hbb03e1e5),
	.w8(32'h3b9ce320),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8de908b),
	.w1(32'hb9b04f8d),
	.w2(32'hbb6e5833),
	.w3(32'h383c7ed8),
	.w4(32'h3b9333a8),
	.w5(32'hbb061b48),
	.w6(32'h3a41f3a8),
	.w7(32'hbafc5a71),
	.w8(32'hbac74dca),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6807bd),
	.w1(32'hbbf63eb1),
	.w2(32'hba5167ec),
	.w3(32'hba2b1baf),
	.w4(32'hbbda7e37),
	.w5(32'h3a1be233),
	.w6(32'hb9fa9240),
	.w7(32'h3b1d4a52),
	.w8(32'h3bac0851),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7652ba),
	.w1(32'hbc046f7c),
	.w2(32'hbbdce164),
	.w3(32'h3b94d809),
	.w4(32'hbc011251),
	.w5(32'h3a7a0f5e),
	.w6(32'hbbd1c8a6),
	.w7(32'hbbbb33cd),
	.w8(32'hbc013525),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d521),
	.w1(32'h3ad188e6),
	.w2(32'hbac33875),
	.w3(32'hbbce008b),
	.w4(32'hbb84ce96),
	.w5(32'hbba8a24e),
	.w6(32'h3840d7c3),
	.w7(32'hb8d2170b),
	.w8(32'hbbae9b9f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb060582),
	.w1(32'hbbb79d85),
	.w2(32'hbc28d87d),
	.w3(32'h38000043),
	.w4(32'h3a60bf51),
	.w5(32'hbc3dbefd),
	.w6(32'hbbbc3abc),
	.w7(32'hbbfd5e1d),
	.w8(32'hbc028074),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6e58e),
	.w1(32'hbb3b82ed),
	.w2(32'hbc20114a),
	.w3(32'hbbdeb278),
	.w4(32'hbb5ed4e0),
	.w5(32'hbbe1f3e7),
	.w6(32'hbafb4cc1),
	.w7(32'hbc04e553),
	.w8(32'hbc00e9a0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b821c),
	.w1(32'h3d02cc13),
	.w2(32'h3e06c247),
	.w3(32'hbbbdf309),
	.w4(32'hbba425e2),
	.w5(32'h3daeed97),
	.w6(32'hbc8a4bea),
	.w7(32'h3d261ead),
	.w8(32'hbb5b3672),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d956524),
	.w1(32'hb9a5267e),
	.w2(32'h39d0b4b4),
	.w3(32'h3cc29fb2),
	.w4(32'h3a7cb566),
	.w5(32'hbb8febe1),
	.w6(32'hbb01f9d4),
	.w7(32'hbab9ea95),
	.w8(32'hbaf7dbfa),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32bb03),
	.w1(32'hbace7ddf),
	.w2(32'hb829b51f),
	.w3(32'hbbda4d88),
	.w4(32'hbb5e80a1),
	.w5(32'hbba04acf),
	.w6(32'h3a2cf1db),
	.w7(32'hbb5f7305),
	.w8(32'hbb87435e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a296e),
	.w1(32'h3a83ea68),
	.w2(32'h3b21a903),
	.w3(32'hbb24084d),
	.w4(32'h3bcd62cc),
	.w5(32'h3b9ed363),
	.w6(32'h3ba819c3),
	.w7(32'h3bc767fb),
	.w8(32'h3b5e1656),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad61177),
	.w1(32'hbc959784),
	.w2(32'hbcb3e2b1),
	.w3(32'h3b93dff2),
	.w4(32'h3b7bbef8),
	.w5(32'h3b2e2e3f),
	.w6(32'hbba425bb),
	.w7(32'hbc69add1),
	.w8(32'h3a93aed9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85513e),
	.w1(32'h3b2855f4),
	.w2(32'h38268264),
	.w3(32'h3c6600ba),
	.w4(32'hbbcaa3a3),
	.w5(32'hbb1bf8ee),
	.w6(32'h3ac4a3cc),
	.w7(32'h3a42816e),
	.w8(32'h3b6535e2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a37cdd),
	.w1(32'h3ccf5cc2),
	.w2(32'h3d1f97e5),
	.w3(32'h3acf0fc5),
	.w4(32'h3ca1d46f),
	.w5(32'h3d06c4fd),
	.w6(32'h3c7f9f08),
	.w7(32'h3cd2e1df),
	.w8(32'h3c8c7842),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cee2c5a),
	.w1(32'hbbf5f147),
	.w2(32'h3bdb0d58),
	.w3(32'h3cb83a96),
	.w4(32'hbb16c905),
	.w5(32'h3c5fe5e6),
	.w6(32'hbb96d851),
	.w7(32'hbaf0399a),
	.w8(32'h3b283ea3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b856586),
	.w1(32'hbb4265af),
	.w2(32'hbbbd3ba6),
	.w3(32'h3ab8a0f9),
	.w4(32'hbb121dc1),
	.w5(32'hbb82f032),
	.w6(32'hb8e230bb),
	.w7(32'hbb6cfaf6),
	.w8(32'hb962ef30),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c4a7c),
	.w1(32'h3ad39596),
	.w2(32'h3a967c55),
	.w3(32'hbba2954d),
	.w4(32'hbbb7e983),
	.w5(32'hbae861c7),
	.w6(32'hba5bf4f1),
	.w7(32'h39d22af6),
	.w8(32'hbb7d3a54),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb194092),
	.w1(32'hbc04d430),
	.w2(32'h3b1685a0),
	.w3(32'hbbc8b2e8),
	.w4(32'h3bbdb4ca),
	.w5(32'h3c7aa74e),
	.w6(32'hbb91bc34),
	.w7(32'hbba4f874),
	.w8(32'h3b9b0635),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c388248),
	.w1(32'hbb8bd9be),
	.w2(32'h3bf552a6),
	.w3(32'h3c8d8a7f),
	.w4(32'hbbe805d1),
	.w5(32'h3b8f7750),
	.w6(32'hbb8589af),
	.w7(32'h3b10e0ad),
	.w8(32'hb9d66f02),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75424c),
	.w1(32'hbc267b04),
	.w2(32'hb8967f5e),
	.w3(32'h37a92134),
	.w4(32'hba55c547),
	.w5(32'h3bb8e4a4),
	.w6(32'hbbc3f86d),
	.w7(32'hbbc40973),
	.w8(32'hbaa99022),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0864),
	.w1(32'hbb5979b0),
	.w2(32'hbb5655da),
	.w3(32'h3c0ae02b),
	.w4(32'hbb0ff80f),
	.w5(32'h3b09dd75),
	.w6(32'hbb83d0e0),
	.w7(32'h3a83f9a9),
	.w8(32'h3bc1ac09),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb875b2f),
	.w1(32'h3bafda92),
	.w2(32'h3b10ddd3),
	.w3(32'h3a08427d),
	.w4(32'h3b1bba33),
	.w5(32'h38ecde19),
	.w6(32'hbb5e954f),
	.w7(32'h3a3652e5),
	.w8(32'hb992a0b3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2d0bd),
	.w1(32'h3a1d3610),
	.w2(32'hbbc7fa92),
	.w3(32'hbaed58ba),
	.w4(32'hbae93c39),
	.w5(32'h3b6e9baf),
	.w6(32'hbb706e80),
	.w7(32'hbbfd62cd),
	.w8(32'h3bb4e8a9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09a501),
	.w1(32'h3abc05f9),
	.w2(32'h3bc3bdf9),
	.w3(32'hbbc5872d),
	.w4(32'h3b0ff341),
	.w5(32'h3b1c5676),
	.w6(32'h3a9eb647),
	.w7(32'hbb0e8173),
	.w8(32'h3b01f92e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a438d),
	.w1(32'hbca246be),
	.w2(32'hbd298058),
	.w3(32'h3b72f124),
	.w4(32'h3bc26266),
	.w5(32'hbc193784),
	.w6(32'hbb8e3ab8),
	.w7(32'hbc9b3f27),
	.w8(32'hbb30721f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ca40a),
	.w1(32'hbabb462f),
	.w2(32'h3b42e9e7),
	.w3(32'h3bf5114c),
	.w4(32'h3b1d9e73),
	.w5(32'h3bcedffa),
	.w6(32'hbba460fd),
	.w7(32'hbbc9ea3d),
	.w8(32'hbb17fb6c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82b226),
	.w1(32'hbbbad5ca),
	.w2(32'hbb921982),
	.w3(32'h3c0feb76),
	.w4(32'hbbf7d8f7),
	.w5(32'hbc15ff14),
	.w6(32'hbb307a7b),
	.w7(32'hb9cd3dd5),
	.w8(32'hbb11b147),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfe22d),
	.w1(32'hba9af1c4),
	.w2(32'hb9f4558c),
	.w3(32'hbc06de97),
	.w4(32'hbaf505d1),
	.w5(32'hbbcfbfa1),
	.w6(32'hbb8f0a89),
	.w7(32'hbba7a6dd),
	.w8(32'hba9290a1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a75cc),
	.w1(32'h38afbc58),
	.w2(32'h3c10026e),
	.w3(32'hbac24108),
	.w4(32'hbb3c196b),
	.w5(32'h3a0afa31),
	.w6(32'hbb86565d),
	.w7(32'hbaaabf98),
	.w8(32'hbb4e6664),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91459b),
	.w1(32'h3b241de8),
	.w2(32'hbbe4131c),
	.w3(32'hbb1f9726),
	.w4(32'h3b6abd23),
	.w5(32'hbbac5b98),
	.w6(32'h3c0a04b5),
	.w7(32'h3a3aa297),
	.w8(32'h3b735e51),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule