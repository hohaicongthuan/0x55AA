module layer_8_featuremap_71(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87c6410),
	.w1(32'h37d9bc95),
	.w2(32'h39298138),
	.w3(32'h37d3d794),
	.w4(32'h395c42dd),
	.w5(32'h39ca311d),
	.w6(32'hb91e1fc1),
	.w7(32'hb7561277),
	.w8(32'hb82f2448),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb762ffa7),
	.w1(32'hb84565b8),
	.w2(32'hb8ddf787),
	.w3(32'h387a9384),
	.w4(32'hb7cdd5aa),
	.w5(32'hb88dd2a1),
	.w6(32'h36123591),
	.w7(32'hb8569020),
	.w8(32'hb88c3f5a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88604d8),
	.w1(32'hb8855996),
	.w2(32'hb89aee5a),
	.w3(32'h36825f26),
	.w4(32'hb843eea2),
	.w5(32'hb89a9977),
	.w6(32'hb4bb9ca3),
	.w7(32'hb85b219a),
	.w8(32'hb8d9a235),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c407a),
	.w1(32'h3869dac0),
	.w2(32'h3973f891),
	.w3(32'h379f1b11),
	.w4(32'h396dcb6e),
	.w5(32'h394eebb1),
	.w6(32'h391ca12a),
	.w7(32'h38e98c06),
	.w8(32'h3839208e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bc6452),
	.w1(32'h383044b4),
	.w2(32'h3863bc60),
	.w3(32'h3887c90c),
	.w4(32'h3855a2ac),
	.w5(32'h389e0188),
	.w6(32'h37953462),
	.w7(32'h37e8c086),
	.w8(32'h38868ec2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e5951a),
	.w1(32'hb8ae8913),
	.w2(32'hb800d23b),
	.w3(32'h37ccaffd),
	.w4(32'h34aec154),
	.w5(32'hb7a72afe),
	.w6(32'h39479b53),
	.w7(32'h3880c800),
	.w8(32'h398a47b0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a1acc9),
	.w1(32'h369baf5a),
	.w2(32'h368a2f3c),
	.w3(32'h363b58eb),
	.w4(32'h3688db7a),
	.w5(32'h36554ca9),
	.w6(32'h361bfeea),
	.w7(32'h36810b1e),
	.w8(32'h363fbf54),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84cf157),
	.w1(32'hb7ea983b),
	.w2(32'hb8d0dcd8),
	.w3(32'hb7c204c2),
	.w4(32'h38420293),
	.w5(32'h38226331),
	.w6(32'h386048a7),
	.w7(32'h385ccccb),
	.w8(32'h38615fe2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e96f67),
	.w1(32'h36b2b165),
	.w2(32'h3600ee7a),
	.w3(32'hb71782d1),
	.w4(32'hb7cd575c),
	.w5(32'hb7824a15),
	.w6(32'hb59fa8cb),
	.w7(32'hb6215781),
	.w8(32'hb7cc6209),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ff8ce),
	.w1(32'hb90cf65b),
	.w2(32'hb9042a83),
	.w3(32'hb5478664),
	.w4(32'h3877e728),
	.w5(32'h3953fe12),
	.w6(32'hb95f4e2c),
	.w7(32'hb9408d52),
	.w8(32'hb9075bc3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8457a84),
	.w1(32'h3880e81c),
	.w2(32'h39804f69),
	.w3(32'h3864eb10),
	.w4(32'h3942dde9),
	.w5(32'h39bba07a),
	.w6(32'h389c0856),
	.w7(32'h391f0b56),
	.w8(32'h392c8352),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955fe65),
	.w1(32'hb8af5cf6),
	.w2(32'h383603e1),
	.w3(32'hb8323fac),
	.w4(32'h3898dc21),
	.w5(32'h3961774d),
	.w6(32'hb93f9a02),
	.w7(32'hb8c1b8b0),
	.w8(32'h37e87354),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89672d7),
	.w1(32'hb7c4fcc9),
	.w2(32'hb6d9ee0c),
	.w3(32'h37c116c5),
	.w4(32'h37838f70),
	.w5(32'h370e5c76),
	.w6(32'hb842dd05),
	.w7(32'hb8c0b650),
	.w8(32'hb8bffad9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373c9382),
	.w1(32'h37452185),
	.w2(32'h3739a0b7),
	.w3(32'h37001f5d),
	.w4(32'h37594fbe),
	.w5(32'h3731ea2a),
	.w6(32'h36efee65),
	.w7(32'h371f32ef),
	.w8(32'h36ff4867),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d7dba9),
	.w1(32'h362b81ed),
	.w2(32'h35f83348),
	.w3(32'h356f6fb6),
	.w4(32'h3600ed8d),
	.w5(32'h35a41220),
	.w6(32'h360e9cd4),
	.w7(32'h362139df),
	.w8(32'h3606b124),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3738f378),
	.w1(32'h3741ed34),
	.w2(32'h36dab00b),
	.w3(32'h3773ed02),
	.w4(32'h37573a18),
	.w5(32'h37420ae1),
	.w6(32'h375f2e84),
	.w7(32'h374394c3),
	.w8(32'h37311180),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389efdb3),
	.w1(32'h3851cdbf),
	.w2(32'h37d2d5bc),
	.w3(32'h38d9cebd),
	.w4(32'h37154601),
	.w5(32'h38b0b2ee),
	.w6(32'h384c4775),
	.w7(32'h38ac4c6c),
	.w8(32'h38b9dea7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9811654),
	.w1(32'hb913a794),
	.w2(32'hb8762749),
	.w3(32'hb81f9976),
	.w4(32'hb73a8cda),
	.w5(32'h388600b0),
	.w6(32'hb9183f50),
	.w7(32'hb94113dc),
	.w8(32'hb917214a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88dd758),
	.w1(32'h3770c309),
	.w2(32'h39d79c94),
	.w3(32'h39bbd8c7),
	.w4(32'h3a736e05),
	.w5(32'h3ab0adf1),
	.w6(32'hb90aa961),
	.w7(32'h3989bb83),
	.w8(32'h397dc634),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb0146),
	.w1(32'h3896a826),
	.w2(32'h3923fe64),
	.w3(32'hb846f316),
	.w4(32'h3897c4ed),
	.w5(32'h3972588d),
	.w6(32'hb9b570d7),
	.w7(32'hb9bebde9),
	.w8(32'hb952a987),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39076d4c),
	.w1(32'hb6a6d118),
	.w2(32'hb8c0379d),
	.w3(32'h396a54ad),
	.w4(32'hb85c5cd5),
	.w5(32'h37e95d2d),
	.w6(32'hb821ce76),
	.w7(32'hb7a45512),
	.w8(32'h3744afbb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aad8e5),
	.w1(32'hb7cf2c02),
	.w2(32'hb88de2b3),
	.w3(32'h3795be59),
	.w4(32'hb838ebbc),
	.w5(32'hb8b77279),
	.w6(32'hb7e5a73c),
	.w7(32'hb857cbdb),
	.w8(32'hb7a6e2c5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382d7f3e),
	.w1(32'h3902bd50),
	.w2(32'h39d2de7b),
	.w3(32'h395722ae),
	.w4(32'h39dd8863),
	.w5(32'h3a3c343d),
	.w6(32'h38ace9f6),
	.w7(32'h3a00c4c5),
	.w8(32'h39d7d920),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a0b5eb),
	.w1(32'hb7baf279),
	.w2(32'hb8153bae),
	.w3(32'h382dcf47),
	.w4(32'hb7ce7ac6),
	.w5(32'hb89d14e5),
	.w6(32'hb7fcdf45),
	.w7(32'hb8f5f9e6),
	.w8(32'hb82f1f60),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a6bf06),
	.w1(32'h37322160),
	.w2(32'hb55d0473),
	.w3(32'h37f05d24),
	.w4(32'h37d0d12f),
	.w5(32'h381cefc4),
	.w6(32'h382704a1),
	.w7(32'h38023725),
	.w8(32'h3828044b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e90a0),
	.w1(32'hb8888856),
	.w2(32'h38da8b30),
	.w3(32'h38b6e5c3),
	.w4(32'h39434d00),
	.w5(32'h39adade4),
	.w6(32'h38b2a03a),
	.w7(32'h3971ae84),
	.w8(32'h3998ea2d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78dfc9d),
	.w1(32'hb774a037),
	.w2(32'hb72cca77),
	.w3(32'hb7b9ebe3),
	.w4(32'hb7baba6e),
	.w5(32'hb76c7b1d),
	.w6(32'hb7b90e52),
	.w7(32'hb7a0fa2b),
	.w8(32'hb78b2b07),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cebf1),
	.w1(32'h3aad0da9),
	.w2(32'h39756e58),
	.w3(32'h3aad44e4),
	.w4(32'hb7cfae25),
	.w5(32'h3af4b2e0),
	.w6(32'h3b454b52),
	.w7(32'h3af7950a),
	.w8(32'h3b41af2e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f02b5),
	.w1(32'hb882c722),
	.w2(32'h3894b0e5),
	.w3(32'h3748f155),
	.w4(32'h390ad55d),
	.w5(32'h39831185),
	.w6(32'h38157302),
	.w7(32'h38f2efe6),
	.w8(32'h39118b23),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7576621),
	.w1(32'hb7d816a2),
	.w2(32'hb73a8531),
	.w3(32'h3759dda5),
	.w4(32'h36927340),
	.w5(32'h379d54de),
	.w6(32'h37e5f2d0),
	.w7(32'h37e6eca5),
	.w8(32'h382c4bda),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb881503a),
	.w1(32'hb8a3195c),
	.w2(32'hb88df4ee),
	.w3(32'hb75f6829),
	.w4(32'hb79146b6),
	.w5(32'hb728b4c4),
	.w6(32'hb79a4380),
	.w7(32'hb77a7538),
	.w8(32'hb79a60df),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88854d3),
	.w1(32'hb87fb93e),
	.w2(32'hb86f4c23),
	.w3(32'hb8381881),
	.w4(32'hb8a0e589),
	.w5(32'hb7a817e0),
	.w6(32'hb8b17fc0),
	.w7(32'hb873d9fa),
	.w8(32'h37097235),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36509433),
	.w1(32'h366474ac),
	.w2(32'h361cd696),
	.w3(32'h361c352f),
	.w4(32'h3694ae35),
	.w5(32'h36428d3d),
	.w6(32'h36adba4e),
	.w7(32'h366a1bd0),
	.w8(32'h365a9654),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367dc2d9),
	.w1(32'h365f8fe7),
	.w2(32'h362ad0aa),
	.w3(32'h3523eef1),
	.w4(32'h36008562),
	.w5(32'h3598e770),
	.w6(32'hb5a061da),
	.w7(32'hb52e6e65),
	.w8(32'hb54eb9b1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f468f),
	.w1(32'h38c9332d),
	.w2(32'h37ea225e),
	.w3(32'h3811a518),
	.w4(32'h386ddc1e),
	.w5(32'hb879550f),
	.w6(32'hb8994b64),
	.w7(32'hb8a1c610),
	.w8(32'hb88d4fc4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c60b1),
	.w1(32'hb91f2569),
	.w2(32'hb918b362),
	.w3(32'h38e131bb),
	.w4(32'h387bfeb7),
	.w5(32'h39222041),
	.w6(32'hb8bb1a17),
	.w7(32'hb828dce6),
	.w8(32'hb8d349c2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370428fa),
	.w1(32'h3634cd60),
	.w2(32'h36a7ac51),
	.w3(32'h36d284aa),
	.w4(32'h368b7016),
	.w5(32'h3700cfd3),
	.w6(32'h36c98a1e),
	.w7(32'h36983c21),
	.w8(32'h36c3209d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83a652d),
	.w1(32'hb81013f4),
	.w2(32'hb7ee5dba),
	.w3(32'h37ba0a32),
	.w4(32'h35ee52d3),
	.w5(32'h35fde343),
	.w6(32'h37d8a852),
	.w7(32'h3789030d),
	.w8(32'h37f96eeb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36112b50),
	.w1(32'h369a9a86),
	.w2(32'h36abb731),
	.w3(32'hb60ea751),
	.w4(32'hb6524ceb),
	.w5(32'hb6995d66),
	.w6(32'hb6223190),
	.w7(32'hb5f42f0e),
	.w8(32'hb58dc0dd),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378ff0e5),
	.w1(32'hb6cef7e2),
	.w2(32'h36e5e5cc),
	.w3(32'h36f03380),
	.w4(32'hb6cf72c4),
	.w5(32'h34ddd32e),
	.w6(32'hb6c7cd98),
	.w7(32'h36890c9d),
	.w8(32'h36e0e504),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b49b2),
	.w1(32'hb9b8d6b4),
	.w2(32'h39710e61),
	.w3(32'h358a54e8),
	.w4(32'h3950cc09),
	.w5(32'h39f8dfcf),
	.w6(32'h38d1772f),
	.w7(32'h38885922),
	.w8(32'hba3b6eff),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5309bc),
	.w1(32'hba2d17f6),
	.w2(32'hb9dab589),
	.w3(32'hb9a41e7d),
	.w4(32'hb88ab974),
	.w5(32'hb9872e6e),
	.w6(32'hb9a31e81),
	.w7(32'hb95509c3),
	.w8(32'h3b721a82),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6593e2),
	.w1(32'hba4ace23),
	.w2(32'h3b2ab28d),
	.w3(32'h3b84a394),
	.w4(32'hbb282e57),
	.w5(32'h3b141351),
	.w6(32'hbb2d23ba),
	.w7(32'h3a7fd851),
	.w8(32'hba3c01c6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cd93a),
	.w1(32'hb9b303dc),
	.w2(32'h35d668f8),
	.w3(32'hb95595db),
	.w4(32'h38eca0a6),
	.w5(32'h388c8671),
	.w6(32'hb92696b2),
	.w7(32'h37d5821d),
	.w8(32'h394476c0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4e24e),
	.w1(32'h397dff58),
	.w2(32'h3a108ab5),
	.w3(32'h3981ea35),
	.w4(32'h3a52ddf7),
	.w5(32'h3a5b912a),
	.w6(32'h3a21ffa7),
	.w7(32'h3a3e5cde),
	.w8(32'hbabc52d9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070f3c),
	.w1(32'hbac10a50),
	.w2(32'hba98a66d),
	.w3(32'hbacc377e),
	.w4(32'hba1901b3),
	.w5(32'hba31fe17),
	.w6(32'hbad06c0d),
	.w7(32'hbab92f1b),
	.w8(32'hba591036),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67f2d1),
	.w1(32'hbad5e45b),
	.w2(32'hb9ecf783),
	.w3(32'hbae8d233),
	.w4(32'hbb939164),
	.w5(32'h39d05efe),
	.w6(32'hbb47eb45),
	.w7(32'hbad0acec),
	.w8(32'hbab451aa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13880b),
	.w1(32'hbab2f070),
	.w2(32'hba99166a),
	.w3(32'hbb141f78),
	.w4(32'hba1568e0),
	.w5(32'hba48c2e7),
	.w6(32'hb9b039ea),
	.w7(32'hba206220),
	.w8(32'h3b2092c6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b5a8f),
	.w1(32'hbab7bcdf),
	.w2(32'hbace4cb4),
	.w3(32'h3b266a35),
	.w4(32'h3938c346),
	.w5(32'hb7f80b65),
	.w6(32'hb9ed1bc0),
	.w7(32'hba4b0db1),
	.w8(32'hb9219bd1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53ce42),
	.w1(32'hb98e86a2),
	.w2(32'h391b4f1e),
	.w3(32'hb9902646),
	.w4(32'h39d0b69a),
	.w5(32'h3a0ccd00),
	.w6(32'h38f7d8b8),
	.w7(32'h399379cd),
	.w8(32'hb9a6e966),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94dc22e),
	.w1(32'hb98501e9),
	.w2(32'hb9b9af17),
	.w3(32'hb88c06ef),
	.w4(32'h393c990d),
	.w5(32'hb9811296),
	.w6(32'h3802d1a2),
	.w7(32'h3827081d),
	.w8(32'hba836275),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ea7fa),
	.w1(32'hb9cb0be8),
	.w2(32'hb98fccc4),
	.w3(32'h38a8a9ef),
	.w4(32'h3a4dc2a3),
	.w5(32'h3895101b),
	.w6(32'h3a493aaf),
	.w7(32'h3a4b9be7),
	.w8(32'h3a3cea41),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21325f),
	.w1(32'hba8927c6),
	.w2(32'h393c8d35),
	.w3(32'hb9c1740a),
	.w4(32'hba01a74c),
	.w5(32'hbad4ba38),
	.w6(32'hba471932),
	.w7(32'hb7f92b0e),
	.w8(32'h3ae32307),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c57be),
	.w1(32'hb9794c28),
	.w2(32'hb979b611),
	.w3(32'h3ae10221),
	.w4(32'h3a45554f),
	.w5(32'h3a8d1f35),
	.w6(32'h392ea4b8),
	.w7(32'hb9aa9f0c),
	.w8(32'hb9a1fc84),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996436f),
	.w1(32'h3bc6c63a),
	.w2(32'h3b877376),
	.w3(32'hba60e61e),
	.w4(32'h3b1b6ae1),
	.w5(32'h3b26e1ec),
	.w6(32'h3aa41f8a),
	.w7(32'h3b282f05),
	.w8(32'hbb4b1962),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78c936),
	.w1(32'hbba663fc),
	.w2(32'hbb3d254b),
	.w3(32'hbb3e53b1),
	.w4(32'hbb43f600),
	.w5(32'hba9608ff),
	.w6(32'hbb73121e),
	.w7(32'hbad442dc),
	.w8(32'hbae6158d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e25bd),
	.w1(32'hb96f40c8),
	.w2(32'h3a5e19fc),
	.w3(32'hba5c482a),
	.w4(32'hbabd9b4b),
	.w5(32'h3972f659),
	.w6(32'hbb4e5fde),
	.w7(32'h392bc8ba),
	.w8(32'h3acf29f3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa7f63),
	.w1(32'hba174e19),
	.w2(32'hba90ce03),
	.w3(32'hba34d1db),
	.w4(32'h39b007b9),
	.w5(32'h3a470f14),
	.w6(32'hb9ebe547),
	.w7(32'hb9051288),
	.w8(32'h3b55715b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2faec5),
	.w1(32'hb92351ac),
	.w2(32'h39ccdb69),
	.w3(32'h3b6d6e9b),
	.w4(32'h3a90fafb),
	.w5(32'h3aa15edc),
	.w6(32'h3a6132cf),
	.w7(32'h3a915b67),
	.w8(32'hba37dfad),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d35f5),
	.w1(32'hb99c3b2b),
	.w2(32'hba8dbc60),
	.w3(32'hbae9058c),
	.w4(32'hbad3df64),
	.w5(32'hbab7c73b),
	.w6(32'hbaf86342),
	.w7(32'hbb189839),
	.w8(32'h3b08b4ac),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e21d8),
	.w1(32'hbb115c6f),
	.w2(32'h3b2bb06d),
	.w3(32'h394ae91d),
	.w4(32'hb867968e),
	.w5(32'h3aa5df08),
	.w6(32'hbb756e86),
	.w7(32'h3a98d174),
	.w8(32'hbb064731),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb371faf),
	.w1(32'hbb1f226d),
	.w2(32'hbaefd90e),
	.w3(32'hbb200187),
	.w4(32'hbb0964e4),
	.w5(32'hbad9d73c),
	.w6(32'hbabfbf88),
	.w7(32'hbaea037d),
	.w8(32'h3ac140ae),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d4f86),
	.w1(32'hba298f3d),
	.w2(32'h39613a58),
	.w3(32'h3ac068c9),
	.w4(32'h3a456a0b),
	.w5(32'h3a72ef79),
	.w6(32'h3a1c229f),
	.w7(32'h3a79cf04),
	.w8(32'hbafbd257),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84686e),
	.w1(32'hbba3c1b4),
	.w2(32'hbb028603),
	.w3(32'hbb4483d4),
	.w4(32'hbba0e518),
	.w5(32'hbb049f5f),
	.w6(32'hbabe19b0),
	.w7(32'hbb068d89),
	.w8(32'hb84b1b40),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3791649c),
	.w1(32'hb7b866e9),
	.w2(32'h3a0c2c3d),
	.w3(32'h39be5ce3),
	.w4(32'h39ba7ffe),
	.w5(32'h39c60a68),
	.w6(32'h39b711a1),
	.w7(32'h3a3382a3),
	.w8(32'hba2b06b6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1177e6),
	.w1(32'hb9db103e),
	.w2(32'hba077d02),
	.w3(32'hb9a66ab5),
	.w4(32'hb95f0536),
	.w5(32'hb9e6253e),
	.w6(32'hb9d49645),
	.w7(32'hb9eaaa04),
	.w8(32'hb9d41c5c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6c454),
	.w1(32'hb999119e),
	.w2(32'hb973317c),
	.w3(32'hb733a06d),
	.w4(32'h38c978a5),
	.w5(32'hb9154f61),
	.w6(32'hb8523bbd),
	.w7(32'hb8d1e881),
	.w8(32'hba6de2ad),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17d96e),
	.w1(32'hbb003207),
	.w2(32'hb97cc097),
	.w3(32'hba8f1062),
	.w4(32'hbb018d07),
	.w5(32'hba374612),
	.w6(32'hba9378b7),
	.w7(32'hba92e49b),
	.w8(32'hb92ea663),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba087a51),
	.w1(32'hb82b46ee),
	.w2(32'h38c7fa58),
	.w3(32'hb91e56e7),
	.w4(32'h399b09ea),
	.w5(32'h39907996),
	.w6(32'h386ebe32),
	.w7(32'h39010abd),
	.w8(32'h3b3bbb84),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49fbf8),
	.w1(32'h3acbc598),
	.w2(32'h3b387068),
	.w3(32'h3b5e937e),
	.w4(32'h3afaf5b4),
	.w5(32'h3b24b6db),
	.w6(32'h3b0c374b),
	.w7(32'h3b4f0c5e),
	.w8(32'h3a02afaf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dcc312),
	.w1(32'hb96c48ff),
	.w2(32'hb7ff2cad),
	.w3(32'h38d388bd),
	.w4(32'h398d86d1),
	.w5(32'h381cd36e),
	.w6(32'hb7949cce),
	.w7(32'h390f0bb4),
	.w8(32'hb9b29cc2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48328c),
	.w1(32'hb908d576),
	.w2(32'hb5fb333d),
	.w3(32'hba031df3),
	.w4(32'h39689be3),
	.w5(32'h39b47fa4),
	.w6(32'hb9242fcb),
	.w7(32'hb7e924b1),
	.w8(32'hba14b5ce),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0493b3),
	.w1(32'h390c1611),
	.w2(32'hb8660e9b),
	.w3(32'hb7290baf),
	.w4(32'h3a0cca8b),
	.w5(32'h378e8d8b),
	.w6(32'h38fdd00e),
	.w7(32'hb6342713),
	.w8(32'hbb39dce4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10eb1b),
	.w1(32'hbaeadef9),
	.w2(32'hba63bef4),
	.w3(32'hbb9cfbf5),
	.w4(32'hbb89aca0),
	.w5(32'hbb3863a5),
	.w6(32'hba259231),
	.w7(32'hb9a67877),
	.w8(32'hba4fb1aa),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90f1ca),
	.w1(32'hba0a277a),
	.w2(32'hb9d03a79),
	.w3(32'hba40a1ce),
	.w4(32'h37f594b9),
	.w5(32'hb915cc5e),
	.w6(32'hb8fb0f2c),
	.w7(32'hb9aaa31e),
	.w8(32'hb9e68c3d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a3040),
	.w1(32'hb7d174f1),
	.w2(32'h3915c0c3),
	.w3(32'h39142c5d),
	.w4(32'h39dc4ae9),
	.w5(32'h3941d658),
	.w6(32'h391a3ba4),
	.w7(32'h39a1dd1c),
	.w8(32'hb94803d1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19b4e6),
	.w1(32'hb9c7aafa),
	.w2(32'hb9c6a1dc),
	.w3(32'hb96b3a39),
	.w4(32'h3836e59f),
	.w5(32'hb89974da),
	.w6(32'hb9267cf0),
	.w7(32'hb9619881),
	.w8(32'h3b79f408),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e1f5b),
	.w1(32'h3ab86736),
	.w2(32'h3b2d0dc8),
	.w3(32'h3b9056ca),
	.w4(32'h3b199d30),
	.w5(32'h3b332289),
	.w6(32'h3b102389),
	.w7(32'h3b419340),
	.w8(32'h3acbe470),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba672d),
	.w1(32'h3a5e5fe5),
	.w2(32'h3aa9ba2b),
	.w3(32'h3aca53a1),
	.w4(32'h3a9dcfdb),
	.w5(32'h3abfc866),
	.w6(32'h3a96be4f),
	.w7(32'h3ace4968),
	.w8(32'hba1084c9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fa2ad),
	.w1(32'h39718639),
	.w2(32'h3830dcdc),
	.w3(32'hb929a534),
	.w4(32'hb89a0fdf),
	.w5(32'h37c336be),
	.w6(32'hb903f061),
	.w7(32'hb9282b7c),
	.w8(32'hbb262488),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9488ca),
	.w1(32'hbb7f5803),
	.w2(32'hba9d1b35),
	.w3(32'hb9a10362),
	.w4(32'hba7a9e80),
	.w5(32'hba85dee5),
	.w6(32'hbb67f783),
	.w7(32'hbb50c4e0),
	.w8(32'hba7c0146),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa44bb0),
	.w1(32'hba62973e),
	.w2(32'hba45365d),
	.w3(32'hba647dbe),
	.w4(32'hb9e332ac),
	.w5(32'hba2e677c),
	.w6(32'hba0dbf26),
	.w7(32'hba49c12c),
	.w8(32'hba8c7525),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacea368),
	.w1(32'h3a5db7e0),
	.w2(32'h398a3e9a),
	.w3(32'hba5553e8),
	.w4(32'h3a931621),
	.w5(32'h3a180a4d),
	.w6(32'hb996e6af),
	.w7(32'hb98adbb1),
	.w8(32'hb946f473),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a779179),
	.w1(32'h3a095148),
	.w2(32'hbac3767f),
	.w3(32'h3a268676),
	.w4(32'hbafdaa01),
	.w5(32'h3a5eecf4),
	.w6(32'hb9b25626),
	.w7(32'hbb2c3ff7),
	.w8(32'h3a4e5940),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bea2ed),
	.w1(32'h39d3922d),
	.w2(32'h3a24d80a),
	.w3(32'h3a8d01fb),
	.w4(32'h3a9c195f),
	.w5(32'h3a991290),
	.w6(32'h3a231a88),
	.w7(32'h3a425c38),
	.w8(32'h3a21492e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c5d19),
	.w1(32'hb96a9140),
	.w2(32'h399c70e4),
	.w3(32'h395a75e7),
	.w4(32'h39bee957),
	.w5(32'h3a2642ea),
	.w6(32'h3a1b2c9e),
	.w7(32'h3a0f019e),
	.w8(32'h3b56ac3a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adba242),
	.w1(32'hbaec4f47),
	.w2(32'hbb072bd4),
	.w3(32'h3b5eb46c),
	.w4(32'h397478e9),
	.w5(32'hb8c5a732),
	.w6(32'hba0a0acc),
	.w7(32'hba813f96),
	.w8(32'hb90ca661),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99532ce),
	.w1(32'h3a2874bb),
	.w2(32'h39ff97af),
	.w3(32'hb99478fc),
	.w4(32'h3a55eecc),
	.w5(32'h37d437e6),
	.w6(32'h3a399d79),
	.w7(32'h398865c4),
	.w8(32'hbaf29517),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6fd2d),
	.w1(32'hba1ce7f2),
	.w2(32'hbadfa76b),
	.w3(32'hbb121aa0),
	.w4(32'hbafff29e),
	.w5(32'hbb03146e),
	.w6(32'hbb224fca),
	.w7(32'hbb51e43a),
	.w8(32'h3b326729),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7ff0e),
	.w1(32'hbad78081),
	.w2(32'hbaef11fa),
	.w3(32'h3b50c71c),
	.w4(32'h39883066),
	.w5(32'hb7a7ea8d),
	.w6(32'hb9f59e98),
	.w7(32'hba597534),
	.w8(32'h3b1d9b4b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae7fb3),
	.w1(32'hbaad4430),
	.w2(32'hbac4bf12),
	.w3(32'h3b38a672),
	.w4(32'h39ac9cd2),
	.w5(32'h389647f8),
	.w6(32'hb98874d7),
	.w7(32'hba1c5821),
	.w8(32'h3a13e48b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904d77f),
	.w1(32'hba5148fe),
	.w2(32'hba34e7ed),
	.w3(32'h39ec8aa5),
	.w4(32'hba37697a),
	.w5(32'hb9e1e956),
	.w6(32'hba407f11),
	.w7(32'hba317ec2),
	.w8(32'hbaa27818),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66b2b3),
	.w1(32'h3a8a9793),
	.w2(32'h3a3f9579),
	.w3(32'hbb0d106b),
	.w4(32'hbafbc14a),
	.w5(32'hb8a43640),
	.w6(32'hba5697ce),
	.w7(32'hb9b14439),
	.w8(32'hb9d95b6b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcc69c),
	.w1(32'hb9c36ee6),
	.w2(32'hb988b5c1),
	.w3(32'hb98d4e09),
	.w4(32'hb5f314f2),
	.w5(32'hb8505649),
	.w6(32'hb924089f),
	.w7(32'hb927a420),
	.w8(32'hbb33ccfd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa356d5),
	.w1(32'hbb25b40c),
	.w2(32'hba8389c9),
	.w3(32'hbb8a370d),
	.w4(32'hbb670c7c),
	.w5(32'hbb31b4ca),
	.w6(32'hbb876ac9),
	.w7(32'hbb6ad515),
	.w8(32'h39991795),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a8e9c),
	.w1(32'hbaa4de44),
	.w2(32'hba685a0b),
	.w3(32'hb782465a),
	.w4(32'hba59964d),
	.w5(32'hba01fafb),
	.w6(32'hb77ff865),
	.w7(32'hb896a7fa),
	.w8(32'h3a926478),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d35ee),
	.w1(32'hbafb8ab9),
	.w2(32'hb9861b1f),
	.w3(32'hba48e3c8),
	.w4(32'h399dd7e6),
	.w5(32'h3a0dc93d),
	.w6(32'h39b18608),
	.w7(32'h39a98776),
	.w8(32'h3aba0be8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a811d5d),
	.w1(32'h395fd7f4),
	.w2(32'h3a0ca232),
	.w3(32'hbada4905),
	.w4(32'hbb5e08f3),
	.w5(32'h39f38a6d),
	.w6(32'h3b3d703f),
	.w7(32'hba72abd9),
	.w8(32'h3b599c88),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b583410),
	.w1(32'h3aa0f53f),
	.w2(32'h3b0d1bf4),
	.w3(32'h3b7108c7),
	.w4(32'h3aeca6cd),
	.w5(32'h3b0242cd),
	.w6(32'h3af7626b),
	.w7(32'h3b1a749c),
	.w8(32'hb9866296),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bda11),
	.w1(32'h3a8007b3),
	.w2(32'h3a46095e),
	.w3(32'h3943cba9),
	.w4(32'h3a6e35dd),
	.w5(32'h39c6b3d1),
	.w6(32'h3a0bb8de),
	.w7(32'h39e03275),
	.w8(32'hba8c65de),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba974fea),
	.w1(32'hbab56ed8),
	.w2(32'hba54324d),
	.w3(32'hbab53077),
	.w4(32'hbadf259a),
	.w5(32'hba36d034),
	.w6(32'hbb20bb7b),
	.w7(32'hbac9c327),
	.w8(32'hb9e43816),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d27bf),
	.w1(32'hb9bda15f),
	.w2(32'hb994a42b),
	.w3(32'hb682c665),
	.w4(32'h3948dd4d),
	.w5(32'hb92603a4),
	.w6(32'hb902509a),
	.w7(32'hb8ce2323),
	.w8(32'h3ae3564b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec9fe4),
	.w1(32'h3a937048),
	.w2(32'h3b19635c),
	.w3(32'h3afc4f60),
	.w4(32'h3ac2523c),
	.w5(32'h3b00a10a),
	.w6(32'h3ad6994b),
	.w7(32'h3b30c0be),
	.w8(32'h3938365d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39781a93),
	.w1(32'h3888f7d0),
	.w2(32'hb8e3efe3),
	.w3(32'h3a29f117),
	.w4(32'hb9769ecd),
	.w5(32'hb956cdbf),
	.w6(32'hba33398c),
	.w7(32'hba114a30),
	.w8(32'h3a675260),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f81cf2),
	.w1(32'hba38ac09),
	.w2(32'hba57f40c),
	.w3(32'h3a8abe2f),
	.w4(32'hb7617290),
	.w5(32'hb8f52655),
	.w6(32'hb9a048af),
	.w7(32'hb9fec046),
	.w8(32'h3a907ba5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e2198),
	.w1(32'hbb978a72),
	.w2(32'h3b6a31d4),
	.w3(32'h39de6bb2),
	.w4(32'hb870f7be),
	.w5(32'h3a59a3be),
	.w6(32'h3ac32c79),
	.w7(32'h3b3b0709),
	.w8(32'hb8d2578a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb011f92),
	.w1(32'hbc4c5db1),
	.w2(32'h3c635e76),
	.w3(32'h3c259c77),
	.w4(32'hbb9527d3),
	.w5(32'hbb030a30),
	.w6(32'hbbce8cb2),
	.w7(32'h3c728799),
	.w8(32'h3b0841b7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad11c7a),
	.w1(32'hbbda9a12),
	.w2(32'hb9841cc7),
	.w3(32'hbaec8f7a),
	.w4(32'hba311841),
	.w5(32'h3a601357),
	.w6(32'h3b6107e0),
	.w7(32'h3b202cf6),
	.w8(32'h3b719649),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cefa12),
	.w1(32'hbbcfc8b2),
	.w2(32'h391d9f7a),
	.w3(32'hba856ae4),
	.w4(32'hbaae7dd6),
	.w5(32'h3a903352),
	.w6(32'h3a9c67f6),
	.w7(32'hbaf9f375),
	.w8(32'hbb9c19f7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f9a842),
	.w1(32'hbc5df684),
	.w2(32'hbc4d585b),
	.w3(32'h3a87708b),
	.w4(32'hbb2ce31c),
	.w5(32'hbb9a3dba),
	.w6(32'hbb63a8e9),
	.w7(32'hbc043271),
	.w8(32'hbb155c8c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbefdc),
	.w1(32'h3c5523bb),
	.w2(32'hbac6a1ec),
	.w3(32'hba954023),
	.w4(32'hba800eb8),
	.w5(32'h3be22ee2),
	.w6(32'hbbdd71e9),
	.w7(32'hbb38349c),
	.w8(32'hba2f2cfc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a853aac),
	.w1(32'hbc931343),
	.w2(32'h3a0abcc4),
	.w3(32'hbb61956d),
	.w4(32'hbba73d75),
	.w5(32'h39815b6c),
	.w6(32'hbc38b8cf),
	.w7(32'hbb51cf92),
	.w8(32'h3bc991d2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc00601),
	.w1(32'h3a84041d),
	.w2(32'hbba81621),
	.w3(32'h3c8f5259),
	.w4(32'h3c32b1be),
	.w5(32'h3bb81e42),
	.w6(32'h3ae746a7),
	.w7(32'h3b8112a8),
	.w8(32'h3b5f7a8a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eec7d),
	.w1(32'hbc5ea0c1),
	.w2(32'hbaae86dd),
	.w3(32'h39f956db),
	.w4(32'hbb3d80d2),
	.w5(32'h395ce9ba),
	.w6(32'hba4617cf),
	.w7(32'hbb2045eb),
	.w8(32'hb9c69817),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba831c9e),
	.w1(32'hba8fe207),
	.w2(32'h392ba9aa),
	.w3(32'hbb2e37ea),
	.w4(32'hba96dabb),
	.w5(32'h3994190e),
	.w6(32'hb65e3dc7),
	.w7(32'h3a0723c6),
	.w8(32'hb890044b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64eb45),
	.w1(32'hbb95147f),
	.w2(32'h39b10e78),
	.w3(32'hbbb0e2fe),
	.w4(32'hbb41bf67),
	.w5(32'hb8424c4d),
	.w6(32'h3b4b7d2d),
	.w7(32'h3b3099dc),
	.w8(32'h399e0315),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cd6e1),
	.w1(32'h3c744009),
	.w2(32'hbc66ed75),
	.w3(32'hbcabb837),
	.w4(32'h3cf27e16),
	.w5(32'hb96b7441),
	.w6(32'hbd3e2676),
	.w7(32'hbc967e5a),
	.w8(32'h3b3a36b0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3ae47),
	.w1(32'hbc0626f3),
	.w2(32'hbc21af9f),
	.w3(32'h3c763226),
	.w4(32'h3afffe0f),
	.w5(32'hbb4f27cd),
	.w6(32'hbbb73209),
	.w7(32'hbb6da24c),
	.w8(32'h3bfc5f75),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb7cd0),
	.w1(32'hbc0083e6),
	.w2(32'h3c892e4a),
	.w3(32'h3c0ca045),
	.w4(32'hbc2cecef),
	.w5(32'hbab0238b),
	.w6(32'h3b7a1d37),
	.w7(32'h3c69decc),
	.w8(32'hbb16b01b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46b202),
	.w1(32'hbc8eb7db),
	.w2(32'hbcade8be),
	.w3(32'h3a06acc1),
	.w4(32'hbc425106),
	.w5(32'hbc1d5124),
	.w6(32'hbc23dead),
	.w7(32'hbabc95c2),
	.w8(32'h3c122f9f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a188b0f),
	.w1(32'h3beff9d1),
	.w2(32'hbbb01f41),
	.w3(32'h3b4bdea3),
	.w4(32'h3c2d55c9),
	.w5(32'hbc256803),
	.w6(32'h3b9c0b9d),
	.w7(32'hba8d067e),
	.w8(32'h3bf019db),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80e75d),
	.w1(32'h3b241f6b),
	.w2(32'hba41af6a),
	.w3(32'h387fed08),
	.w4(32'h3ba95a68),
	.w5(32'hbba9c82f),
	.w6(32'hbab82f7e),
	.w7(32'hba274051),
	.w8(32'h3c089450),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b931cbf),
	.w1(32'h39a3019b),
	.w2(32'h3b42e549),
	.w3(32'h3c0c3911),
	.w4(32'h3bdb9473),
	.w5(32'h3bd1e422),
	.w6(32'h3be83d27),
	.w7(32'h3c0d9eaa),
	.w8(32'h3b3f1dec),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b71f30),
	.w1(32'hbb8f14ba),
	.w2(32'hbb69444c),
	.w3(32'h3b942bb2),
	.w4(32'h3bcf7228),
	.w5(32'hbb26f215),
	.w6(32'hbbea67c1),
	.w7(32'hbc1e1fb5),
	.w8(32'hbc1dda7a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ff625),
	.w1(32'hbc8cd6ff),
	.w2(32'hbbc22288),
	.w3(32'hbb285bc1),
	.w4(32'h3c824cab),
	.w5(32'h3c9aa287),
	.w6(32'hbcc20aa8),
	.w7(32'hbbf1e176),
	.w8(32'hbc27d4f6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa64633),
	.w1(32'hbca1eb68),
	.w2(32'hbc396090),
	.w3(32'hbb37b887),
	.w4(32'hbbfc64d6),
	.w5(32'hbbc87bbe),
	.w6(32'hbc1d001e),
	.w7(32'h39df7fc3),
	.w8(32'h3b45c7f6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8dcf9),
	.w1(32'hbbef5ecf),
	.w2(32'h3a0c186d),
	.w3(32'h397160a7),
	.w4(32'hbb03b03e),
	.w5(32'h3a8d8cef),
	.w6(32'h3b62a981),
	.w7(32'h3bd1284d),
	.w8(32'h3b854e63),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca86ff8),
	.w1(32'h3ca4c72a),
	.w2(32'h3aa9e618),
	.w3(32'hbbae7a2d),
	.w4(32'h3ca837d6),
	.w5(32'h3c7240a9),
	.w6(32'h3be23968),
	.w7(32'hbad26e65),
	.w8(32'h3abb95f7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule