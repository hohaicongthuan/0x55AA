module layer_8_featuremap_164(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca970c5),
	.w1(32'h3bb50401),
	.w2(32'h3b04ef01),
	.w3(32'h3c8d86e3),
	.w4(32'h3c8c7532),
	.w5(32'h3c2d0d18),
	.w6(32'h3c32889b),
	.w7(32'h3bd0bf79),
	.w8(32'h3bb1a314),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fac82),
	.w1(32'hbba3beca),
	.w2(32'hbbe4b95d),
	.w3(32'hbb56627c),
	.w4(32'hba449f3a),
	.w5(32'hbabc90c2),
	.w6(32'hbba60412),
	.w7(32'hbadf7e9c),
	.w8(32'hba235d1c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc231805),
	.w1(32'hbbad341c),
	.w2(32'hbbbe25cf),
	.w3(32'hbbb2880d),
	.w4(32'hbb7962ca),
	.w5(32'hbc32303c),
	.w6(32'hbc5b1f94),
	.w7(32'hbc2dc4dd),
	.w8(32'hbc5f1704),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28c9a5),
	.w1(32'hbb0945bc),
	.w2(32'hbb9f6f40),
	.w3(32'hbc994b37),
	.w4(32'hbb8d5eea),
	.w5(32'hbc2a2f9a),
	.w6(32'h3b4433ac),
	.w7(32'hbc1d884d),
	.w8(32'hbc9f333f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56afde),
	.w1(32'hbb6671f2),
	.w2(32'hbbca3770),
	.w3(32'hbc7185c9),
	.w4(32'h3aed0575),
	.w5(32'hbae2b982),
	.w6(32'h3a5fe7f2),
	.w7(32'h3bae87d2),
	.w8(32'h3bb1c36b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65c248),
	.w1(32'hbc2b140c),
	.w2(32'hbbda2677),
	.w3(32'hbc589819),
	.w4(32'hbbc1dca3),
	.w5(32'h3b73471f),
	.w6(32'hbc5ebfd2),
	.w7(32'hbc2fab13),
	.w8(32'h3a10c068),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb057dc),
	.w1(32'hbabdf90f),
	.w2(32'h3a4f19c7),
	.w3(32'hbb1fc492),
	.w4(32'hba3ce1ad),
	.w5(32'h3a0ad045),
	.w6(32'hbaeee47e),
	.w7(32'hba2f788b),
	.w8(32'h392d1565),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a945b5e),
	.w1(32'h39978e4b),
	.w2(32'h3c092387),
	.w3(32'h3b91e729),
	.w4(32'h3a8bb228),
	.w5(32'h3c262e15),
	.w6(32'h3a3a7d32),
	.w7(32'h3aad13e6),
	.w8(32'h3ab9f285),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083ff8),
	.w1(32'hbb96563a),
	.w2(32'hbbac16de),
	.w3(32'h3986870d),
	.w4(32'h3b4d43bb),
	.w5(32'h3b84889a),
	.w6(32'hbbdfd36a),
	.w7(32'h3ba1c7c9),
	.w8(32'h3b0b2c52),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e42ba),
	.w1(32'h3c07b1aa),
	.w2(32'h3bb246a3),
	.w3(32'h3b4e84be),
	.w4(32'h3b8b348e),
	.w5(32'h3b8c132c),
	.w6(32'hbbdb2ba4),
	.w7(32'h3bddb282),
	.w8(32'h3b92ba2d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5297bc),
	.w1(32'h3acbceaa),
	.w2(32'h3b96bcbf),
	.w3(32'hbb2bb8b6),
	.w4(32'hba382d44),
	.w5(32'h38aea96c),
	.w6(32'h3bd1298e),
	.w7(32'h3c08bcc7),
	.w8(32'h3c507b7c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb288c29),
	.w1(32'hbbcd2df1),
	.w2(32'hbbc287b4),
	.w3(32'hba052e23),
	.w4(32'h3aacebbc),
	.w5(32'hb83d7b2a),
	.w6(32'hbb0621a1),
	.w7(32'hbb41e507),
	.w8(32'h3ab80d5a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8f748),
	.w1(32'hbb0050db),
	.w2(32'h3abaee39),
	.w3(32'hbb2d63c5),
	.w4(32'h3c2f9be7),
	.w5(32'h3bc7d22a),
	.w6(32'hbc0dfa0e),
	.w7(32'hbb30692a),
	.w8(32'hbc2e05d0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9d91f),
	.w1(32'hbb455e83),
	.w2(32'hbbbac828),
	.w3(32'hbc406ae2),
	.w4(32'hba02a1da),
	.w5(32'hbb942c7e),
	.w6(32'hbb8c785d),
	.w7(32'hbc0e13f5),
	.w8(32'hbbe62826),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b53cb),
	.w1(32'hba1e340b),
	.w2(32'h3b3fad86),
	.w3(32'hbc031fd4),
	.w4(32'hba58787e),
	.w5(32'h3af1f6f0),
	.w6(32'hbb3f243a),
	.w7(32'hb841fecf),
	.w8(32'hba19ecb2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38efe34d),
	.w1(32'h3b073e14),
	.w2(32'hba598f96),
	.w3(32'hb9d0d2db),
	.w4(32'h3c6b1580),
	.w5(32'h3b3c93e9),
	.w6(32'h3a87fe89),
	.w7(32'h38e5177d),
	.w8(32'hbc0dae1f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc117698),
	.w1(32'h3aaaaf79),
	.w2(32'hbb627a35),
	.w3(32'hbad26ab9),
	.w4(32'h3ac9eeca),
	.w5(32'hbb82ccb7),
	.w6(32'hbb95066a),
	.w7(32'hbb4f3bc2),
	.w8(32'hbc09eec0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc158ec7),
	.w1(32'hbbab1cd6),
	.w2(32'hbc30e32f),
	.w3(32'hbb0aa2e1),
	.w4(32'h3aeec9d4),
	.w5(32'hbb89e177),
	.w6(32'hbc27a5e7),
	.w7(32'hba0a0f2d),
	.w8(32'hbc10932e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c952d),
	.w1(32'hbcbda0cc),
	.w2(32'hbd02c255),
	.w3(32'hbad86f96),
	.w4(32'hbab28bbb),
	.w5(32'hbbf9a957),
	.w6(32'hbb8eae60),
	.w7(32'h3c0600a6),
	.w8(32'hbb8000c1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdbf2f),
	.w1(32'h3bc51ffa),
	.w2(32'h3bc0ff60),
	.w3(32'h3bf59c73),
	.w4(32'h3c64b970),
	.w5(32'h3bdfbc7a),
	.w6(32'h3ad3e75d),
	.w7(32'h3c204977),
	.w8(32'h3b65b1d2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f61c2f),
	.w1(32'hbb5c69ec),
	.w2(32'hbbf0562c),
	.w3(32'h397f677b),
	.w4(32'h3c0b8e01),
	.w5(32'hbbb2cc37),
	.w6(32'hbbcb1bf2),
	.w7(32'hbb6e0919),
	.w8(32'hbbd4c72d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62f1b9),
	.w1(32'hbbcf74ca),
	.w2(32'hbb8c002c),
	.w3(32'hbc49309a),
	.w4(32'h3c22a44c),
	.w5(32'hb9328456),
	.w6(32'hbbb43504),
	.w7(32'hbb1f0992),
	.w8(32'hbb2885d0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca30694),
	.w1(32'h3c21c9d7),
	.w2(32'h3b6f6ddc),
	.w3(32'h3d04badf),
	.w4(32'h3cbdcf38),
	.w5(32'h3cb89ea5),
	.w6(32'hbaedcd2b),
	.w7(32'h3c7a4f87),
	.w8(32'h3cf0e8d2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a0d20),
	.w1(32'h3b281360),
	.w2(32'hba247e5e),
	.w3(32'h3af978f5),
	.w4(32'h3b66dc23),
	.w5(32'hbac7c38d),
	.w6(32'h3b1405e2),
	.w7(32'hba766be2),
	.w8(32'h3c08a598),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023f16),
	.w1(32'hb9d1af90),
	.w2(32'hbbac0008),
	.w3(32'hbbbbb662),
	.w4(32'hbad9672f),
	.w5(32'hbc277b77),
	.w6(32'hbb47e48c),
	.w7(32'h37d48aee),
	.w8(32'h3a319d09),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4d5f8),
	.w1(32'h3cb9110e),
	.w2(32'h3c234064),
	.w3(32'h3bb4da15),
	.w4(32'h3c9bc8cb),
	.w5(32'h3b0f2cdf),
	.w6(32'h3ca4ca53),
	.w7(32'h3c48d4c3),
	.w8(32'h3c853b49),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12ee70),
	.w1(32'h3b569379),
	.w2(32'hba0381b9),
	.w3(32'hbc2ba4d6),
	.w4(32'h3bcac85c),
	.w5(32'h3a879032),
	.w6(32'h3b906797),
	.w7(32'hbb966b27),
	.w8(32'hbb57aa6a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda4716),
	.w1(32'hbc26073a),
	.w2(32'hbc20d476),
	.w3(32'h3ce44de8),
	.w4(32'h3ce75741),
	.w5(32'h3bd2cd56),
	.w6(32'h3cbc2690),
	.w7(32'h3c31d3c5),
	.w8(32'h3b898588),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20fd07),
	.w1(32'hba35910b),
	.w2(32'h382f9c5c),
	.w3(32'hbb51b180),
	.w4(32'h3c5309ef),
	.w5(32'h3c0a7180),
	.w6(32'hba9f5c9f),
	.w7(32'h3b4edfe6),
	.w8(32'h3c20b766),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c3d02),
	.w1(32'hbafda248),
	.w2(32'hb99f535e),
	.w3(32'h3c17c788),
	.w4(32'h3aa3f528),
	.w5(32'h3a8ae720),
	.w6(32'hbb4ef099),
	.w7(32'h3a804680),
	.w8(32'h3ac307d1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92f452),
	.w1(32'h3a8f4a46),
	.w2(32'h3b9a8e26),
	.w3(32'hbbcf5b47),
	.w4(32'h3c2faf34),
	.w5(32'h3c25c4d2),
	.w6(32'hbbe796ef),
	.w7(32'hba4a78e9),
	.w8(32'hbb13f848),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399839be),
	.w1(32'hbae52927),
	.w2(32'hbbf7a998),
	.w3(32'h3b1250cc),
	.w4(32'hbb5d5c1f),
	.w5(32'hbb5f87c7),
	.w6(32'hbb34c60f),
	.w7(32'h3a9f5f48),
	.w8(32'h3b4430eb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bebd4),
	.w1(32'h3c011a60),
	.w2(32'h3b8494bc),
	.w3(32'h3c556fc9),
	.w4(32'h3b6b099e),
	.w5(32'h3b5098fe),
	.w6(32'h3b8de8c9),
	.w7(32'h3bc5d3c3),
	.w8(32'hbac63d92),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f06d2),
	.w1(32'hbb9c1889),
	.w2(32'hbc0d36b2),
	.w3(32'hbb5e4f29),
	.w4(32'hbbaad615),
	.w5(32'hba3edbb0),
	.w6(32'hbbcfc0d1),
	.w7(32'hbbfe1e25),
	.w8(32'hba640daf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2976a3),
	.w1(32'h3bf98c63),
	.w2(32'h3c289899),
	.w3(32'hbc48892d),
	.w4(32'h3aaa77ba),
	.w5(32'h3b9b7e13),
	.w6(32'hbbb39ad5),
	.w7(32'h397f782e),
	.w8(32'h3a8d75ee),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87625c),
	.w1(32'hba2eeabe),
	.w2(32'hbbe67df7),
	.w3(32'h3c0ff3f0),
	.w4(32'h3ba24126),
	.w5(32'h3b23a865),
	.w6(32'h3b7bae90),
	.w7(32'h3b870f51),
	.w8(32'h3959e026),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b382779),
	.w1(32'h3ba0f9dc),
	.w2(32'h3b6dbbd6),
	.w3(32'h3a451d06),
	.w4(32'h3bd08aa7),
	.w5(32'h3b27d7bd),
	.w6(32'hb9fd3491),
	.w7(32'hb9bc60fd),
	.w8(32'hbb1f5526),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba025667),
	.w1(32'h39a7124f),
	.w2(32'h3a7a60ea),
	.w3(32'hbaafded5),
	.w4(32'h3a91d163),
	.w5(32'h3b81d70a),
	.w6(32'hbb1ad6c9),
	.w7(32'h3b836084),
	.w8(32'hb94670d6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3c398),
	.w1(32'hbaa105be),
	.w2(32'h3c25458b),
	.w3(32'h3b046582),
	.w4(32'hba8687f6),
	.w5(32'h3ba3a2d5),
	.w6(32'hbb08ba30),
	.w7(32'h3b09595a),
	.w8(32'hbb13bde7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a390d5a),
	.w1(32'hbbbbcb69),
	.w2(32'hbbb879b0),
	.w3(32'hb98dbb75),
	.w4(32'hbbddd67b),
	.w5(32'hbbd34bb7),
	.w6(32'hbbad72e8),
	.w7(32'hbbc76ce9),
	.w8(32'hba7cbb11),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec095d),
	.w1(32'hbabc099a),
	.w2(32'hbad0389a),
	.w3(32'h3bbb22f0),
	.w4(32'h3c243b5b),
	.w5(32'h3bdfb1d6),
	.w6(32'h3bfb45f2),
	.w7(32'h3bd765ad),
	.w8(32'h3bbe425f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b416622),
	.w1(32'hbbbe87c9),
	.w2(32'hbb5e2fd7),
	.w3(32'h3a7e3a3f),
	.w4(32'hba3dc0ee),
	.w5(32'h3b3f90cb),
	.w6(32'hbbf65f44),
	.w7(32'hbaa5ad04),
	.w8(32'h3bdfc938),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c266664),
	.w1(32'h38a2b3d9),
	.w2(32'h3b8fbafd),
	.w3(32'h3c348523),
	.w4(32'hbb3ea57a),
	.w5(32'hbaa107b1),
	.w6(32'hbb003ed5),
	.w7(32'h3a968bd8),
	.w8(32'hba072842),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e4780),
	.w1(32'hbbb78487),
	.w2(32'hbb3c12b8),
	.w3(32'hbb3457da),
	.w4(32'hbbe176fd),
	.w5(32'hbba472a6),
	.w6(32'hbafa6077),
	.w7(32'h3b964bb2),
	.w8(32'hbab526da),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaef5f),
	.w1(32'h3b149de3),
	.w2(32'hbbe17877),
	.w3(32'hbbb0ef8b),
	.w4(32'h3b80b355),
	.w5(32'h3b1de4ff),
	.w6(32'hb96d7823),
	.w7(32'hb93df672),
	.w8(32'h3b3a222a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9699af),
	.w1(32'hbc0d4b13),
	.w2(32'hbbb37a48),
	.w3(32'h3b6720d5),
	.w4(32'hbb177479),
	.w5(32'h3b90b983),
	.w6(32'hbbe32ffb),
	.w7(32'hbb3a6354),
	.w8(32'h3b9761be),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab46b1d),
	.w1(32'hbbeeb032),
	.w2(32'hbb9e35af),
	.w3(32'h3a89fcd3),
	.w4(32'hbb87bcee),
	.w5(32'h3a7511b3),
	.w6(32'hbc42a467),
	.w7(32'hbbadce01),
	.w8(32'hbb8bdb64),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafee14),
	.w1(32'h3a95bfd2),
	.w2(32'hbc36fea5),
	.w3(32'h3c8b07b5),
	.w4(32'h3bd23724),
	.w5(32'hbbf4a47d),
	.w6(32'h3bef9996),
	.w7(32'h3a8015f0),
	.w8(32'h3bf76700),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c9df3),
	.w1(32'h3b52e802),
	.w2(32'hbac70b51),
	.w3(32'hbc0f4a36),
	.w4(32'h3c31e744),
	.w5(32'hbae739e8),
	.w6(32'hbbc6bd88),
	.w7(32'hbbc685f7),
	.w8(32'hba86b531),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedffb4),
	.w1(32'hbb6df8aa),
	.w2(32'hbc0175a8),
	.w3(32'hbcb4953c),
	.w4(32'hbbc4ffda),
	.w5(32'hbbd5fbe5),
	.w6(32'h3bb4d25d),
	.w7(32'hbb6cad32),
	.w8(32'hbbdcd0d3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d0ac1),
	.w1(32'hbbff3ce5),
	.w2(32'hbc89fbb6),
	.w3(32'hbc51ddc0),
	.w4(32'h3786fbee),
	.w5(32'hbc263f83),
	.w6(32'hbb470a17),
	.w7(32'hbbaba1b9),
	.w8(32'hbbf01659),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88ec6b),
	.w1(32'hbc1854d9),
	.w2(32'hbcdb979d),
	.w3(32'hba3eb94b),
	.w4(32'hbb86d86e),
	.w5(32'hbc885c02),
	.w6(32'hbbf0fef8),
	.w7(32'h3aa31dbe),
	.w8(32'hbbdc401e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78e927),
	.w1(32'h3a91df86),
	.w2(32'hbb982427),
	.w3(32'h3b843c73),
	.w4(32'h3b7cf6e5),
	.w5(32'hbb2c3084),
	.w6(32'h3ab744e1),
	.w7(32'h3c0c20f4),
	.w8(32'h3a82ec11),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf94549),
	.w1(32'h3aff8f4a),
	.w2(32'h3bfe3b23),
	.w3(32'hba21fbd9),
	.w4(32'h3c008aa3),
	.w5(32'h3c8178df),
	.w6(32'hbb62e455),
	.w7(32'h3c4719ba),
	.w8(32'h3bf48f60),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd460bc),
	.w1(32'h3b22d323),
	.w2(32'h3a240445),
	.w3(32'hbb87d81b),
	.w4(32'hbbb697a1),
	.w5(32'hbb91e2dc),
	.w6(32'h3b71d031),
	.w7(32'hbba1c4d2),
	.w8(32'hbb059929),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bb4ac),
	.w1(32'h3afc0add),
	.w2(32'hbc8e0fe2),
	.w3(32'h3bec930e),
	.w4(32'h3c055d2c),
	.w5(32'hbaabb311),
	.w6(32'hb98712de),
	.w7(32'h3c1b8bf8),
	.w8(32'hba252fb4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f5b51),
	.w1(32'h3afca5ba),
	.w2(32'h3b9b408d),
	.w3(32'hbc289fa7),
	.w4(32'h3c41063a),
	.w5(32'h3a94dafb),
	.w6(32'hbc0e254b),
	.w7(32'hbb1e7e2d),
	.w8(32'hbbc14ef3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2eb0db),
	.w1(32'h3a758890),
	.w2(32'hba0a6e45),
	.w3(32'hbc814179),
	.w4(32'h3b1598f9),
	.w5(32'h3bc53c73),
	.w6(32'hbb40a1e8),
	.w7(32'h3b7554cb),
	.w8(32'h3adfc0e1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81927e),
	.w1(32'hba0fd86e),
	.w2(32'hba61b99e),
	.w3(32'h39f5968f),
	.w4(32'h3a12f85c),
	.w5(32'h3afe5d5c),
	.w6(32'h3aaeba27),
	.w7(32'h3b00cd1b),
	.w8(32'h3bbe8b83),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b812b15),
	.w1(32'hbc1048c2),
	.w2(32'hbbaed94b),
	.w3(32'h3b96b6b8),
	.w4(32'hbba4c21b),
	.w5(32'hbbd46359),
	.w6(32'hbc397e98),
	.w7(32'hbc4f35cb),
	.w8(32'h3a549751),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26fd1f),
	.w1(32'hbbd758fd),
	.w2(32'hbb526760),
	.w3(32'hbc652af3),
	.w4(32'h3b9bbbc9),
	.w5(32'hbaff9d29),
	.w6(32'hbb29aec0),
	.w7(32'hbad1518e),
	.w8(32'h3b120420),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c6971),
	.w1(32'hbb0b5abd),
	.w2(32'hbbd41412),
	.w3(32'hbc1ac4b8),
	.w4(32'hbb461dd7),
	.w5(32'hbb780adc),
	.w6(32'hbc25fa3d),
	.w7(32'hbc32e275),
	.w8(32'hbc13a471),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf134e),
	.w1(32'hbb834003),
	.w2(32'hbc139e0d),
	.w3(32'h3c84ab6d),
	.w4(32'h3aebb7d8),
	.w5(32'h3b05add5),
	.w6(32'hba7a1977),
	.w7(32'h3bcc514a),
	.w8(32'hbb3c3d14),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f40bc2),
	.w1(32'h3bdf7567),
	.w2(32'h3bb5622a),
	.w3(32'h3b16bc3d),
	.w4(32'h3b8f038b),
	.w5(32'h3b560ff9),
	.w6(32'h3ab2770c),
	.w7(32'h3bc1d6bc),
	.w8(32'h3bfec369),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c255d95),
	.w1(32'h378dbda4),
	.w2(32'h3bb49b53),
	.w3(32'h3c04878c),
	.w4(32'h39d08482),
	.w5(32'h3c09f7cd),
	.w6(32'h39cb8916),
	.w7(32'h3ad61821),
	.w8(32'h3bb31e56),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd30ffc),
	.w1(32'hbc189da0),
	.w2(32'hbbf088e5),
	.w3(32'h3c2253d2),
	.w4(32'hbb16a755),
	.w5(32'hbb75b8b3),
	.w6(32'h3786c868),
	.w7(32'h39ada83a),
	.w8(32'hbab9f7cb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2afca7),
	.w1(32'h3b36e0d6),
	.w2(32'hbc8817cc),
	.w3(32'hbb96f40a),
	.w4(32'h384de5a8),
	.w5(32'hbc0fbb9c),
	.w6(32'h3a3fee64),
	.w7(32'h3a1b7940),
	.w8(32'hbb14ddd8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc066650),
	.w1(32'hbb9210bb),
	.w2(32'hbc386a5c),
	.w3(32'h3b77199b),
	.w4(32'h39895081),
	.w5(32'hba5d50c2),
	.w6(32'hbbf57f6b),
	.w7(32'hbbbb5b64),
	.w8(32'hbc0b74ed),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22b7b8),
	.w1(32'h390adbc2),
	.w2(32'hbc08b3a4),
	.w3(32'hbb8dd2cb),
	.w4(32'h3b4c220a),
	.w5(32'h3b04aef3),
	.w6(32'hb9c49320),
	.w7(32'hbb9b1c76),
	.w8(32'hbb9628e2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7a35b),
	.w1(32'h3c5ec26f),
	.w2(32'h3c0d539e),
	.w3(32'h3c4a279c),
	.w4(32'h3c8f97df),
	.w5(32'h3bc872f7),
	.w6(32'h3a68a21c),
	.w7(32'h3b90fa90),
	.w8(32'h3cb97560),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66eefb),
	.w1(32'hbc01bb52),
	.w2(32'hbb51d615),
	.w3(32'hbbe3e4d6),
	.w4(32'hbc44299f),
	.w5(32'hbbaf88a8),
	.w6(32'hbbb2ae96),
	.w7(32'h3a75cd78),
	.w8(32'h3b77e958),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e72b7),
	.w1(32'h39acf36a),
	.w2(32'hbb8648a7),
	.w3(32'h3b8e5820),
	.w4(32'h3b9051ca),
	.w5(32'hbbcaa5ba),
	.w6(32'hbb8e2bb8),
	.w7(32'h3a157c57),
	.w8(32'hbb85b60c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba980ab4),
	.w1(32'hbb8a0af9),
	.w2(32'hbb631128),
	.w3(32'hbae377ec),
	.w4(32'hbb011c8d),
	.w5(32'hbc0bc2cd),
	.w6(32'h3a3d2384),
	.w7(32'hbb8eebc2),
	.w8(32'hbc0d4973),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb7c64),
	.w1(32'hbbf7c916),
	.w2(32'h3b66d2b7),
	.w3(32'hbbfcf9ce),
	.w4(32'h3c05037a),
	.w5(32'h3c0e2ff3),
	.w6(32'hbbbf4852),
	.w7(32'h3b74a77a),
	.w8(32'hbb45d342),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f3ccd),
	.w1(32'hbb714732),
	.w2(32'hbbef5db3),
	.w3(32'hbc15837e),
	.w4(32'hbb3f2f29),
	.w5(32'hbbcc13a8),
	.w6(32'hbbe51cd2),
	.w7(32'hbc0c417e),
	.w8(32'h39deee86),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fc52d),
	.w1(32'h3adddab4),
	.w2(32'h3b4ff3d0),
	.w3(32'hba4a8727),
	.w4(32'h3bcc46f1),
	.w5(32'h38ffe2d8),
	.w6(32'h3b035829),
	.w7(32'h3c68b1d9),
	.w8(32'h3be426cd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a5852),
	.w1(32'hb9b86955),
	.w2(32'h3965df64),
	.w3(32'h3b447b01),
	.w4(32'hbb6bca89),
	.w5(32'hbb6316f2),
	.w6(32'hbbb1ad7d),
	.w7(32'hbac15b6c),
	.w8(32'h3b88dd0c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c55c3),
	.w1(32'h3bf6d4d5),
	.w2(32'hbb2b3d7a),
	.w3(32'h3b2b309e),
	.w4(32'h3c1adc7a),
	.w5(32'h3b801edd),
	.w6(32'h3c0256a5),
	.w7(32'h3c4168ff),
	.w8(32'h3c02f3f3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79ab23),
	.w1(32'hbb11eb53),
	.w2(32'h3b10970e),
	.w3(32'h3ae5b114),
	.w4(32'h3bfe90b7),
	.w5(32'h3c2ac5b4),
	.w6(32'h3c058cb7),
	.w7(32'h3bf2758e),
	.w8(32'h3aacbd50),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecf1b8),
	.w1(32'hbb629a60),
	.w2(32'hbc0e9cdc),
	.w3(32'hbbc0f145),
	.w4(32'hbabc9e8e),
	.w5(32'hbbd5ed0e),
	.w6(32'h3b6f0199),
	.w7(32'hbb7d3b7f),
	.w8(32'hbbc0c824),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9af65b),
	.w1(32'h3be0af9f),
	.w2(32'h3bd09590),
	.w3(32'h3aae2782),
	.w4(32'h3c27962e),
	.w5(32'hbb91134f),
	.w6(32'h3b6de63d),
	.w7(32'hba8ccd61),
	.w8(32'hbc0945a8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a9220),
	.w1(32'hbc3994e2),
	.w2(32'hbc51ee59),
	.w3(32'hbc972550),
	.w4(32'hbc1ff6b7),
	.w5(32'hbc0af8d9),
	.w6(32'hbc837744),
	.w7(32'hbc566800),
	.w8(32'hbc180097),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38a453),
	.w1(32'hbb950b4c),
	.w2(32'hb853093a),
	.w3(32'h3b9f53c7),
	.w4(32'h3c3da2e4),
	.w5(32'h3c0998dd),
	.w6(32'h3b19f3f4),
	.w7(32'h3c2121b8),
	.w8(32'h3c5ae47b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ae485),
	.w1(32'hbcbc0b00),
	.w2(32'hbcdf303a),
	.w3(32'hbc916e62),
	.w4(32'hbcd29ab4),
	.w5(32'hbc851b83),
	.w6(32'hbc82c0c2),
	.w7(32'hbcccd3d6),
	.w8(32'hbd014e65),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95e28),
	.w1(32'h3c4da636),
	.w2(32'h3909bf84),
	.w3(32'h3bf0eab5),
	.w4(32'h3cbe2246),
	.w5(32'h3c091806),
	.w6(32'h3c835813),
	.w7(32'h3c410d2f),
	.w8(32'h3c0b0e3a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc1682),
	.w1(32'h37fcfdd8),
	.w2(32'hbb02ed4d),
	.w3(32'hbac1e8b8),
	.w4(32'h3c2ab540),
	.w5(32'h3b807119),
	.w6(32'h3b9a26e1),
	.w7(32'h3c54ffa3),
	.w8(32'h3bbbf581),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983d2c0),
	.w1(32'h391a8e64),
	.w2(32'h3b207d71),
	.w3(32'hbb0ab79e),
	.w4(32'hba521cdc),
	.w5(32'h3b0dd7dd),
	.w6(32'h3b4d2998),
	.w7(32'h3bd856ea),
	.w8(32'h3ba73cf0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d1690),
	.w1(32'hbb8d3f0c),
	.w2(32'h3a916f2b),
	.w3(32'h3b01c8b4),
	.w4(32'hbb79233c),
	.w5(32'h3aaac2c4),
	.w6(32'hbbe91e08),
	.w7(32'hbb19de70),
	.w8(32'h3b08ed0b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13dff6),
	.w1(32'h3bfe17bd),
	.w2(32'h3bd35425),
	.w3(32'h3ba70c7e),
	.w4(32'h3be57af7),
	.w5(32'h3bc1ac98),
	.w6(32'h3b8c2a68),
	.w7(32'h3bd34f9d),
	.w8(32'h3b3fad67),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5a98e),
	.w1(32'h3bea653e),
	.w2(32'h3be41b01),
	.w3(32'h3b5f35ca),
	.w4(32'h3c98ea6d),
	.w5(32'h3ba3e2f7),
	.w6(32'h3c748f79),
	.w7(32'h3bd2fd7a),
	.w8(32'h3c120758),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2e5f9),
	.w1(32'hbb631901),
	.w2(32'hbb2445e6),
	.w3(32'hbc8aee18),
	.w4(32'h399f39c8),
	.w5(32'hbb2ea1d1),
	.w6(32'h3acad535),
	.w7(32'hbbcafdcb),
	.w8(32'hbb5b88ad),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f7761),
	.w1(32'hbb9b8f8f),
	.w2(32'hbbe8f27b),
	.w3(32'hbbef5f8f),
	.w4(32'h3aee815e),
	.w5(32'hbbb8f95e),
	.w6(32'hbbad2021),
	.w7(32'hbc020939),
	.w8(32'hbba5ae04),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaee4f),
	.w1(32'hbbaf9cb5),
	.w2(32'hbb1d7bea),
	.w3(32'hbbc60e1b),
	.w4(32'hbb9ee7e3),
	.w5(32'hbb45eb8b),
	.w6(32'hbc283c2b),
	.w7(32'hbbbb50bc),
	.w8(32'hbb21f8b6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0f3ce),
	.w1(32'hbab005f5),
	.w2(32'hbbb3cce2),
	.w3(32'h3bc02ebd),
	.w4(32'h3ba07828),
	.w5(32'h3ae288ff),
	.w6(32'hbb66cb69),
	.w7(32'h3a25bf54),
	.w8(32'h39554361),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b533),
	.w1(32'hbbd9e939),
	.w2(32'h3b4d9170),
	.w3(32'h3bc16642),
	.w4(32'hbc0d82d3),
	.w5(32'h3c160a62),
	.w6(32'hbc462a76),
	.w7(32'hbb6a5cd3),
	.w8(32'h392c4e3f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74f9c0),
	.w1(32'h3b1530df),
	.w2(32'hbbb1a9e6),
	.w3(32'hbad731b6),
	.w4(32'h3b93e80b),
	.w5(32'hb86c81cc),
	.w6(32'h3b6dd7ec),
	.w7(32'h3b9bfdca),
	.w8(32'h3b0a5c48),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72ca10),
	.w1(32'h3a0d5b9d),
	.w2(32'hbc16d189),
	.w3(32'h3b6670f5),
	.w4(32'h3c41229c),
	.w5(32'hbaeaad8f),
	.w6(32'h3bec1706),
	.w7(32'h3c888d85),
	.w8(32'h3bd77556),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39c624),
	.w1(32'hbb88b0cb),
	.w2(32'h3b450cfa),
	.w3(32'hbc52fac8),
	.w4(32'hbb37601e),
	.w5(32'hba4d3d8a),
	.w6(32'hbc33730f),
	.w7(32'hbb86cda5),
	.w8(32'hbc0b45f0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc351091),
	.w1(32'hbb93afad),
	.w2(32'hbab0b010),
	.w3(32'hbc15143f),
	.w4(32'hbbde005c),
	.w5(32'hbb5b4a78),
	.w6(32'hbbbcdacf),
	.w7(32'h3b8d676e),
	.w8(32'hbad7f038),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5df47),
	.w1(32'hbbddba7d),
	.w2(32'hbb1b182b),
	.w3(32'h3a5add41),
	.w4(32'hbbf4d41b),
	.w5(32'h3a25e254),
	.w6(32'hbc65a7d2),
	.w7(32'h392425a6),
	.w8(32'h3be2e0ae),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8d011),
	.w1(32'hbb267e7b),
	.w2(32'h3997780f),
	.w3(32'hbb8ade1f),
	.w4(32'hbbd8c9c8),
	.w5(32'hbc074a82),
	.w6(32'hbb0d4fda),
	.w7(32'h3b976b82),
	.w8(32'h3b8e7891),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1c28c),
	.w1(32'h3b0afbcc),
	.w2(32'hbb3c14fa),
	.w3(32'hbc15ee87),
	.w4(32'h3c01d80b),
	.w5(32'hbb2742f7),
	.w6(32'hbb77eb08),
	.w7(32'h3bb228b7),
	.w8(32'h3b5f74aa),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb74918),
	.w1(32'hbc2848fd),
	.w2(32'hbbedc2d0),
	.w3(32'hbb3afe43),
	.w4(32'hbbe6643e),
	.w5(32'hbbaaae01),
	.w6(32'hbbfa97db),
	.w7(32'hbc457c7d),
	.w8(32'hbba2c92a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ec077),
	.w1(32'h3bfda519),
	.w2(32'hbb77e6eb),
	.w3(32'hbbc2d825),
	.w4(32'h3c27b43f),
	.w5(32'hbc2272b3),
	.w6(32'hbc0d0a54),
	.w7(32'hbaa86c1d),
	.w8(32'hbb5f9c0a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f01b5),
	.w1(32'hbaea90ba),
	.w2(32'hbbba96a8),
	.w3(32'hbca7127d),
	.w4(32'h3bba5a87),
	.w5(32'hbb2571bd),
	.w6(32'hbb87eb6a),
	.w7(32'hbc10eeff),
	.w8(32'hbbc8a1db),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d56a8),
	.w1(32'h3ab90430),
	.w2(32'hba94a326),
	.w3(32'h3c9572a5),
	.w4(32'h394bd58e),
	.w5(32'h3b3901a8),
	.w6(32'h3b2e2e20),
	.w7(32'h3baa7d27),
	.w8(32'h3ba1d1c0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b881c37),
	.w1(32'h3c55591d),
	.w2(32'h3c6e2ab8),
	.w3(32'h3ba8e822),
	.w4(32'h3c932b43),
	.w5(32'h3c29b34b),
	.w6(32'h3c54fdb9),
	.w7(32'h3c892e0d),
	.w8(32'h3c8f0f2b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1bc98),
	.w1(32'h3bf36129),
	.w2(32'h3c024410),
	.w3(32'hbbf1b1ec),
	.w4(32'h3bc7ad28),
	.w5(32'h3a3e40af),
	.w6(32'hbac79c88),
	.w7(32'h3b48bb2d),
	.w8(32'hba6e7392),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b394c1c),
	.w1(32'hbaf52aa4),
	.w2(32'hbb1a1f31),
	.w3(32'hbb782d5f),
	.w4(32'hbb81f8aa),
	.w5(32'h3b1cc4d0),
	.w6(32'hbbaaa9ef),
	.w7(32'hbbb1fa32),
	.w8(32'hb9576104),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd607cc),
	.w1(32'hba912c24),
	.w2(32'hbb17707e),
	.w3(32'h3c713113),
	.w4(32'h3bb22d4a),
	.w5(32'h3bed4159),
	.w6(32'hbb02ffe8),
	.w7(32'h3ba1057c),
	.w8(32'h3ba7d041),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ecef1),
	.w1(32'hbc4126ed),
	.w2(32'hbc857a59),
	.w3(32'h3b5c17e3),
	.w4(32'hbbade2d8),
	.w5(32'hbbbe81c4),
	.w6(32'hbc4b96ba),
	.w7(32'hbc34e59d),
	.w8(32'hbc39972d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc882bb8),
	.w1(32'hbba8db04),
	.w2(32'hbba4e7db),
	.w3(32'hbbc6da6a),
	.w4(32'h39f7aa8d),
	.w5(32'h3abcd958),
	.w6(32'hbc354de7),
	.w7(32'hbbb17d60),
	.w8(32'hbb3e5205),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41aa9b),
	.w1(32'hbc469e4f),
	.w2(32'hbc1616d7),
	.w3(32'h3b9f1cf9),
	.w4(32'hbc5dcc65),
	.w5(32'hbbe2a193),
	.w6(32'hbc69fcc7),
	.w7(32'hbc6b7825),
	.w8(32'hbc1b5b90),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50a8e6),
	.w1(32'h3bd1af63),
	.w2(32'hbb886164),
	.w3(32'hbbb6a66e),
	.w4(32'h3b657189),
	.w5(32'hbb72417e),
	.w6(32'h3b22d506),
	.w7(32'hbaee0c30),
	.w8(32'h3988db77),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29a258),
	.w1(32'hba853b5b),
	.w2(32'hbb1995cd),
	.w3(32'hbc6e7c5e),
	.w4(32'h3b49d31d),
	.w5(32'h3b63ef25),
	.w6(32'h3b594703),
	.w7(32'h395cbece),
	.w8(32'hbb8aed4c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa9206),
	.w1(32'hb9b3a476),
	.w2(32'hbacd964d),
	.w3(32'h3a83f25e),
	.w4(32'h3b31588a),
	.w5(32'h3b523af8),
	.w6(32'hba65746f),
	.w7(32'h3a2d5ecc),
	.w8(32'h3976de15),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba14bd7),
	.w1(32'h3af89417),
	.w2(32'hbb3a37b5),
	.w3(32'hbad5ac40),
	.w4(32'h39efa310),
	.w5(32'hbb5a721c),
	.w6(32'hba8c1aeb),
	.w7(32'hbb10b2ca),
	.w8(32'hba8fd143),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb444fba),
	.w1(32'hbc4ac618),
	.w2(32'hbc65fc15),
	.w3(32'hbada384a),
	.w4(32'hbc4449e8),
	.w5(32'hbc7df9c7),
	.w6(32'hbc25ba8d),
	.w7(32'hbc0b0078),
	.w8(32'hbc21f4d2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64466),
	.w1(32'h3add88e9),
	.w2(32'hbb82ff71),
	.w3(32'hbb7da467),
	.w4(32'h3a8ce211),
	.w5(32'h3abb8339),
	.w6(32'h3b8bbec5),
	.w7(32'hba8d0a06),
	.w8(32'hbc14d3bd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc200cd4),
	.w1(32'h3aef23a5),
	.w2(32'hbb8e20f2),
	.w3(32'hbc012d57),
	.w4(32'h3b7fbfdd),
	.w5(32'hbb6b8b66),
	.w6(32'h3b5cf924),
	.w7(32'h3a8065ed),
	.w8(32'h3aaf1ebc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0d634),
	.w1(32'hbbf7b461),
	.w2(32'hbb8eaf16),
	.w3(32'hbabf4506),
	.w4(32'h39d44380),
	.w5(32'h3b2cf46c),
	.w6(32'hbb99d775),
	.w7(32'hbba3f10d),
	.w8(32'hbbf9817d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e2dc5),
	.w1(32'h3afaa5ab),
	.w2(32'h3b0678aa),
	.w3(32'hbab39356),
	.w4(32'h3c249001),
	.w5(32'h3bfdc508),
	.w6(32'hba136f4d),
	.w7(32'h3bed2a5b),
	.w8(32'h3b7d1607),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8344d7),
	.w1(32'hbbf48294),
	.w2(32'hbb266497),
	.w3(32'h3b395000),
	.w4(32'hbb55ba15),
	.w5(32'h395bf07b),
	.w6(32'hbc0ae466),
	.w7(32'hbbbeaf0c),
	.w8(32'hba159ad6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb439d4e),
	.w1(32'hbc2d43cf),
	.w2(32'hbc513d7c),
	.w3(32'hbb0568d4),
	.w4(32'hbc569154),
	.w5(32'hbc6dbc6b),
	.w6(32'hbc9d9e1f),
	.w7(32'hbc692bbb),
	.w8(32'hbc818397),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fc1a1),
	.w1(32'h3ba03d4f),
	.w2(32'hba8d625d),
	.w3(32'hbc0f2241),
	.w4(32'hbc0061a7),
	.w5(32'hbc0b9724),
	.w6(32'h3a5bae1d),
	.w7(32'hbba1929b),
	.w8(32'h396f40e6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22ccea),
	.w1(32'hbc2415c9),
	.w2(32'hbc4df4d8),
	.w3(32'hbb820fd9),
	.w4(32'hb91fc917),
	.w5(32'hbc800253),
	.w6(32'hbc1b1ecb),
	.w7(32'hbc31c0e1),
	.w8(32'hbbf36de3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc061c01),
	.w1(32'hbac39b1c),
	.w2(32'hbbae1be6),
	.w3(32'hbc7d2d43),
	.w4(32'h3b3b5f6c),
	.w5(32'h3b436f4d),
	.w6(32'h38d1d601),
	.w7(32'h3aa39d4b),
	.w8(32'h39df61e2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dbcbc),
	.w1(32'hbbc8dfe6),
	.w2(32'hba185dcc),
	.w3(32'h3a3fadd0),
	.w4(32'hbb944c99),
	.w5(32'hbbc4c407),
	.w6(32'hbc0802b1),
	.w7(32'h3b5296bf),
	.w8(32'hbb93e7d0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule