module layer_10_featuremap_443(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1ed9b),
	.w1(32'hb9353504),
	.w2(32'hba114d52),
	.w3(32'hba53be23),
	.w4(32'hb9b7f9f7),
	.w5(32'h3977c644),
	.w6(32'h39f9a68e),
	.w7(32'hba8e2b7a),
	.w8(32'hba27a121),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f0e1b),
	.w1(32'hbabf91dd),
	.w2(32'hbb516229),
	.w3(32'hba1bf59a),
	.w4(32'hba90b16a),
	.w5(32'hbafe0bbe),
	.w6(32'hba911218),
	.w7(32'hba870d93),
	.w8(32'hbab609bb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95487af),
	.w1(32'hba608242),
	.w2(32'h3884ddb4),
	.w3(32'hb91a5fde),
	.w4(32'hb9e872b3),
	.w5(32'h3ad4cdfd),
	.w6(32'hb994485b),
	.w7(32'hb9ec4010),
	.w8(32'h3abec3c6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a623d2a),
	.w1(32'h3a94258e),
	.w2(32'hb944f48c),
	.w3(32'h39e1a63c),
	.w4(32'h3a19f18c),
	.w5(32'h3a4258a5),
	.w6(32'h3ae7f8be),
	.w7(32'h3ada25aa),
	.w8(32'h3b336327),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3f633),
	.w1(32'h3a6e2105),
	.w2(32'h382b8e1c),
	.w3(32'h3b36cbdd),
	.w4(32'hb8e6e1da),
	.w5(32'h3ac51630),
	.w6(32'h3b2d3334),
	.w7(32'h39c95f48),
	.w8(32'h3a7da7b0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aca3ba),
	.w1(32'h3987b70c),
	.w2(32'h3a224447),
	.w3(32'hb9a8d6ee),
	.w4(32'h3ac9d775),
	.w5(32'h3a3a6095),
	.w6(32'hb954f2ec),
	.w7(32'h3a03745d),
	.w8(32'h391b0c1d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1117d4),
	.w1(32'h39288373),
	.w2(32'hba9cc4c4),
	.w3(32'h3a662410),
	.w4(32'hb9fea29c),
	.w5(32'hbb2c4a9e),
	.w6(32'h3a9f8720),
	.w7(32'hba5f1b6f),
	.w8(32'hbaf0970f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba912146),
	.w1(32'hbad5034b),
	.w2(32'hba456729),
	.w3(32'hbaba8f52),
	.w4(32'hb8b7c0f9),
	.w5(32'h389f102e),
	.w6(32'hba5131e2),
	.w7(32'h39952dc8),
	.w8(32'hbae09728),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba719cd1),
	.w1(32'h3aa90dda),
	.w2(32'h3a229c7c),
	.w3(32'hbaece24f),
	.w4(32'h3938e9bd),
	.w5(32'h3a855af7),
	.w6(32'hba9823a1),
	.w7(32'h38c5dae1),
	.w8(32'h3ab681c7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69b9e1),
	.w1(32'hba409eb1),
	.w2(32'hba09e21a),
	.w3(32'h380a4ccf),
	.w4(32'hba90c270),
	.w5(32'hbabfaf8b),
	.w6(32'h3a3a6b78),
	.w7(32'hba00134c),
	.w8(32'hbac4f754),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84615e),
	.w1(32'hba244100),
	.w2(32'hb9f0f721),
	.w3(32'hbaa3fcd2),
	.w4(32'h38eb8d60),
	.w5(32'h3a43c4ef),
	.w6(32'hbabe8d0a),
	.w7(32'hb942996d),
	.w8(32'hb8c2cda0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c32a1b),
	.w1(32'h3b0c19ac),
	.w2(32'h3b4c758a),
	.w3(32'h3a934186),
	.w4(32'h3b1ea23d),
	.w5(32'h3af15b95),
	.w6(32'h3a3831cc),
	.w7(32'h3b12dd7e),
	.w8(32'h3ab8f4f1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7226bf),
	.w1(32'h3876feaa),
	.w2(32'hba6a60e8),
	.w3(32'h39b3c702),
	.w4(32'hb95b903b),
	.w5(32'hbb7fdda0),
	.w6(32'hb99f27c9),
	.w7(32'hb9c2a10f),
	.w8(32'hbb26a10b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba1d7f),
	.w1(32'hba1bef04),
	.w2(32'hba6d91e9),
	.w3(32'hb9d9ff29),
	.w4(32'hba99d2b7),
	.w5(32'hb9f998d4),
	.w6(32'h3a1b03df),
	.w7(32'hb9fb5776),
	.w8(32'h3a176370),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba857c76),
	.w1(32'hbab381e4),
	.w2(32'h38f49db8),
	.w3(32'hb9db89d4),
	.w4(32'hbb0960bc),
	.w5(32'h3aa1a28e),
	.w6(32'h3a4a0c65),
	.w7(32'hb99fa60e),
	.w8(32'hb872a4b5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7ed4c),
	.w1(32'hba030576),
	.w2(32'h39d9cca7),
	.w3(32'h390e54b9),
	.w4(32'hb90acf87),
	.w5(32'h37de347c),
	.w6(32'hb916d616),
	.w7(32'h3a7dd6ba),
	.w8(32'hb9c9cb18),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8533906),
	.w1(32'hba5f1d42),
	.w2(32'h39f09c9b),
	.w3(32'hba0cf9d0),
	.w4(32'hba6468e1),
	.w5(32'hb986469c),
	.w6(32'hba7fa7d7),
	.w7(32'h3aaeb0d7),
	.w8(32'h3a35f2be),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff6e13),
	.w1(32'hba9989a2),
	.w2(32'hba7a1a88),
	.w3(32'h3a21113a),
	.w4(32'hbab144f9),
	.w5(32'hb9293eea),
	.w6(32'h39d00696),
	.w7(32'hbb1333ca),
	.w8(32'hba940d3a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990f5f2),
	.w1(32'h3901a85d),
	.w2(32'h3ad3f954),
	.w3(32'hba1af9f1),
	.w4(32'hba2c5d4d),
	.w5(32'h3a512f07),
	.w6(32'hbade7301),
	.w7(32'hba571363),
	.w8(32'h38957b01),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395068bd),
	.w1(32'hbaeb0a01),
	.w2(32'hba1815ca),
	.w3(32'hba24f943),
	.w4(32'hbabe7dc2),
	.w5(32'h3a53bfd2),
	.w6(32'hba379c93),
	.w7(32'hb97fd922),
	.w8(32'hb9805aa6),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61e33e),
	.w1(32'h3b138f8d),
	.w2(32'h3b01f087),
	.w3(32'hbac80c06),
	.w4(32'h3afcd52c),
	.w5(32'h3a0061d4),
	.w6(32'hba95113f),
	.w7(32'hb890409f),
	.w8(32'h39a92cfc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86c511),
	.w1(32'hba210d44),
	.w2(32'h39b9df2c),
	.w3(32'h39a27d65),
	.w4(32'h3a88fe66),
	.w5(32'h392e6bda),
	.w6(32'h3ab1f480),
	.w7(32'h3b0b7f8f),
	.w8(32'hba4380af),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadadac8),
	.w1(32'hbab8e37b),
	.w2(32'hbab957b1),
	.w3(32'hbb1a7c46),
	.w4(32'h3a00dff5),
	.w5(32'hba13f241),
	.w6(32'hbb0631e8),
	.w7(32'hba2e5743),
	.w8(32'hb9cf7842),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac794ab),
	.w1(32'h3a0cb613),
	.w2(32'h39a17579),
	.w3(32'hba49ac7d),
	.w4(32'hbaa3a3eb),
	.w5(32'hbb169ae6),
	.w6(32'hb9ec2c0c),
	.w7(32'h39cd8091),
	.w8(32'hba7e4ee6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bdc97),
	.w1(32'hbaaa99f5),
	.w2(32'hba27e50e),
	.w3(32'hbb468a24),
	.w4(32'hbb1664b7),
	.w5(32'h3a5838a5),
	.w6(32'hbae3ac08),
	.w7(32'hbb314eac),
	.w8(32'hba80a82b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6f68d),
	.w1(32'hb87d9d1a),
	.w2(32'h3a515477),
	.w3(32'hba88fd31),
	.w4(32'h3978bf93),
	.w5(32'hb95e0aa1),
	.w6(32'hba79b4de),
	.w7(32'hb990ed3a),
	.w8(32'hbb0aed18),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2004d),
	.w1(32'h3b15872c),
	.w2(32'hb9d7c163),
	.w3(32'hb9abb1ec),
	.w4(32'h3a016ab2),
	.w5(32'hbae4ecae),
	.w6(32'hbb2929c9),
	.w7(32'h394078ac),
	.w8(32'hba9ffdac),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cc1f5),
	.w1(32'hba289dbd),
	.w2(32'hba01ba56),
	.w3(32'hbb04d6ef),
	.w4(32'hba70629d),
	.w5(32'hba31c728),
	.w6(32'hb95e1560),
	.w7(32'hba11d9fd),
	.w8(32'hb9a1e24a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d3d2d6),
	.w1(32'hb8ee02a7),
	.w2(32'hbb11a653),
	.w3(32'hb93f021a),
	.w4(32'hbaa3d9d1),
	.w5(32'hbac00317),
	.w6(32'hb8f877d2),
	.w7(32'hba91cfc3),
	.w8(32'hbb0af6be),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac37d36),
	.w1(32'h3a92192a),
	.w2(32'h3a8fd2f5),
	.w3(32'hb8bc0304),
	.w4(32'h3abb3450),
	.w5(32'h3a7c79a6),
	.w6(32'hb9e9f7cb),
	.w7(32'h3a4625be),
	.w8(32'h3a75a65d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85acda),
	.w1(32'hba0d7852),
	.w2(32'h3a1a0c5f),
	.w3(32'hb98dd34f),
	.w4(32'hba68e73a),
	.w5(32'hbaff458d),
	.w6(32'h3a1ad844),
	.w7(32'hb918cf9d),
	.w8(32'hbb17a658),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6c263),
	.w1(32'hbab0e4b6),
	.w2(32'hba8fa10e),
	.w3(32'hbb016cfb),
	.w4(32'hb9451928),
	.w5(32'h3a5389b1),
	.w6(32'hbb1de2be),
	.w7(32'h393ee898),
	.w8(32'h3a9a7763),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4b47e),
	.w1(32'hbad14c00),
	.w2(32'hb985ad56),
	.w3(32'h3ad291b4),
	.w4(32'h398278dd),
	.w5(32'h39de6587),
	.w6(32'h3ab69795),
	.w7(32'hb9517954),
	.w8(32'h3a056560),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab14777),
	.w1(32'hba83b72f),
	.w2(32'h3986188f),
	.w3(32'hbaf37f13),
	.w4(32'hb98e653d),
	.w5(32'hba31e492),
	.w6(32'hba0c132d),
	.w7(32'hba2a3ba1),
	.w8(32'hb95d85e8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba083d26),
	.w1(32'hbad95c2d),
	.w2(32'h39ba4a0c),
	.w3(32'hb950d8d5),
	.w4(32'hb9920137),
	.w5(32'h3a8b3aa6),
	.w6(32'h37f6643c),
	.w7(32'h3aac8317),
	.w8(32'h3ad11218),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba628727),
	.w1(32'h399d6798),
	.w2(32'h3a2d8a5b),
	.w3(32'hb991e3ae),
	.w4(32'h3992306c),
	.w5(32'h3a2370c2),
	.w6(32'h3a992120),
	.w7(32'h3a37a306),
	.w8(32'h3a421096),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaace739),
	.w1(32'h3a6ea259),
	.w2(32'hbad7eee4),
	.w3(32'hbab18b26),
	.w4(32'hb86f35bb),
	.w5(32'hba38b50a),
	.w6(32'hbaeed679),
	.w7(32'hba6c6d83),
	.w8(32'hba087cc2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20f0d2),
	.w1(32'hbb037758),
	.w2(32'hbad3bffc),
	.w3(32'hba9e8a23),
	.w4(32'h393e4b67),
	.w5(32'h3a83dcfd),
	.w6(32'h3a6681da),
	.w7(32'h3a29d460),
	.w8(32'h3a1bfb2a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a73c0),
	.w1(32'hba82c810),
	.w2(32'hb97aebed),
	.w3(32'h3ae981ed),
	.w4(32'hbb06b201),
	.w5(32'h3a35506b),
	.w6(32'h3a49c5fc),
	.w7(32'hba853997),
	.w8(32'hb9d21de1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfc0d3),
	.w1(32'hbade731c),
	.w2(32'hb95b8594),
	.w3(32'hb8847386),
	.w4(32'hba1dc52e),
	.w5(32'h39d244ad),
	.w6(32'h39d3e398),
	.w7(32'hba31ff71),
	.w8(32'h38ee1c02),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1af427),
	.w1(32'h3a6c1f5f),
	.w2(32'hba213944),
	.w3(32'h3ab99074),
	.w4(32'hba9ebd40),
	.w5(32'hbb0d1d4e),
	.w6(32'h37b65689),
	.w7(32'hb9b67b61),
	.w8(32'hba2762dd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c7bee),
	.w1(32'h3980625f),
	.w2(32'hb9c249ab),
	.w3(32'h3a183566),
	.w4(32'hba826979),
	.w5(32'hbade7c11),
	.w6(32'hba964c6f),
	.w7(32'hba2c90ac),
	.w8(32'hba7158c7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0d6dc),
	.w1(32'hba831613),
	.w2(32'hbb28152a),
	.w3(32'hb9d66d63),
	.w4(32'hbad30c0d),
	.w5(32'hba91332f),
	.w6(32'hb9a937e5),
	.w7(32'hb90daa60),
	.w8(32'h3939fe95),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99503b0),
	.w1(32'h3ac85078),
	.w2(32'h37bbf136),
	.w3(32'h3a97b69e),
	.w4(32'h3ab0ed94),
	.w5(32'h3a0dddb7),
	.w6(32'h39f2f520),
	.w7(32'h39abac6b),
	.w8(32'h3aa95de9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abeeb21),
	.w1(32'h3929cfb8),
	.w2(32'h3a0f6f4b),
	.w3(32'h3b307d99),
	.w4(32'hb93fdea8),
	.w5(32'h3a17af37),
	.w6(32'h3b4c4d44),
	.w7(32'h3847fff6),
	.w8(32'h39a417a7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fca5df),
	.w1(32'hba093b41),
	.w2(32'hbab21816),
	.w3(32'hba537308),
	.w4(32'hb9ff69ea),
	.w5(32'hba505169),
	.w6(32'hba999a5e),
	.w7(32'h396f7d5c),
	.w8(32'hbb006275),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd1c97),
	.w1(32'hb8d0dd6d),
	.w2(32'h39b3b1d5),
	.w3(32'hbb22b6cb),
	.w4(32'hbad90bcf),
	.w5(32'hbac2ad38),
	.w6(32'hbaea1b26),
	.w7(32'hb9aeb928),
	.w8(32'hba7a6838),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc526e),
	.w1(32'hbb1d299c),
	.w2(32'hba8a1c1a),
	.w3(32'h3ad9a153),
	.w4(32'hbb151528),
	.w5(32'hba660bc6),
	.w6(32'h3a8d7b7f),
	.w7(32'hbb26d074),
	.w8(32'hbae717a3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb177521),
	.w1(32'h37749f25),
	.w2(32'h3a1d2721),
	.w3(32'hbacf51d1),
	.w4(32'hb9735617),
	.w5(32'h3a2d95fe),
	.w6(32'hbaa038dc),
	.w7(32'hb90aea3f),
	.w8(32'h39a52ac5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6e0a0),
	.w1(32'hba83f0ff),
	.w2(32'h3a294e00),
	.w3(32'hbb0fd9f6),
	.w4(32'hba3aeeb7),
	.w5(32'h38bda917),
	.w6(32'hbb111f84),
	.w7(32'hba657cc6),
	.w8(32'h38f263be),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afec432),
	.w1(32'h39b0d43d),
	.w2(32'hba376f37),
	.w3(32'h3a779e3e),
	.w4(32'hb9c19e06),
	.w5(32'hba93c2da),
	.w6(32'hba210ae2),
	.w7(32'h3a0f76c2),
	.w8(32'hb97d5f5b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e5692),
	.w1(32'hba3b5f5e),
	.w2(32'hba6dc7ce),
	.w3(32'h3a680a39),
	.w4(32'h3a6fab87),
	.w5(32'hb9817401),
	.w6(32'hb99a4ea7),
	.w7(32'h3a9b2a26),
	.w8(32'h3a630197),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81d61e),
	.w1(32'h39e53918),
	.w2(32'h3ae4241a),
	.w3(32'hba7809af),
	.w4(32'h3adaf0c8),
	.w5(32'h3aa80881),
	.w6(32'hba1d4733),
	.w7(32'h3a80d3b5),
	.w8(32'h399e56af),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89e1c7),
	.w1(32'hb980a9a7),
	.w2(32'h39602309),
	.w3(32'hb9dfd72d),
	.w4(32'h3a96af2d),
	.w5(32'h3ac92fc6),
	.w6(32'hb9fc105c),
	.w7(32'h395a4e1f),
	.w8(32'h3a7eeaf8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38ac15),
	.w1(32'hbafa889b),
	.w2(32'h391a55be),
	.w3(32'hba60eb9b),
	.w4(32'hba6c3023),
	.w5(32'h3aaedd38),
	.w6(32'h393fe6ee),
	.w7(32'hb9512502),
	.w8(32'h378205fb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba163824),
	.w1(32'hbac1f4e7),
	.w2(32'hba9fcef3),
	.w3(32'hb9f2560e),
	.w4(32'hbad63d2e),
	.w5(32'h3a6d17af),
	.w6(32'hba0c3d4e),
	.w7(32'hbac1eb09),
	.w8(32'hbad7d2c9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7a545),
	.w1(32'h3a5f51aa),
	.w2(32'h3892977b),
	.w3(32'hb9aa6020),
	.w4(32'hb8701ea8),
	.w5(32'hba814751),
	.w6(32'hba26c451),
	.w7(32'hba4f9cd4),
	.w8(32'hba477817),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976aa79),
	.w1(32'hb8d01980),
	.w2(32'hbafc07c2),
	.w3(32'hba3499b6),
	.w4(32'h3a967c7f),
	.w5(32'hba809c21),
	.w6(32'h3878bccd),
	.w7(32'h39e1c543),
	.w8(32'hbae431e1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac39d6f),
	.w1(32'h388f8a4e),
	.w2(32'hbb1291bf),
	.w3(32'hba82b3a1),
	.w4(32'hb91f58fd),
	.w5(32'hbabad9b2),
	.w6(32'hbae6ed23),
	.w7(32'h38813d8d),
	.w8(32'hbac3102d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa0444),
	.w1(32'hbad96435),
	.w2(32'h3a8cfff3),
	.w3(32'h388c4abd),
	.w4(32'hbaeaeb7b),
	.w5(32'h3aa01d50),
	.w6(32'h39390119),
	.w7(32'hb8c0d4f6),
	.w8(32'hba60174e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80002a),
	.w1(32'h37e2c59c),
	.w2(32'hba469749),
	.w3(32'h39fe7b42),
	.w4(32'hbaece023),
	.w5(32'hba799f73),
	.w6(32'hba777a43),
	.w7(32'hb8a43afc),
	.w8(32'hba1c3598),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaac78f),
	.w1(32'hbaa6da61),
	.w2(32'hba50b9f2),
	.w3(32'hbac9d5d2),
	.w4(32'hbad82467),
	.w5(32'hb8e98c15),
	.w6(32'hba896bf4),
	.w7(32'hbaa38ecf),
	.w8(32'hba3f35d6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24b93a),
	.w1(32'hbb1738c5),
	.w2(32'hbb39c10d),
	.w3(32'hb9dfc680),
	.w4(32'hbb720f9a),
	.w5(32'hbafbc24a),
	.w6(32'hba77ad08),
	.w7(32'hbad4e70c),
	.w8(32'hbaaa5840),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7c1e7),
	.w1(32'h3b06edb0),
	.w2(32'h3ad78e7b),
	.w3(32'hba33375b),
	.w4(32'h3a88acf0),
	.w5(32'h3ab4eb8b),
	.w6(32'hbad958c4),
	.w7(32'h398085fb),
	.w8(32'h3a851333),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af74904),
	.w1(32'h3ad70cc5),
	.w2(32'h3b07b17e),
	.w3(32'h3a58f7b7),
	.w4(32'h3b04ed9b),
	.w5(32'h3b0af680),
	.w6(32'hba59bbd1),
	.w7(32'h3b1ec6d1),
	.w8(32'h3b357232),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b271653),
	.w1(32'h3a894025),
	.w2(32'h39c5d401),
	.w3(32'h3b1eae98),
	.w4(32'hb9f2b8bd),
	.w5(32'hba9ab207),
	.w6(32'h3b09453a),
	.w7(32'hba1e18d0),
	.w8(32'hbad720c7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba562fe7),
	.w1(32'hb7c7cd98),
	.w2(32'h3ad403ee),
	.w3(32'hba5cd6cd),
	.w4(32'h39af6b24),
	.w5(32'h39ddabad),
	.w6(32'hb9eb7c7f),
	.w7(32'hb37af2c0),
	.w8(32'hb855cee7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41db87),
	.w1(32'hba977252),
	.w2(32'hbad1a2b6),
	.w3(32'hba825931),
	.w4(32'hbb42a323),
	.w5(32'hbb392d46),
	.w6(32'hba6e3569),
	.w7(32'hbb1de86e),
	.w8(32'hbb2225fb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad97dd6),
	.w1(32'hbaf24a41),
	.w2(32'hbb23a3fd),
	.w3(32'hbb10359d),
	.w4(32'hbb1acdbf),
	.w5(32'hba83bd04),
	.w6(32'hbb082ba5),
	.w7(32'hba67b405),
	.w8(32'hb9e1bf16),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53cc07),
	.w1(32'h3b6077fb),
	.w2(32'hbb87a022),
	.w3(32'hbaf15bbf),
	.w4(32'hbae71012),
	.w5(32'hbaa4c087),
	.w6(32'hba446790),
	.w7(32'h392fbcc8),
	.w8(32'hbb0e3a2a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6caf0),
	.w1(32'hbb6b549c),
	.w2(32'h3a803a0d),
	.w3(32'hbb42c2eb),
	.w4(32'hbc507ad9),
	.w5(32'hbb744c16),
	.w6(32'h3b096659),
	.w7(32'hbbe4bae3),
	.w8(32'hbaa8e645),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7a8e0),
	.w1(32'hbb897617),
	.w2(32'hbbb36295),
	.w3(32'hbb8dbce9),
	.w4(32'hb9d57462),
	.w5(32'hbbfca44c),
	.w6(32'hbb9757c4),
	.w7(32'hbb641bd5),
	.w8(32'hba812054),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8b283),
	.w1(32'h3bbdd18a),
	.w2(32'h3a5d84af),
	.w3(32'hbbd27116),
	.w4(32'h3baa4101),
	.w5(32'h3be7b7b7),
	.w6(32'hbbb96148),
	.w7(32'hbb453dd6),
	.w8(32'h3ae43836),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40142a),
	.w1(32'hbb1dd30d),
	.w2(32'hbb23f479),
	.w3(32'hbb65492a),
	.w4(32'h3a3d8f55),
	.w5(32'hbb64085f),
	.w6(32'h3ae5b0e0),
	.w7(32'hba0d5742),
	.w8(32'hb8120386),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9878e6),
	.w1(32'hbb51216b),
	.w2(32'hbb788f13),
	.w3(32'h3ba46864),
	.w4(32'hbaf85551),
	.w5(32'hbb4b5689),
	.w6(32'h3a409385),
	.w7(32'hbb73f1e1),
	.w8(32'hbb331bfe),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babb389),
	.w1(32'hba8f8639),
	.w2(32'hbb281e43),
	.w3(32'hbbbb24db),
	.w4(32'h3b0eee27),
	.w5(32'hbaa52370),
	.w6(32'hbaa60363),
	.w7(32'h3a52c27f),
	.w8(32'h3b70429e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b9ddb),
	.w1(32'hbbc07db5),
	.w2(32'hbb9bfaaa),
	.w3(32'hba9c542e),
	.w4(32'hbc0e0fcf),
	.w5(32'hbbbbd256),
	.w6(32'h3b86defb),
	.w7(32'hbae994b2),
	.w8(32'hba9ebf1b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea5f50),
	.w1(32'hbb9052cd),
	.w2(32'h3c1a87ef),
	.w3(32'h3baa8d08),
	.w4(32'h3b07010e),
	.w5(32'h3b2ecddb),
	.w6(32'h3be5383b),
	.w7(32'h3b46e3ca),
	.w8(32'h3c58a144),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80cc89),
	.w1(32'hba7f9eba),
	.w2(32'h3b11f708),
	.w3(32'h3a007586),
	.w4(32'hbbb9656b),
	.w5(32'h3b8528bb),
	.w6(32'hbb20d15c),
	.w7(32'hbbb4b9e6),
	.w8(32'hbb0e1137),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97d980),
	.w1(32'h3b39aa89),
	.w2(32'h39caca49),
	.w3(32'hbba31b9d),
	.w4(32'h3b89e0f5),
	.w5(32'h3a92d758),
	.w6(32'hbb12a1e8),
	.w7(32'h3bdb865e),
	.w8(32'h3ad590e6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26ea27),
	.w1(32'h3b57cb7a),
	.w2(32'h3a1281bb),
	.w3(32'h3c4d700a),
	.w4(32'hbb2a8838),
	.w5(32'hbb48ce49),
	.w6(32'h3aea7208),
	.w7(32'h3a9332fa),
	.w8(32'h3a57b646),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc4e2f),
	.w1(32'h3ba21251),
	.w2(32'h3c264e40),
	.w3(32'h3b60b71d),
	.w4(32'h3ae0920e),
	.w5(32'h3bc6f078),
	.w6(32'h3bd34b5c),
	.w7(32'h3b5f3386),
	.w8(32'h3be0a913),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f5512),
	.w1(32'h3ade67a2),
	.w2(32'h3b7968c7),
	.w3(32'h3bb9cc66),
	.w4(32'h396c2787),
	.w5(32'h3b990677),
	.w6(32'h3af8993b),
	.w7(32'hbace5998),
	.w8(32'h3b3c699b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1d383),
	.w1(32'hba80217f),
	.w2(32'hbbd065a1),
	.w3(32'h3bbdb23b),
	.w4(32'hbb56aacc),
	.w5(32'hbbd89714),
	.w6(32'h3b75af76),
	.w7(32'hb90bf9b2),
	.w8(32'hbb79fd9c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb128c54),
	.w1(32'h3b00cb00),
	.w2(32'h3c2cf0ae),
	.w3(32'hbbf7685c),
	.w4(32'h3b59c447),
	.w5(32'h3c22d9e5),
	.w6(32'hbb147088),
	.w7(32'hba920709),
	.w8(32'h3c468eee),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad33d14),
	.w1(32'hba7147f4),
	.w2(32'h3bbbdb96),
	.w3(32'h3ab5cc44),
	.w4(32'h34b642e5),
	.w5(32'h39ca6525),
	.w6(32'hba3dc1b7),
	.w7(32'hbb038f4d),
	.w8(32'hbc4e7d13),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb131e66),
	.w1(32'hbb0c0b7b),
	.w2(32'hbacd12f8),
	.w3(32'hbbd861e5),
	.w4(32'hbb78dbd6),
	.w5(32'h3a930942),
	.w6(32'hbbbb2b5d),
	.w7(32'h3a81d48e),
	.w8(32'hb958fa8a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b667deb),
	.w1(32'h3b0e7f95),
	.w2(32'h3a44cbe0),
	.w3(32'h3bf59076),
	.w4(32'hbb8c4daa),
	.w5(32'h3c02ea61),
	.w6(32'h3b391923),
	.w7(32'hbb7e97ac),
	.w8(32'h3a92d6f7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43e898),
	.w1(32'hbbdea449),
	.w2(32'hbbfed6e5),
	.w3(32'h3a032b04),
	.w4(32'hbbef06cd),
	.w5(32'hbc075280),
	.w6(32'hba56cd0b),
	.w7(32'hbb57dde5),
	.w8(32'hbb9c4ed2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13c3c2),
	.w1(32'h3bb11099),
	.w2(32'h3b5733c4),
	.w3(32'hbb477e9e),
	.w4(32'hba8d5c94),
	.w5(32'hbbb467dd),
	.w6(32'h39ec4ad9),
	.w7(32'h3c1bd498),
	.w8(32'hbb9bbbb2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb225f9b),
	.w1(32'hbae43456),
	.w2(32'hbb8862ae),
	.w3(32'hbaa01072),
	.w4(32'h3af6fe61),
	.w5(32'h3b0d0617),
	.w6(32'hbbced2e7),
	.w7(32'h3bf74940),
	.w8(32'h3c054918),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b136ef3),
	.w1(32'h3c2e066c),
	.w2(32'h3b4aa92c),
	.w3(32'h3bb82854),
	.w4(32'h3b8fd0fc),
	.w5(32'hbac5668f),
	.w6(32'h3be72b48),
	.w7(32'h3c1d36fc),
	.w8(32'h3b248061),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9331901),
	.w1(32'hbb4c4082),
	.w2(32'hbb8fcbd2),
	.w3(32'h3a0bde45),
	.w4(32'hbb8f7fc5),
	.w5(32'hbbc20118),
	.w6(32'h3b9c8080),
	.w7(32'hbbd83271),
	.w8(32'hbc1352f6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc08f9c),
	.w1(32'hb8c4b7e7),
	.w2(32'hbb4ae74f),
	.w3(32'hbbab4f57),
	.w4(32'h3b34500c),
	.w5(32'h38d59732),
	.w6(32'hbb71c97a),
	.w7(32'hbb28030e),
	.w8(32'hbb4126b5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3ca52),
	.w1(32'hba141685),
	.w2(32'hbb9b151d),
	.w3(32'hbbaca668),
	.w4(32'h3abefb54),
	.w5(32'hbb99f981),
	.w6(32'hb9e866ee),
	.w7(32'hbb6fb147),
	.w8(32'hbb152d73),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d7f16),
	.w1(32'hbbc1bd1d),
	.w2(32'hbc79d3e7),
	.w3(32'hbb11db5a),
	.w4(32'hbb22acc3),
	.w5(32'hbc3e5135),
	.w6(32'hbbaf0543),
	.w7(32'hbac9e70b),
	.w8(32'hbbf94dd0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40da1f),
	.w1(32'h3b247342),
	.w2(32'h3bcae41f),
	.w3(32'h3b196921),
	.w4(32'h39a03d49),
	.w5(32'h3bad8cad),
	.w6(32'h3ab71284),
	.w7(32'h3ade0de6),
	.w8(32'h3b71048b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8621d6),
	.w1(32'h3bea0f16),
	.w2(32'h3b692cc7),
	.w3(32'h3a92191a),
	.w4(32'h3ae5b3c5),
	.w5(32'hbb827045),
	.w6(32'hbac99d2d),
	.w7(32'h3a93dd65),
	.w8(32'h3b4d27dd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd24b65),
	.w1(32'h3943026e),
	.w2(32'hbbbd3461),
	.w3(32'h3c3fc598),
	.w4(32'h3b2d80e7),
	.w5(32'hbb9eb541),
	.w6(32'h3ad97507),
	.w7(32'h3c2fa09d),
	.w8(32'hba7ee035),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5af54),
	.w1(32'hbb2f38fa),
	.w2(32'h3c0f9361),
	.w3(32'hbab29833),
	.w4(32'h3aaa0c9c),
	.w5(32'h3ba913a4),
	.w6(32'hbacf9299),
	.w7(32'hbb920e36),
	.w8(32'h3b2b1538),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4565d2),
	.w1(32'hbb45668a),
	.w2(32'hbb99c3af),
	.w3(32'h3bdb0d6a),
	.w4(32'h380a0369),
	.w5(32'hbb43baf9),
	.w6(32'h3b627681),
	.w7(32'hba64a7f0),
	.w8(32'h3a7c56e2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a029dcf),
	.w1(32'hbaaef7b3),
	.w2(32'h3bc6ae9d),
	.w3(32'h3a86b890),
	.w4(32'hba0104da),
	.w5(32'h3b7279f5),
	.w6(32'h3b9a3156),
	.w7(32'hba3aa66f),
	.w8(32'h3afb2fca),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e4aff),
	.w1(32'hb89fc480),
	.w2(32'hbba2a8d0),
	.w3(32'hbaa4eaa4),
	.w4(32'h3b3a413b),
	.w5(32'hbbe9cb48),
	.w6(32'hbbc4273b),
	.w7(32'h3adb65e0),
	.w8(32'h3b65d0bd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4977f),
	.w1(32'hba74afd0),
	.w2(32'h3c23104c),
	.w3(32'h3bb7d8ae),
	.w4(32'h39926103),
	.w5(32'h3c1432d7),
	.w6(32'h3b205909),
	.w7(32'h3b5517f9),
	.w8(32'h3c234e8c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9b208),
	.w1(32'hbb93a70d),
	.w2(32'hb9af0263),
	.w3(32'hbacabd86),
	.w4(32'hbbf911ec),
	.w5(32'h3a01f179),
	.w6(32'h3ac21766),
	.w7(32'hbbe6d624),
	.w8(32'hbb7aac2d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4a2ec),
	.w1(32'h3b39280b),
	.w2(32'h3b8b0f67),
	.w3(32'h390c4312),
	.w4(32'h3b1ced56),
	.w5(32'h3bb3f02d),
	.w6(32'h3802f8fc),
	.w7(32'h3b21f719),
	.w8(32'h3b4efcb3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc1d99),
	.w1(32'h3b11088f),
	.w2(32'h3bfae0b2),
	.w3(32'h3bc04c18),
	.w4(32'hbbe1f3b3),
	.w5(32'hbab169d7),
	.w6(32'h3b9dd546),
	.w7(32'hbb459492),
	.w8(32'hbada5ab6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eec87),
	.w1(32'h3b30ebd4),
	.w2(32'hbbb07f79),
	.w3(32'hbb9210c0),
	.w4(32'h3b3a7365),
	.w5(32'h3a4497f5),
	.w6(32'hbb3a5e21),
	.w7(32'h3aab0b7d),
	.w8(32'hbb86334e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e89cfc),
	.w1(32'h3a2bb6a3),
	.w2(32'h3b25e121),
	.w3(32'hbb857ea0),
	.w4(32'h3b5eb30d),
	.w5(32'h3ab2a65b),
	.w6(32'hba90f6c4),
	.w7(32'h3bd746e2),
	.w8(32'h3b731e49),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c54d1),
	.w1(32'h3b9a68cb),
	.w2(32'hbb30ea81),
	.w3(32'h3be5ad6c),
	.w4(32'h3b30f873),
	.w5(32'hbaf2bf3b),
	.w6(32'h3bdc58df),
	.w7(32'hbb194c47),
	.w8(32'hbb42ee1e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad191b7),
	.w1(32'h3b807a56),
	.w2(32'hbad06588),
	.w3(32'h3bdf79e5),
	.w4(32'h3bb90f00),
	.w5(32'h3afbb871),
	.w6(32'hb956ae08),
	.w7(32'h3bc1d4c9),
	.w8(32'hbaff4565),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dc7bf),
	.w1(32'h3ba7b041),
	.w2(32'h3c50f6db),
	.w3(32'hba807ab1),
	.w4(32'h3c25e90d),
	.w5(32'h3a7be673),
	.w6(32'hbb265fef),
	.w7(32'h3c25b8e1),
	.w8(32'h3be6a45c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07dbc),
	.w1(32'h3b77cbf2),
	.w2(32'h3af6cfec),
	.w3(32'h3b5ff9c7),
	.w4(32'h3b07e45f),
	.w5(32'h3abcba15),
	.w6(32'h3b05acad),
	.w7(32'hba77c4fa),
	.w8(32'h3ae89667),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91218e),
	.w1(32'hbb708766),
	.w2(32'h3c033ca9),
	.w3(32'h3bfbe629),
	.w4(32'h3a93097d),
	.w5(32'hba8a0f72),
	.w6(32'h3b39ad55),
	.w7(32'h3af92fec),
	.w8(32'h3b90cf18),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64ed10),
	.w1(32'hbb69149d),
	.w2(32'hbb300928),
	.w3(32'h3b38a27f),
	.w4(32'hbb19c47e),
	.w5(32'hbb8df664),
	.w6(32'h3beb5b2a),
	.w7(32'hbb9a276a),
	.w8(32'hba9c178f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c090a68),
	.w1(32'h390a901a),
	.w2(32'h3bd106fa),
	.w3(32'h3bf9bba8),
	.w4(32'h39787e5c),
	.w5(32'h3c5f8f64),
	.w6(32'h38333474),
	.w7(32'h3ba4ab72),
	.w8(32'h3c1990e6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4b916),
	.w1(32'h3b42df2e),
	.w2(32'hbac6d63e),
	.w3(32'h3b3c3fcf),
	.w4(32'h3b0e758a),
	.w5(32'h3a469d82),
	.w6(32'h3b8c7958),
	.w7(32'hb9ea01ed),
	.w8(32'hbac140ed),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c138606),
	.w1(32'h39df0a8c),
	.w2(32'h3b81109e),
	.w3(32'h3c35daf4),
	.w4(32'h3c2075a4),
	.w5(32'hba31b570),
	.w6(32'h3b74494e),
	.w7(32'h3be9dffd),
	.w8(32'h3c0ce5fb),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdd041),
	.w1(32'hbada2bc6),
	.w2(32'hbc05656a),
	.w3(32'h3bf275a2),
	.w4(32'hbb885667),
	.w5(32'hbbe7124e),
	.w6(32'h3c3cf828),
	.w7(32'hbb511e84),
	.w8(32'hbba651c1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29c573),
	.w1(32'hba63fef0),
	.w2(32'hbba00f83),
	.w3(32'hbb9b9343),
	.w4(32'h3ab1e3f3),
	.w5(32'hbbf893f7),
	.w6(32'hbbb9e973),
	.w7(32'hbb098e99),
	.w8(32'hbb8a4ef6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1ddb6),
	.w1(32'hbb82e67a),
	.w2(32'hbb3dda53),
	.w3(32'hba0438a3),
	.w4(32'hbbe73098),
	.w5(32'h3b001904),
	.w6(32'hba03ec1f),
	.w7(32'hbbabc661),
	.w8(32'h3b52a96b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b6f9a),
	.w1(32'hbc248fef),
	.w2(32'hbbea9f94),
	.w3(32'h3ad01981),
	.w4(32'hbc0b0a7f),
	.w5(32'hbb82c885),
	.w6(32'h3a074fcd),
	.w7(32'h3a7f9d66),
	.w8(32'hbb592ac1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac9d29),
	.w1(32'h3acd931f),
	.w2(32'h3bf3ebf9),
	.w3(32'hbbc46bc4),
	.w4(32'hbbb165a5),
	.w5(32'h3b931954),
	.w6(32'hba910bb7),
	.w7(32'hbb028961),
	.w8(32'h3bf47393),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2edb8d),
	.w1(32'hbb59ce14),
	.w2(32'h3992898f),
	.w3(32'h3c0ea037),
	.w4(32'hbb8d22ea),
	.w5(32'hbb917dc9),
	.w6(32'h3bdfbd70),
	.w7(32'hbba4a05e),
	.w8(32'hbb319cc4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8002d),
	.w1(32'hbba7c663),
	.w2(32'h3adf23f0),
	.w3(32'hbb4ef60f),
	.w4(32'h3bb1cf7e),
	.w5(32'hbb80657a),
	.w6(32'hbb27f863),
	.w7(32'h3a569054),
	.w8(32'h3bd2c7b6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48b668),
	.w1(32'hbad57f4e),
	.w2(32'h3a4972aa),
	.w3(32'hbb1e7147),
	.w4(32'hbbd282f1),
	.w5(32'hbaec4ac9),
	.w6(32'h39959a22),
	.w7(32'hbba98de2),
	.w8(32'hbaa77b44),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13667e),
	.w1(32'hbaf60136),
	.w2(32'hbc046b60),
	.w3(32'hbad38198),
	.w4(32'h3b5f1078),
	.w5(32'hbb6b1ff7),
	.w6(32'h3a613c72),
	.w7(32'h3bdea40f),
	.w8(32'h3bda528e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b5cfc),
	.w1(32'hbb6d7c6a),
	.w2(32'hbb5fef31),
	.w3(32'hb9c53d3f),
	.w4(32'hbaaf0c8f),
	.w5(32'hba815b2b),
	.w6(32'h3b4e2b96),
	.w7(32'h39ce392c),
	.w8(32'hbbcefcee),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd82713),
	.w1(32'hbb7bf473),
	.w2(32'hbbb741a1),
	.w3(32'hbb85228a),
	.w4(32'hbb077d09),
	.w5(32'hbaf8a7c4),
	.w6(32'hbb8e55b0),
	.w7(32'hba26a906),
	.w8(32'hbb80cc16),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46c4d8),
	.w1(32'h3a807959),
	.w2(32'h3b96d86f),
	.w3(32'h3b7d4811),
	.w4(32'hbb02eb4c),
	.w5(32'hb9dfad16),
	.w6(32'h3b2b4b8f),
	.w7(32'hba8f04c4),
	.w8(32'h3b752745),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc373c6),
	.w1(32'h38673b2b),
	.w2(32'hba1d72c3),
	.w3(32'hbbd581b3),
	.w4(32'h3b3ab7fc),
	.w5(32'h3a20a98c),
	.w6(32'hbb8f0e1d),
	.w7(32'hb9703a89),
	.w8(32'h3b4cecab),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f270d),
	.w1(32'hbb5b01f4),
	.w2(32'hb9b2d727),
	.w3(32'h3afc178b),
	.w4(32'hbb839e65),
	.w5(32'h3985dd83),
	.w6(32'h39da9c94),
	.w7(32'h3abcebf3),
	.w8(32'h3b8e5a91),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dfa8d),
	.w1(32'h3a604bcf),
	.w2(32'hbab0df4d),
	.w3(32'hbb51e3bc),
	.w4(32'hb99a027b),
	.w5(32'hbb5a7265),
	.w6(32'h3b97182c),
	.w7(32'h3b25f390),
	.w8(32'hbb02d0a9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f4867),
	.w1(32'hba804bbd),
	.w2(32'h3b4020b9),
	.w3(32'hbb20bb1d),
	.w4(32'h3be7d32b),
	.w5(32'hbb09a04b),
	.w6(32'hbba88fa7),
	.w7(32'hbb420e3c),
	.w8(32'h3bd0ca1f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2348de),
	.w1(32'hbbf2ab7a),
	.w2(32'hbbf3d5b6),
	.w3(32'h3af8a90b),
	.w4(32'hbadb6ebb),
	.w5(32'hbb883819),
	.w6(32'h3aa4d790),
	.w7(32'hbbb5ae5f),
	.w8(32'hbbc79611),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6484865),
	.w1(32'h3b41e641),
	.w2(32'hbb2d35cf),
	.w3(32'hba4cc400),
	.w4(32'h3bbe9023),
	.w5(32'h3a6d1ea0),
	.w6(32'hbb39283b),
	.w7(32'h3a55a534),
	.w8(32'h3b13e30c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f828),
	.w1(32'hbb0bb258),
	.w2(32'h3b90e4d6),
	.w3(32'hbb0bd317),
	.w4(32'hba143a78),
	.w5(32'hba0242c1),
	.w6(32'h39be2bf1),
	.w7(32'h39a7cde3),
	.w8(32'hba1750a2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf10e41),
	.w1(32'hba332606),
	.w2(32'h3ab34029),
	.w3(32'h3c024b35),
	.w4(32'h3badee46),
	.w5(32'h3b3b0e72),
	.w6(32'h3be561d2),
	.w7(32'h3a834a13),
	.w8(32'h3b8e7f02),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0c274),
	.w1(32'h3b057232),
	.w2(32'h3aea5302),
	.w3(32'hba49bef4),
	.w4(32'h3b167e33),
	.w5(32'h3ba767b3),
	.w6(32'h3b3eb734),
	.w7(32'hba91e9e9),
	.w8(32'h3b01a7db),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa0bb6),
	.w1(32'hb9a57dae),
	.w2(32'h3b1fd5fc),
	.w3(32'h3b0844db),
	.w4(32'hbba2fe78),
	.w5(32'hbaffc2da),
	.w6(32'h3b89958a),
	.w7(32'hbb82dbc6),
	.w8(32'h3a88c2ff),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b211a40),
	.w1(32'h3b1223c7),
	.w2(32'h3c869353),
	.w3(32'h3a2eb481),
	.w4(32'hbbb73b44),
	.w5(32'h3c766b7f),
	.w6(32'hbab022bd),
	.w7(32'hbb1395fd),
	.w8(32'h3c4588d8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f4d19),
	.w1(32'h3a63b034),
	.w2(32'h3ad4ff25),
	.w3(32'h3b61e24d),
	.w4(32'h3b50f6af),
	.w5(32'h3b0dab49),
	.w6(32'h3bbbab35),
	.w7(32'h3b210fa4),
	.w8(32'h3b94ba05),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922a163),
	.w1(32'hbab570b3),
	.w2(32'h3c6693da),
	.w3(32'h3bbe54ac),
	.w4(32'h3a335454),
	.w5(32'h3bcc633f),
	.w6(32'h3bb2dd7d),
	.w7(32'hbb3bc829),
	.w8(32'h3c0758c5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca6f66),
	.w1(32'h3a00fbd4),
	.w2(32'h3c3776f1),
	.w3(32'h3baf6a70),
	.w4(32'hbb2ebae7),
	.w5(32'h3c1b29a6),
	.w6(32'h3abc9b35),
	.w7(32'hb9c3fb62),
	.w8(32'h3bf1c6a2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25ff92),
	.w1(32'hbba1146d),
	.w2(32'h3ab08e41),
	.w3(32'h3b3871fe),
	.w4(32'hbbbea96a),
	.w5(32'hbbff9760),
	.w6(32'h3b38175b),
	.w7(32'h3ae473c8),
	.w8(32'hbba48a5f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68338b),
	.w1(32'hbb3aed3e),
	.w2(32'hbc1fe278),
	.w3(32'hbb140d7c),
	.w4(32'h3a384080),
	.w5(32'hbb8fb569),
	.w6(32'hbbb91ef4),
	.w7(32'h3b16ad0f),
	.w8(32'hbae55a19),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38944e99),
	.w1(32'hbaac16d6),
	.w2(32'h3bb4737e),
	.w3(32'hbb0f64f2),
	.w4(32'h3a044d3b),
	.w5(32'h39a77838),
	.w6(32'h3bcc14d6),
	.w7(32'h3a9dfd64),
	.w8(32'h3ba1fcad),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e3c1a),
	.w1(32'h3ab251d0),
	.w2(32'h3bac20f4),
	.w3(32'hb9504f51),
	.w4(32'hbb618360),
	.w5(32'h3c669fed),
	.w6(32'hbaeba490),
	.w7(32'h3a3d9e20),
	.w8(32'h3be10b33),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96eb0f),
	.w1(32'hbb4035b7),
	.w2(32'h3b754392),
	.w3(32'h3b5b3113),
	.w4(32'hbbd9d418),
	.w5(32'hbbd3c0b9),
	.w6(32'h3c342a98),
	.w7(32'hbbf24403),
	.w8(32'hbbaadbf1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53cc5b),
	.w1(32'hbab42add),
	.w2(32'h3c4a9bf3),
	.w3(32'hbba36c66),
	.w4(32'hbb843516),
	.w5(32'h3c4fca90),
	.w6(32'hbbb12914),
	.w7(32'hba60aa6b),
	.w8(32'h3c6bcc9f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba1276),
	.w1(32'hbb263f54),
	.w2(32'h3b791a72),
	.w3(32'h3aa2d966),
	.w4(32'h3b2a1d4d),
	.w5(32'h3b0f1842),
	.w6(32'hbbd44354),
	.w7(32'hbba31fca),
	.w8(32'hbb1f1559),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d2660),
	.w1(32'hbac6b1fc),
	.w2(32'hbbbbb77b),
	.w3(32'hbbf1c966),
	.w4(32'hbbbb1625),
	.w5(32'hbc5a8eb1),
	.w6(32'hbbdcb811),
	.w7(32'h39c4b73f),
	.w8(32'hbb4ba1ad),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db78d),
	.w1(32'h3b1f7dca),
	.w2(32'hbc15ef00),
	.w3(32'hbc000ef2),
	.w4(32'h3b55c739),
	.w5(32'hbb63cd70),
	.w6(32'h3ab2b63d),
	.w7(32'h3aa0d53c),
	.w8(32'hbb53568a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee4e1c),
	.w1(32'h3bdcf62a),
	.w2(32'h3b9e06fa),
	.w3(32'hba18e0b8),
	.w4(32'hbb3621b0),
	.w5(32'h3b3f18fb),
	.w6(32'h3a2836df),
	.w7(32'h3ade1ff5),
	.w8(32'h3983e368),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959c3e2),
	.w1(32'hbbf1cdee),
	.w2(32'h3b81200b),
	.w3(32'hbb32208e),
	.w4(32'hbb128f32),
	.w5(32'h3b48a48d),
	.w6(32'h3aadb973),
	.w7(32'hbb7013fe),
	.w8(32'h381909f9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79326b),
	.w1(32'h3b34430e),
	.w2(32'hbb854c04),
	.w3(32'h3ba18d48),
	.w4(32'h3b95a7ad),
	.w5(32'hbb3964e6),
	.w6(32'h3918d00e),
	.w7(32'hbb09b002),
	.w8(32'hbbd1a2e6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5b878),
	.w1(32'hbc32eda5),
	.w2(32'hbb99338b),
	.w3(32'hbb9df6ab),
	.w4(32'hbb9e6656),
	.w5(32'hbba11fff),
	.w6(32'hbb787e03),
	.w7(32'hbbf060a4),
	.w8(32'hbafad25e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b2375),
	.w1(32'h3bb55a9f),
	.w2(32'h3b9c4c35),
	.w3(32'hbb4522b7),
	.w4(32'h3aaf3691),
	.w5(32'hb9a4458a),
	.w6(32'hbad8ccab),
	.w7(32'h3abdf33a),
	.w8(32'h3a0cc7a4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74d609),
	.w1(32'hbb4d0705),
	.w2(32'h3a1d5cd4),
	.w3(32'hbb8b665e),
	.w4(32'h3b3dea14),
	.w5(32'h3bf3cef3),
	.w6(32'hbaa20f62),
	.w7(32'hbb355ebf),
	.w8(32'hbbc92f0b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958fe95),
	.w1(32'h385aa04e),
	.w2(32'h3b8f2e0e),
	.w3(32'h3b9a97a1),
	.w4(32'hbb260e3c),
	.w5(32'h3ab1b207),
	.w6(32'hba78f2d5),
	.w7(32'hbacfd6ef),
	.w8(32'h3bbde52c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d1bb9),
	.w1(32'hba5b3285),
	.w2(32'h3b7be2b1),
	.w3(32'h3ab1de7e),
	.w4(32'h38feb0e4),
	.w5(32'h39586e92),
	.w6(32'h3ac83d5f),
	.w7(32'h3a249b6e),
	.w8(32'h3b7047bf),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1615c3),
	.w1(32'hbb6f07ed),
	.w2(32'h3b5fc7de),
	.w3(32'h3adaa37c),
	.w4(32'h3b474736),
	.w5(32'h3ba46c49),
	.w6(32'h3baa5e0c),
	.w7(32'h3a2476bc),
	.w8(32'h3a94bbac),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31793e),
	.w1(32'hbaf82618),
	.w2(32'hb990fb7f),
	.w3(32'h3b9cbc21),
	.w4(32'h3ae43697),
	.w5(32'hbb42b417),
	.w6(32'h3bd0f153),
	.w7(32'h39f183e5),
	.w8(32'h39a4f6b2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74e151),
	.w1(32'hbba576ae),
	.w2(32'hbbae5b10),
	.w3(32'h3b8dee46),
	.w4(32'hbb60dc05),
	.w5(32'hbbb4e7d6),
	.w6(32'h3b1b6199),
	.w7(32'hbb6a8f53),
	.w8(32'hbba7b4a0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9194719),
	.w1(32'h3b5b885d),
	.w2(32'h3b0399fc),
	.w3(32'hbaddd320),
	.w4(32'h3be08035),
	.w5(32'h3c36585d),
	.w6(32'hbb344243),
	.w7(32'h3b0714f1),
	.w8(32'h3bb1259c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5332b6),
	.w1(32'h3a9bb07d),
	.w2(32'h3bd8df37),
	.w3(32'hbb945e80),
	.w4(32'hba9dd548),
	.w5(32'h3bb3a2c6),
	.w6(32'hba900546),
	.w7(32'hba80c261),
	.w8(32'h3bbdcf24),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae81129),
	.w1(32'hbbaf4769),
	.w2(32'hbc54a406),
	.w3(32'hb9d31e43),
	.w4(32'hbb1a1bad),
	.w5(32'hbc0e978d),
	.w6(32'hbb0a1cea),
	.w7(32'hbbaf2d37),
	.w8(32'hbbf4e1ea),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dbe02),
	.w1(32'hbb7e3dad),
	.w2(32'hbb66de38),
	.w3(32'h3bef6af3),
	.w4(32'hbbb66924),
	.w5(32'h3713b55d),
	.w6(32'hbadd6d4c),
	.w7(32'hbbc270c5),
	.w8(32'hbb1f73d8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb06de),
	.w1(32'h3a9859f6),
	.w2(32'h3be0e6c3),
	.w3(32'hbba59793),
	.w4(32'h3ae7accd),
	.w5(32'h3abf7f30),
	.w6(32'hbb20e7f6),
	.w7(32'hbaf070de),
	.w8(32'h3b40cad0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affd5bf),
	.w1(32'hb952fd0c),
	.w2(32'h3be16011),
	.w3(32'h3b83b81d),
	.w4(32'h3a91327b),
	.w5(32'h3b88c518),
	.w6(32'h3b888f9b),
	.w7(32'hbba5e60c),
	.w8(32'hb9963ef3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba285129),
	.w1(32'hba52b59b),
	.w2(32'h3be679df),
	.w3(32'h3a9de99f),
	.w4(32'hbb7fda6b),
	.w5(32'h3bca8dc3),
	.w6(32'hbab3b7fd),
	.w7(32'h3b5c10f3),
	.w8(32'h3b4d10d5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba202608),
	.w1(32'hbbdf24e4),
	.w2(32'hbbc70367),
	.w3(32'hbb091e39),
	.w4(32'hbb016089),
	.w5(32'hbba295cc),
	.w6(32'hbb10dd92),
	.w7(32'hbac5e9d3),
	.w8(32'hbb30dd20),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b902b99),
	.w1(32'h3ac61c9d),
	.w2(32'hbafad684),
	.w3(32'h3bf82d60),
	.w4(32'hb84a56f3),
	.w5(32'h3a525599),
	.w6(32'h3c066851),
	.w7(32'hbb55663c),
	.w8(32'hbb7878eb),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89e7f5),
	.w1(32'h3a6e798b),
	.w2(32'hba42be06),
	.w3(32'hbb97bb15),
	.w4(32'hbb668d7c),
	.w5(32'hbb7f93d1),
	.w6(32'hbb48a801),
	.w7(32'h3a5dbb6a),
	.w8(32'hba90d851),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4c0f6),
	.w1(32'h3abf1329),
	.w2(32'hbabb1437),
	.w3(32'hbb38177b),
	.w4(32'hbb7686c8),
	.w5(32'h3b27865d),
	.w6(32'hbb1fb360),
	.w7(32'hbbff069c),
	.w8(32'hbbef588f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7084c4),
	.w1(32'hbb4daf57),
	.w2(32'hbbcbc908),
	.w3(32'hbb652f72),
	.w4(32'h399ee6c8),
	.w5(32'hbb1b860b),
	.w6(32'hbbd4cf50),
	.w7(32'h3a81f94b),
	.w8(32'hbb273062),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f6dd0),
	.w1(32'hbb4e8272),
	.w2(32'hbbb283b5),
	.w3(32'h3b29bcce),
	.w4(32'hbbb83edd),
	.w5(32'hbbeb991c),
	.w6(32'h3b3eab59),
	.w7(32'hbb03a6ac),
	.w8(32'hbbea7949),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb95f8),
	.w1(32'hbabbdc2e),
	.w2(32'hbb99fa58),
	.w3(32'hbbb671e5),
	.w4(32'hbacb6da8),
	.w5(32'hbb9945cc),
	.w6(32'hbbc2b1e5),
	.w7(32'hbb66f171),
	.w8(32'hbb5772ef),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91185d),
	.w1(32'hba9c08c7),
	.w2(32'h3b31b583),
	.w3(32'hbbac1186),
	.w4(32'hbb55bba7),
	.w5(32'hb92912e0),
	.w6(32'hbb9ea25e),
	.w7(32'h3b35c9dd),
	.w8(32'h3ac18b6f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e99ac),
	.w1(32'hbad1be59),
	.w2(32'h3bcdb5aa),
	.w3(32'h3c1ec2ef),
	.w4(32'hbb02255c),
	.w5(32'h3b28e8ae),
	.w6(32'h3b829618),
	.w7(32'hbb7bc14b),
	.w8(32'h3a173d9e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c38b1),
	.w1(32'h38a738ae),
	.w2(32'hbbaee4f9),
	.w3(32'h3c4272d1),
	.w4(32'h3b11f969),
	.w5(32'hbb6224f1),
	.w6(32'h3abee9c8),
	.w7(32'hbb8df72b),
	.w8(32'hbbd635bb),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccfe0d),
	.w1(32'hb9f23902),
	.w2(32'h3b2f33c0),
	.w3(32'hba241af5),
	.w4(32'h39608230),
	.w5(32'h3b97ec49),
	.w6(32'hb98234f6),
	.w7(32'hbb7acb1f),
	.w8(32'h378a8bd5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5298a9),
	.w1(32'hb9a83a60),
	.w2(32'hba25d812),
	.w3(32'hb975a5e2),
	.w4(32'hb917a394),
	.w5(32'h3c2d7c92),
	.w6(32'h3b3d11f5),
	.w7(32'h3aa0432a),
	.w8(32'h3c39ba6e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaa213),
	.w1(32'hba081380),
	.w2(32'h3b478390),
	.w3(32'hbb7f311d),
	.w4(32'hbbb56e2d),
	.w5(32'hba2fe741),
	.w6(32'hbb89aeba),
	.w7(32'hbb88d90b),
	.w8(32'h39c22788),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e74bb),
	.w1(32'h3b02aee2),
	.w2(32'h3b8fa1c5),
	.w3(32'hb99ec07e),
	.w4(32'h3ab22fb0),
	.w5(32'hbb6bb996),
	.w6(32'h3b2de656),
	.w7(32'h3b8f1dfc),
	.w8(32'h3af9b2c0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9c4f4),
	.w1(32'h3be35fca),
	.w2(32'h3c2fc4d2),
	.w3(32'h3b97dfc4),
	.w4(32'h3b7afc31),
	.w5(32'h3b69bd6d),
	.w6(32'h3a901800),
	.w7(32'h3b3b1923),
	.w8(32'h3c31c074),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d132f),
	.w1(32'hbb6308ac),
	.w2(32'h3aa1cb81),
	.w3(32'h3b872895),
	.w4(32'hbb94ff62),
	.w5(32'h3bbe9183),
	.w6(32'h3baf5034),
	.w7(32'h3b53c65a),
	.w8(32'h36cdaae1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7971ac),
	.w1(32'h3bc035b8),
	.w2(32'hbc0aa3a1),
	.w3(32'hb9b57bf7),
	.w4(32'h3b81f69b),
	.w5(32'hbb4c41c0),
	.w6(32'hbb3dd10e),
	.w7(32'hbb500d73),
	.w8(32'hba025b30),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03beba),
	.w1(32'h3b84c604),
	.w2(32'hbb1ad823),
	.w3(32'hbb104801),
	.w4(32'hba19ef40),
	.w5(32'hbb4c48bf),
	.w6(32'hbc15ae77),
	.w7(32'h3a2e8f65),
	.w8(32'hbb1a9e2d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa59a0e),
	.w1(32'h3a797654),
	.w2(32'hbb3bc439),
	.w3(32'hbb8d5c69),
	.w4(32'h382d828d),
	.w5(32'hbb80be0d),
	.w6(32'hbba225bf),
	.w7(32'hbb2e546e),
	.w8(32'h3a6aa319),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39d73f),
	.w1(32'hbbb4343a),
	.w2(32'hbc22bc65),
	.w3(32'hbaa26e17),
	.w4(32'hbb7f9d98),
	.w5(32'hbbb3af8c),
	.w6(32'hba809c17),
	.w7(32'hba0cd9e7),
	.w8(32'hba90bf2c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf52cf5),
	.w1(32'h398ddb63),
	.w2(32'h3b5a2510),
	.w3(32'hbbe51c09),
	.w4(32'hbb5ab639),
	.w5(32'h3b41a08a),
	.w6(32'hbb1066c4),
	.w7(32'hbb0c371f),
	.w8(32'h3b37f812),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfa680),
	.w1(32'h3bc506e7),
	.w2(32'h3c0b3e9c),
	.w3(32'h3bcb8c4d),
	.w4(32'h3b06b1ed),
	.w5(32'h3a5d428b),
	.w6(32'h3b8e1c7b),
	.w7(32'h3b85f4a3),
	.w8(32'h3b8aab9f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f4c18),
	.w1(32'hbb9d5c4b),
	.w2(32'hbc2de58a),
	.w3(32'h3bde28eb),
	.w4(32'hbb90a779),
	.w5(32'hbc0c4546),
	.w6(32'h3c11743e),
	.w7(32'hbb7cf072),
	.w8(32'hbc17fb5c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52e58),
	.w1(32'h3b67f42e),
	.w2(32'hbaa80d3f),
	.w3(32'hbb9bab1e),
	.w4(32'h3bb4153c),
	.w5(32'h3bb15269),
	.w6(32'hbc0af11f),
	.w7(32'h3c0b6810),
	.w8(32'h3b0fb360),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91120c),
	.w1(32'h3aa8f5f9),
	.w2(32'hbbc8ff62),
	.w3(32'h3c4558fe),
	.w4(32'hbad07d0b),
	.w5(32'hb9bae64b),
	.w6(32'h3bec568c),
	.w7(32'h3c1d2eb2),
	.w8(32'h3b385703),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d1161),
	.w1(32'hbc265416),
	.w2(32'hbbc386a5),
	.w3(32'h3c002fc1),
	.w4(32'hbb5bc5c2),
	.w5(32'hbb24d6ff),
	.w6(32'h3c1bfed5),
	.w7(32'hbad131dd),
	.w8(32'hbb1d67ac),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8adfda),
	.w1(32'h3b0b7f94),
	.w2(32'h3b788880),
	.w3(32'h3b31b85f),
	.w4(32'hbaa2d095),
	.w5(32'h3b0bd0c9),
	.w6(32'hb6a38d91),
	.w7(32'h3ab50b54),
	.w8(32'hbc0c0de0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936c225),
	.w1(32'hbb680442),
	.w2(32'hbbc5825b),
	.w3(32'h3a919029),
	.w4(32'hbb69edd3),
	.w5(32'hba38794d),
	.w6(32'hbb6f8059),
	.w7(32'hbb81e54d),
	.w8(32'hb91739d0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade38ef),
	.w1(32'hb91e0d27),
	.w2(32'hbb807f08),
	.w3(32'hbb2fe796),
	.w4(32'hbc05d530),
	.w5(32'hbc016cb3),
	.w6(32'h398a7837),
	.w7(32'hbb2412fc),
	.w8(32'h3a315e0b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb282108),
	.w1(32'hbbf234bf),
	.w2(32'hbb3c3ff0),
	.w3(32'hbb009286),
	.w4(32'hbb568609),
	.w5(32'hbb865396),
	.w6(32'hbb1abd9c),
	.w7(32'h39a296bd),
	.w8(32'hbc0784aa),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b05c3),
	.w1(32'h399b0d90),
	.w2(32'hbb4bf265),
	.w3(32'h3b6b74bf),
	.w4(32'hbb37e9e9),
	.w5(32'hbb622b93),
	.w6(32'hbb6e923b),
	.w7(32'hbaca1425),
	.w8(32'hbad0e999),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62afbc),
	.w1(32'hbbb33223),
	.w2(32'hbad551cb),
	.w3(32'h39ea5ab7),
	.w4(32'hba020406),
	.w5(32'hbb1478b0),
	.w6(32'hbb55c593),
	.w7(32'hbb2b9d5b),
	.w8(32'hbaf9db2c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b4337),
	.w1(32'hbada86ab),
	.w2(32'hbbba4261),
	.w3(32'hbba50ec2),
	.w4(32'hba8fd3b3),
	.w5(32'hbb2a59e8),
	.w6(32'hbae35aa6),
	.w7(32'h3a497daa),
	.w8(32'h3b04a759),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884e0e1),
	.w1(32'h3a6dcddc),
	.w2(32'h3b8a4e94),
	.w3(32'h3b6d6f84),
	.w4(32'h3a940626),
	.w5(32'hb9125f00),
	.w6(32'h3a6c033c),
	.w7(32'h3a9a2be1),
	.w8(32'h3b16f3ee),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d21b0),
	.w1(32'hbbad5f48),
	.w2(32'hbb561c90),
	.w3(32'h3a2c1161),
	.w4(32'hbb322658),
	.w5(32'hbb1d7399),
	.w6(32'hbbdb39d2),
	.w7(32'hbbf9dc98),
	.w8(32'hbc247225),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3b924),
	.w1(32'hbb626d98),
	.w2(32'h3ab3c15a),
	.w3(32'hbb94e845),
	.w4(32'h3903436e),
	.w5(32'h3b23d5e8),
	.w6(32'hbbb4faa7),
	.w7(32'h3b17c2b5),
	.w8(32'h3bc7b9a0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06940b),
	.w1(32'hbbb89a92),
	.w2(32'hbbbd4280),
	.w3(32'h3b4d53cd),
	.w4(32'hbbd627b9),
	.w5(32'hb9c89bc3),
	.w6(32'hbb3d47b8),
	.w7(32'hbaf78740),
	.w8(32'hbb8015aa),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaacfae),
	.w1(32'h3c11a17b),
	.w2(32'h3bb1cc57),
	.w3(32'hbb1d4870),
	.w4(32'h3ad9932d),
	.w5(32'h3b9bf635),
	.w6(32'hbb3c04ce),
	.w7(32'h3c0b7e56),
	.w8(32'h3c36b245),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b591726),
	.w1(32'h3a8c3511),
	.w2(32'h39ea88c9),
	.w3(32'h3c162d96),
	.w4(32'hba69d7fb),
	.w5(32'h3bcdd29f),
	.w6(32'h3bdfa809),
	.w7(32'h3b1f55df),
	.w8(32'h3ba5f7ee),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e2f88),
	.w1(32'h3b3d402d),
	.w2(32'h3a5275d7),
	.w3(32'h3b485930),
	.w4(32'hbb11c370),
	.w5(32'hbb868eb3),
	.w6(32'h3b09dac3),
	.w7(32'hbb0ed491),
	.w8(32'h3972a687),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44cce4),
	.w1(32'hba381ee5),
	.w2(32'h3b857d96),
	.w3(32'hbb53aa1f),
	.w4(32'h3a9a6763),
	.w5(32'h3c6f4e0f),
	.w6(32'hbb6ee6b9),
	.w7(32'h3ad5da75),
	.w8(32'hba2e8d44),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bd9f0),
	.w1(32'hbb8d598f),
	.w2(32'hbb363207),
	.w3(32'hbb43287e),
	.w4(32'hbb4eef95),
	.w5(32'hbb4c955f),
	.w6(32'h3b8865b9),
	.w7(32'hbb1d9520),
	.w8(32'hbaf5464f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e2ada),
	.w1(32'hbb44594d),
	.w2(32'h3becd43b),
	.w3(32'hbb2262ee),
	.w4(32'h3be0ec75),
	.w5(32'hbc2fd216),
	.w6(32'hbb2a2263),
	.w7(32'h3b381bcf),
	.w8(32'hbad76b53),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48a083),
	.w1(32'hbbcf896f),
	.w2(32'hbbc916eb),
	.w3(32'hbaf21213),
	.w4(32'h3ad471e5),
	.w5(32'hbb50fcf9),
	.w6(32'hba3358dc),
	.w7(32'hbb464028),
	.w8(32'hbb93b192),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb78d),
	.w1(32'hbb115078),
	.w2(32'hbb8c41f2),
	.w3(32'hbbc99b95),
	.w4(32'h38b84980),
	.w5(32'hbb6f03e7),
	.w6(32'hbb8596e8),
	.w7(32'hbb383479),
	.w8(32'hba728bed),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2782f4),
	.w1(32'h3b4e62b6),
	.w2(32'h3b5fe5c9),
	.w3(32'hbb0069e0),
	.w4(32'h3a49192b),
	.w5(32'h3b262c72),
	.w6(32'h3b5c7d00),
	.w7(32'hbb79350f),
	.w8(32'h3a1a4f56),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967618),
	.w1(32'hbac9e533),
	.w2(32'hbb33616a),
	.w3(32'hbb052ff4),
	.w4(32'hbadd9394),
	.w5(32'hbb028068),
	.w6(32'hbb86023f),
	.w7(32'hbb5b4dcf),
	.w8(32'hbb980da0),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba871b09),
	.w1(32'h3917cf51),
	.w2(32'hbb0fda59),
	.w3(32'hb8b799bb),
	.w4(32'hbb04d08e),
	.w5(32'hbb1c4bb5),
	.w6(32'hb970eb4f),
	.w7(32'h3b17862d),
	.w8(32'h3b848aa4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6be283),
	.w1(32'h3b62e79f),
	.w2(32'h3bc684ca),
	.w3(32'hbafca8cc),
	.w4(32'h3c2e87ac),
	.w5(32'hbb7630a1),
	.w6(32'hbaeb692c),
	.w7(32'hbb950b41),
	.w8(32'h3a6fdba2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc308d),
	.w1(32'h3b399ce0),
	.w2(32'h3b1fc397),
	.w3(32'hbb710f19),
	.w4(32'h3b1faa10),
	.w5(32'h3afb1b17),
	.w6(32'hb8ff8a18),
	.w7(32'h3bc54d2b),
	.w8(32'h3b721d04),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b164f11),
	.w1(32'h3a0a0f3b),
	.w2(32'h3b2b9728),
	.w3(32'h3ba1debb),
	.w4(32'hbb3d4cbd),
	.w5(32'h3a249628),
	.w6(32'h3995ea70),
	.w7(32'h3a58b5df),
	.w8(32'h3ad5d681),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc9cce),
	.w1(32'hbb666bba),
	.w2(32'hbbf9cde6),
	.w3(32'h3b350c33),
	.w4(32'h3b771e70),
	.w5(32'h3b9d0983),
	.w6(32'h3b4275d5),
	.w7(32'hbc0292a7),
	.w8(32'hbb8c1458),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3104e),
	.w1(32'hbbe7baa2),
	.w2(32'hbbda60da),
	.w3(32'hbb46700f),
	.w4(32'hbbbe0077),
	.w5(32'hbbf8165c),
	.w6(32'hbbaec127),
	.w7(32'hbbba5b45),
	.w8(32'hbbc3bbb3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd556),
	.w1(32'h3ae2f31e),
	.w2(32'h3ae8e672),
	.w3(32'h3a1311da),
	.w4(32'hba4a39e7),
	.w5(32'h3a05d28b),
	.w6(32'hbb579821),
	.w7(32'hba79b90c),
	.w8(32'hbb05c344),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a7173),
	.w1(32'hb89ef5a9),
	.w2(32'hbb8a3955),
	.w3(32'h3b261352),
	.w4(32'hbb09f399),
	.w5(32'hbaa6a4f6),
	.w6(32'hbab4e6fb),
	.w7(32'hba346ee2),
	.w8(32'h3af18cea),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11f5d8),
	.w1(32'hbb12f0d5),
	.w2(32'hbbc0d3f2),
	.w3(32'h3c152002),
	.w4(32'hbc009d37),
	.w5(32'h3b6b3b34),
	.w6(32'h3c0b58ac),
	.w7(32'hb9d1203a),
	.w8(32'h3b8092c9),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03315d),
	.w1(32'hbb524ed7),
	.w2(32'hbb7c1f78),
	.w3(32'hbb32f6ca),
	.w4(32'hbb2cc5ef),
	.w5(32'hbb8958e4),
	.w6(32'hbc50080c),
	.w7(32'hb8c9dc31),
	.w8(32'h3a3e4686),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba679dd9),
	.w1(32'h3a28655d),
	.w2(32'h3ae64a31),
	.w3(32'hbbc56947),
	.w4(32'h3ba5ee7e),
	.w5(32'h3be2ffbd),
	.w6(32'hbb87e0b2),
	.w7(32'h3b6a7936),
	.w8(32'h3b99cffc),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab17f32),
	.w1(32'hba9b84e3),
	.w2(32'hb9fde90f),
	.w3(32'h3c050a68),
	.w4(32'hbb82845d),
	.w5(32'hbb0c8dac),
	.w6(32'h3a5b752b),
	.w7(32'hbb28a30c),
	.w8(32'hbb081405),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8906b6),
	.w1(32'hba48d58b),
	.w2(32'hbb16b00b),
	.w3(32'h3a92768a),
	.w4(32'hbb2efce2),
	.w5(32'hbb51c004),
	.w6(32'h3a8448f6),
	.w7(32'hbb3f2df5),
	.w8(32'h3a9bbcf7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb6abe),
	.w1(32'hbb592b4c),
	.w2(32'hb9b69b7b),
	.w3(32'h3ab5c748),
	.w4(32'hbb60b377),
	.w5(32'hbb7b3988),
	.w6(32'hb9a41029),
	.w7(32'hbba11f99),
	.w8(32'hbb50db0a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55f1ba),
	.w1(32'h3b007930),
	.w2(32'h3af3a8b3),
	.w3(32'h3b15f3d7),
	.w4(32'hbacd26af),
	.w5(32'h3a4b25fe),
	.w6(32'hbba8ad6b),
	.w7(32'hb90f3976),
	.w8(32'h3b8d62ad),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba85b43),
	.w1(32'h3a8ce60b),
	.w2(32'h3b86ed03),
	.w3(32'h39981731),
	.w4(32'h3b93ef1c),
	.w5(32'h3bc7843e),
	.w6(32'hbb24eff0),
	.w7(32'h3be448db),
	.w8(32'h3bcf6981),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02cc74),
	.w1(32'h3b4ed245),
	.w2(32'h39847374),
	.w3(32'h3b15b0d8),
	.w4(32'h3b18a27e),
	.w5(32'hbb10b0d7),
	.w6(32'h3b223b8b),
	.w7(32'hb98e8863),
	.w8(32'hbabfaff2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb140765),
	.w1(32'hbaa42cf8),
	.w2(32'hbb39c19e),
	.w3(32'hbb71344b),
	.w4(32'hbb23b478),
	.w5(32'hbb07dddc),
	.w6(32'hbb201c7c),
	.w7(32'hbb914514),
	.w8(32'hbb8d441f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54035b),
	.w1(32'h3b80ab29),
	.w2(32'h3b1f80a8),
	.w3(32'hbbd2fb50),
	.w4(32'hbb6ed3f9),
	.w5(32'hbb1be464),
	.w6(32'hbbc17d16),
	.w7(32'h3bac41b4),
	.w8(32'h39850688),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b622950),
	.w1(32'hbb4a1a5e),
	.w2(32'hbb916fff),
	.w3(32'h3b84ec7e),
	.w4(32'h3ae1a597),
	.w5(32'hba6b41f4),
	.w6(32'h3acacb39),
	.w7(32'hbb94e41e),
	.w8(32'hbbd16905),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9715a4),
	.w1(32'h3be79c31),
	.w2(32'hba48fc9b),
	.w3(32'hbb5837f3),
	.w4(32'h3b1b3871),
	.w5(32'hba118d2e),
	.w6(32'hbb92e6ad),
	.w7(32'hbb45c9a9),
	.w8(32'hbb8c09ad),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff87d0),
	.w1(32'h3782db02),
	.w2(32'h3b822895),
	.w3(32'h3b01ce87),
	.w4(32'hbb9db42d),
	.w5(32'hbaf7608b),
	.w6(32'hbb060003),
	.w7(32'hbb775c8f),
	.w8(32'h3b17704a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b177abe),
	.w1(32'hb98c7657),
	.w2(32'hbb5aa593),
	.w3(32'h3b64bb0c),
	.w4(32'hbaa8dbb1),
	.w5(32'hbad67da6),
	.w6(32'h3ab0553d),
	.w7(32'hba2df2b8),
	.w8(32'h3a6a9d1b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f8582),
	.w1(32'hbab65bcb),
	.w2(32'h39296d57),
	.w3(32'h3be149ef),
	.w4(32'h3b17c7c7),
	.w5(32'hbb88899f),
	.w6(32'h3b90ec4c),
	.w7(32'h39d9d4f2),
	.w8(32'h3aa6d515),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d4339),
	.w1(32'h3a321452),
	.w2(32'h3899b936),
	.w3(32'h3b623f8a),
	.w4(32'h3b7126d9),
	.w5(32'hbb733494),
	.w6(32'h39e1feb7),
	.w7(32'hbac19f0a),
	.w8(32'h3b1f3836),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83a42b),
	.w1(32'hbbf150e2),
	.w2(32'hbb1eede3),
	.w3(32'h3a457794),
	.w4(32'hbbfb6916),
	.w5(32'h3b6d262a),
	.w6(32'hbb042183),
	.w7(32'hbab81a23),
	.w8(32'hba9ac2e4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf92066),
	.w1(32'hbada6a13),
	.w2(32'h3b39ebd7),
	.w3(32'hbae2cf39),
	.w4(32'h3ba05b27),
	.w5(32'hbb07cd96),
	.w6(32'hbb990c7a),
	.w7(32'h3bbdfff2),
	.w8(32'hba9df312),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ac45c),
	.w1(32'hbb4225b9),
	.w2(32'h3a6bf4dc),
	.w3(32'hbb932ce4),
	.w4(32'hbb9e6aa8),
	.w5(32'hb98b3c0b),
	.w6(32'hbb637603),
	.w7(32'hba428c82),
	.w8(32'h3be85b84),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908ec48),
	.w1(32'hbb8de5e8),
	.w2(32'hbbf2d8ce),
	.w3(32'h3b538ea0),
	.w4(32'hbb7b295b),
	.w5(32'hbbdad358),
	.w6(32'h3b9b100a),
	.w7(32'hbb2e95e0),
	.w8(32'hbbb2bea1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8140cb),
	.w1(32'h3a54a1f0),
	.w2(32'hbb405c62),
	.w3(32'hbbaf5c2d),
	.w4(32'hb952fa27),
	.w5(32'hbb1cbc44),
	.w6(32'hbbab9007),
	.w7(32'hba8e2513),
	.w8(32'hbb616961),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9b65f),
	.w1(32'hbadc9a7f),
	.w2(32'h3b01dff0),
	.w3(32'hba7ae5d2),
	.w4(32'hb9d6fd33),
	.w5(32'hbb4cbf91),
	.w6(32'hbabee68f),
	.w7(32'hbb428729),
	.w8(32'hba1764aa),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac79de),
	.w1(32'h3b78001c),
	.w2(32'hbaa59956),
	.w3(32'hbb572612),
	.w4(32'hbadb0475),
	.w5(32'h3b088c1c),
	.w6(32'hbbc40b60),
	.w7(32'h3b9bb745),
	.w8(32'hbba07078),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5649e),
	.w1(32'hbaa5e711),
	.w2(32'hbb2c6ab2),
	.w3(32'hbafe4a1c),
	.w4(32'hbbb3e7bc),
	.w5(32'hb9f304f4),
	.w6(32'hbbc6e5d8),
	.w7(32'hbb8f8e2d),
	.w8(32'hbac4a79a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40a631),
	.w1(32'hbb24c807),
	.w2(32'hbba95ad7),
	.w3(32'hbb6a5561),
	.w4(32'hbc0584af),
	.w5(32'hbad8134d),
	.w6(32'hbb2c29f3),
	.w7(32'hba8a2349),
	.w8(32'hbb0d8a52),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd67496),
	.w1(32'hbb6dfe97),
	.w2(32'hbbb36432),
	.w3(32'h3b2c4122),
	.w4(32'hbbd9e5d4),
	.w5(32'hbbe1e2db),
	.w6(32'h390f04c0),
	.w7(32'h39a90a98),
	.w8(32'hbb252772),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e6ff0),
	.w1(32'hbb0d00b7),
	.w2(32'hbba5d409),
	.w3(32'hbbba259b),
	.w4(32'hbb096d6d),
	.w5(32'hbace9e5a),
	.w6(32'hbb610dca),
	.w7(32'hbae359fb),
	.w8(32'h3b4ef0da),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabef020),
	.w1(32'h3ab10ee3),
	.w2(32'hbb7c7954),
	.w3(32'h3ba4b74b),
	.w4(32'h3afe8283),
	.w5(32'hbbf5336f),
	.w6(32'hbaa43da4),
	.w7(32'h38ba3d99),
	.w8(32'hbb1458f6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6a0d5),
	.w1(32'h3b865421),
	.w2(32'h3c371305),
	.w3(32'hbbf7fc56),
	.w4(32'h3beba50b),
	.w5(32'h3bf53a63),
	.w6(32'hbb633b7e),
	.w7(32'h3c17c961),
	.w8(32'h3b31157c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule