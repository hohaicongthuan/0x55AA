module layer_8_featuremap_35(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb226a7f),
	.w1(32'hba4cba85),
	.w2(32'h3c094a67),
	.w3(32'hbbfa77c2),
	.w4(32'hbbd90bac),
	.w5(32'h3bc4bf53),
	.w6(32'hbb86b5ad),
	.w7(32'hbb843012),
	.w8(32'h3b0b61ea),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac12e6),
	.w1(32'hba752718),
	.w2(32'hbaea8e2e),
	.w3(32'hba9ed2f2),
	.w4(32'hba9c034d),
	.w5(32'hbb15eb03),
	.w6(32'hba984b81),
	.w7(32'hba20bf98),
	.w8(32'hbb3c61e1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919fe7d),
	.w1(32'h3a380cb2),
	.w2(32'hb9d9a2a1),
	.w3(32'hb83ec748),
	.w4(32'hb9b7086a),
	.w5(32'hbabfbe76),
	.w6(32'h3a8a30e0),
	.w7(32'h3a71736b),
	.w8(32'hba8c748c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f96a7),
	.w1(32'hbafba1ab),
	.w2(32'h3ac67c63),
	.w3(32'hbbe397ab),
	.w4(32'hbb80a113),
	.w5(32'h39df69ec),
	.w6(32'hbb8b822c),
	.w7(32'h3b0e2235),
	.w8(32'h3abb4685),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a20f4),
	.w1(32'hb59e3f04),
	.w2(32'h377e5134),
	.w3(32'h3aa5127d),
	.w4(32'hba88d163),
	.w5(32'hbaae257f),
	.w6(32'h3abcfb77),
	.w7(32'hbabf301c),
	.w8(32'hba8c4a52),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce088c),
	.w1(32'h3b8e5035),
	.w2(32'hbbd8bfbd),
	.w3(32'h3bd990ff),
	.w4(32'h3b486948),
	.w5(32'hbbacddc5),
	.w6(32'h3b9c1fcd),
	.w7(32'hb9ca8756),
	.w8(32'hbbf10052),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ebc04),
	.w1(32'hb966b802),
	.w2(32'h396cfd76),
	.w3(32'hba541bf0),
	.w4(32'hba251913),
	.w5(32'hb945ef7f),
	.w6(32'hba03c475),
	.w7(32'hb98c1ffd),
	.w8(32'h3903ca83),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac0526),
	.w1(32'h38cc0442),
	.w2(32'h3bc8b863),
	.w3(32'hbb928ec5),
	.w4(32'h3958ec9a),
	.w5(32'h3bd3d97d),
	.w6(32'hbb51de60),
	.w7(32'h3916800f),
	.w8(32'h3b8a2b7b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b63d4),
	.w1(32'h3717df6c),
	.w2(32'hba939e16),
	.w3(32'h3927423b),
	.w4(32'hb93b0073),
	.w5(32'hba4ef55b),
	.w6(32'h39c7054c),
	.w7(32'hb9833f11),
	.w8(32'hbaf146f7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb58d66),
	.w1(32'h3b8e13d5),
	.w2(32'h3c500c5c),
	.w3(32'hbc12476c),
	.w4(32'hbad64001),
	.w5(32'h3c627d99),
	.w6(32'hba0580d1),
	.w7(32'h3b15c7c7),
	.w8(32'h3b94eae5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394cec62),
	.w1(32'h3b6d0131),
	.w2(32'h3c1309d2),
	.w3(32'hbba174ed),
	.w4(32'hbafcf776),
	.w5(32'h3bebe8b7),
	.w6(32'hbb979fa3),
	.w7(32'hbb1474b1),
	.w8(32'h3b53c8d8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d8349),
	.w1(32'hb886afa2),
	.w2(32'h3af0093f),
	.w3(32'hbbe1e3d1),
	.w4(32'hbb7bf45a),
	.w5(32'h39b33bb1),
	.w6(32'hba9d60ed),
	.w7(32'hbb32d5f7),
	.w8(32'hbb61942c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5db992),
	.w1(32'hba455c27),
	.w2(32'hba8823eb),
	.w3(32'hba73cf58),
	.w4(32'hbb1f68fb),
	.w5(32'hbb53797a),
	.w6(32'h3ab1e1fc),
	.w7(32'hb8745f63),
	.w8(32'hbace5ac5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98357c7),
	.w1(32'hba0d6a0d),
	.w2(32'hb89a0aed),
	.w3(32'h396e7eb4),
	.w4(32'hb99ac32c),
	.w5(32'h3a41c5a1),
	.w6(32'h3a43c524),
	.w7(32'hb9471f25),
	.w8(32'h3a2590bd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4f6f2),
	.w1(32'hb9c88d9a),
	.w2(32'hb9b33685),
	.w3(32'hb9dfd511),
	.w4(32'hbaa5bd5c),
	.w5(32'hb93c62bb),
	.w6(32'h398f0de1),
	.w7(32'hb9132d92),
	.w8(32'hb87a8dfc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eab631),
	.w1(32'h3a19cf9d),
	.w2(32'h3a19cead),
	.w3(32'h39fc2a67),
	.w4(32'h373c9455),
	.w5(32'h3a2573cc),
	.w6(32'h37be6ee9),
	.w7(32'hb997f7b2),
	.w8(32'h3abb175e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c8013),
	.w1(32'hbb6aa2fd),
	.w2(32'h3aa81b86),
	.w3(32'hbbaded4f),
	.w4(32'hbc0af556),
	.w5(32'hbaca5f10),
	.w6(32'hbab8c227),
	.w7(32'hbb17684e),
	.w8(32'h3a66099a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dc18c),
	.w1(32'h3b0e413d),
	.w2(32'h3b8d0932),
	.w3(32'hbb2bcc0f),
	.w4(32'hbaaada85),
	.w5(32'h3ae4bfb4),
	.w6(32'h3ab99009),
	.w7(32'h3a6a206a),
	.w8(32'h3a881ed3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80994e),
	.w1(32'h3bd47832),
	.w2(32'h3d061665),
	.w3(32'hbcc15a2a),
	.w4(32'hbc354079),
	.w5(32'h3cf5d430),
	.w6(32'hbc87a9b3),
	.w7(32'hbb1f3800),
	.w8(32'h3c993f7c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7a22e),
	.w1(32'hbbbfe82b),
	.w2(32'hbb9ea0f2),
	.w3(32'hbab03140),
	.w4(32'hbbee583b),
	.w5(32'hbc259f8a),
	.w6(32'h3b946fc8),
	.w7(32'hbae8ca72),
	.w8(32'hbb8f24ab),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ee5cd),
	.w1(32'hb8ea95b4),
	.w2(32'hbb4b2c92),
	.w3(32'hb7b5f05a),
	.w4(32'hbbf826bc),
	.w5(32'hbbb105a8),
	.w6(32'h3b0b0d78),
	.w7(32'hbc0bec72),
	.w8(32'hbbadd66c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4c25a),
	.w1(32'hba83ec73),
	.w2(32'hbb5cdcf6),
	.w3(32'hba02fd3c),
	.w4(32'hbac62f86),
	.w5(32'hbb635fd5),
	.w6(32'hb82963de),
	.w7(32'h39c16b2d),
	.w8(32'hbb633bbf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeafa2),
	.w1(32'h39df660d),
	.w2(32'h3cb0cb49),
	.w3(32'hbc743ddc),
	.w4(32'hbbd490e6),
	.w5(32'h3cc28afa),
	.w6(32'hbc7168ec),
	.w7(32'hbc0d9113),
	.w8(32'h3c420e62),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00e03b),
	.w1(32'hba5fc458),
	.w2(32'hbb4acf65),
	.w3(32'hb9810b71),
	.w4(32'hba2b406a),
	.w5(32'hbb214ee9),
	.w6(32'h3aaea4c3),
	.w7(32'hba5f0242),
	.w8(32'hbbd45cb1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb411e19),
	.w1(32'hbb552278),
	.w2(32'hbb5f17dc),
	.w3(32'h3a0c853b),
	.w4(32'h3b09781f),
	.w5(32'hba465167),
	.w6(32'hbba053dd),
	.w7(32'hbba01def),
	.w8(32'hba190668),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e28c1),
	.w1(32'h3ade238c),
	.w2(32'h3ba13a74),
	.w3(32'hbb4bb046),
	.w4(32'hbb6fc278),
	.w5(32'h3b35b436),
	.w6(32'hbb1f19c3),
	.w7(32'hbbc14cb4),
	.w8(32'hba2fa8c0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c523a7),
	.w1(32'hb9cb47cd),
	.w2(32'hb902d444),
	.w3(32'hb9c5ee41),
	.w4(32'hb938f04b),
	.w5(32'hba15e802),
	.w6(32'hb9faafef),
	.w7(32'h3945986e),
	.w8(32'hba51b1fe),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0257e0),
	.w1(32'h3d30809f),
	.w2(32'hbcc255a6),
	.w3(32'hbce60fc3),
	.w4(32'h3bc71d0e),
	.w5(32'hbd285230),
	.w6(32'hbd49c602),
	.w7(32'hbcf5d457),
	.w8(32'hbbfd85fe),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1c1e7),
	.w1(32'hbae6f79c),
	.w2(32'h3c080609),
	.w3(32'hbbea0e8a),
	.w4(32'hba90b637),
	.w5(32'h3c12104e),
	.w6(32'hbbcc1bd1),
	.w7(32'hbb1d0735),
	.w8(32'h3b0c2611),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba145990),
	.w1(32'hb994a8a4),
	.w2(32'hba1bd888),
	.w3(32'hba311509),
	.w4(32'hba437e07),
	.w5(32'hba4a0664),
	.w6(32'hba384717),
	.w7(32'hba411d18),
	.w8(32'h3a99cb18),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b93332),
	.w1(32'h3ae28424),
	.w2(32'h3a89f063),
	.w3(32'hbaad0242),
	.w4(32'hbba490cc),
	.w5(32'hbb136cf8),
	.w6(32'h3a8e75bd),
	.w7(32'hbaf7676b),
	.w8(32'hb91dc2ce),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e52bd),
	.w1(32'hbac192bd),
	.w2(32'hbb98b9ad),
	.w3(32'h3b06fec0),
	.w4(32'hb98601e9),
	.w5(32'hbb97875d),
	.w6(32'hbae6ff4e),
	.w7(32'hbb6725b6),
	.w8(32'hbb015eee),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39828bf1),
	.w1(32'h37d8c0a6),
	.w2(32'hba5b19aa),
	.w3(32'hbb53b0e9),
	.w4(32'hbbb50d34),
	.w5(32'hbba7abb8),
	.w6(32'h39ae7178),
	.w7(32'hba451b1c),
	.w8(32'h399dc307),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb700493),
	.w1(32'hbb732631),
	.w2(32'hbb3bbd85),
	.w3(32'h3ae59f42),
	.w4(32'h3ace833d),
	.w5(32'h3b598423),
	.w6(32'h3acb17ee),
	.w7(32'hbb36409e),
	.w8(32'h3a9f79bb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fb02f),
	.w1(32'hbb17bb6a),
	.w2(32'hbba39a9d),
	.w3(32'hba31da66),
	.w4(32'h3a30afab),
	.w5(32'hbb89674d),
	.w6(32'h3aee7b21),
	.w7(32'h3b1b6d04),
	.w8(32'hbaf68180),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9087a9),
	.w1(32'hba51c798),
	.w2(32'h3bcc065f),
	.w3(32'hbc110611),
	.w4(32'hbbd490dd),
	.w5(32'h3b6ce03c),
	.w6(32'hbbb371bd),
	.w7(32'hbb896640),
	.w8(32'hb9a5179a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a480f38),
	.w1(32'h39c6a26b),
	.w2(32'hba2d04cd),
	.w3(32'h3a64c485),
	.w4(32'h3a0cd9ba),
	.w5(32'hb9373a72),
	.w6(32'hbabdd441),
	.w7(32'hbac0cacd),
	.w8(32'hba240b4e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dc1fd),
	.w1(32'hb9a560b3),
	.w2(32'hb95a9e8a),
	.w3(32'hbac8955b),
	.w4(32'hba6c824a),
	.w5(32'hba3530a6),
	.w6(32'hba5cd99d),
	.w7(32'h38be48bb),
	.w8(32'h3aa1cd70),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab7b7b),
	.w1(32'hba3f0880),
	.w2(32'hba219ee8),
	.w3(32'hba45d5c2),
	.w4(32'hbb4a6471),
	.w5(32'hba082aba),
	.w6(32'h39926234),
	.w7(32'h38bdd292),
	.w8(32'hba9fcedf),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e506f2),
	.w1(32'h3a27450c),
	.w2(32'h396967a5),
	.w3(32'h3a1cb283),
	.w4(32'h39c4b8cd),
	.w5(32'hb8ba3536),
	.w6(32'hbad0ae16),
	.w7(32'hbaa16602),
	.w8(32'h39938e18),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef0d68),
	.w1(32'h3c45c224),
	.w2(32'h3ad7926a),
	.w3(32'hbaa829aa),
	.w4(32'h3c0b277e),
	.w5(32'h39d43366),
	.w6(32'hbb0ddc18),
	.w7(32'h3b897909),
	.w8(32'hbc511b98),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8827f6),
	.w1(32'hbb1c4776),
	.w2(32'h3ac72a67),
	.w3(32'hbbccfa68),
	.w4(32'hbb5c754d),
	.w5(32'h3b0c03b9),
	.w6(32'hbba26a8f),
	.w7(32'hbb1c63cf),
	.w8(32'hba7f0390),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a5dac),
	.w1(32'hbac21125),
	.w2(32'hbb0ec0f6),
	.w3(32'hba768fe4),
	.w4(32'h3a2c9c45),
	.w5(32'hbab6d3e7),
	.w6(32'hbb34af74),
	.w7(32'hbb21099a),
	.w8(32'hba66aeea),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bd8a20),
	.w1(32'h392f98ac),
	.w2(32'h39f6dc20),
	.w3(32'hbab8682d),
	.w4(32'hbaa89554),
	.w5(32'h3ae5f660),
	.w6(32'hbb70f3bb),
	.w7(32'hbb683c1b),
	.w8(32'h3a52fcc4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba414a84),
	.w1(32'hb92b7b1a),
	.w2(32'h3c43a3f7),
	.w3(32'hbbd1001f),
	.w4(32'hbb6be721),
	.w5(32'h3c556118),
	.w6(32'hbc095674),
	.w7(32'hbb9bca28),
	.w8(32'h3c082492),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4db78),
	.w1(32'hbb77446e),
	.w2(32'h3bf99290),
	.w3(32'hbc2b0552),
	.w4(32'hbb73ceab),
	.w5(32'h3be4b364),
	.w6(32'hbbd91b36),
	.w7(32'hba1fb212),
	.w8(32'h3a8b530f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c828d),
	.w1(32'h3b91d73f),
	.w2(32'h3a1241c1),
	.w3(32'h3ac57d7d),
	.w4(32'h3b21fb10),
	.w5(32'hba3d02c7),
	.w6(32'hb97afc79),
	.w7(32'hbacedb85),
	.w8(32'hba87aca5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc063d51),
	.w1(32'hbc117488),
	.w2(32'h3ba68650),
	.w3(32'hbbf7fd64),
	.w4(32'hbc2706e7),
	.w5(32'h3ba79d5c),
	.w6(32'hbc07d5f2),
	.w7(32'hbbf1b308),
	.w8(32'h3ba0c90d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c6add),
	.w1(32'h3a8c2567),
	.w2(32'h3977f9f3),
	.w3(32'hbaa013a4),
	.w4(32'h3a9dceff),
	.w5(32'h3a0773c0),
	.w6(32'hba17d89f),
	.w7(32'h3a070f04),
	.w8(32'hb86cf7e7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a552b4),
	.w1(32'h3acd79b9),
	.w2(32'h3bfb4082),
	.w3(32'hbb8d7c82),
	.w4(32'hba02a257),
	.w5(32'h3bfc93f4),
	.w6(32'hbb667299),
	.w7(32'h3955ec93),
	.w8(32'h3b3f07d7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92a67a),
	.w1(32'hbb4a008c),
	.w2(32'hbbcc45e7),
	.w3(32'h3b9f3d43),
	.w4(32'hbb5e77ad),
	.w5(32'hbc0dda54),
	.w6(32'h3c03db4e),
	.w7(32'h3a5944ec),
	.w8(32'hbc190725),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8257d0),
	.w1(32'h3c5e5162),
	.w2(32'h3c8f345d),
	.w3(32'hbb6d842d),
	.w4(32'h3c0e674e),
	.w5(32'h3cbb90cc),
	.w6(32'hbc50aa3e),
	.w7(32'hbb20aa26),
	.w8(32'h3c888b59),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32416d),
	.w1(32'hbb634d8b),
	.w2(32'hba117ce3),
	.w3(32'hbad76d8a),
	.w4(32'hbace5dea),
	.w5(32'h3b34bcb6),
	.w6(32'hbbaafe16),
	.w7(32'hbc082bc0),
	.w8(32'h3a143de2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0fbd3),
	.w1(32'hbb94116a),
	.w2(32'h3c26f883),
	.w3(32'hbc21f888),
	.w4(32'hbbc026a5),
	.w5(32'h3c1d82e8),
	.w6(32'hbac5d0fb),
	.w7(32'h3aff988c),
	.w8(32'h3b6ab894),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4b34c),
	.w1(32'h38752f7d),
	.w2(32'h380239dc),
	.w3(32'hba0356fc),
	.w4(32'h3b3e4bf7),
	.w5(32'h3b046b83),
	.w6(32'hbb5230a0),
	.w7(32'hbb422856),
	.w8(32'hba6186eb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc915756),
	.w1(32'hbc406661),
	.w2(32'h3c6573ae),
	.w3(32'hbc81f013),
	.w4(32'hbc596e3f),
	.w5(32'h3c373555),
	.w6(32'hbc415653),
	.w7(32'hbbf9a239),
	.w8(32'h3bb04fa6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86440b),
	.w1(32'hbb829f6a),
	.w2(32'h3a5ad59c),
	.w3(32'hba816884),
	.w4(32'hba4fd1a1),
	.w5(32'h3b966fed),
	.w6(32'hbade7ecf),
	.w7(32'hbb054c12),
	.w8(32'h3a48af3d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab740f8),
	.w1(32'h3bc697e6),
	.w2(32'h3bf30edc),
	.w3(32'hbbf9adec),
	.w4(32'h3b90c250),
	.w5(32'h3c14335b),
	.w6(32'hbbeb06e7),
	.w7(32'h3a02a267),
	.w8(32'h3bcd18d1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb355ab5),
	.w1(32'hbb63aa60),
	.w2(32'h3b05154f),
	.w3(32'hbaec339f),
	.w4(32'hbb20c52b),
	.w5(32'h3ba093ff),
	.w6(32'hbba9cf6c),
	.w7(32'hbbc85258),
	.w8(32'h3aa91350),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee39a6),
	.w1(32'h394d876c),
	.w2(32'hb9bea89e),
	.w3(32'hbb382dcc),
	.w4(32'hba62b492),
	.w5(32'hba42aa37),
	.w6(32'hbb8e2ac3),
	.w7(32'hba2e488a),
	.w8(32'hbaf26dbb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab03540),
	.w1(32'h39bff8a0),
	.w2(32'hba8498fe),
	.w3(32'h39c96826),
	.w4(32'h3ae049b6),
	.w5(32'h3aadcc8b),
	.w6(32'hbab421c7),
	.w7(32'hbacd8d10),
	.w8(32'hba00c48a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0da543),
	.w1(32'h39446c4b),
	.w2(32'h38c15e45),
	.w3(32'hbab2d552),
	.w4(32'hba9b1710),
	.w5(32'hb9571c75),
	.w6(32'hba19975b),
	.w7(32'hba25f64e),
	.w8(32'h3ab67286),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacc37a),
	.w1(32'h3b19cc45),
	.w2(32'h3bc38488),
	.w3(32'hbbcb0c7d),
	.w4(32'h3a05f387),
	.w5(32'h3bc7016c),
	.w6(32'hba5b5c36),
	.w7(32'h3b0bcacc),
	.w8(32'h3a6bb48f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18d96a),
	.w1(32'h3b1170bc),
	.w2(32'hb8da32e0),
	.w3(32'hbb007614),
	.w4(32'hb9b3cdce),
	.w5(32'hbb4a1a46),
	.w6(32'hbae7cc3c),
	.w7(32'hba8c1d54),
	.w8(32'h3a9b30b6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381aef08),
	.w1(32'hb999abde),
	.w2(32'hb97e2df1),
	.w3(32'h39707a68),
	.w4(32'hb9b5aa80),
	.w5(32'hb9dce3e6),
	.w6(32'hb94cb06a),
	.w7(32'hb95406b4),
	.w8(32'hba0357e0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea7544),
	.w1(32'h3a91da3f),
	.w2(32'h3a75d0ad),
	.w3(32'hbb364c0c),
	.w4(32'hbb14de6d),
	.w5(32'hba90f6e6),
	.w6(32'hbb1e3b65),
	.w7(32'hbb00a919),
	.w8(32'hba3e8ca8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bcac4),
	.w1(32'hba0a1122),
	.w2(32'hbb4b23ff),
	.w3(32'h3b052ab4),
	.w4(32'hb94582e8),
	.w5(32'hbb1dee53),
	.w6(32'h3a36a862),
	.w7(32'hb9fcedff),
	.w8(32'hbb02730c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07a1b0),
	.w1(32'hbb13528e),
	.w2(32'h3997e50c),
	.w3(32'hbb8c80f4),
	.w4(32'hbbd1910e),
	.w5(32'hbb26ae81),
	.w6(32'h39c72415),
	.w7(32'hbb6babe7),
	.w8(32'hbb09f214),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fdebeb),
	.w1(32'h396de904),
	.w2(32'h3a14945a),
	.w3(32'h3a050df1),
	.w4(32'h3966d942),
	.w5(32'h39939e6d),
	.w6(32'h3a0c88ea),
	.w7(32'h3a26416f),
	.w8(32'h3a8a52a4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81f782),
	.w1(32'hba999082),
	.w2(32'h3c02e92c),
	.w3(32'hbacf6e6a),
	.w4(32'hbc2f5ccf),
	.w5(32'h3c0816f3),
	.w6(32'hbc7cf44a),
	.w7(32'hbca6398b),
	.w8(32'h3be95b70),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ada203),
	.w1(32'hba270663),
	.w2(32'hb9db9569),
	.w3(32'hb93035dd),
	.w4(32'hba46e7eb),
	.w5(32'hba55079c),
	.w6(32'hb8d8401c),
	.w7(32'hb8269d0c),
	.w8(32'h3a3e53a5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a46d5),
	.w1(32'hba203c16),
	.w2(32'hbaea176a),
	.w3(32'hba915625),
	.w4(32'hb98c3c26),
	.w5(32'hba9594dc),
	.w6(32'hbb662664),
	.w7(32'hbb07a475),
	.w8(32'hbb19e987),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29c136),
	.w1(32'hb92f47ef),
	.w2(32'hba362947),
	.w3(32'hba46e974),
	.w4(32'hb9c5cf7a),
	.w5(32'hbabfbdb8),
	.w6(32'hba2ae45a),
	.w7(32'h3982c327),
	.w8(32'h3b875d4a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb617562),
	.w1(32'h3c032408),
	.w2(32'h3c1e6504),
	.w3(32'hbbd17a47),
	.w4(32'h39db076e),
	.w5(32'h3b3de726),
	.w6(32'h3b1a9743),
	.w7(32'hbaadd3ca),
	.w8(32'hb9f4ba83),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cb5c0),
	.w1(32'h3a73fcba),
	.w2(32'h3a2ee348),
	.w3(32'h3a07b9b1),
	.w4(32'h393537d5),
	.w5(32'h38209c09),
	.w6(32'h3a8e3038),
	.w7(32'h3a6c24ac),
	.w8(32'hb90c49bb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23c382),
	.w1(32'h3abc8ca9),
	.w2(32'h3b714168),
	.w3(32'h3aa6804b),
	.w4(32'h3a184948),
	.w5(32'h3ba0cce7),
	.w6(32'hbac6de9b),
	.w7(32'hbac17dc2),
	.w8(32'h3b2ffa92),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0353f),
	.w1(32'hb97888f5),
	.w2(32'hb98bb975),
	.w3(32'hb9660e65),
	.w4(32'hba12e231),
	.w5(32'hba3caabe),
	.w6(32'h394e5910),
	.w7(32'h38ed649e),
	.w8(32'h3a9d71e3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f63e6),
	.w1(32'h3b712bc2),
	.w2(32'h3bca19ca),
	.w3(32'hb7497cf1),
	.w4(32'hbb5ab567),
	.w5(32'h3b8db65c),
	.w6(32'hbbae4175),
	.w7(32'hbb986690),
	.w8(32'h3adedb9f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8f7e1),
	.w1(32'hbb34ca27),
	.w2(32'h3c25aba6),
	.w3(32'hbc12e0a7),
	.w4(32'hbaee284c),
	.w5(32'h3c15b0a7),
	.w6(32'hbb9a95c5),
	.w7(32'h3a0359a4),
	.w8(32'h3c0cfd6d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf551b),
	.w1(32'h391456a0),
	.w2(32'h39d4e8c7),
	.w3(32'h38f82cd0),
	.w4(32'hb9a38425),
	.w5(32'hb97c4900),
	.w6(32'h39fcd5eb),
	.w7(32'h3a2f3e05),
	.w8(32'h381b24d8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cc047),
	.w1(32'h3b7daaa6),
	.w2(32'h3aa73ab7),
	.w3(32'h3acf3e4a),
	.w4(32'h3b5e1498),
	.w5(32'h3ad62cd0),
	.w6(32'h3a10d33e),
	.w7(32'hba98f845),
	.w8(32'h389910f0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a316dd1),
	.w1(32'h3b4dee7c),
	.w2(32'hbabdc986),
	.w3(32'hba4a566c),
	.w4(32'h3a9f3645),
	.w5(32'hba047507),
	.w6(32'hbb9ab27e),
	.w7(32'hbba5e414),
	.w8(32'h3a97c795),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10ce22),
	.w1(32'h3ae50320),
	.w2(32'h3b3da137),
	.w3(32'hbb51fd5c),
	.w4(32'hbad6211b),
	.w5(32'h3b747ee7),
	.w6(32'hbb84b74a),
	.w7(32'hbb41d072),
	.w8(32'hbb7b4204),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18845b),
	.w1(32'h3b0ced4a),
	.w2(32'hba9b0b2f),
	.w3(32'hb94ac6fc),
	.w4(32'h3b02b9ff),
	.w5(32'hbc0dbfa4),
	.w6(32'hb9cece04),
	.w7(32'h3b8c7518),
	.w8(32'hbc88fb37),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62c946),
	.w1(32'h3a1782b1),
	.w2(32'h3c2eef23),
	.w3(32'hbc4d275e),
	.w4(32'hbbf1b600),
	.w5(32'h3c2f4249),
	.w6(32'hbc2cc6a2),
	.w7(32'hbc0dcda8),
	.w8(32'h3aeabfce),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe8fd5),
	.w1(32'h3bb0a144),
	.w2(32'h3aef22e4),
	.w3(32'h3aa002f9),
	.w4(32'h3bd121ee),
	.w5(32'h3babd1d1),
	.w6(32'hba5da89e),
	.w7(32'hbabe28c4),
	.w8(32'h3b3945e0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3898f8af),
	.w1(32'h385f94a4),
	.w2(32'hb9b80461),
	.w3(32'hb8a592ce),
	.w4(32'h39fa194b),
	.w5(32'h3a750580),
	.w6(32'hb98cdf28),
	.w7(32'hb884bcee),
	.w8(32'h38dabced),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bf0ac6),
	.w1(32'h392235ad),
	.w2(32'h3a2532be),
	.w3(32'h3a269da2),
	.w4(32'h3a02e89b),
	.w5(32'h3a63784b),
	.w6(32'hb998e503),
	.w7(32'h393c2aee),
	.w8(32'hb9fc1c38),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0aa1c),
	.w1(32'h38e3bc5d),
	.w2(32'hba3b21a8),
	.w3(32'hbaf744fa),
	.w4(32'hbad84027),
	.w5(32'hbaf3565a),
	.w6(32'hb96195df),
	.w7(32'hba84dcf5),
	.w8(32'hb9849067),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8a3d6),
	.w1(32'hba1b7783),
	.w2(32'h3980ea71),
	.w3(32'hbae1e1ab),
	.w4(32'h39b60fd0),
	.w5(32'h3b1fe50f),
	.w6(32'hbb27cad4),
	.w7(32'hbac3ae9f),
	.w8(32'h3a085799),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f32bf),
	.w1(32'h3b208c25),
	.w2(32'h3a1fe103),
	.w3(32'hbb2def99),
	.w4(32'h3b02d15f),
	.w5(32'h3ae5d2e4),
	.w6(32'hba8a19e1),
	.w7(32'hba8f7912),
	.w8(32'hba827b17),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f1b17),
	.w1(32'h392f5695),
	.w2(32'h39ae232a),
	.w3(32'hba1ca472),
	.w4(32'hb7c65b5a),
	.w5(32'h39c54c80),
	.w6(32'hb85c9f23),
	.w7(32'hb8b700cc),
	.w8(32'hbb4ea35e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8acd1),
	.w1(32'h3965cdd0),
	.w2(32'hbb653cf2),
	.w3(32'h3bd59642),
	.w4(32'h3b70cdca),
	.w5(32'h38cf86d5),
	.w6(32'hbad215d8),
	.w7(32'hba8ad62e),
	.w8(32'hba3a7b90),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47a21d),
	.w1(32'h3aa1509e),
	.w2(32'h3b39b271),
	.w3(32'hbb00dca9),
	.w4(32'hb9384c6f),
	.w5(32'h3b0c0392),
	.w6(32'hba4875aa),
	.w7(32'h38673cfa),
	.w8(32'hbb0aa892),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d21df),
	.w1(32'h3a63414c),
	.w2(32'hba9747a9),
	.w3(32'hbb3eebcc),
	.w4(32'hba003ce6),
	.w5(32'hbacc44ea),
	.w6(32'hba9cddf5),
	.w7(32'hbb60cab0),
	.w8(32'hbb905bd8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0df875),
	.w1(32'hbbc35dda),
	.w2(32'h3b12b51d),
	.w3(32'hbb512847),
	.w4(32'hbc0136fb),
	.w5(32'h3b02144b),
	.w6(32'hbb1cc7dc),
	.w7(32'hbb917d08),
	.w8(32'h3ba29020),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2ffa0),
	.w1(32'h3b305898),
	.w2(32'h3ba11334),
	.w3(32'hbac3f4ed),
	.w4(32'h3a8568c8),
	.w5(32'h3be7f037),
	.w6(32'hbb9413a2),
	.w7(32'hbba0b004),
	.w8(32'h3a9db0c9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95cac0),
	.w1(32'h3bf60585),
	.w2(32'h3bac9725),
	.w3(32'h3a518a29),
	.w4(32'h3b1caa04),
	.w5(32'h39f949f3),
	.w6(32'h39e78124),
	.w7(32'h3a644052),
	.w8(32'h3a9533f9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d4af0f),
	.w1(32'hb982fc1a),
	.w2(32'h398382d2),
	.w3(32'h3adad5bc),
	.w4(32'h3a35ecc8),
	.w5(32'h3a453769),
	.w6(32'h3a73034c),
	.w7(32'h3a8f74ac),
	.w8(32'h3838c272),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383895ac),
	.w1(32'hb9c390ec),
	.w2(32'h396c6529),
	.w3(32'h3992c722),
	.w4(32'hb997f87c),
	.w5(32'h37b23782),
	.w6(32'hb9412f8a),
	.w7(32'h383a312c),
	.w8(32'hba721256),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc8724),
	.w1(32'h3a4467eb),
	.w2(32'hb89584e1),
	.w3(32'hb955d4c7),
	.w4(32'h396e5200),
	.w5(32'hb9fd4d37),
	.w6(32'hba44ff06),
	.w7(32'hba4f5fe4),
	.w8(32'h39aac05b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97597e5),
	.w1(32'h3a1e20dd),
	.w2(32'h3a307ba3),
	.w3(32'hb9a3e762),
	.w4(32'hba37d2c5),
	.w5(32'h38049bbe),
	.w6(32'hb91c5f12),
	.w7(32'hb9ae0ef6),
	.w8(32'hb9a55770),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cacc07),
	.w1(32'hba1c2d91),
	.w2(32'h3a6b56f6),
	.w3(32'h3b0151b5),
	.w4(32'h3a7b8689),
	.w5(32'h3aa707f4),
	.w6(32'h3a3c5b13),
	.w7(32'h3a758d37),
	.w8(32'hba414c59),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b70fa),
	.w1(32'h3b1fa1c0),
	.w2(32'hbb8e24f8),
	.w3(32'h39f5fcd5),
	.w4(32'h3b01be51),
	.w5(32'hbba7b6c2),
	.w6(32'h3a8cfe77),
	.w7(32'h3a08b362),
	.w8(32'hbb27138b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c608e),
	.w1(32'hb81dcf07),
	.w2(32'hbaa4570c),
	.w3(32'h392d04fe),
	.w4(32'h3a9e608e),
	.w5(32'hba283650),
	.w6(32'h39fc0eca),
	.w7(32'h3aa017f6),
	.w8(32'h382b42ad),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba389987),
	.w1(32'h3b479fad),
	.w2(32'h3bc407f7),
	.w3(32'hbb8fcdbe),
	.w4(32'hbb4b318e),
	.w5(32'h3b7418fd),
	.w6(32'hbbcedda2),
	.w7(32'hbc1bb24b),
	.w8(32'hba85c148),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8fad5),
	.w1(32'h3c43664d),
	.w2(32'hb8ecbadc),
	.w3(32'hba93f172),
	.w4(32'h3bab0f8b),
	.w5(32'hba52621c),
	.w6(32'h3ab62b55),
	.w7(32'hbbb26f62),
	.w8(32'hb99c1f7b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e8feb),
	.w1(32'hbb48dedb),
	.w2(32'hbb7b054a),
	.w3(32'h3a711195),
	.w4(32'hba01dcf2),
	.w5(32'hbad08d6e),
	.w6(32'h3a79d039),
	.w7(32'hb9f4a1e3),
	.w8(32'hba6a550c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96adbc),
	.w1(32'hb9a67e8f),
	.w2(32'h3837579c),
	.w3(32'hb9cd4a2f),
	.w4(32'h39fd2e9f),
	.w5(32'h3a0d1fe1),
	.w6(32'hb9dc7560),
	.w7(32'h3a1a81cb),
	.w8(32'hb91c0a5a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10e0ec),
	.w1(32'hb9c1fd5d),
	.w2(32'h3ad59237),
	.w3(32'hbaf76c97),
	.w4(32'h3a63be0e),
	.w5(32'h3b023dc3),
	.w6(32'hbae6bfb6),
	.w7(32'hbad5dcba),
	.w8(32'hbb0402e6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5e4ce),
	.w1(32'hbba1ea87),
	.w2(32'hbbeb8c15),
	.w3(32'h391cb2c3),
	.w4(32'hbb843c49),
	.w5(32'hbbc388d9),
	.w6(32'h3b4a0520),
	.w7(32'hbafddfc5),
	.w8(32'hbbf67ee6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fd417),
	.w1(32'hbb4cd0e3),
	.w2(32'hbaf1bedb),
	.w3(32'hbac95099),
	.w4(32'hbb2b1368),
	.w5(32'hbbdc5605),
	.w6(32'hbb0996cc),
	.w7(32'hba17588b),
	.w8(32'hbb134906),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d5371),
	.w1(32'h3aa1ca80),
	.w2(32'h39ff9c69),
	.w3(32'h3a925128),
	.w4(32'h3b218069),
	.w5(32'h3a79f0df),
	.w6(32'hba4117bd),
	.w7(32'h3a4b6314),
	.w8(32'h3a9f1c57),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b2200),
	.w1(32'hba4de9b3),
	.w2(32'hb9039885),
	.w3(32'hba998e01),
	.w4(32'h3846c28b),
	.w5(32'hb9b1c270),
	.w6(32'hba21d25f),
	.w7(32'hba3734b9),
	.w8(32'h39baaa83),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba628bf1),
	.w1(32'hb91e7c0c),
	.w2(32'h3aaa3ae6),
	.w3(32'hbaa859fc),
	.w4(32'hb9a212c8),
	.w5(32'h3ad79c4d),
	.w6(32'hbae39b22),
	.w7(32'h3a3597c9),
	.w8(32'h3ad32070),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f3156),
	.w1(32'hb909ccb9),
	.w2(32'hba10eaa5),
	.w3(32'hba6f92bd),
	.w4(32'h37a17121),
	.w5(32'hb7709ba3),
	.w6(32'hba74d616),
	.w7(32'hba92f3b1),
	.w8(32'h388c14a1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0b276),
	.w1(32'h3b87f573),
	.w2(32'hbb51db7e),
	.w3(32'h3aa02a68),
	.w4(32'h3b829623),
	.w5(32'hbb35e9d2),
	.w6(32'hbb025a8c),
	.w7(32'hbad4ca74),
	.w8(32'h3bc8fb9e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ec16a),
	.w1(32'h3b59d0d2),
	.w2(32'h3bbf5dd3),
	.w3(32'h38b0bb1f),
	.w4(32'h3a99f6ac),
	.w5(32'h3be7fc46),
	.w6(32'hbb05c84c),
	.w7(32'hbb070d9c),
	.w8(32'h3a8f7e17),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f4714),
	.w1(32'hbb2f29d5),
	.w2(32'hbb007bee),
	.w3(32'h39361bc0),
	.w4(32'hbb808c7e),
	.w5(32'hbb1db49b),
	.w6(32'hbba29a06),
	.w7(32'h3a8432ac),
	.w8(32'hbb7195d6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7702d5),
	.w1(32'hba84f43b),
	.w2(32'hba4d5b1b),
	.w3(32'hbb466e1c),
	.w4(32'hb9bf71fe),
	.w5(32'hba860971),
	.w6(32'hbacb1d03),
	.w7(32'hbb0bb2f1),
	.w8(32'hba690713),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6d55b),
	.w1(32'hbbf3dce2),
	.w2(32'hba25dce2),
	.w3(32'hbbae17e5),
	.w4(32'h39e1bd5b),
	.w5(32'h3b30b517),
	.w6(32'hbba3eb34),
	.w7(32'hbb74c82e),
	.w8(32'hbb170746),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c039d6b),
	.w1(32'h3be197d9),
	.w2(32'hbaac5cce),
	.w3(32'h3a5d6461),
	.w4(32'h3b88573b),
	.w5(32'h3b000d2c),
	.w6(32'hbb606e82),
	.w7(32'h3b55b551),
	.w8(32'h3a790227),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e9094),
	.w1(32'h38b8fbd4),
	.w2(32'h3a1ebf17),
	.w3(32'h3a847511),
	.w4(32'h3a50919a),
	.w5(32'h3abd2eb9),
	.w6(32'h3864611b),
	.w7(32'h3a3b73b5),
	.w8(32'hbb6527a0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90ce5b),
	.w1(32'hbb1b5e77),
	.w2(32'hbb89ca20),
	.w3(32'hbb7bf20b),
	.w4(32'hbb8f693c),
	.w5(32'hbb98f89c),
	.w6(32'hbb4d3a4a),
	.w7(32'hbba4417d),
	.w8(32'hbb4859fb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaf0e7),
	.w1(32'h3b364a6a),
	.w2(32'h398a7f40),
	.w3(32'h3b807205),
	.w4(32'h3c20a080),
	.w5(32'hbab5d523),
	.w6(32'hbae4b6b7),
	.w7(32'hba0df6cf),
	.w8(32'hba6a3e86),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aee709),
	.w1(32'hbba8c5e7),
	.w2(32'hbb8c5258),
	.w3(32'hbaed8f03),
	.w4(32'hbbb16c5a),
	.w5(32'hbb863d5e),
	.w6(32'hba7e6fd2),
	.w7(32'hbb3236f6),
	.w8(32'h3a171976),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13a09c),
	.w1(32'h3b0c7320),
	.w2(32'h3b82105d),
	.w3(32'hbb4f0642),
	.w4(32'h3adbd04d),
	.w5(32'h3b8803fc),
	.w6(32'hb96c5889),
	.w7(32'h395ea3ad),
	.w8(32'h3b2aaf41),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1f2f3),
	.w1(32'h3bcc56ef),
	.w2(32'h3a8bcf3b),
	.w3(32'hbbdbc804),
	.w4(32'hbbfeb57c),
	.w5(32'h3bee97dc),
	.w6(32'hbbfc0a1e),
	.w7(32'hbc26d140),
	.w8(32'h3b2ee53a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule