module layer_8_featuremap_197(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd722bb),
	.w1(32'h39a7c00d),
	.w2(32'hbb787368),
	.w3(32'h3b3582a4),
	.w4(32'hbcb00ac1),
	.w5(32'hbba6580d),
	.w6(32'hba01f3e9),
	.w7(32'h3a962811),
	.w8(32'h3b7694a9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbee328),
	.w1(32'h3b2cbeca),
	.w2(32'h3bc40e51),
	.w3(32'h3c8f57d0),
	.w4(32'h3b3c28b6),
	.w5(32'h39b0baea),
	.w6(32'h3bc632cd),
	.w7(32'h3c0139ff),
	.w8(32'h3b80371e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c452e79),
	.w1(32'hbaf928e9),
	.w2(32'h3a616d3a),
	.w3(32'h3c392daa),
	.w4(32'h3bbcb142),
	.w5(32'h3b086d41),
	.w6(32'h3c2f4e48),
	.w7(32'h3c50a164),
	.w8(32'h3a945c9d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06e03b),
	.w1(32'hbc599962),
	.w2(32'h3b2857ef),
	.w3(32'hbc8fb730),
	.w4(32'hbc7690b6),
	.w5(32'hbcaf72b7),
	.w6(32'h3c49eb1b),
	.w7(32'h3c4cc5c8),
	.w8(32'h3bf0e862),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b4d6f),
	.w1(32'h3b44a7d9),
	.w2(32'h3b3422ff),
	.w3(32'hbbc84a11),
	.w4(32'h3b50f1d5),
	.w5(32'h3b10f894),
	.w6(32'hba5067b3),
	.w7(32'hbb5cf56b),
	.w8(32'hbbd38352),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17d1b9),
	.w1(32'hbb2561d4),
	.w2(32'hbbdcd3d0),
	.w3(32'h3c052692),
	.w4(32'hbab3dc91),
	.w5(32'hbbe58a0d),
	.w6(32'hbabc6c69),
	.w7(32'hbbebecc5),
	.w8(32'hbb59bf5e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc223872),
	.w1(32'h3bbc4d80),
	.w2(32'h3ba8bd27),
	.w3(32'h3bdf7ba1),
	.w4(32'h3b828d58),
	.w5(32'h3bc29c36),
	.w6(32'hba812a50),
	.w7(32'hbb987e47),
	.w8(32'hbb822873),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafcdd8),
	.w1(32'h3a683171),
	.w2(32'hb9fde736),
	.w3(32'h3b696edc),
	.w4(32'hba866081),
	.w5(32'hbb9e9ec5),
	.w6(32'hbb3328f0),
	.w7(32'hbb96ac8a),
	.w8(32'hbb81d240),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0eade),
	.w1(32'h3c32ccde),
	.w2(32'h3c84c814),
	.w3(32'h3a94b80f),
	.w4(32'hba869b8a),
	.w5(32'h3c20475c),
	.w6(32'h3ad35173),
	.w7(32'hbb8072f8),
	.w8(32'hbbb04733),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390697),
	.w1(32'h3d19cb36),
	.w2(32'h3cb979bd),
	.w3(32'h3c41675c),
	.w4(32'h3ccc5c19),
	.w5(32'h3d2adc9b),
	.w6(32'h3a5fbdd1),
	.w7(32'hbc8b9f5c),
	.w8(32'hbc70e689),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ee0d4),
	.w1(32'hbd3f8d43),
	.w2(32'h39b14105),
	.w3(32'h3b83cf08),
	.w4(32'hbcd1b99e),
	.w5(32'hbd1785ed),
	.w6(32'hbc4c3659),
	.w7(32'h3ca64c52),
	.w8(32'h3cc1341c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d485e04),
	.w1(32'hbadeb1f6),
	.w2(32'hbbdf9e0c),
	.w3(32'h3c740d37),
	.w4(32'h3bbbe7dd),
	.w5(32'hba456c77),
	.w6(32'hb9063bce),
	.w7(32'h3ad55cac),
	.w8(32'h3b12b693),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c328dc0),
	.w1(32'h3c4f7cd0),
	.w2(32'h3b3d44af),
	.w3(32'h3c3c158b),
	.w4(32'h3c8c4870),
	.w5(32'h3bcbb329),
	.w6(32'h3c0649b7),
	.w7(32'h3b943626),
	.w8(32'hbb490fd3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c1001),
	.w1(32'hbac7f856),
	.w2(32'hbca2a07e),
	.w3(32'hbb9f4c39),
	.w4(32'h3c2f5b64),
	.w5(32'h3bc92a28),
	.w6(32'hbc1a4e26),
	.w7(32'h3aca4df1),
	.w8(32'h395de529),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc949476),
	.w1(32'h3bc3b8f7),
	.w2(32'h3ba6ebe5),
	.w3(32'hbc426326),
	.w4(32'h3b11bb6e),
	.w5(32'h3bf024cb),
	.w6(32'hbb47ccec),
	.w7(32'hbbe47825),
	.w8(32'hbc0d718a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e3b1b),
	.w1(32'hbb8bef35),
	.w2(32'h3961c4d9),
	.w3(32'hbbb447a6),
	.w4(32'hbcb165b5),
	.w5(32'hba51baa6),
	.w6(32'hbb8b7f70),
	.w7(32'h3b845200),
	.w8(32'h3c75f3d1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33a889),
	.w1(32'h3c201dc8),
	.w2(32'h3c80a437),
	.w3(32'h3c1addd5),
	.w4(32'hbb75f968),
	.w5(32'h3b9137c0),
	.w6(32'h3bb3143d),
	.w7(32'h3c102db9),
	.w8(32'hbb249f93),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59df72),
	.w1(32'h3bf1be97),
	.w2(32'hbc920202),
	.w3(32'h3bf412e1),
	.w4(32'h3c6c3571),
	.w5(32'hbaf17c5a),
	.w6(32'hbc01aa5e),
	.w7(32'hbc33be3c),
	.w8(32'h3bf9d10f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f668b),
	.w1(32'hbc3b08e1),
	.w2(32'hbca35697),
	.w3(32'hbc959aaf),
	.w4(32'hbb4398e0),
	.w5(32'h3c0478c2),
	.w6(32'h3b03f6c2),
	.w7(32'hbcbb33a3),
	.w8(32'hbb87271f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd23262),
	.w1(32'hbafc2dcc),
	.w2(32'hba68fd61),
	.w3(32'hbb838e4c),
	.w4(32'hbac4008c),
	.w5(32'h3b675143),
	.w6(32'hbb804eab),
	.w7(32'hbc104403),
	.w8(32'hbc4e93e3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc9873),
	.w1(32'hbb827979),
	.w2(32'hbcfa2148),
	.w3(32'h3a785f4e),
	.w4(32'h3cbddb6b),
	.w5(32'h3c165b1e),
	.w6(32'hbb5cb149),
	.w7(32'hbbaa6286),
	.w8(32'h3bfe29ec),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2744a4),
	.w1(32'h3c8eaf71),
	.w2(32'h3ca801a3),
	.w3(32'hbc31881e),
	.w4(32'h3c2e2b7d),
	.w5(32'h3c9c1e03),
	.w6(32'h3c1dbea3),
	.w7(32'h3be74be1),
	.w8(32'h39e4cdae),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd39eec),
	.w1(32'h3c64bd50),
	.w2(32'hbb357eab),
	.w3(32'hbbb507f8),
	.w4(32'h39589b67),
	.w5(32'hbc126e2e),
	.w6(32'hbbcc9011),
	.w7(32'hbc8bae89),
	.w8(32'hbbe579fa),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58263e),
	.w1(32'h3b8b9bf7),
	.w2(32'h3b8a4854),
	.w3(32'hbb6eea95),
	.w4(32'h3ae82317),
	.w5(32'h3bc127bc),
	.w6(32'hba7b22c5),
	.w7(32'h3a969f1b),
	.w8(32'hbbbec061),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc8e1a),
	.w1(32'hbb195c7e),
	.w2(32'h3b01edef),
	.w3(32'hb79c5f39),
	.w4(32'hba5377b8),
	.w5(32'hb9790637),
	.w6(32'hbbbabc27),
	.w7(32'hb988b59e),
	.w8(32'hbc355b27),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01faf7),
	.w1(32'h3c04f3b4),
	.w2(32'h3b75cf0c),
	.w3(32'hbb733c1c),
	.w4(32'h3a73f67d),
	.w5(32'h3ad2a48d),
	.w6(32'hbad3fdde),
	.w7(32'hbc55bf80),
	.w8(32'hbc45d1f2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00fc65),
	.w1(32'hbb730ba1),
	.w2(32'h3c50f85c),
	.w3(32'hba87b2fc),
	.w4(32'h3b1ffc42),
	.w5(32'h3b696a4e),
	.w6(32'hba8486e8),
	.w7(32'h3c341f9e),
	.w8(32'h3bdbd77f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d14e807),
	.w1(32'hbd03a1f8),
	.w2(32'hbd3c8dcc),
	.w3(32'hbd3ce906),
	.w4(32'hbd5aa661),
	.w5(32'hbd86a9ee),
	.w6(32'hbd5d6b0b),
	.w7(32'h3c1900ac),
	.w8(32'hbbdabaf1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5209b3),
	.w1(32'hbb9b91a4),
	.w2(32'h3bba2522),
	.w3(32'h3a6037c2),
	.w4(32'hbb90661f),
	.w5(32'h3bcfadf4),
	.w6(32'hbb096c88),
	.w7(32'h3badf04a),
	.w8(32'hbaeb03ac),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f20d5),
	.w1(32'h3a90bfd0),
	.w2(32'h3b629c72),
	.w3(32'h3c033121),
	.w4(32'hbb603be0),
	.w5(32'hba1d676b),
	.w6(32'hbb469190),
	.w7(32'hbb2cf26e),
	.w8(32'h3bf28228),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a822b),
	.w1(32'hbc1e4193),
	.w2(32'hbce282f3),
	.w3(32'h3c06fa2d),
	.w4(32'h3c2131a0),
	.w5(32'hbb553666),
	.w6(32'hbc739851),
	.w7(32'hbc5dcdd1),
	.w8(32'hbb6d6791),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e8513),
	.w1(32'h3ba98d8d),
	.w2(32'h3b864788),
	.w3(32'hbca9741c),
	.w4(32'hbbb17e66),
	.w5(32'hbb289e0a),
	.w6(32'h3c489932),
	.w7(32'h3c30cdeb),
	.w8(32'h3bab0da4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaf2b9),
	.w1(32'h3c352581),
	.w2(32'h3c074d8c),
	.w3(32'h3b8569ff),
	.w4(32'h3c8754c1),
	.w5(32'h3c5711a0),
	.w6(32'hbc5700a8),
	.w7(32'h3be1c6d0),
	.w8(32'h3a05f8c3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af735a5),
	.w1(32'hbbe885e8),
	.w2(32'hbc7b6ba8),
	.w3(32'h3b928fa0),
	.w4(32'h3bae2fdb),
	.w5(32'hbbb3c6cc),
	.w6(32'hbc250812),
	.w7(32'h3a1a7f65),
	.w8(32'h3bca1baa),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9f72e),
	.w1(32'hbb820ea1),
	.w2(32'hbbea11e3),
	.w3(32'hbc23743c),
	.w4(32'h3a81bb92),
	.w5(32'hba8b8ff0),
	.w6(32'hbbfa1bef),
	.w7(32'hbc23642c),
	.w8(32'hbba3aeaa),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc521cb4),
	.w1(32'hbc4295db),
	.w2(32'hbc21da9d),
	.w3(32'hbbe4ae30),
	.w4(32'hbc78ee04),
	.w5(32'hbbf8aae4),
	.w6(32'hba8d4b0a),
	.w7(32'hbbce1e08),
	.w8(32'hbc2ba847),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde079c),
	.w1(32'h3ac26e44),
	.w2(32'h3c0ee5e4),
	.w3(32'hbb57ad70),
	.w4(32'hbc10a49e),
	.w5(32'h3b08cc04),
	.w6(32'h3adb8504),
	.w7(32'h3bd07e19),
	.w8(32'hb9ba1a49),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c337383),
	.w1(32'h3c5fcd68),
	.w2(32'h3c57d580),
	.w3(32'h3bb28f2d),
	.w4(32'h3c157b24),
	.w5(32'h3c117a85),
	.w6(32'h3c0add63),
	.w7(32'h3b789c41),
	.w8(32'h3a3a8a11),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec39c),
	.w1(32'hbbce20ff),
	.w2(32'hbc487db8),
	.w3(32'h3a955ad2),
	.w4(32'hbb8cb47d),
	.w5(32'hbc4d8af6),
	.w6(32'hbbc11a95),
	.w7(32'hbc09a1c7),
	.w8(32'hbc42b89e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc781460),
	.w1(32'h3aa19f24),
	.w2(32'h3c068402),
	.w3(32'hbc3b8e30),
	.w4(32'hbaa79483),
	.w5(32'h3aef01b9),
	.w6(32'hbb2b9b0c),
	.w7(32'hbb8993ab),
	.w8(32'hbb6c2529),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2c978),
	.w1(32'h3b98d1f5),
	.w2(32'hbb3fedbd),
	.w3(32'hb9dda88c),
	.w4(32'h3b3f54b2),
	.w5(32'hbb4d06e3),
	.w6(32'h3c223db4),
	.w7(32'h3b9aed5b),
	.w8(32'h3a2ae894),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1a379),
	.w1(32'h3b5c3a72),
	.w2(32'hbd0a0764),
	.w3(32'h3ba78949),
	.w4(32'h3cbde972),
	.w5(32'hbc16fa3c),
	.w6(32'hbc20e24d),
	.w7(32'hbc8b6cfc),
	.w8(32'h3bfff04e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012558),
	.w1(32'hbc0ee33a),
	.w2(32'h3c047c69),
	.w3(32'hbc2659a0),
	.w4(32'hbc4ae09e),
	.w5(32'hbba2084d),
	.w6(32'hbb4b7d68),
	.w7(32'h3c4bf6f7),
	.w8(32'h3b4a8a3e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c488f06),
	.w1(32'h3b687c1d),
	.w2(32'hbc90e669),
	.w3(32'hbb74fa10),
	.w4(32'h3bd6c918),
	.w5(32'hbbf8d636),
	.w6(32'hbae208fb),
	.w7(32'hbc8db7da),
	.w8(32'hbbae31d8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8187e4),
	.w1(32'hbc593904),
	.w2(32'h39264c1b),
	.w3(32'hbb434dc5),
	.w4(32'hbc72244d),
	.w5(32'hbb5fe9de),
	.w6(32'hbbb337f7),
	.w7(32'hb6dffb6d),
	.w8(32'hbc14b2ec),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec7512),
	.w1(32'h3bd93edc),
	.w2(32'h3bac6763),
	.w3(32'hbc1a7e32),
	.w4(32'h3b9101c3),
	.w5(32'h3b67e8e0),
	.w6(32'h3b90aff3),
	.w7(32'h3abaf1c1),
	.w8(32'hbb02298e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf809c0),
	.w1(32'h3b978789),
	.w2(32'hbbf1a5d8),
	.w3(32'h3aab2175),
	.w4(32'h3c6bea21),
	.w5(32'h3bf975f4),
	.w6(32'hbb88581f),
	.w7(32'hbc8235e3),
	.w8(32'hbc96e1fb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad4f34),
	.w1(32'h3c372013),
	.w2(32'h3bc1a42a),
	.w3(32'hbc6a030e),
	.w4(32'hbbce31e7),
	.w5(32'h3aff0510),
	.w6(32'h3c012e58),
	.w7(32'hbbc05580),
	.w8(32'hbb9cc265),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15bbe8),
	.w1(32'h3c0a9bc4),
	.w2(32'h3c410cda),
	.w3(32'h3bb3632c),
	.w4(32'hba871c74),
	.w5(32'h3c233318),
	.w6(32'h3bd96ae8),
	.w7(32'h3a94d527),
	.w8(32'h3aea55dc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acef4ce),
	.w1(32'hbbcad9e2),
	.w2(32'hbc2a0f58),
	.w3(32'h397eb878),
	.w4(32'h3c0111ce),
	.w5(32'hbcbd3f4e),
	.w6(32'hbc09c31b),
	.w7(32'hbb9091ab),
	.w8(32'h3bbde1f5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76e2ea),
	.w1(32'h3c6d836d),
	.w2(32'h3ac306d4),
	.w3(32'hbbaac6f8),
	.w4(32'h3c1d2b18),
	.w5(32'h389fe652),
	.w6(32'h3c3f7950),
	.w7(32'h3c0f5834),
	.w8(32'h3c062ba3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84b290),
	.w1(32'hbc81fe30),
	.w2(32'hbc8f1e99),
	.w3(32'hbc3ab449),
	.w4(32'hbc0b69e9),
	.w5(32'hbbfbb824),
	.w6(32'hbbf1bba7),
	.w7(32'hbcb2c229),
	.w8(32'hbbc7f95f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc377b86),
	.w1(32'hbb554386),
	.w2(32'hb95f32dc),
	.w3(32'hbc191bb3),
	.w4(32'hbc10c830),
	.w5(32'hbc09b646),
	.w6(32'hbb8f9705),
	.w7(32'hbb5edbd7),
	.w8(32'hbba92959),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1d766),
	.w1(32'hbb5e8b39),
	.w2(32'hbc21c861),
	.w3(32'hbb6bee8c),
	.w4(32'h3ca018bb),
	.w5(32'h3c064af2),
	.w6(32'hbb8ce5ba),
	.w7(32'hbb0f63a7),
	.w8(32'h3c201148),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc26443),
	.w1(32'h3d18b0f3),
	.w2(32'h3c53d68e),
	.w3(32'h3b3742ff),
	.w4(32'h3c5af70c),
	.w5(32'h3d42b595),
	.w6(32'h3c0da1ae),
	.w7(32'hbc7f8a3c),
	.w8(32'hbb41499c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe390a1),
	.w1(32'h3b90d5d9),
	.w2(32'hbcd375ce),
	.w3(32'h3c33f16c),
	.w4(32'h3c1f7017),
	.w5(32'hbc6fe500),
	.w6(32'hbc0b21b1),
	.w7(32'hbc46a941),
	.w8(32'h3c1068b0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b52fe),
	.w1(32'hbc49d2e2),
	.w2(32'h3c0fc6c6),
	.w3(32'hbc29b157),
	.w4(32'hbbd2281e),
	.w5(32'h398504e9),
	.w6(32'hbc0d17c4),
	.w7(32'h3ba53083),
	.w8(32'h3b9d4b03),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d1db3),
	.w1(32'hb96ae51a),
	.w2(32'h3c0f2b3b),
	.w3(32'hbb820733),
	.w4(32'hbc3562fb),
	.w5(32'h3a037b72),
	.w6(32'h3a3b1e61),
	.w7(32'h3b548859),
	.w8(32'h3c1488c8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa13ee),
	.w1(32'hbbb2317e),
	.w2(32'hbbdf34ef),
	.w3(32'hba93d1d2),
	.w4(32'hbb57d9a7),
	.w5(32'hbba57906),
	.w6(32'hbbf429c6),
	.w7(32'hbc0bf9d4),
	.w8(32'hbc2ecb2f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba17fc7),
	.w1(32'h3bac1c9b),
	.w2(32'h3c0953b7),
	.w3(32'hbb64c43d),
	.w4(32'h3b8e26f4),
	.w5(32'h3c320777),
	.w6(32'h3b5aca0c),
	.w7(32'h3bb75f09),
	.w8(32'h3aa9de9e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa10023),
	.w1(32'h3c4d96f1),
	.w2(32'h3c83e99e),
	.w3(32'h3b2281cd),
	.w4(32'h3ba93cce),
	.w5(32'h3c2acb7f),
	.w6(32'h3bc53929),
	.w7(32'h3b5f60f7),
	.w8(32'hbbf0f7c2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2613a0),
	.w1(32'h3b0cd817),
	.w2(32'h3c9fcb65),
	.w3(32'h3978647c),
	.w4(32'hbc587cec),
	.w5(32'hba33217a),
	.w6(32'h3adf92ed),
	.w7(32'h3b581c83),
	.w8(32'hbbcbcfbb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf26b69),
	.w1(32'hbc074137),
	.w2(32'hbb4d5bca),
	.w3(32'h3ba5217d),
	.w4(32'hbc472f75),
	.w5(32'hbc2705f0),
	.w6(32'h3c320a9e),
	.w7(32'h3c3f783f),
	.w8(32'h3c4c3c98),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cb1ef),
	.w1(32'h3981255d),
	.w2(32'hb8bb7644),
	.w3(32'h3c899edf),
	.w4(32'h3be2bcfa),
	.w5(32'h3ba1b861),
	.w6(32'h3bd4aec0),
	.w7(32'h3b6fe827),
	.w8(32'h3aa4c7a2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8490ac),
	.w1(32'hbbeab2a7),
	.w2(32'hbc6440b4),
	.w3(32'h3ba1b051),
	.w4(32'hbb7558c3),
	.w5(32'hbc44efbf),
	.w6(32'hbbaea77c),
	.w7(32'hbbaba590),
	.w8(32'hbbd90fd8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1fee),
	.w1(32'h3bdb3541),
	.w2(32'h3a6e9594),
	.w3(32'hbbc32837),
	.w4(32'h3be6cb42),
	.w5(32'h3c509342),
	.w6(32'h3b5711e0),
	.w7(32'hbb32f71a),
	.w8(32'h3af52ccc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01b103),
	.w1(32'hbc65de50),
	.w2(32'hbbcac424),
	.w3(32'h3b848811),
	.w4(32'hbc33010e),
	.w5(32'hbc29f47f),
	.w6(32'h3b9bcccd),
	.w7(32'h3c5cf9fa),
	.w8(32'h3bd1161a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7ec7a),
	.w1(32'h3bf2945a),
	.w2(32'hbcb8b307),
	.w3(32'hbc02e55b),
	.w4(32'h3c9709ca),
	.w5(32'hbbbbc6ec),
	.w6(32'hbae816fc),
	.w7(32'hbc3b75aa),
	.w8(32'hbc06495c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83c334),
	.w1(32'hbb2430f4),
	.w2(32'hbcf09589),
	.w3(32'hbb99ad48),
	.w4(32'hbade4f15),
	.w5(32'hbba22522),
	.w6(32'hbcc1b602),
	.w7(32'hbbcb1503),
	.w8(32'hb892a08f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b461b),
	.w1(32'hbc7d83d3),
	.w2(32'hbc75ba9e),
	.w3(32'hbcf303ff),
	.w4(32'hbc9f099d),
	.w5(32'hbb965569),
	.w6(32'hbbf1a3ca),
	.w7(32'hbc97eebc),
	.w8(32'hbcbe9a43),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f1f81),
	.w1(32'h3c2e7e26),
	.w2(32'h3b64d8db),
	.w3(32'hbc3b19dc),
	.w4(32'h3c1b9457),
	.w5(32'h3c162fde),
	.w6(32'h3b2b418a),
	.w7(32'hbbb39262),
	.w8(32'hbb66a8b6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ef70a),
	.w1(32'h39f9416b),
	.w2(32'hbb639dbd),
	.w3(32'hbb5fe2ad),
	.w4(32'h3b72a124),
	.w5(32'h3c1b4991),
	.w6(32'h3aba1284),
	.w7(32'h3bd5ae28),
	.w8(32'h3b18fdb6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc373d5e),
	.w1(32'h3b9777b2),
	.w2(32'h39cc983a),
	.w3(32'h3c016932),
	.w4(32'h3b36f9a9),
	.w5(32'h3c17fe10),
	.w6(32'h3ba490d0),
	.w7(32'hbb5d805d),
	.w8(32'h3abbe2cc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fb430),
	.w1(32'h3c0d6e09),
	.w2(32'h3c0b3594),
	.w3(32'h3ba6e81b),
	.w4(32'h3b8a8c5c),
	.w5(32'h3b60df5a),
	.w6(32'hb9f7e65e),
	.w7(32'h3bdc6ae0),
	.w8(32'h3b8ff10a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb769499),
	.w1(32'hbbea909a),
	.w2(32'hbaadefcf),
	.w3(32'hba9d31ef),
	.w4(32'hbb4cd758),
	.w5(32'hba281c54),
	.w6(32'hbc53d18f),
	.w7(32'hbc606728),
	.w8(32'h3a8ea571),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91e8bb),
	.w1(32'hbbe1714c),
	.w2(32'hbcaccee8),
	.w3(32'hbbb901d2),
	.w4(32'hbc00f433),
	.w5(32'hbc6dfc35),
	.w6(32'hbc434d1e),
	.w7(32'hbc611fc6),
	.w8(32'h3ad4fad8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd288d1),
	.w1(32'h3b817c4e),
	.w2(32'h3c0e9e54),
	.w3(32'hbaf3e1d9),
	.w4(32'h3b58103b),
	.w5(32'hbb27c45e),
	.w6(32'h3b3bd03d),
	.w7(32'h3c02f863),
	.w8(32'h3c0027ec),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf614e7),
	.w1(32'h37c42794),
	.w2(32'hb84e1a70),
	.w3(32'hbbc68986),
	.w4(32'hbbac9cad),
	.w5(32'hbc0ce28b),
	.w6(32'hbb961f0a),
	.w7(32'hbb89d748),
	.w8(32'h3bb606c7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf25f2),
	.w1(32'h3c0657b7),
	.w2(32'hbc860020),
	.w3(32'hbb475536),
	.w4(32'h3c7fb702),
	.w5(32'h3c38367c),
	.w6(32'hb99bcc2a),
	.w7(32'hbbe3c2a8),
	.w8(32'h3c0abe53),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f4e7d),
	.w1(32'hba711a5a),
	.w2(32'hbc908aa2),
	.w3(32'hbb66d74f),
	.w4(32'h3b85121b),
	.w5(32'hbc93f11b),
	.w6(32'hbc87f9b5),
	.w7(32'h3a90baab),
	.w8(32'h3c2e9983),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8955c2),
	.w1(32'h3aacf7dd),
	.w2(32'hbc31f606),
	.w3(32'h3bace17c),
	.w4(32'h3c6a3dd1),
	.w5(32'h3b1cc467),
	.w6(32'hbb1354b9),
	.w7(32'h3b06eadc),
	.w8(32'h39e667cd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2122ec),
	.w1(32'hbc061095),
	.w2(32'hbc76614c),
	.w3(32'hbc959086),
	.w4(32'h3ab12811),
	.w5(32'h3ace74e1),
	.w6(32'hbca3ae4f),
	.w7(32'hbc2986b6),
	.w8(32'h3b15cd8b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26f03e),
	.w1(32'hbc2a57d4),
	.w2(32'hbca5eb91),
	.w3(32'hbc88639a),
	.w4(32'hbc2119d9),
	.w5(32'hbca179da),
	.w6(32'hbc7caeb1),
	.w7(32'hbc9da42a),
	.w8(32'hbb5e9d54),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56ee95),
	.w1(32'h3b73fb38),
	.w2(32'hbc31072d),
	.w3(32'hbc169fd4),
	.w4(32'h3c2e3f2d),
	.w5(32'h3bca9f16),
	.w6(32'h3ad72904),
	.w7(32'hb9de9587),
	.w8(32'h3c4f9424),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad92e1e),
	.w1(32'hbc797feb),
	.w2(32'hbd0059c1),
	.w3(32'hbbcd5297),
	.w4(32'hbbd23a45),
	.w5(32'hbc3009ad),
	.w6(32'hbc4b86cb),
	.w7(32'hb954153f),
	.w8(32'h3c40c8dd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc850625),
	.w1(32'hbbe3d458),
	.w2(32'hbbee3b09),
	.w3(32'hbca6ad94),
	.w4(32'h3bf4156f),
	.w5(32'h3a4dea9d),
	.w6(32'h3ba42b96),
	.w7(32'hba9eb229),
	.w8(32'hbc24dc8c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68cd40),
	.w1(32'h3c113312),
	.w2(32'hbb1bfca9),
	.w3(32'hbbe3a6fe),
	.w4(32'h3bd8e77a),
	.w5(32'h3bc714c5),
	.w6(32'hbbad6688),
	.w7(32'hbc3ed742),
	.w8(32'hbb891920),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66339b),
	.w1(32'h3b88f901),
	.w2(32'h3c26dede),
	.w3(32'h3b82629e),
	.w4(32'hbbc6a829),
	.w5(32'hba12d1ea),
	.w6(32'h3c57f180),
	.w7(32'h3c91d2d9),
	.w8(32'h3b3eb741),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8432b7),
	.w1(32'hba851d64),
	.w2(32'hbc0430d9),
	.w3(32'h3c359cc5),
	.w4(32'h3b2672dd),
	.w5(32'hbaa24e4b),
	.w6(32'hbbdfcb6c),
	.w7(32'hbbc8c041),
	.w8(32'hba1457c7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea0fc5),
	.w1(32'hbbb7fbec),
	.w2(32'hbc8ff1a8),
	.w3(32'hbbb6b94f),
	.w4(32'hbba41a2f),
	.w5(32'hba932f41),
	.w6(32'hbb899da6),
	.w7(32'hbbc09838),
	.w8(32'hbbf00e50),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5daa5b),
	.w1(32'h3c2964df),
	.w2(32'hba8c9ec0),
	.w3(32'hbbddd2ae),
	.w4(32'h3bcc53d9),
	.w5(32'h3c258312),
	.w6(32'h3b2a779b),
	.w7(32'h3c197938),
	.w8(32'h3beba2d5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0d22),
	.w1(32'hba603e62),
	.w2(32'hbbae9230),
	.w3(32'h3b2c591d),
	.w4(32'hbb5c282f),
	.w5(32'h3b8291a1),
	.w6(32'hbbf858fd),
	.w7(32'h3bb4a54d),
	.w8(32'h3a344c09),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41b18a),
	.w1(32'h3a35d58d),
	.w2(32'h3b6db007),
	.w3(32'hbbeb2d04),
	.w4(32'h3aea8d3a),
	.w5(32'h3bda9bc9),
	.w6(32'hbadb27ac),
	.w7(32'h389659ee),
	.w8(32'h3a587b9f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb380de),
	.w1(32'h3b915659),
	.w2(32'h39f17e6a),
	.w3(32'h3baa8be9),
	.w4(32'h3bb66742),
	.w5(32'h3b298a5b),
	.w6(32'h3a8faf71),
	.w7(32'h3a771a11),
	.w8(32'hbae002e4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fa254),
	.w1(32'h3cb095db),
	.w2(32'h3cf16c41),
	.w3(32'h3b8f2486),
	.w4(32'h3b36aa3d),
	.w5(32'h3cd3abe9),
	.w6(32'h3c1d9628),
	.w7(32'h3a4a480a),
	.w8(32'hbbb49ea6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab17802),
	.w1(32'hbbbce0d6),
	.w2(32'hbb7382d5),
	.w3(32'h3b8cfc07),
	.w4(32'hbc24499c),
	.w5(32'hbbf8a3cb),
	.w6(32'h3b965bb8),
	.w7(32'h3b1886f9),
	.w8(32'h399d79ca),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c301c),
	.w1(32'h3b0aabae),
	.w2(32'hbbc63bcc),
	.w3(32'hbb8435fb),
	.w4(32'h3a865322),
	.w5(32'hbbc0f5d8),
	.w6(32'hbc0c63b4),
	.w7(32'hbc45e512),
	.w8(32'hbbb9fe3d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a8562),
	.w1(32'h3b9c4a9b),
	.w2(32'h3aa37949),
	.w3(32'hbb7cffba),
	.w4(32'h3ab16ef7),
	.w5(32'hbbc7cf45),
	.w6(32'h3b9e8923),
	.w7(32'hbc2395fe),
	.w8(32'h3bac402a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826893),
	.w1(32'h3be9b45f),
	.w2(32'hbc628fa9),
	.w3(32'hb9cd2be9),
	.w4(32'h3be63cf0),
	.w5(32'hbbb48d7a),
	.w6(32'hb7931b16),
	.w7(32'hbc00f06e),
	.w8(32'hbbb257b4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80f2f6),
	.w1(32'hbc2a84ad),
	.w2(32'h3c3b6abf),
	.w3(32'hbbf60bf7),
	.w4(32'hbc57b84a),
	.w5(32'hbc484a19),
	.w6(32'hbaca0458),
	.w7(32'h3c9f3a56),
	.w8(32'h3c01a326),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb01fa4),
	.w1(32'hbc190ae1),
	.w2(32'hbd002492),
	.w3(32'h3bde7fb5),
	.w4(32'h3ce9a32d),
	.w5(32'hbb0024ed),
	.w6(32'hbc631aba),
	.w7(32'h3b41f35d),
	.w8(32'h3bb57535),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ac0d1),
	.w1(32'h3bcf42ac),
	.w2(32'h3c6337ce),
	.w3(32'hbc0fc5f0),
	.w4(32'hbc2e5e96),
	.w5(32'h3bc1310f),
	.w6(32'h3b9f2be8),
	.w7(32'hbb436a5f),
	.w8(32'hbc3af9ef),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a975e6),
	.w1(32'hbbbbc0b8),
	.w2(32'hbc9c82b6),
	.w3(32'h3ba10b27),
	.w4(32'h3c953eb2),
	.w5(32'h3b34456f),
	.w6(32'hbbe62fc1),
	.w7(32'h3b62108e),
	.w8(32'h3c4d3ab8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72a725),
	.w1(32'h3c8b6f93),
	.w2(32'h3c3a6398),
	.w3(32'hbc0c02b9),
	.w4(32'h3bc11abc),
	.w5(32'h3c757d6c),
	.w6(32'hba3403a0),
	.w7(32'h3a8d6ca5),
	.w8(32'hbb9e7b18),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934df3),
	.w1(32'h3b678c1c),
	.w2(32'hbad35524),
	.w3(32'h3b22bcf9),
	.w4(32'h3bef78b0),
	.w5(32'hbb1b6524),
	.w6(32'hbc236d52),
	.w7(32'h3beb2efc),
	.w8(32'h3c4fd9da),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae7a5e),
	.w1(32'hbb805c95),
	.w2(32'hbc048135),
	.w3(32'hbc07f4e9),
	.w4(32'hbbbf19f3),
	.w5(32'hbbd8c188),
	.w6(32'hbc3e91eb),
	.w7(32'hbc7d89e0),
	.w8(32'hbc6597c6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbade622),
	.w1(32'h3af2fb45),
	.w2(32'hbc5a6231),
	.w3(32'hbbc4d3ef),
	.w4(32'hbbc85e4e),
	.w5(32'hbb5af98a),
	.w6(32'hbc0e8bc8),
	.w7(32'hbc804d5d),
	.w8(32'hbbdeb247),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b6b6a),
	.w1(32'hbb64a61f),
	.w2(32'h3b4c3c42),
	.w3(32'hbc0dad97),
	.w4(32'hbc990b84),
	.w5(32'hbbd4de80),
	.w6(32'hbc3ad6f0),
	.w7(32'h3a67391c),
	.w8(32'hb90be318),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fae0f),
	.w1(32'hbb8235e1),
	.w2(32'hbc0df5aa),
	.w3(32'hbbcde9ce),
	.w4(32'hbc0c3461),
	.w5(32'hbbdabe0b),
	.w6(32'hba46e379),
	.w7(32'hbc1ef346),
	.w8(32'hbc3274a6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb0f0),
	.w1(32'h3ac6407a),
	.w2(32'hb9e31d07),
	.w3(32'hbabc9a3f),
	.w4(32'h3ac5210c),
	.w5(32'hbb6eff21),
	.w6(32'h3aecbdf8),
	.w7(32'h3b855ca7),
	.w8(32'h3b3fec19),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba845c4d),
	.w1(32'hbc9656d4),
	.w2(32'hbb625d85),
	.w3(32'hbb79fd51),
	.w4(32'h3bf4455f),
	.w5(32'hbc114aaa),
	.w6(32'h3c074b2c),
	.w7(32'h3c091799),
	.w8(32'h3b03a1e5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92f2de),
	.w1(32'hbb557236),
	.w2(32'hbb5bedca),
	.w3(32'hbc5c3864),
	.w4(32'hba6b9660),
	.w5(32'hbac2cf16),
	.w6(32'hb9cf0c7d),
	.w7(32'hba44f617),
	.w8(32'hbabdc35d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ea12),
	.w1(32'h3b387694),
	.w2(32'h3b3c2070),
	.w3(32'h3b7a997b),
	.w4(32'h3b6761c0),
	.w5(32'h3b3e9f9d),
	.w6(32'h39c31604),
	.w7(32'hbae772a0),
	.w8(32'h39f48940),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb057f93),
	.w1(32'h3b0c2af4),
	.w2(32'hbb06bcde),
	.w3(32'hbb6f24a2),
	.w4(32'hbb03d6da),
	.w5(32'h3a0590af),
	.w6(32'h3aacd634),
	.w7(32'h3b977599),
	.w8(32'h3aad4b73),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f1a17),
	.w1(32'hbb48f2ce),
	.w2(32'hbcac9b62),
	.w3(32'hbc57949e),
	.w4(32'h3c20fb7e),
	.w5(32'hb9f69569),
	.w6(32'hbc0bbb05),
	.w7(32'hbc3e8afe),
	.w8(32'h3aab1b3b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb873aa6),
	.w1(32'hba03631f),
	.w2(32'hbb4a9ef1),
	.w3(32'hbb901ac6),
	.w4(32'hbb4eeee5),
	.w5(32'hbbb6e12a),
	.w6(32'h399a14e3),
	.w7(32'h3b872a40),
	.w8(32'h3ba1745f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b937398),
	.w1(32'hbaad8b37),
	.w2(32'hba80f7e4),
	.w3(32'hb8439b3a),
	.w4(32'hbc3d5a82),
	.w5(32'hbbcbb898),
	.w6(32'h3af600a1),
	.w7(32'hba91c025),
	.w8(32'hbb965457),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e7912),
	.w1(32'hb9fbb7df),
	.w2(32'h3a52188e),
	.w3(32'hbaeeace1),
	.w4(32'hbaca639b),
	.w5(32'hbc20bac2),
	.w6(32'hbbae7da6),
	.w7(32'hbbb09772),
	.w8(32'hbae92b0c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b893d77),
	.w1(32'hbb4df200),
	.w2(32'hbca477a1),
	.w3(32'hbb90d2fb),
	.w4(32'hba40038f),
	.w5(32'hbbb74ab7),
	.w6(32'hbc5e662c),
	.w7(32'hbb9de28e),
	.w8(32'hbbd2b124),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc41863),
	.w1(32'hba0ec665),
	.w2(32'hbb56c768),
	.w3(32'hbc8626e3),
	.w4(32'h3b85a4ff),
	.w5(32'hbad99359),
	.w6(32'hbb9d8dbb),
	.w7(32'hbc2ae39a),
	.w8(32'h3ad67a77),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb856073),
	.w1(32'h3a70da3e),
	.w2(32'hbd0f56c2),
	.w3(32'hbb5fa15d),
	.w4(32'h3b970057),
	.w5(32'hbb953ffe),
	.w6(32'hbca5baaf),
	.w7(32'hbc797f58),
	.w8(32'h3b043550),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73c101),
	.w1(32'h3bfb927a),
	.w2(32'hbc853cec),
	.w3(32'hbc8f522b),
	.w4(32'h3b4f89b1),
	.w5(32'h3bc294ba),
	.w6(32'hbb54f43c),
	.w7(32'h3b827ee3),
	.w8(32'hbadac186),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb820f202),
	.w1(32'hbb939ea7),
	.w2(32'hbb3a57b1),
	.w3(32'h39696f8e),
	.w4(32'hb9cf0b51),
	.w5(32'hbb7a0ed4),
	.w6(32'hbb35c7f1),
	.w7(32'hbb5cb47b),
	.w8(32'hbbcbce04),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c99d9),
	.w1(32'h3a034511),
	.w2(32'h3b33b3a0),
	.w3(32'h3b958c0e),
	.w4(32'h3956ec0c),
	.w5(32'hbbe9da94),
	.w6(32'hbb6817ac),
	.w7(32'hb9b5c7ab),
	.w8(32'hbb6bcdae),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3db21),
	.w1(32'h3cafdefa),
	.w2(32'h3c3e1858),
	.w3(32'h3b2eca4a),
	.w4(32'h3c05b65c),
	.w5(32'h3c798e9f),
	.w6(32'h3c18ab94),
	.w7(32'hbbbc00cd),
	.w8(32'h3b0bf055),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd89179),
	.w1(32'h3c744620),
	.w2(32'h3c5a0fed),
	.w3(32'h3be3e481),
	.w4(32'h3b8b267d),
	.w5(32'h3c049462),
	.w6(32'h3c024ec0),
	.w7(32'h3bc60e19),
	.w8(32'h3ba21cde),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ecfef),
	.w1(32'h3841e883),
	.w2(32'hb9ba6aa2),
	.w3(32'hb9fd1cee),
	.w4(32'h3a9e74f4),
	.w5(32'hbacb315d),
	.w6(32'hbb04de17),
	.w7(32'h3a096f3b),
	.w8(32'hba03d456),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a696de),
	.w1(32'hbb9fdeb8),
	.w2(32'hbc57a920),
	.w3(32'hba155db9),
	.w4(32'hbbc44a1d),
	.w5(32'hbb3e5639),
	.w6(32'h3aa864e8),
	.w7(32'h39f21859),
	.w8(32'h3c2b6d99),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule