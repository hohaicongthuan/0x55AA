module layer_10_featuremap_80(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd1949),
	.w1(32'h3acb1f24),
	.w2(32'hbb6646cc),
	.w3(32'h3871c2f0),
	.w4(32'h3b83e3d0),
	.w5(32'h3b5fbbf4),
	.w6(32'hbd5abde1),
	.w7(32'hbad65b5c),
	.w8(32'hbaba734f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ed77f),
	.w1(32'h3a89d249),
	.w2(32'hbae94758),
	.w3(32'h3b1f7ed0),
	.w4(32'h3be9309a),
	.w5(32'hbae9ceaa),
	.w6(32'hbbecc084),
	.w7(32'hbb0c3bac),
	.w8(32'h3ba2703b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818f27),
	.w1(32'hbb65b3cf),
	.w2(32'hbc4b7a93),
	.w3(32'h3bbaaed4),
	.w4(32'hbc063eed),
	.w5(32'hbae5c3e2),
	.w6(32'hbbc9fdc2),
	.w7(32'hbba03e01),
	.w8(32'hbbd5f8e6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23240d),
	.w1(32'hba8d2761),
	.w2(32'hba8b9a1d),
	.w3(32'hb8b7d23b),
	.w4(32'h3b34c57f),
	.w5(32'hbbba9f68),
	.w6(32'hba841d5f),
	.w7(32'hbbb55fd2),
	.w8(32'h3c123aea),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b120d91),
	.w1(32'hbb8a1006),
	.w2(32'hbb8984a2),
	.w3(32'h3aa13333),
	.w4(32'hbbf2e6e1),
	.w5(32'hbb2dbefb),
	.w6(32'h3ba7b7ca),
	.w7(32'h3baaf999),
	.w8(32'h3cf7c3ab),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0258a3),
	.w1(32'hbb2cce2f),
	.w2(32'h3af364ab),
	.w3(32'hbb7b8cb5),
	.w4(32'hbc3280c0),
	.w5(32'hbb0ffbcf),
	.w6(32'hbce29e38),
	.w7(32'hbaca6b59),
	.w8(32'hbad567a8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7fbb9),
	.w1(32'hb9e126d3),
	.w2(32'hb8dfa9df),
	.w3(32'h3b671714),
	.w4(32'hbbfacbdc),
	.w5(32'hbcff13a8),
	.w6(32'hb9b3aa77),
	.w7(32'h3b311ee4),
	.w8(32'h3d5d086a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe34c),
	.w1(32'hba9737a4),
	.w2(32'hbc69a7c5),
	.w3(32'hbc5800f7),
	.w4(32'hbbfb0e6d),
	.w5(32'h3ab9295c),
	.w6(32'hbc692cee),
	.w7(32'hbac9ba5e),
	.w8(32'hbbc76c7f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44501d),
	.w1(32'hba9d5a12),
	.w2(32'hbc0bd177),
	.w3(32'hbb8bb4ed),
	.w4(32'hbbcf0c4c),
	.w5(32'h3b69c3da),
	.w6(32'h3a2fdd7a),
	.w7(32'hbb168c7c),
	.w8(32'h3a20d569),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e9e67),
	.w1(32'h3a7b37cf),
	.w2(32'hbbeb8325),
	.w3(32'hbb7fb9c5),
	.w4(32'h39778bad),
	.w5(32'hbc131deb),
	.w6(32'hbb8dbcba),
	.w7(32'h3c4aeed4),
	.w8(32'hbc1ad495),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b48cc),
	.w1(32'hb999157a),
	.w2(32'h3ae10755),
	.w3(32'h3ab9cdeb),
	.w4(32'h3d66bdf8),
	.w5(32'hbd50bbc8),
	.w6(32'h3bd1be6f),
	.w7(32'hb802d467),
	.w8(32'hbb22d815),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2b6092),
	.w1(32'h3b1ad1fc),
	.w2(32'h3c3bfd00),
	.w3(32'h37e46a5a),
	.w4(32'h3caaa1d5),
	.w5(32'hbb119d30),
	.w6(32'h3ae632a8),
	.w7(32'h3a52b6be),
	.w8(32'hbb1c207f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb991f6e),
	.w1(32'hbbb72b66),
	.w2(32'hbba91092),
	.w3(32'hbb65e94f),
	.w4(32'hbbc6f716),
	.w5(32'hbbac8a56),
	.w6(32'h3a5e25c0),
	.w7(32'hbb7daade),
	.w8(32'hba874ac4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c350b83),
	.w1(32'h3c50b88c),
	.w2(32'hbaea0891),
	.w3(32'hbb8eed14),
	.w4(32'hbaa65aff),
	.w5(32'h3b15d2ac),
	.w6(32'h3bf15ab2),
	.w7(32'h3d895150),
	.w8(32'hbb37c287),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896a4c),
	.w1(32'hbb54a5de),
	.w2(32'hbb1a1d5b),
	.w3(32'hbbaec405),
	.w4(32'h390dbf90),
	.w5(32'hb9b2b3ef),
	.w6(32'h3c42d7ec),
	.w7(32'h3c40bd17),
	.w8(32'hbc778e22),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4150e9),
	.w1(32'hbb0f4b06),
	.w2(32'h3949044c),
	.w3(32'hbd12f049),
	.w4(32'hbb9d7779),
	.w5(32'hbb159bf5),
	.w6(32'hbb1533ce),
	.w7(32'hbb9bea04),
	.w8(32'hbb93253f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962799a),
	.w1(32'h3cf98f74),
	.w2(32'hbb275f8b),
	.w3(32'hb9a3f7ff),
	.w4(32'hb7d742d7),
	.w5(32'h3b844643),
	.w6(32'h3aead6bf),
	.w7(32'hbbc8b4f2),
	.w8(32'hbb360455),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb576c88),
	.w1(32'hbd4229f8),
	.w2(32'hbc94f133),
	.w3(32'hbb72efce),
	.w4(32'hba10cf61),
	.w5(32'hbb343492),
	.w6(32'hbc435750),
	.w7(32'h3c6b08e2),
	.w8(32'hbbad5684),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab1d0e),
	.w1(32'hbd8da7a6),
	.w2(32'hbba53953),
	.w3(32'hb9b84205),
	.w4(32'h3b6624cc),
	.w5(32'h37982d7f),
	.w6(32'hb9995f67),
	.w7(32'hbadd3de6),
	.w8(32'hbbc578ec),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9873b6),
	.w1(32'hbbb13c66),
	.w2(32'h3b43dcff),
	.w3(32'h3b75ce06),
	.w4(32'h3ba04dab),
	.w5(32'h3b98ef97),
	.w6(32'h39e8ba24),
	.w7(32'hbb19760d),
	.w8(32'hbb991694),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a582275),
	.w1(32'hb9ef59c0),
	.w2(32'hbc3cb953),
	.w3(32'hbb6af3ee),
	.w4(32'hbb6cb58a),
	.w5(32'h3b969fb5),
	.w6(32'hbd0c4665),
	.w7(32'hbbc87098),
	.w8(32'h3b866709),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfbc65a),
	.w1(32'h3b9f331e),
	.w2(32'hba1ea300),
	.w3(32'hba002b1a),
	.w4(32'hb98b6aa8),
	.w5(32'hb99af0f9),
	.w6(32'hbba97443),
	.w7(32'h3ab573b2),
	.w8(32'h39c348a2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b6fda),
	.w1(32'hbabf97cb),
	.w2(32'hbc25e8ac),
	.w3(32'hbbae0a16),
	.w4(32'hbb97c3ac),
	.w5(32'hbd0fc24a),
	.w6(32'hbc04821f),
	.w7(32'h3a862a3e),
	.w8(32'hbc79765d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96920bb),
	.w1(32'h3bda50ee),
	.w2(32'hbbb5b4c3),
	.w3(32'h3ba1dbef),
	.w4(32'h3be8c5cb),
	.w5(32'hbaaf67e7),
	.w6(32'hbb002c95),
	.w7(32'h3a833c12),
	.w8(32'hbb974648),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a3e82),
	.w1(32'h39ade9ed),
	.w2(32'hbbd47db3),
	.w3(32'h3aee3fe2),
	.w4(32'hbbe9b707),
	.w5(32'hbbef8b68),
	.w6(32'hbc03525d),
	.w7(32'h3bca46d7),
	.w8(32'hbc5934ca),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ff472),
	.w1(32'h3c27443f),
	.w2(32'h3a8c5f1a),
	.w3(32'hbb8f45da),
	.w4(32'h3c807fa7),
	.w5(32'hb989bc05),
	.w6(32'h3d1b921c),
	.w7(32'hba839363),
	.w8(32'hbb9a9832),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32e6f5),
	.w1(32'h3a9a8cf0),
	.w2(32'hbca8e983),
	.w3(32'hbc0b8237),
	.w4(32'hbb3d141b),
	.w5(32'hba27bbce),
	.w6(32'h3aded8e5),
	.w7(32'hba96066b),
	.w8(32'h39c74b0f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4759a),
	.w1(32'hbbcab563),
	.w2(32'h3b2e1d41),
	.w3(32'hbbd8c875),
	.w4(32'h3bab4753),
	.w5(32'h3ba7e2c0),
	.w6(32'h3c039449),
	.w7(32'hbc8252a2),
	.w8(32'h3b2248e3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27a5ef),
	.w1(32'h3badf411),
	.w2(32'h3b6f0b7c),
	.w3(32'hb92a8592),
	.w4(32'h3b369298),
	.w5(32'h3a1255fe),
	.w6(32'h3b809c39),
	.w7(32'hbb0901c9),
	.w8(32'h3ba3477d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d8d52),
	.w1(32'hbb775d42),
	.w2(32'hbc0dbe61),
	.w3(32'hbbbcf030),
	.w4(32'h3c1d6282),
	.w5(32'hbb25647b),
	.w6(32'h3bc73aec),
	.w7(32'h3c4ab2d7),
	.w8(32'hb6adf226),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955d72),
	.w1(32'h3914f65b),
	.w2(32'hbd6aa1b1),
	.w3(32'h3acbbbc0),
	.w4(32'h393b620b),
	.w5(32'hb92b378e),
	.w6(32'hbb21ea6e),
	.w7(32'hbba13cc7),
	.w8(32'hbc66b213),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdf6f0),
	.w1(32'h3bc9e566),
	.w2(32'h3ad967da),
	.w3(32'h3bbea7be),
	.w4(32'hbbca7b09),
	.w5(32'h3bb9a6ad),
	.w6(32'h3a805773),
	.w7(32'hbbb37deb),
	.w8(32'hbb4daa70),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedb0b3),
	.w1(32'hbb348a1e),
	.w2(32'h3bab03e0),
	.w3(32'hba134da5),
	.w4(32'hbbb73c3a),
	.w5(32'h3a9b0be2),
	.w6(32'hbbccd264),
	.w7(32'hbb96dbb7),
	.w8(32'h3b950324),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb235128),
	.w1(32'hbcee6708),
	.w2(32'hba4fc933),
	.w3(32'h3bc4e60f),
	.w4(32'h3b9bc519),
	.w5(32'hbb740eb6),
	.w6(32'h3a1c06fe),
	.w7(32'h3c1b5764),
	.w8(32'h3903dc4c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09403c),
	.w1(32'hbb697d03),
	.w2(32'h3b3884ba),
	.w3(32'hbbb96ac7),
	.w4(32'hbb322ab6),
	.w5(32'h3b4d3c29),
	.w6(32'h3b8b4328),
	.w7(32'h3bd1bfdd),
	.w8(32'h3baf5ab1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf21978),
	.w1(32'h3af74a2e),
	.w2(32'hbc06fd27),
	.w3(32'h394bfb06),
	.w4(32'h3b04fa05),
	.w5(32'hbadd430b),
	.w6(32'h3bd7f3e4),
	.w7(32'h3bacf3fb),
	.w8(32'hbbf3f41e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfd07c),
	.w1(32'hbac9093b),
	.w2(32'hbc10c002),
	.w3(32'hbb3e02ea),
	.w4(32'h3b2714a5),
	.w5(32'h3b5943f1),
	.w6(32'hb9d10507),
	.w7(32'h3ab3c200),
	.w8(32'h3b994afa),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc113fed),
	.w1(32'h3b920a5f),
	.w2(32'hbc5a2d04),
	.w3(32'hbc83918f),
	.w4(32'h3d4953e0),
	.w5(32'h3ace4ab9),
	.w6(32'hbb951891),
	.w7(32'h3bf38e0c),
	.w8(32'hb8aa5b1d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49c4e7),
	.w1(32'hbc0bba57),
	.w2(32'h3b3d73fd),
	.w3(32'hbc0f2a65),
	.w4(32'h3bb20b44),
	.w5(32'hbc4f1570),
	.w6(32'hbc3cdf84),
	.w7(32'hbb9ff019),
	.w8(32'hb98f4fd1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb25f92),
	.w1(32'hbb01f07f),
	.w2(32'h3949db5f),
	.w3(32'h39fc9832),
	.w4(32'h3b27cfe8),
	.w5(32'h39b03539),
	.w6(32'hbb1ff0d4),
	.w7(32'hbb8330a7),
	.w8(32'h3cca7c32),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37af0c14),
	.w1(32'hbb9166ec),
	.w2(32'h3c0381eb),
	.w3(32'h3d4e32c3),
	.w4(32'hbaf9cb94),
	.w5(32'h39ba3b07),
	.w6(32'hb880210a),
	.w7(32'hbc4c5df2),
	.w8(32'hbb83177f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b0fc4),
	.w1(32'hbb2e10da),
	.w2(32'hbc02a166),
	.w3(32'hbb164b1b),
	.w4(32'h3ba02b6d),
	.w5(32'h3cd010b3),
	.w6(32'h3b42f45c),
	.w7(32'h3a0c87f0),
	.w8(32'hbdb67047),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7d293),
	.w1(32'h3b4d2550),
	.w2(32'hbbfbcb16),
	.w3(32'h3b994f7d),
	.w4(32'h3c18f38a),
	.w5(32'hba408c25),
	.w6(32'hb963faf3),
	.w7(32'h3b0db410),
	.w8(32'hbbd709e9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc351e),
	.w1(32'hbb357543),
	.w2(32'hbc80e969),
	.w3(32'hbc14d309),
	.w4(32'hbb885917),
	.w5(32'hbba34a19),
	.w6(32'h3c2325f6),
	.w7(32'hbb448a28),
	.w8(32'hbc375254),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a40f7),
	.w1(32'h3c0aa2c3),
	.w2(32'hbbbe9704),
	.w3(32'hbbba7aca),
	.w4(32'h39ef7d18),
	.w5(32'h3af5f5f0),
	.w6(32'h3b567867),
	.w7(32'h3b82c2b5),
	.w8(32'hbae6325e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8baf97),
	.w1(32'h3b3b93cb),
	.w2(32'hbc1a1f77),
	.w3(32'hbb7789ae),
	.w4(32'h3a2cb2d9),
	.w5(32'hbc46303e),
	.w6(32'hbabe3946),
	.w7(32'h3c19d975),
	.w8(32'hbbb8cd6f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfcceb9),
	.w1(32'hbbb806af),
	.w2(32'hbc34397c),
	.w3(32'hbbbb661a),
	.w4(32'hbb6cd4c1),
	.w5(32'hbbf4644c),
	.w6(32'h3af80522),
	.w7(32'h3afeb9db),
	.w8(32'hbb7c9fd4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba091d93),
	.w1(32'hbbccd0f3),
	.w2(32'hbb64c571),
	.w3(32'hbc0d942b),
	.w4(32'hbc4ef055),
	.w5(32'hbc48932b),
	.w6(32'hbc1f4670),
	.w7(32'hbcba074b),
	.w8(32'hbafe4cbd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdefdda),
	.w1(32'hba7ecc63),
	.w2(32'hbba4558f),
	.w3(32'hbbeb8a5a),
	.w4(32'hbbd932d9),
	.w5(32'hbc1174a3),
	.w6(32'h3ba23fd6),
	.w7(32'hb9f7ce1d),
	.w8(32'hbb8f77b2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6f08d),
	.w1(32'hba6a0ebc),
	.w2(32'hbb2ffc11),
	.w3(32'h3c0b8baf),
	.w4(32'hbc75717c),
	.w5(32'h3ab54f1c),
	.w6(32'h3a2690b8),
	.w7(32'h3a561a4b),
	.w8(32'hb7d65860),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ab4ff),
	.w1(32'h3b34ab23),
	.w2(32'hbaf4c490),
	.w3(32'h3ad46f8d),
	.w4(32'h3a8e369a),
	.w5(32'hb8213a5a),
	.w6(32'h3b378ed6),
	.w7(32'h3acebe76),
	.w8(32'hbb303152),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d3952),
	.w1(32'hb91e550f),
	.w2(32'h3bb72462),
	.w3(32'hbce03dfd),
	.w4(32'h3a628ec1),
	.w5(32'hbb6d709a),
	.w6(32'h3c231e35),
	.w7(32'h3a991f1a),
	.w8(32'h3ae217d9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace8d37),
	.w1(32'h3c4da67c),
	.w2(32'hbbbdd548),
	.w3(32'h3afb0c6e),
	.w4(32'hbc23c87f),
	.w5(32'h3ba13296),
	.w6(32'hbb416bd3),
	.w7(32'hbac9a743),
	.w8(32'h3b90bb39),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03051d),
	.w1(32'h3a424494),
	.w2(32'h3a16cf54),
	.w3(32'hbc161cb9),
	.w4(32'hbc32a693),
	.w5(32'hbc14db51),
	.w6(32'hbc0130b9),
	.w7(32'h3a1e06cb),
	.w8(32'hbc49d9ef),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26f36d),
	.w1(32'h3997f8db),
	.w2(32'hbafd1489),
	.w3(32'h3c3c1134),
	.w4(32'hbc826efd),
	.w5(32'hb7e85403),
	.w6(32'hb9fbe5f1),
	.w7(32'h3bd66f6b),
	.w8(32'h3be9dee7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ccbe7),
	.w1(32'hbb6695d4),
	.w2(32'hbaba1a5b),
	.w3(32'h3a2a7d73),
	.w4(32'h3b2f9f3e),
	.w5(32'hbba009f2),
	.w6(32'h3b74e73b),
	.w7(32'h3ac56e85),
	.w8(32'hbbcff576),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91924f),
	.w1(32'hba9428ea),
	.w2(32'h3a77c343),
	.w3(32'h39fb4416),
	.w4(32'hbac24c63),
	.w5(32'h3b37f5b5),
	.w6(32'h39a9f2e6),
	.w7(32'hbb882035),
	.w8(32'hba763760),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cb202),
	.w1(32'h3ba3074b),
	.w2(32'hbb020d8e),
	.w3(32'h3b28fbeb),
	.w4(32'hbb5bd5d5),
	.w5(32'hb9a13b35),
	.w6(32'hbab9bc17),
	.w7(32'hbb41436a),
	.w8(32'h3c042e9f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9dfa3),
	.w1(32'hba7e3582),
	.w2(32'hbb4ac5b8),
	.w3(32'h3a14e875),
	.w4(32'h3bbb781a),
	.w5(32'h38da2ab3),
	.w6(32'hbb239b79),
	.w7(32'h3b07bfe2),
	.w8(32'hba8a57db),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca4d3c),
	.w1(32'h3ba11695),
	.w2(32'hb90168c0),
	.w3(32'hbbdbc4df),
	.w4(32'h3b0e6008),
	.w5(32'hba53ee30),
	.w6(32'hbaf95149),
	.w7(32'h3b8dddca),
	.w8(32'h3b2dab08),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8438f),
	.w1(32'h399e4de1),
	.w2(32'hbb4b301c),
	.w3(32'h3b83cd6d),
	.w4(32'h3a60d2d0),
	.w5(32'h37db3672),
	.w6(32'h3bc342a0),
	.w7(32'h39af72ba),
	.w8(32'h3a9e6150),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad352c),
	.w1(32'hbb8aca66),
	.w2(32'hbae08461),
	.w3(32'h3aff0581),
	.w4(32'hbb3cb69a),
	.w5(32'hb9986018),
	.w6(32'hbb3bb574),
	.w7(32'h38c14069),
	.w8(32'hbaea1a8c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55619b),
	.w1(32'h3b1614ce),
	.w2(32'hb9687e12),
	.w3(32'h3b26ee40),
	.w4(32'hbb019bad),
	.w5(32'hba0d7369),
	.w6(32'hbad84481),
	.w7(32'hbb93de8d),
	.w8(32'h3a140909),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f5c89),
	.w1(32'hbc1217a1),
	.w2(32'h3d0227ae),
	.w3(32'hba2d12db),
	.w4(32'hbb8f8f81),
	.w5(32'h3ae36760),
	.w6(32'hbb5d17aa),
	.w7(32'hb975076b),
	.w8(32'hbbbdd2da),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d6530),
	.w1(32'h3a725054),
	.w2(32'h398a0cac),
	.w3(32'h3a0537d8),
	.w4(32'h3aa03c78),
	.w5(32'h3af645be),
	.w6(32'hba4f8775),
	.w7(32'hbb02a410),
	.w8(32'hbb161e93),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96f95e),
	.w1(32'hbb1f7818),
	.w2(32'h3a1c8dc4),
	.w3(32'hba7af95b),
	.w4(32'hba8efea7),
	.w5(32'h38c207fc),
	.w6(32'h3c90c439),
	.w7(32'h3c0831ae),
	.w8(32'h3bfa178a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05eadc),
	.w1(32'hb9392ffd),
	.w2(32'hba45fd61),
	.w3(32'hbaec662a),
	.w4(32'hbc7292f7),
	.w5(32'h3b58bb97),
	.w6(32'hbb25be8a),
	.w7(32'hb9262df4),
	.w8(32'h3b7902ae),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe82084),
	.w1(32'hbbd420a1),
	.w2(32'hbc04d5ed),
	.w3(32'hbb177960),
	.w4(32'h3b719f72),
	.w5(32'hbb53c160),
	.w6(32'hb96c4470),
	.w7(32'h3b8cf953),
	.w8(32'hbb59c58a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1df1a),
	.w1(32'h3a76d657),
	.w2(32'hbb348836),
	.w3(32'hbb784445),
	.w4(32'h3b8947e8),
	.w5(32'h3b804647),
	.w6(32'hbaa1ab7d),
	.w7(32'h3c64e0e3),
	.w8(32'h3b510781),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc056bff),
	.w1(32'hba7c941d),
	.w2(32'hbba009cb),
	.w3(32'h39e6e174),
	.w4(32'h3b61d0bc),
	.w5(32'hbbb13e19),
	.w6(32'hb9f4f781),
	.w7(32'h3be6e638),
	.w8(32'h3ba6f218),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c74e8),
	.w1(32'hbbe9710a),
	.w2(32'hbad97a6d),
	.w3(32'h3af8a21d),
	.w4(32'hbb2d58ae),
	.w5(32'hbb841267),
	.w6(32'hbb93f23d),
	.w7(32'h3ba3d94e),
	.w8(32'hbba44da9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a272a61),
	.w1(32'h3b28399a),
	.w2(32'h39a933bb),
	.w3(32'h3b02e360),
	.w4(32'hba9285b1),
	.w5(32'h3b655010),
	.w6(32'hbb7c45e8),
	.w7(32'hbb637327),
	.w8(32'h3b2b4e31),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce3b500),
	.w1(32'hba0c11f9),
	.w2(32'h3b323ca2),
	.w3(32'h3ba630c2),
	.w4(32'h39bb1fdb),
	.w5(32'h3c8666f8),
	.w6(32'h389a5f9d),
	.w7(32'hbaa2c5ff),
	.w8(32'h39ed977c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4c00a),
	.w1(32'hb8ccdfe9),
	.w2(32'hbc65e439),
	.w3(32'hb8c6dd3b),
	.w4(32'h3a70bddf),
	.w5(32'h3ab74eac),
	.w6(32'h3bd7f168),
	.w7(32'h3b09c92f),
	.w8(32'hbb8ca5e5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb250c41),
	.w1(32'h3962db85),
	.w2(32'h3a1c23cb),
	.w3(32'hbb303d51),
	.w4(32'h3c14d3f0),
	.w5(32'hba34f957),
	.w6(32'hbb921725),
	.w7(32'hba08ad0d),
	.w8(32'h3b0ca981),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a311dc9),
	.w1(32'hbb2d6808),
	.w2(32'hbac8a04c),
	.w3(32'hbba603c9),
	.w4(32'hbbb2c097),
	.w5(32'h39205318),
	.w6(32'h3b1dfa3c),
	.w7(32'h3b82916a),
	.w8(32'h3b678439),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06fba7),
	.w1(32'hbb82816d),
	.w2(32'hbbb62309),
	.w3(32'h3acb024c),
	.w4(32'h3a03b813),
	.w5(32'hba2851a8),
	.w6(32'h3adb16eb),
	.w7(32'h388fa721),
	.w8(32'hbb34606b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c773d),
	.w1(32'hbbc1c8e8),
	.w2(32'hbb07506d),
	.w3(32'h3c055fc5),
	.w4(32'hbbf8adf3),
	.w5(32'hbc089723),
	.w6(32'hbbea998a),
	.w7(32'hbc521077),
	.w8(32'hbc7a0b4e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0f4bf),
	.w1(32'hba9325b9),
	.w2(32'hbb113112),
	.w3(32'h3aa69ff9),
	.w4(32'h39c94535),
	.w5(32'hbbaf5fb5),
	.w6(32'h3a180275),
	.w7(32'hb9e45d31),
	.w8(32'hbb340ae8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41811c),
	.w1(32'hb9ede3a9),
	.w2(32'hbc3b86d0),
	.w3(32'hbb0b32ca),
	.w4(32'hb92c7a7e),
	.w5(32'hbb82b1db),
	.w6(32'hba327399),
	.w7(32'h3a0db610),
	.w8(32'hbaa8ae0d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b6f25),
	.w1(32'hbb47ecab),
	.w2(32'hbbaa48b9),
	.w3(32'hbb0035c2),
	.w4(32'h3a4bbd47),
	.w5(32'hbb26671f),
	.w6(32'hbb825654),
	.w7(32'h3b7fc594),
	.w8(32'h3a9cc805),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24e8f2),
	.w1(32'h37f22cce),
	.w2(32'hbacafeaf),
	.w3(32'hbb606d74),
	.w4(32'hbba4c004),
	.w5(32'hbb1de55e),
	.w6(32'hbb13c4d4),
	.w7(32'hba3cd0b4),
	.w8(32'hbb12d6ac),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b790897),
	.w1(32'hbbd2514b),
	.w2(32'hb9894be2),
	.w3(32'hbbf99076),
	.w4(32'hbaafcfbb),
	.w5(32'hbace29f3),
	.w6(32'h3a94ba05),
	.w7(32'hba7ce529),
	.w8(32'hbb31aac0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3abad6),
	.w1(32'hbb051f2c),
	.w2(32'h3ad301c5),
	.w3(32'hbbb92a54),
	.w4(32'h3a1dea17),
	.w5(32'h3c32f2e8),
	.w6(32'h3b0630bd),
	.w7(32'hbbb0ebd4),
	.w8(32'h3b8bcb6b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c3739),
	.w1(32'h3ba1f5e5),
	.w2(32'h3c505e4f),
	.w3(32'hba7cf91c),
	.w4(32'hbbb0a2c7),
	.w5(32'h3ad28b1a),
	.w6(32'h3c88c2e3),
	.w7(32'hbba502f4),
	.w8(32'hbb0554ac),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a8af3),
	.w1(32'hbb1ad1ba),
	.w2(32'h3b32efc1),
	.w3(32'hbb8b17d9),
	.w4(32'hbb5e90b7),
	.w5(32'hba870879),
	.w6(32'hbaf0ff34),
	.w7(32'hbb6f0a6f),
	.w8(32'h3bb4861b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18de8a),
	.w1(32'h3b33a9b5),
	.w2(32'h3a82a99e),
	.w3(32'h3b1cce6f),
	.w4(32'h3bd8083e),
	.w5(32'hbacb706b),
	.w6(32'hbb2ff1d7),
	.w7(32'hbb25b9e9),
	.w8(32'h3c1f9b2f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad19fb7),
	.w1(32'hbbd7ae15),
	.w2(32'hbb2429c5),
	.w3(32'hba046050),
	.w4(32'h3c3e241c),
	.w5(32'hbc824a6c),
	.w6(32'h3bcbbe41),
	.w7(32'h3c404cbc),
	.w8(32'h3b9d13e3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16bac0),
	.w1(32'hba061405),
	.w2(32'hba22a7c1),
	.w3(32'hbaef0772),
	.w4(32'hbbb507b9),
	.w5(32'hbab749fa),
	.w6(32'h3b93bb5f),
	.w7(32'h399015dd),
	.w8(32'h3b6072c9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f9333),
	.w1(32'hbad66748),
	.w2(32'h3c4a4697),
	.w3(32'hba5bcb74),
	.w4(32'hbc0ee03c),
	.w5(32'hbb615318),
	.w6(32'h3b5d33e4),
	.w7(32'h3812d615),
	.w8(32'h3ab36134),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabdf8d),
	.w1(32'h3b6ed5e0),
	.w2(32'hbc2d16cc),
	.w3(32'h3a98a783),
	.w4(32'h3a464d4b),
	.w5(32'hb9c79666),
	.w6(32'hbbb2a74b),
	.w7(32'hbc194bfe),
	.w8(32'hbb8a3cc5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae352dd),
	.w1(32'hb9c8a2ff),
	.w2(32'hbba6628c),
	.w3(32'hbbabfd67),
	.w4(32'h3ba6dcde),
	.w5(32'hbb73ca5e),
	.w6(32'hbbe73635),
	.w7(32'h3c3df458),
	.w8(32'h3c072aed),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2beff0),
	.w1(32'h3ca7bf1f),
	.w2(32'hbbf4d642),
	.w3(32'h3bc17a2c),
	.w4(32'h3c2b8211),
	.w5(32'hbbda57a7),
	.w6(32'h3c39b827),
	.w7(32'h39888630),
	.w8(32'h39f3caa2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85b599),
	.w1(32'hbaaf23d2),
	.w2(32'h3a41b5ea),
	.w3(32'hba75507f),
	.w4(32'h3c311908),
	.w5(32'hbb4fcf4c),
	.w6(32'h3c134285),
	.w7(32'h3b9b6368),
	.w8(32'h3adea27f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c860c84),
	.w1(32'hbbf5ce3d),
	.w2(32'hba6fab0b),
	.w3(32'hbb1db1b4),
	.w4(32'h3c0a3b8c),
	.w5(32'h3c437545),
	.w6(32'hb9afcd8b),
	.w7(32'hbb4190a5),
	.w8(32'h3b9dd31a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75c1f1),
	.w1(32'hbb2da45e),
	.w2(32'hbaf13c1f),
	.w3(32'hbc1ec11d),
	.w4(32'h39c8265a),
	.w5(32'h3ace9ac8),
	.w6(32'h39f423d4),
	.w7(32'hbb82fb95),
	.w8(32'h3a67295f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6348a),
	.w1(32'hbb95da59),
	.w2(32'h3bcbc4bd),
	.w3(32'hbba84b1b),
	.w4(32'hbc2f3229),
	.w5(32'h3b1af7d4),
	.w6(32'h3b46488d),
	.w7(32'h3a823608),
	.w8(32'h38ad62e3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31712c),
	.w1(32'h3ad4875e),
	.w2(32'hbbedc88a),
	.w3(32'h385b3455),
	.w4(32'hba17eed4),
	.w5(32'hbbc52c43),
	.w6(32'hbb9fc099),
	.w7(32'h3c113db7),
	.w8(32'hbc3308ac),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd2a91),
	.w1(32'hba6a3db2),
	.w2(32'hba4c756b),
	.w3(32'h3b461387),
	.w4(32'hbb8ea106),
	.w5(32'h3be2d813),
	.w6(32'hbb0445d7),
	.w7(32'h3c3eccf4),
	.w8(32'h3a2c7545),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84519f),
	.w1(32'hbbcbc78f),
	.w2(32'h3c3091eb),
	.w3(32'hbbe68420),
	.w4(32'hbbbe9408),
	.w5(32'hbbd29b41),
	.w6(32'hbba3009b),
	.w7(32'hbc99b457),
	.w8(32'hbbdbfbaf),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c9502),
	.w1(32'h3b4a6671),
	.w2(32'hbb74f875),
	.w3(32'hbb40651f),
	.w4(32'h3c49e256),
	.w5(32'h37199536),
	.w6(32'hbb2aed8c),
	.w7(32'h3cdb7481),
	.w8(32'h3c64e25f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04f3b4),
	.w1(32'hbb881cf0),
	.w2(32'h3b4cec88),
	.w3(32'h3b5391ea),
	.w4(32'hba462757),
	.w5(32'hbbb9aa00),
	.w6(32'hbc1218db),
	.w7(32'h3bcd8b70),
	.w8(32'hbc0f2b1f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e9b4f),
	.w1(32'hbb3c517a),
	.w2(32'h3ba2d5f9),
	.w3(32'hbbf62602),
	.w4(32'h3b70dc36),
	.w5(32'hbbec6b37),
	.w6(32'hbb53e971),
	.w7(32'hbb4c97ef),
	.w8(32'hbc6b022f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87792d),
	.w1(32'h3bef0f73),
	.w2(32'h3b93325c),
	.w3(32'h3885c1e6),
	.w4(32'hbafc3cbd),
	.w5(32'h3c5e5db3),
	.w6(32'hbab1a109),
	.w7(32'hbba90c2f),
	.w8(32'hbbc76c89),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16360a),
	.w1(32'hbaad8d78),
	.w2(32'h3ca1f1fa),
	.w3(32'hbc175a1d),
	.w4(32'hbb8803d2),
	.w5(32'h3c357ab6),
	.w6(32'hbb670479),
	.w7(32'hbc15c19b),
	.w8(32'hbc26ac6f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfe0b3),
	.w1(32'hbc007195),
	.w2(32'hbbb33615),
	.w3(32'hbc244516),
	.w4(32'hbbd03181),
	.w5(32'hbc4ef140),
	.w6(32'h3bb0a86c),
	.w7(32'hbb4a4119),
	.w8(32'hbb5c4604),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43386),
	.w1(32'hb948a44f),
	.w2(32'h3be4442f),
	.w3(32'hbb237a2e),
	.w4(32'hbae343c9),
	.w5(32'h3b96242a),
	.w6(32'hbb9929d3),
	.w7(32'hbada10a4),
	.w8(32'hb822b403),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b2a17),
	.w1(32'hb9ee7320),
	.w2(32'hba416557),
	.w3(32'hbbae461f),
	.w4(32'hba19d7e0),
	.w5(32'hbaf3fdb0),
	.w6(32'hbaf8e3fb),
	.w7(32'h3bb65ea4),
	.w8(32'h3a6084b7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bbb0d),
	.w1(32'h3baaef72),
	.w2(32'hbbeba373),
	.w3(32'hb9d5ec4a),
	.w4(32'hbb8a81ed),
	.w5(32'hbbbd7939),
	.w6(32'hbc3ca4da),
	.w7(32'hbc4a80e2),
	.w8(32'hbb9fc743),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba6eb8),
	.w1(32'hbbbe3f4d),
	.w2(32'h3a8f55be),
	.w3(32'hbb7f9367),
	.w4(32'h39ddeb9f),
	.w5(32'h3aa31ea0),
	.w6(32'h3a9f8bae),
	.w7(32'h3ab45409),
	.w8(32'hbbe24dad),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97205c),
	.w1(32'hbbbdb342),
	.w2(32'h3bbcdcc9),
	.w3(32'hbb57f94e),
	.w4(32'h3ac1842f),
	.w5(32'h3c124716),
	.w6(32'hbc21f1b5),
	.w7(32'h3b2cfbf2),
	.w8(32'h3aaa6b3d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99bab8),
	.w1(32'h3c63910a),
	.w2(32'hba898248),
	.w3(32'hbb96f2f5),
	.w4(32'h3b62c45b),
	.w5(32'h3b34a1b4),
	.w6(32'hbb8ab22a),
	.w7(32'hbbc2e9e2),
	.w8(32'h3a95c6ce),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12c717),
	.w1(32'h3a0cb0f0),
	.w2(32'hbb81a682),
	.w3(32'hba55ad02),
	.w4(32'h3b599e29),
	.w5(32'h3b14dbc7),
	.w6(32'hb9f00913),
	.w7(32'h3b094fae),
	.w8(32'h3cf6595f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a0799),
	.w1(32'h3acc68b5),
	.w2(32'hbb82a56f),
	.w3(32'hbd2469b6),
	.w4(32'hba32d5f2),
	.w5(32'h3a997168),
	.w6(32'hbb81250d),
	.w7(32'h39a6e63d),
	.w8(32'hbbb570d1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2ca8b0),
	.w1(32'hbb02f1fe),
	.w2(32'hbb4efd05),
	.w3(32'hbab0c110),
	.w4(32'hba83dc48),
	.w5(32'h3d395de4),
	.w6(32'h3b5ee786),
	.w7(32'hba2b2e8e),
	.w8(32'hbbf194c5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ac8b2),
	.w1(32'hba0830d5),
	.w2(32'hbb9a82a7),
	.w3(32'h3b1012c5),
	.w4(32'hbb50d321),
	.w5(32'hbb92311d),
	.w6(32'hbc249afe),
	.w7(32'h3ba99a37),
	.w8(32'h3a154ed7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f8f6d),
	.w1(32'h3b347276),
	.w2(32'h3b66cccb),
	.w3(32'hb9e20ee9),
	.w4(32'h3b551341),
	.w5(32'h3b821a86),
	.w6(32'h3c7f3f81),
	.w7(32'hba69be3f),
	.w8(32'h3b0514b6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb225981),
	.w1(32'h3a39ead9),
	.w2(32'hba8aee89),
	.w3(32'h3a535af4),
	.w4(32'hbadffa0b),
	.w5(32'h3b15d684),
	.w6(32'h3b2cfebf),
	.w7(32'h3b1e5e29),
	.w8(32'hbbeb8f48),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb526fe7),
	.w1(32'hbb2f97f7),
	.w2(32'hbc3fe96b),
	.w3(32'hbb28f027),
	.w4(32'h3b2d0bfa),
	.w5(32'hbbd671ec),
	.w6(32'hbaa72f34),
	.w7(32'h391691ee),
	.w8(32'hb96f36b6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc405fb8),
	.w1(32'hba69b272),
	.w2(32'hbb81f171),
	.w3(32'hbaec24b3),
	.w4(32'hba8a806c),
	.w5(32'hbae9ff27),
	.w6(32'h3b65f470),
	.w7(32'h3bb71e6a),
	.w8(32'hbb2b48fd),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57328a),
	.w1(32'hbbc61397),
	.w2(32'hbc54263d),
	.w3(32'h3b7c16bc),
	.w4(32'hbb6c7407),
	.w5(32'hbbbde8de),
	.w6(32'hbc046e61),
	.w7(32'hbcd16ef0),
	.w8(32'h3a9f7aa3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd0476),
	.w1(32'h3a2fb78f),
	.w2(32'h3a9b32da),
	.w3(32'hbb4c68d2),
	.w4(32'h3b99d109),
	.w5(32'h3c406b5e),
	.w6(32'hbbe8d1c9),
	.w7(32'hbb32b116),
	.w8(32'h3b263c62),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc798b),
	.w1(32'hbb4e79f6),
	.w2(32'hbb41f1d7),
	.w3(32'hbd067672),
	.w4(32'h3b3744c3),
	.w5(32'h3a0595ce),
	.w6(32'h3b99b089),
	.w7(32'h397559f7),
	.w8(32'h3a891a97),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11e1c1),
	.w1(32'h3cee7324),
	.w2(32'h3b9cb019),
	.w3(32'h38d445bf),
	.w4(32'h3b82df1d),
	.w5(32'h3aaa8f4f),
	.w6(32'hbbbf1315),
	.w7(32'h3bfdb910),
	.w8(32'h39b11d8b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5f7b6),
	.w1(32'h3a2f2fca),
	.w2(32'hbb88ec82),
	.w3(32'hbab4c671),
	.w4(32'h3a8b2227),
	.w5(32'h3d0963dd),
	.w6(32'hbc883966),
	.w7(32'h3d27424e),
	.w8(32'hba7d40d8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b016d89),
	.w1(32'h37822f13),
	.w2(32'h3b9235e9),
	.w3(32'h3b8661be),
	.w4(32'h3b3c1dea),
	.w5(32'hbadac3a2),
	.w6(32'hbad231dc),
	.w7(32'h38bb2903),
	.w8(32'hb8da5fd8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb890924),
	.w1(32'h3c32a4af),
	.w2(32'hbaf7f090),
	.w3(32'hbb630dd7),
	.w4(32'h3b3998a6),
	.w5(32'hbd174d0f),
	.w6(32'hbaac6634),
	.w7(32'h3a6726c3),
	.w8(32'hba847822),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddcf75),
	.w1(32'hbcf97c4b),
	.w2(32'hbb7062be),
	.w3(32'hbbbbbfd1),
	.w4(32'hbb6a784d),
	.w5(32'h3a02a83d),
	.w6(32'hbbd6e536),
	.w7(32'hba7fd24e),
	.w8(32'hba20d60f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace7e74),
	.w1(32'hba380762),
	.w2(32'hbc242559),
	.w3(32'h3b712403),
	.w4(32'h3b358d2c),
	.w5(32'hbaacd6ac),
	.w6(32'h3b7b3b6a),
	.w7(32'hbb2cb504),
	.w8(32'hbcf1f3d3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1073a),
	.w1(32'h3af0925d),
	.w2(32'hbce1d622),
	.w3(32'hbaf5a7b5),
	.w4(32'hbbb06069),
	.w5(32'h3a86a166),
	.w6(32'h396486ae),
	.w7(32'h3b0dcf27),
	.w8(32'h3ac4c289),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0eb3),
	.w1(32'h3b68aa49),
	.w2(32'hbb865208),
	.w3(32'hbcb31f15),
	.w4(32'hbb8c52ae),
	.w5(32'hba5d8f75),
	.w6(32'hba1fbb84),
	.w7(32'h3c99e666),
	.w8(32'hbb56fd39),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a781f71),
	.w1(32'hbbee9390),
	.w2(32'hbb8eaeeb),
	.w3(32'h3d13ebc7),
	.w4(32'h3ccfc61e),
	.w5(32'hba360345),
	.w6(32'h39d08842),
	.w7(32'hba708896),
	.w8(32'hbbba43bc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78cf07),
	.w1(32'h3b375ddf),
	.w2(32'h3b501e69),
	.w3(32'h3caf8f22),
	.w4(32'hbad224fb),
	.w5(32'h3cda1ed5),
	.w6(32'hbad17966),
	.w7(32'h3b9b15cd),
	.w8(32'hbb935b5f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48fa48),
	.w1(32'hbace56b5),
	.w2(32'hbbea177a),
	.w3(32'h3b873b05),
	.w4(32'hbaaeac53),
	.w5(32'h3be30d6f),
	.w6(32'hbb8978b5),
	.w7(32'h3bba6438),
	.w8(32'h3b9352a0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc6bf6),
	.w1(32'hbb8ae118),
	.w2(32'h3a539c6e),
	.w3(32'hbb5243b6),
	.w4(32'hbbe30b9b),
	.w5(32'h3c39319b),
	.w6(32'hbb053bec),
	.w7(32'hbb8d834a),
	.w8(32'hbb5a2f6a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf34a4a),
	.w1(32'h3a3256ac),
	.w2(32'hbb800853),
	.w3(32'h3bbb360f),
	.w4(32'h3a9d947a),
	.w5(32'hb99fe3ce),
	.w6(32'h3b33d4ca),
	.w7(32'h3aad032e),
	.w8(32'h39653ce8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c3bae),
	.w1(32'h3a536fdc),
	.w2(32'hbbac5bf5),
	.w3(32'hbb1c6300),
	.w4(32'h3c0a4166),
	.w5(32'hbad251d1),
	.w6(32'hbb31e65a),
	.w7(32'h3c189f93),
	.w8(32'hbba572d2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb856aeb),
	.w1(32'h3b9f3a41),
	.w2(32'hba9fa626),
	.w3(32'hbc290e39),
	.w4(32'hbb4c2bef),
	.w5(32'hbaa3eebf),
	.w6(32'hbae1fbd6),
	.w7(32'h3aa51f9c),
	.w8(32'hbb50c042),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h353362ae),
	.w1(32'h3b646b3d),
	.w2(32'hbb86ee2b),
	.w3(32'hbb99d234),
	.w4(32'h3b97ab06),
	.w5(32'h3c07c32c),
	.w6(32'h3ba87a5a),
	.w7(32'h3990d493),
	.w8(32'hbb97fee6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5c574),
	.w1(32'hbb0246d5),
	.w2(32'hbbb218ab),
	.w3(32'hbb993411),
	.w4(32'hba816de7),
	.w5(32'hbc0f5b0e),
	.w6(32'hba950c48),
	.w7(32'h3bda84db),
	.w8(32'h3a778073),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28fcd1),
	.w1(32'h3a7f74c4),
	.w2(32'hbb37df8a),
	.w3(32'hbb8147f7),
	.w4(32'h38c06a01),
	.w5(32'hb9e25229),
	.w6(32'h3b24877b),
	.w7(32'h3a4a221b),
	.w8(32'h3a5c0b70),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba619338),
	.w1(32'h3bf92c4f),
	.w2(32'hbbb2928c),
	.w3(32'hbb58ccec),
	.w4(32'h3a73799c),
	.w5(32'hbbfec0f5),
	.w6(32'hbc0ae2bd),
	.w7(32'hbb8fcaf0),
	.w8(32'hbb896317),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eb775),
	.w1(32'hbb825958),
	.w2(32'hba2c621d),
	.w3(32'hbb983a53),
	.w4(32'h3c641308),
	.w5(32'hba609557),
	.w6(32'hbb7fac03),
	.w7(32'h3b0027c2),
	.w8(32'h3b0005fc),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cfad0),
	.w1(32'h3b9bbf02),
	.w2(32'h3a555995),
	.w3(32'h3b7f5a9c),
	.w4(32'h3ad01040),
	.w5(32'hb8bc8f8c),
	.w6(32'h3c764689),
	.w7(32'h393383d3),
	.w8(32'hba09c665),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f4ae0),
	.w1(32'hba3101c1),
	.w2(32'h3bc0886b),
	.w3(32'h39bdd157),
	.w4(32'hbb883d25),
	.w5(32'h3b80d432),
	.w6(32'h3a5d0f76),
	.w7(32'hbb880d3d),
	.w8(32'h3b3407a2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8085ec),
	.w1(32'hbb3edb09),
	.w2(32'h3b465b06),
	.w3(32'h3a6b9dac),
	.w4(32'hb985a8b7),
	.w5(32'hb99e0388),
	.w6(32'h3b599b73),
	.w7(32'h3b1c8113),
	.w8(32'hbacf6872),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb263d37),
	.w1(32'hbb5d26d2),
	.w2(32'hbbc2c427),
	.w3(32'h3a3ad39b),
	.w4(32'h3a5bbd66),
	.w5(32'hbb37b426),
	.w6(32'hba7e3794),
	.w7(32'h3a07b2fc),
	.w8(32'hbaa99bf3),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd3781),
	.w1(32'h3a887c9f),
	.w2(32'h3afb0793),
	.w3(32'hbbd09e54),
	.w4(32'hbaecbd85),
	.w5(32'h3a886666),
	.w6(32'hbc033ba1),
	.w7(32'hbbd445eb),
	.w8(32'hbbab21f1),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad64e5a),
	.w1(32'h3bb11455),
	.w2(32'h3be37d18),
	.w3(32'h3ad3ad4c),
	.w4(32'h3b510ca9),
	.w5(32'hba98d0bc),
	.w6(32'h39692013),
	.w7(32'hbab8b88b),
	.w8(32'h39a5ef2f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ef790),
	.w1(32'hbb2e0558),
	.w2(32'hbb8c2bc2),
	.w3(32'hba91be4a),
	.w4(32'hbae252b0),
	.w5(32'hbbc95106),
	.w6(32'h3b292197),
	.w7(32'h3b2d6459),
	.w8(32'h3acb27e6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38c5c8),
	.w1(32'hbaf0aaad),
	.w2(32'h39a252c9),
	.w3(32'hbb134a56),
	.w4(32'hbb1cacb2),
	.w5(32'h3b2481b5),
	.w6(32'h3bbff719),
	.w7(32'hbbffa58f),
	.w8(32'h3b971d32),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa92cc),
	.w1(32'h3ba730c1),
	.w2(32'hbb928bd2),
	.w3(32'hbb413140),
	.w4(32'h3ac41af5),
	.w5(32'h3a265881),
	.w6(32'hb98730b0),
	.w7(32'hbabdf051),
	.w8(32'hbae56419),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae4ff5),
	.w1(32'hbc09180a),
	.w2(32'hbbf45537),
	.w3(32'h3b687a03),
	.w4(32'h3a37a0e9),
	.w5(32'hbad329cb),
	.w6(32'h3b451b03),
	.w7(32'h3b07094c),
	.w8(32'hbafdaf99),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14e3e9),
	.w1(32'hba4744f7),
	.w2(32'h3ac66bdb),
	.w3(32'hbb5590bb),
	.w4(32'hba5cfcbb),
	.w5(32'h3a1a2210),
	.w6(32'h3c017f5d),
	.w7(32'h3b26588a),
	.w8(32'hbb016fd2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357e6e86),
	.w1(32'hba4772b3),
	.w2(32'h3b1c32f6),
	.w3(32'hbba0b228),
	.w4(32'hbb713776),
	.w5(32'h3a83224a),
	.w6(32'h3b0fa107),
	.w7(32'h392fbebb),
	.w8(32'h3b315257),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90830c6),
	.w1(32'h39a12e7a),
	.w2(32'hba416972),
	.w3(32'h3a578d85),
	.w4(32'h3bef6051),
	.w5(32'hbc5660c1),
	.w6(32'hbb7356b2),
	.w7(32'h3b362a09),
	.w8(32'h3b6fb932),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f413a),
	.w1(32'hb99f73a1),
	.w2(32'h3bcea98d),
	.w3(32'hbb60456c),
	.w4(32'h3bca9700),
	.w5(32'h3bfc5bc0),
	.w6(32'hbb0fccd2),
	.w7(32'h3b3ac12c),
	.w8(32'h3a5e3e6b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b67a0),
	.w1(32'hbb4dae8f),
	.w2(32'hbaf5267f),
	.w3(32'hbaec7eca),
	.w4(32'h3b8cbe89),
	.w5(32'hba1dc202),
	.w6(32'hb983efaf),
	.w7(32'h3ab5fc50),
	.w8(32'h39e21eff),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3b6d8),
	.w1(32'hba855936),
	.w2(32'hb9b15e16),
	.w3(32'hbc2198dd),
	.w4(32'h3b635b10),
	.w5(32'h38036944),
	.w6(32'h3adf25c5),
	.w7(32'hbb88f5f5),
	.w8(32'h3b28ced5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dda4a),
	.w1(32'h3a942d8a),
	.w2(32'h3b21d74e),
	.w3(32'hba75ea74),
	.w4(32'hbb816c6e),
	.w5(32'h3bc90978),
	.w6(32'hbb89e566),
	.w7(32'h3ca34fce),
	.w8(32'h3c8b3543),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47a2a2),
	.w1(32'h3a553a2e),
	.w2(32'h3a805ccd),
	.w3(32'hb9e0470a),
	.w4(32'hbb125c56),
	.w5(32'h3b366178),
	.w6(32'hbb02ba50),
	.w7(32'h3c4c6b77),
	.w8(32'h3a91b23c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2479ed),
	.w1(32'h3a8810c2),
	.w2(32'h3b66db29),
	.w3(32'h3b0ef913),
	.w4(32'hb9c91f05),
	.w5(32'hbaf9871b),
	.w6(32'h3c713bbf),
	.w7(32'hba7fb58a),
	.w8(32'hbad433e9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b25ff),
	.w1(32'h3b3fc0de),
	.w2(32'hbb28628c),
	.w3(32'h3a33cd4d),
	.w4(32'h3993c7c6),
	.w5(32'hbb613aa0),
	.w6(32'h3bb299f7),
	.w7(32'h3bcc552b),
	.w8(32'hbb0c152b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fbeece),
	.w1(32'hb8d5e267),
	.w2(32'hb9634609),
	.w3(32'hba0be792),
	.w4(32'h3a0585a6),
	.w5(32'h390c3853),
	.w6(32'h3b6b48fc),
	.w7(32'h3b79afd6),
	.w8(32'h3a628365),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62c3a9),
	.w1(32'hba238e65),
	.w2(32'hbbc4314b),
	.w3(32'hbae4be0e),
	.w4(32'hbb4e711f),
	.w5(32'hbba79ee4),
	.w6(32'hba422554),
	.w7(32'hbae6926b),
	.w8(32'hbc140d04),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce3f39),
	.w1(32'hb9b1c901),
	.w2(32'h3b658862),
	.w3(32'h3a8e786c),
	.w4(32'hba683372),
	.w5(32'hba57c111),
	.w6(32'h3a54aef8),
	.w7(32'h3b0b5a91),
	.w8(32'hbac19557),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3b36a),
	.w1(32'h3b300938),
	.w2(32'h3a307700),
	.w3(32'hba056371),
	.w4(32'h397fa1c0),
	.w5(32'hbb734646),
	.w6(32'h3afe8996),
	.w7(32'hbb123c30),
	.w8(32'h3a8aeb9a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc3ae0),
	.w1(32'h3a70709e),
	.w2(32'hbb2520e3),
	.w3(32'h3c14a2b4),
	.w4(32'hbb272991),
	.w5(32'h3980e8d8),
	.w6(32'h3bb3ed1a),
	.w7(32'h3be9fdae),
	.w8(32'hbba509e9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b6bec),
	.w1(32'h39e4d192),
	.w2(32'hbbc7f5a3),
	.w3(32'h3b20020b),
	.w4(32'h3a0f2da2),
	.w5(32'hbba89d55),
	.w6(32'h3c0c47c4),
	.w7(32'h3b17ee85),
	.w8(32'hbb9d4bed),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91017a),
	.w1(32'h3b4b1059),
	.w2(32'hbba78fff),
	.w3(32'hbad7d5c5),
	.w4(32'hba8b68bf),
	.w5(32'hbc6ce6d5),
	.w6(32'hbacbb979),
	.w7(32'hb9f7db49),
	.w8(32'hbac745fa),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba328b),
	.w1(32'hbad2611d),
	.w2(32'hbb88d451),
	.w3(32'hbb58633b),
	.w4(32'h3af7b7b8),
	.w5(32'hbb81d0fd),
	.w6(32'h3aac4901),
	.w7(32'h3a14bd4e),
	.w8(32'hbb517474),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a4cd),
	.w1(32'hba2e2600),
	.w2(32'h3b9a1577),
	.w3(32'h39927e30),
	.w4(32'hb889b5f9),
	.w5(32'h39660672),
	.w6(32'hbb100360),
	.w7(32'hba8304c1),
	.w8(32'h391a5965),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca0726),
	.w1(32'h39b9ed38),
	.w2(32'h3b17f0f9),
	.w3(32'h3ba4184f),
	.w4(32'h3b4ec4f0),
	.w5(32'hb97f388e),
	.w6(32'h3b4d8a8a),
	.w7(32'h3b7799c4),
	.w8(32'hbbaf4f09),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6ee05),
	.w1(32'h3a013122),
	.w2(32'hb8ae29ef),
	.w3(32'h3b62659b),
	.w4(32'hba89d7b1),
	.w5(32'hbb6256f7),
	.w6(32'hbb245513),
	.w7(32'h3bdccad6),
	.w8(32'hbac5b78c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9d9c8),
	.w1(32'hbad48b37),
	.w2(32'hbb4b753a),
	.w3(32'h3a221962),
	.w4(32'hba749a92),
	.w5(32'h3b99a3d3),
	.w6(32'hba47cfc2),
	.w7(32'h3ad11fe1),
	.w8(32'h38c3cb70),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab914cb),
	.w1(32'hbaa962a2),
	.w2(32'hb8494aeb),
	.w3(32'hba8006c4),
	.w4(32'h39387da3),
	.w5(32'h3ab9152e),
	.w6(32'h3a48155a),
	.w7(32'h3c2e5201),
	.w8(32'hbaa6fdd4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dde72),
	.w1(32'hbb296721),
	.w2(32'h3ab2e6b7),
	.w3(32'h3aac83ef),
	.w4(32'hbb1e0eed),
	.w5(32'hbba7356f),
	.w6(32'h37d7a9ee),
	.w7(32'h3b356448),
	.w8(32'h3b895a4d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143e29),
	.w1(32'h3baa07bf),
	.w2(32'hbbc8fe76),
	.w3(32'hbbbf9cd5),
	.w4(32'h3cb65616),
	.w5(32'hba959bab),
	.w6(32'hbbaf8bf4),
	.w7(32'h3b00a369),
	.w8(32'hba94e658),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6fb8c),
	.w1(32'h390ce397),
	.w2(32'hbb28eb7e),
	.w3(32'h3af8c85b),
	.w4(32'h3938e09e),
	.w5(32'hbb17ce3d),
	.w6(32'hbb3b6e6a),
	.w7(32'hbb10fdca),
	.w8(32'hbb05c598),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c365af8),
	.w1(32'h3c22530b),
	.w2(32'h3b738849),
	.w3(32'h378014f9),
	.w4(32'hba01e84f),
	.w5(32'hbb3458de),
	.w6(32'h3b08e1eb),
	.w7(32'hb913b071),
	.w8(32'h3b9ea460),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09ebf7),
	.w1(32'hbbbe775a),
	.w2(32'h3aba92e1),
	.w3(32'hbb976cf5),
	.w4(32'hbb99dd00),
	.w5(32'hbbe42c20),
	.w6(32'hbc3ad290),
	.w7(32'hba9207ff),
	.w8(32'hbba47a44),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8857022),
	.w1(32'hba860d89),
	.w2(32'hbabae586),
	.w3(32'hbb4bf08f),
	.w4(32'hbbddb26a),
	.w5(32'hbaee4de9),
	.w6(32'h3a592438),
	.w7(32'hbb04eeb1),
	.w8(32'hba6aec85),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15d488),
	.w1(32'h3ba9cd3a),
	.w2(32'hba89419c),
	.w3(32'hba3cd108),
	.w4(32'h3882908a),
	.w5(32'h392e2b71),
	.w6(32'h372f9e25),
	.w7(32'hbb171fba),
	.w8(32'hbac19fd1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07327b),
	.w1(32'h3aa7ef3a),
	.w2(32'h3c144719),
	.w3(32'h3a391a6c),
	.w4(32'hbb8e8d22),
	.w5(32'hbb0188d6),
	.w6(32'hbac13033),
	.w7(32'hba0a8dcf),
	.w8(32'hbb8ee379),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb507702),
	.w1(32'h3b8720b9),
	.w2(32'hbb99b117),
	.w3(32'hbb893f8d),
	.w4(32'h3b91fb61),
	.w5(32'h38626649),
	.w6(32'hbabf227f),
	.w7(32'hbb0bbf67),
	.w8(32'h393d89d2),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d468b9),
	.w1(32'hbb654c97),
	.w2(32'hba9b0aed),
	.w3(32'h3a311abd),
	.w4(32'h3a0c903c),
	.w5(32'h3c8df039),
	.w6(32'hb9d7967f),
	.w7(32'h3b1afcff),
	.w8(32'h3b244f84),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c298a),
	.w1(32'h3b2f87ce),
	.w2(32'h3a863e35),
	.w3(32'h3aa2aef4),
	.w4(32'hba037f89),
	.w5(32'hbb18b937),
	.w6(32'h3a02a149),
	.w7(32'h3c877921),
	.w8(32'h3b09d7cc),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c896c3a),
	.w1(32'h3b880a4a),
	.w2(32'hb9d08fcc),
	.w3(32'h3c8b815e),
	.w4(32'h3abb0a1d),
	.w5(32'h3bce8e93),
	.w6(32'h3ca3b486),
	.w7(32'h3c9148f3),
	.w8(32'h3c31fb6c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9462cb),
	.w1(32'hba661f79),
	.w2(32'hba148996),
	.w3(32'h3b3bf1fa),
	.w4(32'h3b921710),
	.w5(32'h3aa778df),
	.w6(32'h3c40fc08),
	.w7(32'h3bda01d6),
	.w8(32'h3b6c0f10),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48dda3),
	.w1(32'h3ba89c45),
	.w2(32'hba65c7c5),
	.w3(32'hb977d8ae),
	.w4(32'hba85f3c9),
	.w5(32'h3aeb472a),
	.w6(32'hb8447a32),
	.w7(32'h3afe01d1),
	.w8(32'hbb5d32d9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1534d),
	.w1(32'hb9ebbc82),
	.w2(32'hbabcb06e),
	.w3(32'hbaee9a89),
	.w4(32'hbb630bc2),
	.w5(32'hbae1c6dd),
	.w6(32'h3a9a1504),
	.w7(32'h3a90b184),
	.w8(32'h3c414ff9),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedd176),
	.w1(32'hbc06ed3b),
	.w2(32'h393a94d5),
	.w3(32'h3a0038b6),
	.w4(32'hbb0885a6),
	.w5(32'h3896be72),
	.w6(32'h3ab2d532),
	.w7(32'hba667c4a),
	.w8(32'h39a376fa),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43e377),
	.w1(32'hba2f15e2),
	.w2(32'hb93edba3),
	.w3(32'h3a5597e2),
	.w4(32'h3a476626),
	.w5(32'h3b26d39a),
	.w6(32'hb917d728),
	.w7(32'hbb0583fe),
	.w8(32'hba80deba),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b6b8c),
	.w1(32'h3c29fac4),
	.w2(32'h3b0f9fc2),
	.w3(32'hba6a2e43),
	.w4(32'hbc6916ee),
	.w5(32'h3a416194),
	.w6(32'h3a36be0f),
	.w7(32'h3a4c9154),
	.w8(32'hba94853f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db627),
	.w1(32'h3a4d61b0),
	.w2(32'h3b04166a),
	.w3(32'hbb1f1ef7),
	.w4(32'hbb42ffb5),
	.w5(32'hbb22b520),
	.w6(32'hba1182f3),
	.w7(32'hbab7141e),
	.w8(32'hbb4dd1ea),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa795a),
	.w1(32'hba8bcbd7),
	.w2(32'hba01a95c),
	.w3(32'hbb7d05fb),
	.w4(32'hba51416c),
	.w5(32'hbad71372),
	.w6(32'hbbc71be7),
	.w7(32'hba3d8788),
	.w8(32'hbc224b79),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58706d),
	.w1(32'hbbdcdbfa),
	.w2(32'h3aed4da9),
	.w3(32'hbbb0aabd),
	.w4(32'hba129f4b),
	.w5(32'hbab085b6),
	.w6(32'hba8ecc56),
	.w7(32'h3b0db60f),
	.w8(32'hbb230e43),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b5ccd),
	.w1(32'h3a98e1bd),
	.w2(32'hbbb78ec0),
	.w3(32'hbab3b93c),
	.w4(32'hba0a5a21),
	.w5(32'hbbdfbb55),
	.w6(32'h3a220c6c),
	.w7(32'hbb0a416f),
	.w8(32'hbb9d9aff),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db98d),
	.w1(32'h3aa381f5),
	.w2(32'h3a99ac4c),
	.w3(32'h3b008058),
	.w4(32'h3c9b27bf),
	.w5(32'hbabdc431),
	.w6(32'h3b901e99),
	.w7(32'hbb6a5b15),
	.w8(32'hbb20c23a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394afe9b),
	.w1(32'hbc0695bf),
	.w2(32'hbbbd6c96),
	.w3(32'hbaab8798),
	.w4(32'h3b787b10),
	.w5(32'h3b71e2e9),
	.w6(32'h39581e3a),
	.w7(32'hba9c04fa),
	.w8(32'h3aaa9dd0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaac476),
	.w1(32'hbb82fd8e),
	.w2(32'hb920d09c),
	.w3(32'hbc2e5d15),
	.w4(32'hbb2eccbd),
	.w5(32'h3a939647),
	.w6(32'h3a6f6b2d),
	.w7(32'hbb5dca5b),
	.w8(32'h3be92863),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb581a83),
	.w1(32'hbbbdd368),
	.w2(32'h3a059ded),
	.w3(32'hbbaf3aac),
	.w4(32'h39bd81ee),
	.w5(32'hbbe76e86),
	.w6(32'h3adb95b1),
	.w7(32'h3ccb2188),
	.w8(32'h39e8a659),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd21f5),
	.w1(32'hbbd38b0e),
	.w2(32'hbb6bc5f9),
	.w3(32'hbbb51692),
	.w4(32'hbb4d58a9),
	.w5(32'hbad36be5),
	.w6(32'hbab09e81),
	.w7(32'hbbfcb95d),
	.w8(32'hbbbfb215),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98faa6),
	.w1(32'hba8e0589),
	.w2(32'hbb4a77e9),
	.w3(32'hb995c80f),
	.w4(32'hba25f665),
	.w5(32'hba6a1f25),
	.w6(32'hbbbdfb7e),
	.w7(32'h3b0895fb),
	.w8(32'h3a63f89a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a955647),
	.w1(32'hbc4209ac),
	.w2(32'hbb935741),
	.w3(32'hbb9597e2),
	.w4(32'h3abd5a70),
	.w5(32'hbb0e2954),
	.w6(32'hba564a7b),
	.w7(32'h3a1331eb),
	.w8(32'h3afea24e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91e4cd),
	.w1(32'hb7ce9fb3),
	.w2(32'hba4306a8),
	.w3(32'hbb1f3104),
	.w4(32'hbb926be6),
	.w5(32'h3a239717),
	.w6(32'hba76d5b8),
	.w7(32'hbb439cc8),
	.w8(32'h3c422e30),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d3fb4),
	.w1(32'hb9f9e636),
	.w2(32'h3bea2cba),
	.w3(32'h3bb98106),
	.w4(32'h3ba79601),
	.w5(32'hbc04dab2),
	.w6(32'hba417730),
	.w7(32'h3b3b7bd6),
	.w8(32'hbb03bb28),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a049ad1),
	.w1(32'h39124534),
	.w2(32'hbbb3850e),
	.w3(32'hbb82c4b7),
	.w4(32'h3bb99448),
	.w5(32'hbbf554d1),
	.w6(32'hbb69841c),
	.w7(32'hbaf1f1b2),
	.w8(32'h3a2bd109),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09b4a7),
	.w1(32'hbbbd14c5),
	.w2(32'hbbcf472b),
	.w3(32'hbb873383),
	.w4(32'hbbc9aa8a),
	.w5(32'hbc2ca06f),
	.w6(32'hbc20684c),
	.w7(32'hbc07dca0),
	.w8(32'hba80920f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61993d),
	.w1(32'hb9be7133),
	.w2(32'h39e1b470),
	.w3(32'hbba0ec25),
	.w4(32'h3a2c8015),
	.w5(32'hba6d6d67),
	.w6(32'h3a13a59d),
	.w7(32'h3c0a7eea),
	.w8(32'hbc3ca2e4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4ff7),
	.w1(32'h3b2be1ae),
	.w2(32'hb9022541),
	.w3(32'hbb766c8d),
	.w4(32'h3b9eede2),
	.w5(32'h3a9ba358),
	.w6(32'hba204d69),
	.w7(32'h3b07d796),
	.w8(32'hb90336ce),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63418e),
	.w1(32'h3bb3ba7e),
	.w2(32'hbb89ee29),
	.w3(32'h3ad06ef4),
	.w4(32'h3a326b5e),
	.w5(32'h3b9f8c2d),
	.w6(32'h3aec0339),
	.w7(32'h38fa651f),
	.w8(32'hbb7a967d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbababf83),
	.w1(32'hbab8c5a6),
	.w2(32'h3c5d893f),
	.w3(32'h3d1a41db),
	.w4(32'h3b3a823e),
	.w5(32'hbbcc15ca),
	.w6(32'h3b0144f2),
	.w7(32'hbb35beec),
	.w8(32'hbabbd06e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef2225),
	.w1(32'hbbf167f7),
	.w2(32'h3afd2390),
	.w3(32'h3aee931c),
	.w4(32'h3bf633d0),
	.w5(32'hbb94b5bb),
	.w6(32'h3bc0b560),
	.w7(32'hb93185f0),
	.w8(32'h39c383e4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb737110),
	.w1(32'hb8fd6e42),
	.w2(32'hbb923e3b),
	.w3(32'h3b96ed60),
	.w4(32'hbaa92eb1),
	.w5(32'hbba3fdb4),
	.w6(32'hbb3a9dba),
	.w7(32'h3a2428f8),
	.w8(32'hbacf78c3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cca518a),
	.w1(32'hba0346a1),
	.w2(32'hba87e345),
	.w3(32'h3a91c3b8),
	.w4(32'h3cce2f65),
	.w5(32'hbb9033ba),
	.w6(32'hbaf82985),
	.w7(32'hb8248c52),
	.w8(32'hbbf22efc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0bcba),
	.w1(32'h3b763287),
	.w2(32'h3b71dc2d),
	.w3(32'hbb46e347),
	.w4(32'hbca039fd),
	.w5(32'hba0d4728),
	.w6(32'h3bb76683),
	.w7(32'hbb5af2cc),
	.w8(32'hb7f57742),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae378ad),
	.w1(32'h3a5da047),
	.w2(32'hbaceac5f),
	.w3(32'h3cc733e3),
	.w4(32'hbc34dd6e),
	.w5(32'hbb679aab),
	.w6(32'h3a8b78ea),
	.w7(32'hbb748125),
	.w8(32'hbbc0a887),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edfe49),
	.w1(32'hbb6eed22),
	.w2(32'hbb8e888c),
	.w3(32'hbb11fde2),
	.w4(32'h39963dcd),
	.w5(32'hbbbd1a47),
	.w6(32'hbaeffb63),
	.w7(32'h39f46f54),
	.w8(32'h3b9f2d74),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1e797),
	.w1(32'hbb992843),
	.w2(32'hbb7157f0),
	.w3(32'hbb2037ec),
	.w4(32'hbc109d47),
	.w5(32'hbb7fc974),
	.w6(32'hbb9d8ddd),
	.w7(32'h3a3d1015),
	.w8(32'h39cf2636),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa46137),
	.w1(32'hbadd3598),
	.w2(32'hbac3cada),
	.w3(32'h3c36eb5a),
	.w4(32'h3b530bbf),
	.w5(32'hbb5feff3),
	.w6(32'hbb172282),
	.w7(32'h3a50007a),
	.w8(32'hbae561ef),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba16384),
	.w1(32'hba12c89b),
	.w2(32'hbbe8b2a1),
	.w3(32'hbba9b728),
	.w4(32'h3b29f667),
	.w5(32'hbbe5013b),
	.w6(32'h3bda7adf),
	.w7(32'h3ba020f6),
	.w8(32'hbb7eaa70),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe8a9c),
	.w1(32'h3b5e115e),
	.w2(32'hbb7590cb),
	.w3(32'h38b5b4c0),
	.w4(32'hbaec248c),
	.w5(32'h3c0a2929),
	.w6(32'hbbd50d31),
	.w7(32'hbb13ad78),
	.w8(32'hbac301da),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a583d),
	.w1(32'h3a6909ea),
	.w2(32'h39e41a27),
	.w3(32'h3b14155c),
	.w4(32'hbba0e9bb),
	.w5(32'h3c3fbba5),
	.w6(32'h3a332f53),
	.w7(32'h3a023144),
	.w8(32'h39093139),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1b450),
	.w1(32'h3b42acc2),
	.w2(32'h3bd251a9),
	.w3(32'hbaa6724f),
	.w4(32'h3b2c3789),
	.w5(32'h3a2b5b5b),
	.w6(32'hbb81b84b),
	.w7(32'h3d0d66d2),
	.w8(32'hbba93320),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a17a1),
	.w1(32'h3b2ce82d),
	.w2(32'h3a7987d3),
	.w3(32'h3b90808c),
	.w4(32'hba71f9d6),
	.w5(32'h3c24ba10),
	.w6(32'h3b7d9899),
	.w7(32'hbb32e38e),
	.w8(32'hbafb326d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05da20),
	.w1(32'h3c06e931),
	.w2(32'h3bc55097),
	.w3(32'hbb7ec88d),
	.w4(32'h3b69998a),
	.w5(32'hbbbd682f),
	.w6(32'hbb35f36b),
	.w7(32'h3b3c3c59),
	.w8(32'h3b877a4e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b280118),
	.w1(32'hbc75be20),
	.w2(32'hbbd2f6fa),
	.w3(32'hbbd67a1a),
	.w4(32'hbbc908bf),
	.w5(32'h3b812692),
	.w6(32'h3bc7a4e4),
	.w7(32'h3c0bb1ff),
	.w8(32'hbb88cd96),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba12d94),
	.w1(32'h3a84ee04),
	.w2(32'hbc8e0822),
	.w3(32'h388dd4c8),
	.w4(32'h3b42396c),
	.w5(32'hbb2b7bd4),
	.w6(32'h3a427773),
	.w7(32'h3c905e6f),
	.w8(32'h3aa6115a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c77b3),
	.w1(32'h3acc8390),
	.w2(32'h3a96def0),
	.w3(32'hbc3518ed),
	.w4(32'h39c21a5b),
	.w5(32'h3d63f75a),
	.w6(32'h3a262016),
	.w7(32'hbab412b5),
	.w8(32'h3a0f3e44),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c876be5),
	.w1(32'h3a7f9311),
	.w2(32'h3c4a670d),
	.w3(32'hbc5bd061),
	.w4(32'hbc34c55f),
	.w5(32'hbc4d7dd9),
	.w6(32'h3bb4b81a),
	.w7(32'hbb5a9c2c),
	.w8(32'hbc42fb54),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39126d65),
	.w1(32'hba4ee011),
	.w2(32'hbba56717),
	.w3(32'hbc434273),
	.w4(32'h3c199a53),
	.w5(32'hb809bba5),
	.w6(32'hbc342277),
	.w7(32'hbc194a66),
	.w8(32'hbb2a0e93),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4953ab),
	.w1(32'h3aceaaa2),
	.w2(32'hbb0c4cf2),
	.w3(32'h3b1006a5),
	.w4(32'h3c04a623),
	.w5(32'h3bc0a93e),
	.w6(32'h3b97807e),
	.w7(32'h3aa7fd51),
	.w8(32'h3bf80754),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbe907),
	.w1(32'h3b96e751),
	.w2(32'hbad2cefd),
	.w3(32'h3b98fbce),
	.w4(32'hbc114a91),
	.w5(32'hbbac3bcd),
	.w6(32'hbbf857f6),
	.w7(32'h3a60b370),
	.w8(32'h3a674672),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedbffd),
	.w1(32'h3c44d91d),
	.w2(32'hbbad6b6b),
	.w3(32'h3b1f19f1),
	.w4(32'h3b85bcd8),
	.w5(32'hb8c34545),
	.w6(32'hbb55eb4b),
	.w7(32'h3bea5c63),
	.w8(32'hbb96eb56),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5299e9),
	.w1(32'h3aa19ea6),
	.w2(32'h3aa4a341),
	.w3(32'hbb1b4dd4),
	.w4(32'h3b068431),
	.w5(32'hbc34acf0),
	.w6(32'h3bfd8ba3),
	.w7(32'hba0e7224),
	.w8(32'h3c2123e6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b182a31),
	.w1(32'hbc44fa0e),
	.w2(32'h3c14acd3),
	.w3(32'hbb525d5e),
	.w4(32'h3787ff8a),
	.w5(32'hbc202461),
	.w6(32'h3b0c9f25),
	.w7(32'hbd63c610),
	.w8(32'h38625c80),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a577fed),
	.w1(32'hbc8214c8),
	.w2(32'h3a1215bf),
	.w3(32'h3b9f21ea),
	.w4(32'hbc97da14),
	.w5(32'h39c0e0e6),
	.w6(32'h3c521fa3),
	.w7(32'hbbf6ad04),
	.w8(32'hba928161),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9103869),
	.w1(32'hbc8d2455),
	.w2(32'hbb4cb8f5),
	.w3(32'h3a983e8c),
	.w4(32'hbc16ac50),
	.w5(32'hbc6502d1),
	.w6(32'h3b407bc1),
	.w7(32'hb94804b7),
	.w8(32'hbb6b180a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cb6d3),
	.w1(32'hba44bc87),
	.w2(32'hbc6c82bd),
	.w3(32'h39116809),
	.w4(32'hbb114cb4),
	.w5(32'h3b17fe11),
	.w6(32'hbce087cb),
	.w7(32'h3ba2d957),
	.w8(32'h3b669f06),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4a13),
	.w1(32'hbbbc5463),
	.w2(32'h3c4b4810),
	.w3(32'h3c1bfcd4),
	.w4(32'h3c0c5581),
	.w5(32'hbbc76d53),
	.w6(32'h3bb52b48),
	.w7(32'hbbe16b90),
	.w8(32'hbc6b6aeb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3de9d07d),
	.w1(32'hbbbc2fce),
	.w2(32'hbc254aa9),
	.w3(32'h39ecd5f8),
	.w4(32'h3950f73b),
	.w5(32'hbc0bdaae),
	.w6(32'h3ad24d3f),
	.w7(32'h3cf54355),
	.w8(32'h38254cc2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf839c9),
	.w1(32'hbb459c51),
	.w2(32'hbc30141a),
	.w3(32'h3c064f82),
	.w4(32'hbb363974),
	.w5(32'hba3e870e),
	.w6(32'h3ad705fa),
	.w7(32'h3bf56fc4),
	.w8(32'h3b4c83f0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1f981),
	.w1(32'hbc36093e),
	.w2(32'hbb4b612c),
	.w3(32'hba568bef),
	.w4(32'hbc216248),
	.w5(32'h3b5eb549),
	.w6(32'h3b55f781),
	.w7(32'hbbfe6087),
	.w8(32'h3c223760),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ceb054),
	.w1(32'hbbbfc7f6),
	.w2(32'h3be550c4),
	.w3(32'hbbf1d783),
	.w4(32'hbbce0e38),
	.w5(32'h3bd16baa),
	.w6(32'hbbb9e644),
	.w7(32'hbc085687),
	.w8(32'h3bf12ee7),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dd0ba),
	.w1(32'hb963fa7e),
	.w2(32'hba2d6a29),
	.w3(32'hbcaf4ea0),
	.w4(32'hbbb13d9b),
	.w5(32'hbbb28250),
	.w6(32'h3b1e7c07),
	.w7(32'hbbb92913),
	.w8(32'hbc932183),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7061b5),
	.w1(32'h3d06b872),
	.w2(32'hbbcc899b),
	.w3(32'hbb16076b),
	.w4(32'h3babf3b7),
	.w5(32'hbb650b35),
	.w6(32'h3bd4b58c),
	.w7(32'h3ab86e6c),
	.w8(32'h3b9f0a6c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b6165),
	.w1(32'h3c3f2884),
	.w2(32'hbbbb3b96),
	.w3(32'hbb336446),
	.w4(32'h3a96217d),
	.w5(32'hbc024b1c),
	.w6(32'hbac37a02),
	.w7(32'hb9931343),
	.w8(32'hbba09c9f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcd815),
	.w1(32'hbc0994ca),
	.w2(32'h3b50f37f),
	.w3(32'h3bf2ca53),
	.w4(32'h3ba178e8),
	.w5(32'hbaa76f48),
	.w6(32'h3a721d4e),
	.w7(32'h3c7e6ae2),
	.w8(32'h3bd2d2bf),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb8864),
	.w1(32'hbbbb9053),
	.w2(32'hbbd76783),
	.w3(32'hba207fd9),
	.w4(32'h3bb706da),
	.w5(32'h3ba45539),
	.w6(32'h3b71f3cf),
	.w7(32'hba6c17f3),
	.w8(32'hb981885c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7dd06),
	.w1(32'hbc320605),
	.w2(32'hbbd5c62e),
	.w3(32'h3b953f9e),
	.w4(32'h3c1c2d88),
	.w5(32'hbb848a8c),
	.w6(32'h3ced47f0),
	.w7(32'h3b97a889),
	.w8(32'h3aea70ff),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59c597),
	.w1(32'h3b9cc5eb),
	.w2(32'hbc25393a),
	.w3(32'h3c6ed8df),
	.w4(32'hbbb369ee),
	.w5(32'hb598a6b2),
	.w6(32'hb9bb37fa),
	.w7(32'hb9c0a0d0),
	.w8(32'hbbcfa541),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7ce2f),
	.w1(32'hbba9f25d),
	.w2(32'hbb5e3362),
	.w3(32'h3be34cc8),
	.w4(32'hbc85bee3),
	.w5(32'h3a8913fc),
	.w6(32'hbbb7127a),
	.w7(32'hbb77bec7),
	.w8(32'h3b6c83b6),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bdb0e),
	.w1(32'hbc18c4fc),
	.w2(32'hbba260eb),
	.w3(32'h3af5ba17),
	.w4(32'h3b0d741d),
	.w5(32'h3bab17c7),
	.w6(32'hbb02ca14),
	.w7(32'h3b97116a),
	.w8(32'h3b006f42),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33a025),
	.w1(32'hba20e2a8),
	.w2(32'h3b996ac9),
	.w3(32'h3945a2f3),
	.w4(32'h3b11aa14),
	.w5(32'h3aaf15a0),
	.w6(32'h3b83d3ca),
	.w7(32'h3c0137e5),
	.w8(32'h3b20e9d1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafcb23),
	.w1(32'h3bf5516a),
	.w2(32'h3bde8415),
	.w3(32'hbb7ade35),
	.w4(32'h3af1c3dd),
	.w5(32'hbbc7ab1c),
	.w6(32'hbc9d9e94),
	.w7(32'hbbe8411f),
	.w8(32'hbc1edace),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule