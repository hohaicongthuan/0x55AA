module layer_10_featuremap_65(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5f880),
	.w1(32'hbd12486c),
	.w2(32'h3c2699cb),
	.w3(32'h3c020f58),
	.w4(32'hbcda3e93),
	.w5(32'hbc0fad8c),
	.w6(32'h3cbeffa2),
	.w7(32'hbac64c58),
	.w8(32'hbc78188e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd66247),
	.w1(32'h3bc2f231),
	.w2(32'h3c2fd1b5),
	.w3(32'h3cc9099e),
	.w4(32'h3ceb02f8),
	.w5(32'h3ba2d808),
	.w6(32'hbbde0fd2),
	.w7(32'h3cb9880f),
	.w8(32'h3bf600ed),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11af81),
	.w1(32'hbba0f51d),
	.w2(32'hbc081b02),
	.w3(32'hbc4cbd6c),
	.w4(32'hbbf89339),
	.w5(32'hbc458cc5),
	.w6(32'hbbfe0ce0),
	.w7(32'hbaaf5698),
	.w8(32'h39fb2a0b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5509e6),
	.w1(32'hbb66b0be),
	.w2(32'hbb2942da),
	.w3(32'hbba8db24),
	.w4(32'h3a4317b7),
	.w5(32'hbc1a7cf4),
	.w6(32'hbc10ebef),
	.w7(32'hbc3341ed),
	.w8(32'hbb7c9060),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c394d8c),
	.w1(32'hbb9bb8a2),
	.w2(32'hbc881c5a),
	.w3(32'hbc0ce640),
	.w4(32'h39deb5b2),
	.w5(32'hbc456583),
	.w6(32'h3a59546e),
	.w7(32'h3aaf77e4),
	.w8(32'hbc55a0dd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95798f),
	.w1(32'hbc22eeac),
	.w2(32'hb9925d75),
	.w3(32'hbc0e69e9),
	.w4(32'hbc15ec0b),
	.w5(32'hbb6806ed),
	.w6(32'hbc69aed5),
	.w7(32'hbc2436f8),
	.w8(32'hbb259fd4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cba88),
	.w1(32'hbd394372),
	.w2(32'hbd404476),
	.w3(32'hbcbb660d),
	.w4(32'hbd432203),
	.w5(32'hbd099f26),
	.w6(32'hbd0ab2bb),
	.w7(32'hbd4c684d),
	.w8(32'hbcf71436),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc845260),
	.w1(32'h3b5205ea),
	.w2(32'h3d3fd214),
	.w3(32'hbc2b2fee),
	.w4(32'h3ca8d2d6),
	.w5(32'h3cce80a7),
	.w6(32'h3c2341ad),
	.w7(32'h3a7e86dd),
	.w8(32'h3d338ddb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9635ce),
	.w1(32'hbcb7dae8),
	.w2(32'hbb855876),
	.w3(32'h3c199063),
	.w4(32'hbc76a509),
	.w5(32'h3bc5d336),
	.w6(32'h3c3e808d),
	.w7(32'h3af690b9),
	.w8(32'h3c1b0204),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37dac4),
	.w1(32'hbbb54398),
	.w2(32'h3ca3be8a),
	.w3(32'h3c05454f),
	.w4(32'hbc3b00c6),
	.w5(32'h3c5e7729),
	.w6(32'h3c3a5c4d),
	.w7(32'hbca72ff1),
	.w8(32'h3be4f093),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29ba76),
	.w1(32'hbb47bfd0),
	.w2(32'hbba31e2e),
	.w3(32'h3a5ad523),
	.w4(32'hb9faadc2),
	.w5(32'hbb68d856),
	.w6(32'hbb617358),
	.w7(32'h3a23ae9c),
	.w8(32'hbb4ac391),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d032d73),
	.w1(32'hbd183f5b),
	.w2(32'hbd0bb41d),
	.w3(32'h3b4d16b7),
	.w4(32'hbd5ea3c8),
	.w5(32'hbcf03489),
	.w6(32'hbccaa59f),
	.w7(32'hbd8bef1b),
	.w8(32'hbc3a87ec),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26f2e5),
	.w1(32'hbc8d07f1),
	.w2(32'h3abc7493),
	.w3(32'hbbd1a41f),
	.w4(32'hbcac0507),
	.w5(32'h3b4f338c),
	.w6(32'hbc0873e5),
	.w7(32'hbca27511),
	.w8(32'h3b7e77f5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd88072),
	.w1(32'hbb1cb71f),
	.w2(32'h3cb200bf),
	.w3(32'hbcaebc01),
	.w4(32'hbb8d9010),
	.w5(32'h3c91b80c),
	.w6(32'hbbbc1a24),
	.w7(32'hbba84f0d),
	.w8(32'h3ca095db),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be9b7c),
	.w1(32'hbc3f237f),
	.w2(32'h3be61100),
	.w3(32'hbb9c43bc),
	.w4(32'hbc00a2bf),
	.w5(32'hbbbaa7b7),
	.w6(32'h3bb0bffb),
	.w7(32'hbc67d263),
	.w8(32'h3b64ffa4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e8ae5),
	.w1(32'h3bd09de0),
	.w2(32'h3d21bd57),
	.w3(32'h3cb34f79),
	.w4(32'h3ccd590b),
	.w5(32'h3d44a493),
	.w6(32'h3c171319),
	.w7(32'h3cfe6bd0),
	.w8(32'h3d107d43),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b022916),
	.w1(32'hbb92d467),
	.w2(32'h3c108c2c),
	.w3(32'h3babd8cd),
	.w4(32'hb91b492a),
	.w5(32'h3bd9942f),
	.w6(32'hbb189056),
	.w7(32'h398968c0),
	.w8(32'h3c737679),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81abec),
	.w1(32'hbca7ded5),
	.w2(32'h3c8cc611),
	.w3(32'h3bdb12b1),
	.w4(32'hbc8d39e8),
	.w5(32'h3cd697af),
	.w6(32'h3b513b6a),
	.w7(32'hbbada450),
	.w8(32'h3d083465),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31731a),
	.w1(32'hbcb58e99),
	.w2(32'h3c484410),
	.w3(32'hbbbc64ca),
	.w4(32'hbcbb6c46),
	.w5(32'h3bbd33e9),
	.w6(32'hbc28732d),
	.w7(32'hbc5a796a),
	.w8(32'hbc529919),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9194a),
	.w1(32'h3c2b4057),
	.w2(32'h3b3d7b66),
	.w3(32'h3c2ca680),
	.w4(32'h3c817a9e),
	.w5(32'hb9fe1e53),
	.w6(32'h3a3236b2),
	.w7(32'h3c74ac6d),
	.w8(32'h3b1f699e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc54780),
	.w1(32'h3bb25ec8),
	.w2(32'hbb8f979b),
	.w3(32'hbbe4eb59),
	.w4(32'hbb15dc7e),
	.w5(32'hbb80951c),
	.w6(32'hbc37d981),
	.w7(32'hbbef4c33),
	.w8(32'hbad15232),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad55993),
	.w1(32'hbc6249f4),
	.w2(32'h3c1dbb96),
	.w3(32'hbb7cd1de),
	.w4(32'h3bcc2dec),
	.w5(32'h3baf092f),
	.w6(32'h3b1e5c61),
	.w7(32'h3b40f8b0),
	.w8(32'h3a394d1c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d565f3e),
	.w1(32'hbd3566ba),
	.w2(32'hbb78ac42),
	.w3(32'h3d966cdf),
	.w4(32'hbc664526),
	.w5(32'h3d1888c9),
	.w6(32'h3c876567),
	.w7(32'hbcdf5204),
	.w8(32'h3d25eec4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c868762),
	.w1(32'hbc0bbc60),
	.w2(32'h3b60fd63),
	.w3(32'h3bd71718),
	.w4(32'hbc5b29de),
	.w5(32'hba4d9c6e),
	.w6(32'h3c960c13),
	.w7(32'hbbfb0a9f),
	.w8(32'h3c09fccf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7408f0),
	.w1(32'hbcafd13e),
	.w2(32'h3c8deaac),
	.w3(32'h3c396628),
	.w4(32'hbc48ad6b),
	.w5(32'h3d06a90a),
	.w6(32'h3cba1f37),
	.w7(32'hba9b9ae3),
	.w8(32'h3d0f9fd6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a7285),
	.w1(32'h3ac10fe9),
	.w2(32'hbc0bc6f1),
	.w3(32'h3b85ed1b),
	.w4(32'h3c591cf8),
	.w5(32'hbbb5f2be),
	.w6(32'h3c88c940),
	.w7(32'h3bc9286d),
	.w8(32'hbb9b6ae9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae16f6d),
	.w1(32'hbb7780b6),
	.w2(32'h37db974a),
	.w3(32'hbbccb4a0),
	.w4(32'hbb60aefa),
	.w5(32'hb9a69810),
	.w6(32'hbc5d5f7f),
	.w7(32'hbc148934),
	.w8(32'hbad46659),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55793d),
	.w1(32'hbcb26c27),
	.w2(32'hbc5131ed),
	.w3(32'hbbc168df),
	.w4(32'hbc01d7c1),
	.w5(32'hb9eda63e),
	.w6(32'hbc545994),
	.w7(32'hbad7696f),
	.w8(32'h3b82dd7b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb867cda),
	.w1(32'hbb0e3a13),
	.w2(32'hbc3425df),
	.w3(32'h3c24fe61),
	.w4(32'h3c1d4a11),
	.w5(32'h3c5e313d),
	.w6(32'h3c455544),
	.w7(32'h3b4c2333),
	.w8(32'h3b4be6a2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54f7b2),
	.w1(32'hbc998121),
	.w2(32'h3b8bb1e1),
	.w3(32'h3c2409fc),
	.w4(32'hbc9c72ed),
	.w5(32'h3c250d07),
	.w6(32'h3b8fd1f7),
	.w7(32'hbcfdc5a1),
	.w8(32'h3c04eb7a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e4a5b),
	.w1(32'h3aa86221),
	.w2(32'h39e1ba5c),
	.w3(32'h3bd91a0c),
	.w4(32'h3b8f46da),
	.w5(32'hbbe0619d),
	.w6(32'h3b8daec8),
	.w7(32'h3b156fb2),
	.w8(32'hbca3eecb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb961f0),
	.w1(32'hbb7bce9e),
	.w2(32'hb9232efd),
	.w3(32'hbc8df7db),
	.w4(32'hbc9fd776),
	.w5(32'h3bd57616),
	.w6(32'hbba90010),
	.w7(32'hbbd5d9a1),
	.w8(32'hbc001aa3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03925a),
	.w1(32'h3b142d71),
	.w2(32'h3bcd396b),
	.w3(32'h3b876a9b),
	.w4(32'hbc2cae8d),
	.w5(32'h3ada6af9),
	.w6(32'hbc6ef18e),
	.w7(32'hbc63d312),
	.w8(32'h3b8bbb05),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ab3a),
	.w1(32'hbb99211d),
	.w2(32'hbb2af3c5),
	.w3(32'h3b8c19d0),
	.w4(32'h3a2396aa),
	.w5(32'h3c0d2922),
	.w6(32'h3b14d282),
	.w7(32'h39b16f46),
	.w8(32'hbbfa093d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff674f),
	.w1(32'hbc01b03d),
	.w2(32'h3b5f5c75),
	.w3(32'hbba6b478),
	.w4(32'hbc7278d7),
	.w5(32'h3b967131),
	.w6(32'hbc18647e),
	.w7(32'h3c461a6a),
	.w8(32'h3b78abff),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87dabce),
	.w1(32'hbc7672b5),
	.w2(32'hbca1c431),
	.w3(32'hbb509115),
	.w4(32'hbcabbb2a),
	.w5(32'h3c569974),
	.w6(32'hbc0d823b),
	.w7(32'hbc9cd77c),
	.w8(32'hbcfdac78),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8b5ff6),
	.w1(32'h3c8f1aa3),
	.w2(32'hbd90f24c),
	.w3(32'h3dc0fe5b),
	.w4(32'hbc0e3e82),
	.w5(32'hbd39d2dc),
	.w6(32'hbc570461),
	.w7(32'hbd525c9a),
	.w8(32'hbc7fb7ac),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b886fd9),
	.w1(32'hbcb3380c),
	.w2(32'h3c568439),
	.w3(32'h3c82e29d),
	.w4(32'hbb1847e4),
	.w5(32'hbb513f41),
	.w6(32'h3cf47cf4),
	.w7(32'h39a78c39),
	.w8(32'h3d07c27d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9963e3),
	.w1(32'hbd18a019),
	.w2(32'h3bf6ea5b),
	.w3(32'hbc3546f7),
	.w4(32'hbcab2863),
	.w5(32'h3c4f5fcb),
	.w6(32'h3c8c3f9b),
	.w7(32'hbc9d8836),
	.w8(32'h3c85fd5a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe95f3d),
	.w1(32'hbbb6edfc),
	.w2(32'hbb3feaad),
	.w3(32'hbbe07c61),
	.w4(32'h3ba0175c),
	.w5(32'hbb30ac29),
	.w6(32'hbc09ebcf),
	.w7(32'h3b2d5d6c),
	.w8(32'h3a29380a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034869),
	.w1(32'hbbb25f9b),
	.w2(32'hbba605ea),
	.w3(32'hbbe828c4),
	.w4(32'hbb360b7e),
	.w5(32'hbb59e550),
	.w6(32'hbbfa941e),
	.w7(32'hbb115a1b),
	.w8(32'hba88fd37),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc873226),
	.w1(32'hbb6c23ef),
	.w2(32'h3a88caa8),
	.w3(32'h3c079cb1),
	.w4(32'h3c1e5c38),
	.w5(32'hbc21e7f6),
	.w6(32'hbbc1b9bc),
	.w7(32'hbc215d64),
	.w8(32'h3901f55b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e76ca),
	.w1(32'hbbf773af),
	.w2(32'h3b5e601b),
	.w3(32'hbc3ba667),
	.w4(32'hbca7def6),
	.w5(32'h3b90076c),
	.w6(32'h3c2cb772),
	.w7(32'hbbc3e069),
	.w8(32'h3bee070f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01761c),
	.w1(32'hbc83ae85),
	.w2(32'h3d17dbd0),
	.w3(32'h3c619cd1),
	.w4(32'hbc097f48),
	.w5(32'h3d1ff92d),
	.w6(32'h3cbfc88b),
	.w7(32'h3b83c080),
	.w8(32'h3ca4d879),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3cb5b),
	.w1(32'hbcd09af2),
	.w2(32'hbc99ec4c),
	.w3(32'h3cc08549),
	.w4(32'h3b761c58),
	.w5(32'hb6681bb0),
	.w6(32'h3c626a20),
	.w7(32'hbc854b29),
	.w8(32'h3c2c4419),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bed79),
	.w1(32'hbc3442dc),
	.w2(32'h39ac4856),
	.w3(32'h3d5e16db),
	.w4(32'h3cc51bef),
	.w5(32'h3bf9975c),
	.w6(32'h3d510d3a),
	.w7(32'hbcc92fdf),
	.w8(32'h3d0a6867),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c756178),
	.w1(32'h3c0f873b),
	.w2(32'h3ae1e138),
	.w3(32'h3d69c16e),
	.w4(32'h3cc76f3b),
	.w5(32'h3b9eb46d),
	.w6(32'h3d0c2c44),
	.w7(32'hbc6a8671),
	.w8(32'h3c1ab22f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82709a),
	.w1(32'hbd166831),
	.w2(32'hbc97ee41),
	.w3(32'hbb5a7c02),
	.w4(32'hbd0a6b72),
	.w5(32'hbac1d9e6),
	.w6(32'hbcfedb5c),
	.w7(32'hbd24a7f4),
	.w8(32'h3bcb4caa),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d88d4),
	.w1(32'hbadc3708),
	.w2(32'hbc00b37c),
	.w3(32'hbb43bb89),
	.w4(32'hbb7ae6b7),
	.w5(32'hbb436a44),
	.w6(32'hbaa2fb2c),
	.w7(32'hbb991c49),
	.w8(32'h3b9bc6c0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843754),
	.w1(32'hbc0601eb),
	.w2(32'h3c30d314),
	.w3(32'h3c9bc440),
	.w4(32'h3c026ea7),
	.w5(32'hbc0200eb),
	.w6(32'h3c83dabf),
	.w7(32'h3b52643c),
	.w8(32'hbc0a93ac),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4221b8),
	.w1(32'hbbd83e23),
	.w2(32'h3c5f5030),
	.w3(32'hbc54df63),
	.w4(32'h3b435928),
	.w5(32'hbcb5b1e2),
	.w6(32'hbc009632),
	.w7(32'h3c475ccf),
	.w8(32'h3bc6d4be),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09717e),
	.w1(32'hbbeb2af3),
	.w2(32'h3cdc7a00),
	.w3(32'hbc52deea),
	.w4(32'h3b58eca9),
	.w5(32'h3cb42373),
	.w6(32'h3c1ae0ea),
	.w7(32'h3b14e112),
	.w8(32'hbc2c8283),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6f025),
	.w1(32'hbb316b90),
	.w2(32'h3c03bc20),
	.w3(32'h3a48cd5c),
	.w4(32'h3c02f033),
	.w5(32'h3a0f1041),
	.w6(32'h3b9129b8),
	.w7(32'h3c843e32),
	.w8(32'h3b6f318e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42245b),
	.w1(32'hbce2aff0),
	.w2(32'h3d02ea87),
	.w3(32'hbbe9b122),
	.w4(32'hbcc139fb),
	.w5(32'h3c3c596a),
	.w6(32'hbb67a918),
	.w7(32'hbc8b769e),
	.w8(32'h3c87be69),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8d561),
	.w1(32'hbbf007ff),
	.w2(32'h3bf5e162),
	.w3(32'hbc092573),
	.w4(32'hbbf38bd7),
	.w5(32'h3d1b50a8),
	.w6(32'h3c398140),
	.w7(32'h3ba9a03a),
	.w8(32'hbc3f0f92),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb49b40),
	.w1(32'h3cc668fd),
	.w2(32'hbc0d5d45),
	.w3(32'h3cf2b41f),
	.w4(32'h3b8567b5),
	.w5(32'h3b97595c),
	.w6(32'hbc9b7830),
	.w7(32'h39eecf26),
	.w8(32'h3c673bc8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5599),
	.w1(32'h3c6ca8d5),
	.w2(32'hbbfa5752),
	.w3(32'h3c5f89bf),
	.w4(32'h3c6174d9),
	.w5(32'hb9e8ee84),
	.w6(32'hbbf9db31),
	.w7(32'h3a871f4b),
	.w8(32'hbb7c109b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0b9d2),
	.w1(32'hbc045738),
	.w2(32'hb7e9e264),
	.w3(32'hbacea414),
	.w4(32'hbc0b9c13),
	.w5(32'hbadbd3fe),
	.w6(32'hbbb622f9),
	.w7(32'hbc39d6cf),
	.w8(32'h3b124d30),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e1e68),
	.w1(32'hbb0a7c75),
	.w2(32'h3b36e0c3),
	.w3(32'hbb8378e5),
	.w4(32'hbbb4fa68),
	.w5(32'h3a015d77),
	.w6(32'h3b1dbecb),
	.w7(32'h3b576546),
	.w8(32'h38d33272),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f5095),
	.w1(32'hbb85df05),
	.w2(32'hbbb3d601),
	.w3(32'hbada2d6e),
	.w4(32'hbb7e8c53),
	.w5(32'hbb5449cd),
	.w6(32'hbb39c484),
	.w7(32'hb8f704d9),
	.w8(32'hbb14a177),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8de65),
	.w1(32'hbc395c81),
	.w2(32'hb984932a),
	.w3(32'h3c168df0),
	.w4(32'h3abe4906),
	.w5(32'h3c5bdc5f),
	.w6(32'h3a06843e),
	.w7(32'hbbf56041),
	.w8(32'h3ce983f4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87b379),
	.w1(32'h3951117c),
	.w2(32'h3c3b0db4),
	.w3(32'h3c956a98),
	.w4(32'h3c58d4f8),
	.w5(32'h3c8fcba4),
	.w6(32'hba936a28),
	.w7(32'hbc025e87),
	.w8(32'h3d0a4c86),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef4425),
	.w1(32'h3c869e25),
	.w2(32'h3b5cd6b8),
	.w3(32'h3c5915ec),
	.w4(32'h3c0ed0bf),
	.w5(32'hb8acd71e),
	.w6(32'h3a7972bb),
	.w7(32'hbc910d04),
	.w8(32'hbb39e46e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb142a25),
	.w1(32'hbbb152b1),
	.w2(32'h3c35b3c4),
	.w3(32'hbb2000f1),
	.w4(32'hbbe7ef49),
	.w5(32'h3cd36ccd),
	.w6(32'hb96c6436),
	.w7(32'h3babe9af),
	.w8(32'hbc0b7dc7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46745d),
	.w1(32'h3c35801b),
	.w2(32'h3ad619ef),
	.w3(32'h3c2db3b7),
	.w4(32'hbbb2a10a),
	.w5(32'h3ad41c3f),
	.w6(32'hbab88229),
	.w7(32'h3c2d3843),
	.w8(32'hbb5dc39c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d9b2a),
	.w1(32'hbb7eea97),
	.w2(32'hba1bb578),
	.w3(32'h3933a84d),
	.w4(32'h39d96196),
	.w5(32'h3acdc79d),
	.w6(32'hbb49602b),
	.w7(32'h3ad95283),
	.w8(32'h3a9f0fc1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff461),
	.w1(32'hbb840f86),
	.w2(32'h3d6a65b0),
	.w3(32'h3bfd1cca),
	.w4(32'hb92c0a72),
	.w5(32'h3d31c9ea),
	.w6(32'hbcd1be69),
	.w7(32'hbc21e08d),
	.w8(32'h3cc09f96),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aeee2a),
	.w1(32'hbc94ee3a),
	.w2(32'h3c8a241d),
	.w3(32'h3bf33819),
	.w4(32'h378fb468),
	.w5(32'h3c6256f5),
	.w6(32'h3cbf7495),
	.w7(32'h3ca15dc8),
	.w8(32'h3d5e0d6b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a1f3f),
	.w1(32'hbc97586c),
	.w2(32'h3ca63733),
	.w3(32'h3bd60ace),
	.w4(32'hbc88f948),
	.w5(32'h3c9ebcf2),
	.w6(32'h3c8abebc),
	.w7(32'h3bd395a7),
	.w8(32'h3ce9e26c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae631de),
	.w1(32'hbd0a5ded),
	.w2(32'h3c22236c),
	.w3(32'h3bb55962),
	.w4(32'hbce2d347),
	.w5(32'h3c3b43a1),
	.w6(32'h3cef3d8e),
	.w7(32'hbb085d1b),
	.w8(32'h3d01f417),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1941c2),
	.w1(32'h3a46484d),
	.w2(32'h3b131407),
	.w3(32'h3b738030),
	.w4(32'h3ba55447),
	.w5(32'hba957a61),
	.w6(32'hbbb9ce20),
	.w7(32'hbb859d26),
	.w8(32'h3a68f129),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf4731),
	.w1(32'hb9ece6f0),
	.w2(32'hbbbe1fd8),
	.w3(32'h3b3aa4a6),
	.w4(32'h3b58a33c),
	.w5(32'h3c8eeb62),
	.w6(32'hbab00412),
	.w7(32'h3a0805aa),
	.w8(32'h3c05e48e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87db35),
	.w1(32'h3c46a25c),
	.w2(32'h3c52b01a),
	.w3(32'h3cf135e5),
	.w4(32'h3cad87a3),
	.w5(32'hbcceac41),
	.w6(32'h3b6d1eaf),
	.w7(32'hbc79af64),
	.w8(32'h3af18a7a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce61ac1),
	.w1(32'h3a2233f3),
	.w2(32'h3ac0afe2),
	.w3(32'hbd090e00),
	.w4(32'hbcf91e8a),
	.w5(32'h3b006f36),
	.w6(32'h3cd3597c),
	.w7(32'h3cd8f3ce),
	.w8(32'h3b58e6c2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e7ff7),
	.w1(32'hbbc4d718),
	.w2(32'hbabe215a),
	.w3(32'hbaceac99),
	.w4(32'hbb85c103),
	.w5(32'hbbecec91),
	.w6(32'hbb0c45bc),
	.w7(32'hbbbbcf01),
	.w8(32'hbc1b2c7e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b393b21),
	.w1(32'hbc1645f1),
	.w2(32'hbb513df7),
	.w3(32'h3b712d3c),
	.w4(32'hbbb98fe2),
	.w5(32'h3b803ba2),
	.w6(32'hbcbe8216),
	.w7(32'hbcf17a3a),
	.w8(32'hbc462b9b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a29e0),
	.w1(32'h3af426b8),
	.w2(32'h3ba1f14f),
	.w3(32'h3b2b8862),
	.w4(32'hbc7fd861),
	.w5(32'hbb1a0292),
	.w6(32'h3cd745af),
	.w7(32'h3c4dc12e),
	.w8(32'h3c93c5b2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce757ca),
	.w1(32'hbb42f38a),
	.w2(32'h3b8a0e8b),
	.w3(32'h3c24fb05),
	.w4(32'hbc5dd881),
	.w5(32'h3c863402),
	.w6(32'h3ca2ab11),
	.w7(32'h3b8caffc),
	.w8(32'h3b7768c6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2319ee),
	.w1(32'h3c2fa11b),
	.w2(32'h3cafc9cf),
	.w3(32'h3cafde70),
	.w4(32'h3b568b3d),
	.w5(32'h3c8f77dc),
	.w6(32'h3b77ab7f),
	.w7(32'hbab1148a),
	.w8(32'h3c6ae037),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bf936),
	.w1(32'hbc830ede),
	.w2(32'h3c1392f2),
	.w3(32'h39eb8746),
	.w4(32'hbc798a7d),
	.w5(32'hbb917b6e),
	.w6(32'hbbd517b2),
	.w7(32'hbc9fa814),
	.w8(32'h3bf69ecf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a943ad1),
	.w1(32'hbb87c9d4),
	.w2(32'h3bb48df9),
	.w3(32'h3c0e93e3),
	.w4(32'h3b9a4f03),
	.w5(32'h3bf8ecb7),
	.w6(32'h3b87d1dc),
	.w7(32'hbaa66b67),
	.w8(32'hbb591a6f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34f808),
	.w1(32'hbc8bcd53),
	.w2(32'hbc9b1f58),
	.w3(32'hba018757),
	.w4(32'hbc70dfcc),
	.w5(32'h3c3b3d32),
	.w6(32'hbc2eb157),
	.w7(32'hbcb883f5),
	.w8(32'h3bc1aed7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48bdf9),
	.w1(32'hbc58b0ea),
	.w2(32'h3aa1a97a),
	.w3(32'h3ce51afc),
	.w4(32'h3c91defb),
	.w5(32'h3c30408d),
	.w6(32'hbad33879),
	.w7(32'hbc188208),
	.w8(32'h3be45c03),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15351c),
	.w1(32'h3c0084e0),
	.w2(32'hbc8460fe),
	.w3(32'h3c59b072),
	.w4(32'h3b850e79),
	.w5(32'h3c2d55b0),
	.w6(32'hbb583b58),
	.w7(32'hbbc0d866),
	.w8(32'h3c95df1d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba964c16),
	.w1(32'h3ba72801),
	.w2(32'hbbc95657),
	.w3(32'h3d06c90b),
	.w4(32'h3c827d3d),
	.w5(32'hbb9c0fae),
	.w6(32'h3bb13d21),
	.w7(32'hbc220dc1),
	.w8(32'hbc23a97d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d327a),
	.w1(32'h3b7eb3be),
	.w2(32'h3b1eead4),
	.w3(32'hbc2c6b41),
	.w4(32'h3b684ae1),
	.w5(32'h3b9f531b),
	.w6(32'hbbdd70e1),
	.w7(32'hbb841fe7),
	.w8(32'h3b309ad3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b5021),
	.w1(32'h3c087d1a),
	.w2(32'hbc74be8b),
	.w3(32'h3cf77b65),
	.w4(32'h3cbb07fc),
	.w5(32'hbc7893c2),
	.w6(32'h3cd7866d),
	.w7(32'h3c2e7fb6),
	.w8(32'hbc231ae1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ebf4f),
	.w1(32'hbb4ab9bf),
	.w2(32'h3c8efdf7),
	.w3(32'hbbf83f64),
	.w4(32'hbbb9ca83),
	.w5(32'hbc1c87df),
	.w6(32'hba9bdd3d),
	.w7(32'hb99b0bfe),
	.w8(32'hbc448653),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6180f0),
	.w1(32'h3b126712),
	.w2(32'h3bc3166e),
	.w3(32'h3c5f2480),
	.w4(32'h3cc14375),
	.w5(32'h3c23b8ab),
	.w6(32'h3cd9fb40),
	.w7(32'h3cef2c6a),
	.w8(32'h3c1bb27b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cd422),
	.w1(32'hbc5c816f),
	.w2(32'h3bfb7937),
	.w3(32'h3c4cff19),
	.w4(32'hbc03f074),
	.w5(32'h3c928653),
	.w6(32'h3b961231),
	.w7(32'hbb327530),
	.w8(32'h3c891d9a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab572b6),
	.w1(32'hbc80f5de),
	.w2(32'hbc568a8a),
	.w3(32'h3bda94b9),
	.w4(32'hbc111c4a),
	.w5(32'h3b6dc6b4),
	.w6(32'hbb404996),
	.w7(32'hbcda7923),
	.w8(32'hb97e8756),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd3b2a5),
	.w1(32'hbcd805d4),
	.w2(32'hbbb96078),
	.w3(32'h3d13e8e2),
	.w4(32'hbcbcbf48),
	.w5(32'h3c68f628),
	.w6(32'hbb9408f8),
	.w7(32'hbd2457c2),
	.w8(32'h3bf308d2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab61081),
	.w1(32'hbbc04b3c),
	.w2(32'hbb9bd604),
	.w3(32'h3adf290b),
	.w4(32'hbc06ea28),
	.w5(32'hba8705c6),
	.w6(32'hba8c6f59),
	.w7(32'hbbb92ebe),
	.w8(32'h3aeff726),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb350794),
	.w1(32'hbc2b8ab2),
	.w2(32'h3d73b887),
	.w3(32'h3c3c4aa6),
	.w4(32'h3a9d3ff7),
	.w5(32'h3d4d97d6),
	.w6(32'h3c9ce44f),
	.w7(32'h3cba7c74),
	.w8(32'h3d58aa94),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e750c),
	.w1(32'hbc082a81),
	.w2(32'h3ca4b090),
	.w3(32'h3c6a355c),
	.w4(32'h3c252b8e),
	.w5(32'h3be5fc9b),
	.w6(32'h3c4f3c56),
	.w7(32'h3b9165b0),
	.w8(32'h3ce1fe85),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50b563),
	.w1(32'hbc930cb7),
	.w2(32'h3af66189),
	.w3(32'h3d1108c3),
	.w4(32'h3cfd7bc7),
	.w5(32'h3c8cf8ce),
	.w6(32'h3d4ac49e),
	.w7(32'hbac9c1f3),
	.w8(32'h3c1425f2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831dac),
	.w1(32'h3bc55c96),
	.w2(32'hbc72e1e6),
	.w3(32'h3b82234f),
	.w4(32'h3b2b85fa),
	.w5(32'hbb258824),
	.w6(32'hbb289aba),
	.w7(32'hbbaaeca9),
	.w8(32'h3c1bcfb7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3925cf),
	.w1(32'hbc594922),
	.w2(32'h3cae3774),
	.w3(32'h3ca5f7ee),
	.w4(32'hbca13226),
	.w5(32'h3bf5c4fe),
	.w6(32'h3b8ac17e),
	.w7(32'hbca353ac),
	.w8(32'h3aff254d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfdfeed),
	.w1(32'hbd0899bd),
	.w2(32'hbc43637f),
	.w3(32'h3c4218b3),
	.w4(32'hbd260278),
	.w5(32'hbc874a96),
	.w6(32'hbcb9423f),
	.w7(32'hbd1b73e3),
	.w8(32'hbc9d4dc1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e85ec),
	.w1(32'h3bfcc11b),
	.w2(32'hbd283872),
	.w3(32'h3d6dfee4),
	.w4(32'h3bd9a2fa),
	.w5(32'hbcccfca8),
	.w6(32'h3bb9af25),
	.w7(32'hbd038de3),
	.w8(32'h3c49298f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d29da33),
	.w1(32'h3b83992b),
	.w2(32'h3bd7020e),
	.w3(32'h3bb277f0),
	.w4(32'hbb63ef35),
	.w5(32'h3be5c482),
	.w6(32'h3d39499f),
	.w7(32'h3d0edd8d),
	.w8(32'h3cb34d87),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb29d20),
	.w1(32'hba7771d4),
	.w2(32'h3b6e1165),
	.w3(32'hb9c0cc70),
	.w4(32'hbcdb7def),
	.w5(32'h3b5429a4),
	.w6(32'h3ce67de3),
	.w7(32'h3c14f305),
	.w8(32'h3c6be59b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ac658),
	.w1(32'hbc747567),
	.w2(32'hbcf2fab0),
	.w3(32'h3ce33266),
	.w4(32'hbd37a64f),
	.w5(32'hbca26ede),
	.w6(32'hbb91d21a),
	.w7(32'hbd8fd23d),
	.w8(32'hbca0e0e3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b301fb3),
	.w1(32'h3a81b5b6),
	.w2(32'h3b9b9d72),
	.w3(32'hbbc99b46),
	.w4(32'h3b06974a),
	.w5(32'h3c534a34),
	.w6(32'h3bb2ada2),
	.w7(32'hb993ad30),
	.w8(32'h3a15955f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810132),
	.w1(32'h3ce99849),
	.w2(32'hbd08c7cc),
	.w3(32'h3d474095),
	.w4(32'h3d0acfc0),
	.w5(32'hbc9f3c7f),
	.w6(32'hbc1e4797),
	.w7(32'hbd923b1a),
	.w8(32'hbc503dde),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa6e7f),
	.w1(32'h3b545904),
	.w2(32'hbcfeeeac),
	.w3(32'h3baae52e),
	.w4(32'hbc812e2c),
	.w5(32'hbd0019be),
	.w6(32'h3ba11f6f),
	.w7(32'hbce50aea),
	.w8(32'hbd2bbcd3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6824e),
	.w1(32'h3b53210e),
	.w2(32'h3b5ca7c7),
	.w3(32'h3b7f377a),
	.w4(32'h3b02bb91),
	.w5(32'h3c078f99),
	.w6(32'h3acbe42f),
	.w7(32'hba845d89),
	.w8(32'h3bd4d711),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf408fd),
	.w1(32'hbc098afe),
	.w2(32'hbc3022ca),
	.w3(32'h3be2ffb4),
	.w4(32'h3ba87f3f),
	.w5(32'h3d02cf7a),
	.w6(32'h3ba9bb3a),
	.w7(32'h3b8e8767),
	.w8(32'h3cc3e2a2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2df4c4),
	.w1(32'h3a49c2cd),
	.w2(32'h3be60353),
	.w3(32'h3cceb9d3),
	.w4(32'hbb7d7e37),
	.w5(32'hbc0f63dd),
	.w6(32'h3b2e384d),
	.w7(32'hbc7bc698),
	.w8(32'hbb12da58),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb504b01),
	.w1(32'hbc490ea3),
	.w2(32'hbc2ca259),
	.w3(32'hbc81ae3e),
	.w4(32'hbccf9d47),
	.w5(32'h3a58894e),
	.w6(32'h3c619755),
	.w7(32'hbae4fdc0),
	.w8(32'h3c06cae3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95bcbb),
	.w1(32'hbbd25b1a),
	.w2(32'h3bc2800b),
	.w3(32'h3c17f49f),
	.w4(32'hbc283fb7),
	.w5(32'h3b1b0a89),
	.w6(32'h3ab2fc7f),
	.w7(32'hbc478628),
	.w8(32'h3cbea06d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa5b6e),
	.w1(32'h3b745060),
	.w2(32'h3aeda436),
	.w3(32'h3cbdd8e6),
	.w4(32'h3c81d24d),
	.w5(32'h3c8196aa),
	.w6(32'h3c74e947),
	.w7(32'h3bb51417),
	.w8(32'h3c5e5aa2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2774a),
	.w1(32'hbcdfae5d),
	.w2(32'hbd2c5c76),
	.w3(32'h3ba22001),
	.w4(32'hbcb13772),
	.w5(32'hbd1d5878),
	.w6(32'h3c5e953c),
	.w7(32'h3b2d686f),
	.w8(32'h3bfc8210),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc299671),
	.w1(32'hbb398b4b),
	.w2(32'h3cd9e0bb),
	.w3(32'h3b437c3a),
	.w4(32'hbb83e5d6),
	.w5(32'h3d59f8f5),
	.w6(32'h3ca54c24),
	.w7(32'h3be65937),
	.w8(32'h3cef9b12),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c842e4e),
	.w1(32'h3c54a890),
	.w2(32'hbb1622a0),
	.w3(32'h3ce385c6),
	.w4(32'hbb0794e0),
	.w5(32'hba344e7b),
	.w6(32'hb9c51961),
	.w7(32'hba8f04bc),
	.w8(32'h3bbf1250),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e5ca3),
	.w1(32'h3abf86b8),
	.w2(32'hbbe6e265),
	.w3(32'h3b195a8a),
	.w4(32'h3bb0e7bc),
	.w5(32'hbb751af2),
	.w6(32'h3a5a63b7),
	.w7(32'h3a9d36ea),
	.w8(32'hbb497937),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46d94d),
	.w1(32'hbb96c67a),
	.w2(32'h3bd93014),
	.w3(32'hbb254de5),
	.w4(32'hba9f217e),
	.w5(32'h3b6d1077),
	.w6(32'hbbdcd6da),
	.w7(32'hbb2e9673),
	.w8(32'h3ac4fcab),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4e8ba),
	.w1(32'h3abaa2d6),
	.w2(32'h3bd54c7d),
	.w3(32'hbb084835),
	.w4(32'h39ae1d0a),
	.w5(32'hbc8accc5),
	.w6(32'h3b4dc101),
	.w7(32'h3b92b4a3),
	.w8(32'hbc1df145),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c296c20),
	.w1(32'hbaa2eb24),
	.w2(32'h3c32427e),
	.w3(32'hbd019c44),
	.w4(32'hbcc0018e),
	.w5(32'hbb923b38),
	.w6(32'h39290806),
	.w7(32'h3c173d0b),
	.w8(32'hbb9f75b5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb421af),
	.w1(32'h3c3b9fc1),
	.w2(32'hbb1c86e9),
	.w3(32'hb9f1dac1),
	.w4(32'hbc73eb8c),
	.w5(32'hbb1e1994),
	.w6(32'h3cd1f9de),
	.w7(32'h3be8cfd4),
	.w8(32'h3c560899),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b266591),
	.w1(32'h3bacd7ab),
	.w2(32'hbaa5cd9d),
	.w3(32'h394a6534),
	.w4(32'h3bb5d769),
	.w5(32'hbb457816),
	.w6(32'h3c37501a),
	.w7(32'hbc0de0d7),
	.w8(32'hbb5577ec),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2c0fb),
	.w1(32'hbc9857fa),
	.w2(32'hbc51ccc7),
	.w3(32'hbc04d221),
	.w4(32'hbc8b5414),
	.w5(32'hbc43a4aa),
	.w6(32'hbc94f9d3),
	.w7(32'hbcf0222c),
	.w8(32'hbc236936),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fdbb9),
	.w1(32'hbad0cf8e),
	.w2(32'h3cc8ec5a),
	.w3(32'h3c7b822c),
	.w4(32'h3c14ab11),
	.w5(32'h3cfd8c53),
	.w6(32'h3c73331d),
	.w7(32'h3bf0cc10),
	.w8(32'h3d051e9f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bf756),
	.w1(32'h3b323ce8),
	.w2(32'h3ab6fa2e),
	.w3(32'h3ba5868e),
	.w4(32'h3b89c9d2),
	.w5(32'h3bad897d),
	.w6(32'h3b1f683a),
	.w7(32'hbbd149a6),
	.w8(32'h3bdc5f99),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa62db4),
	.w1(32'h3ac5d413),
	.w2(32'h3c1c5417),
	.w3(32'h3bb54482),
	.w4(32'h3ba3fae0),
	.w5(32'hbabe1341),
	.w6(32'h3b8bd58b),
	.w7(32'hb9dc850c),
	.w8(32'hbbbcd546),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44caed),
	.w1(32'h3ad35953),
	.w2(32'hbb19eb47),
	.w3(32'hbac12a63),
	.w4(32'h3baaa9fe),
	.w5(32'h3c9a55ad),
	.w6(32'h3c00f185),
	.w7(32'h3c944971),
	.w8(32'h3bbd0b41),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99784a5),
	.w1(32'h3ba5a7b5),
	.w2(32'hbb542dc3),
	.w3(32'h3cc0ea77),
	.w4(32'h3c9dbff0),
	.w5(32'h3c851ab1),
	.w6(32'hbbcaf1a6),
	.w7(32'hbc08db9f),
	.w8(32'h3b9ef0f2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc45437),
	.w1(32'hbd74a0b7),
	.w2(32'hbd1fa2d5),
	.w3(32'hbc61b257),
	.w4(32'hbcd2c513),
	.w5(32'hbbe017c0),
	.w6(32'h3c1e5b33),
	.w7(32'hbc46473d),
	.w8(32'h3d4c867e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b167f),
	.w1(32'hbc857343),
	.w2(32'h3c8e916d),
	.w3(32'hbbc70a32),
	.w4(32'hbc80f31c),
	.w5(32'h3c257574),
	.w6(32'hbc324fb3),
	.w7(32'hbc0206aa),
	.w8(32'h3c1d3759),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1035de),
	.w1(32'h3a820af1),
	.w2(32'hbc8a92e9),
	.w3(32'h3b790337),
	.w4(32'hbc1935e1),
	.w5(32'hbc5b473e),
	.w6(32'hbc592e03),
	.w7(32'hbc80644c),
	.w8(32'h39cfe03a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f809c),
	.w1(32'hbadcdca3),
	.w2(32'h3c4cd18d),
	.w3(32'hbba33d6f),
	.w4(32'hbc12cfef),
	.w5(32'hbb9d9886),
	.w6(32'hbac9e99a),
	.w7(32'hbacc0a77),
	.w8(32'h3cbca4c5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c096605),
	.w1(32'h3c22ae5c),
	.w2(32'h3c1d8185),
	.w3(32'h3bbe6d8c),
	.w4(32'h3b6b9cec),
	.w5(32'hbc82e44b),
	.w6(32'h3c532a1d),
	.w7(32'hbc485c85),
	.w8(32'h3c933f87),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ab39b),
	.w1(32'hbc5da0da),
	.w2(32'h3c899bfe),
	.w3(32'h3c70f26c),
	.w4(32'h3cad33d3),
	.w5(32'h3cf6154d),
	.w6(32'h3d34828d),
	.w7(32'h3c892436),
	.w8(32'h3c1fce69),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a0b6a),
	.w1(32'hbba36d58),
	.w2(32'h3c5a0d50),
	.w3(32'h3c6107c2),
	.w4(32'h3c36f4e1),
	.w5(32'h3c852cb3),
	.w6(32'hbbb99562),
	.w7(32'hbaab436e),
	.w8(32'h3c08cccb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c6b9a),
	.w1(32'hbce693ab),
	.w2(32'h3c19868f),
	.w3(32'h3b873c00),
	.w4(32'hbcbfa2c8),
	.w5(32'h3ba5cc57),
	.w6(32'hbcd7b6f3),
	.w7(32'hbcf53b26),
	.w8(32'h3bcdd8c9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c330846),
	.w1(32'hbbabb929),
	.w2(32'h3c023ea8),
	.w3(32'hbbdd710b),
	.w4(32'h3b771d1d),
	.w5(32'h3c9b2a61),
	.w6(32'h3c6aabf9),
	.w7(32'h3c9b108a),
	.w8(32'h3c6134b9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8189b5),
	.w1(32'h3b87292a),
	.w2(32'h3ad21798),
	.w3(32'h3c6f4098),
	.w4(32'hbb2319f7),
	.w5(32'h3c18b99d),
	.w6(32'hbb22fc24),
	.w7(32'hbc229612),
	.w8(32'h3bdfd154),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a3130),
	.w1(32'hbcfceea7),
	.w2(32'hba91622a),
	.w3(32'h3bcae899),
	.w4(32'hbcfcedc7),
	.w5(32'h3c0af981),
	.w6(32'hbc982cf6),
	.w7(32'hbd2025ef),
	.w8(32'h3c6fd646),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53a19a),
	.w1(32'h3bbe5840),
	.w2(32'hbbed1b82),
	.w3(32'h3c9219f0),
	.w4(32'h3c4af94c),
	.w5(32'hbc6df85e),
	.w6(32'h3cce3a2c),
	.w7(32'h3c745940),
	.w8(32'h3c2f8c82),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb10021),
	.w1(32'h3b8ccc88),
	.w2(32'h3bf8f7e8),
	.w3(32'h3bd040fa),
	.w4(32'hbae03fa0),
	.w5(32'h3b2d8ccc),
	.w6(32'h3be6d794),
	.w7(32'hbbc2296f),
	.w8(32'h3c1d81e0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba061a6e),
	.w1(32'hbb2f1930),
	.w2(32'h3b738afd),
	.w3(32'hbb921859),
	.w4(32'hbbd3fc4a),
	.w5(32'h3c541236),
	.w6(32'h3a9cad73),
	.w7(32'hbb4cbae6),
	.w8(32'h3b9d21ef),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e0b5b),
	.w1(32'hbd08826c),
	.w2(32'h3c9e54bb),
	.w3(32'h3ca9f9d9),
	.w4(32'hbc749472),
	.w5(32'h3a9ac37a),
	.w6(32'h3cea6b40),
	.w7(32'hbc218ae7),
	.w8(32'h3d4dd3fa),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c314542),
	.w1(32'hbb84497e),
	.w2(32'hbab32c86),
	.w3(32'h3c379800),
	.w4(32'h3d044f24),
	.w5(32'h3c04b95a),
	.w6(32'h3d15a6d4),
	.w7(32'h3be74666),
	.w8(32'h3b108972),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac31ec3),
	.w1(32'hbae5a7e6),
	.w2(32'hb9e5c9e0),
	.w3(32'hba24dbd9),
	.w4(32'h39a51349),
	.w5(32'hba7bc3cd),
	.w6(32'h3b6da409),
	.w7(32'h3c20dd7f),
	.w8(32'h39c89990),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80c97c),
	.w1(32'hbaedf659),
	.w2(32'hbb1068a8),
	.w3(32'h3ab585b7),
	.w4(32'h3a18d535),
	.w5(32'hbc2c90c9),
	.w6(32'hb9be65fa),
	.w7(32'h38b47b71),
	.w8(32'hb83f6082),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a94ef),
	.w1(32'h3b4d2521),
	.w2(32'hbb9d0dca),
	.w3(32'hbba2adfe),
	.w4(32'hbbdb3a11),
	.w5(32'hbaf7ca12),
	.w6(32'h3bb8cd61),
	.w7(32'h3b67798a),
	.w8(32'h3b1a21fe),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3c3cf),
	.w1(32'h3b0335ab),
	.w2(32'hbcbe83b5),
	.w3(32'h3cfe68f3),
	.w4(32'h3c5b3d6f),
	.w5(32'hbc94152b),
	.w6(32'h3c9274c7),
	.w7(32'hbbae4903),
	.w8(32'hbc10280d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80fe55),
	.w1(32'hbc34a326),
	.w2(32'h3c82e514),
	.w3(32'h3b79b412),
	.w4(32'hbcaee868),
	.w5(32'h3c137d43),
	.w6(32'h3c01ec0a),
	.w7(32'hbc6bac77),
	.w8(32'h3c49eca6),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadfdbd),
	.w1(32'h3a313918),
	.w2(32'hbc8d7524),
	.w3(32'hbbb9d6b9),
	.w4(32'h3b3ea067),
	.w5(32'h3b5a4e95),
	.w6(32'h3c0b979d),
	.w7(32'h3bc60c9e),
	.w8(32'h3c242fab),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a40ca),
	.w1(32'hbadfb3cf),
	.w2(32'h3c8b4c16),
	.w3(32'h3c91ac69),
	.w4(32'hbaddcf7e),
	.w5(32'hb8bc5215),
	.w6(32'h3bcfd021),
	.w7(32'hbcaa9f0d),
	.w8(32'h3c493c56),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc40d0),
	.w1(32'hbc07eaf9),
	.w2(32'hbb2e5c24),
	.w3(32'hbc06eb36),
	.w4(32'hbc427ab5),
	.w5(32'hbae18678),
	.w6(32'h3c170e86),
	.w7(32'hbb395440),
	.w8(32'hb8d52128),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05cbc2),
	.w1(32'hbd1c22ff),
	.w2(32'hba557b6a),
	.w3(32'h3bae7fdd),
	.w4(32'hbd0d6649),
	.w5(32'h3c4314d2),
	.w6(32'hbcc447a4),
	.w7(32'hbd4b6f47),
	.w8(32'hbb6bd7fd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb005b0a),
	.w1(32'hbce02053),
	.w2(32'hbc0d938d),
	.w3(32'h3cba3dc7),
	.w4(32'hbba0878f),
	.w5(32'hbbd36b5d),
	.w6(32'h3bf48dad),
	.w7(32'hbce766eb),
	.w8(32'hbc04c7c2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af112dd),
	.w1(32'h3b18c8d3),
	.w2(32'h3c408fd4),
	.w3(32'h3cdbf041),
	.w4(32'h3b3476e6),
	.w5(32'h3c71364c),
	.w6(32'h3cdeebc2),
	.w7(32'h3a764f0c),
	.w8(32'h3c91cacf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e4295),
	.w1(32'h3a6d1ff8),
	.w2(32'hbb07e71b),
	.w3(32'hbc508442),
	.w4(32'hba0aad18),
	.w5(32'hbb5da7fe),
	.w6(32'h3c9a2536),
	.w7(32'h3c8e12ca),
	.w8(32'hbafcfd69),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c310934),
	.w1(32'hbb954e97),
	.w2(32'hba986078),
	.w3(32'h3c2d88e7),
	.w4(32'hba95f8df),
	.w5(32'hb99525b6),
	.w6(32'h3ca31ba7),
	.w7(32'hbb13f2a7),
	.w8(32'hbc0b25c7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07c6cf),
	.w1(32'h3b16783e),
	.w2(32'h3bcc4556),
	.w3(32'h3c9f4fb0),
	.w4(32'h3bb97a65),
	.w5(32'hbb5d5f69),
	.w6(32'h3cbba371),
	.w7(32'h3c1d813c),
	.w8(32'hbc50b9db),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e9313),
	.w1(32'hbbe30295),
	.w2(32'h37f1906c),
	.w3(32'h3bc2ccdb),
	.w4(32'hbc6e0319),
	.w5(32'h3b90cb47),
	.w6(32'h3c23b3a8),
	.w7(32'hbc439082),
	.w8(32'h3bfefb98),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a956a97),
	.w1(32'hbc05426c),
	.w2(32'h3b152669),
	.w3(32'h3adb8bd3),
	.w4(32'hbbdf5ae5),
	.w5(32'hba85c9fe),
	.w6(32'hbb9e151b),
	.w7(32'hbc474ad4),
	.w8(32'hbbe80330),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba31248),
	.w1(32'hbb4f7524),
	.w2(32'h3acf21d4),
	.w3(32'hbadc0716),
	.w4(32'hbc688e28),
	.w5(32'h3bb31124),
	.w6(32'h3c32d96d),
	.w7(32'hbc425e06),
	.w8(32'h3b0a86e6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf560fd),
	.w1(32'hbb54c7c9),
	.w2(32'h3c033689),
	.w3(32'hbc916266),
	.w4(32'hbd1b8cf2),
	.w5(32'h3ac3f5f0),
	.w6(32'h3be353f7),
	.w7(32'hbca8960d),
	.w8(32'h3c9d2035),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1a639),
	.w1(32'hbbd67928),
	.w2(32'h3b2c6a9e),
	.w3(32'hbb80dfa0),
	.w4(32'hbc488015),
	.w5(32'h3b0ff4cc),
	.w6(32'h3bab6d3d),
	.w7(32'hbbe48298),
	.w8(32'h3b28b5f6),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c164b7c),
	.w1(32'hbc3c5731),
	.w2(32'h3bdacbfe),
	.w3(32'h3cb71853),
	.w4(32'hbbb4124c),
	.w5(32'h3c06e146),
	.w6(32'h3d08473c),
	.w7(32'h385a3ad4),
	.w8(32'h3c1548d2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a8ba6),
	.w1(32'h3b918d32),
	.w2(32'hbb6b8898),
	.w3(32'h3a52ba15),
	.w4(32'h3b2affe5),
	.w5(32'h3b5ad150),
	.w6(32'h3bab2584),
	.w7(32'hb9bb2363),
	.w8(32'h3bbf0513),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97d77e),
	.w1(32'hbb7b5f34),
	.w2(32'h3bb2d0c1),
	.w3(32'hbd163bf8),
	.w4(32'hbca585fa),
	.w5(32'h3c08daa6),
	.w6(32'hbceab2f8),
	.w7(32'hbcb45e14),
	.w8(32'h3c74105d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7904c),
	.w1(32'h3af4e50f),
	.w2(32'hba51154e),
	.w3(32'hbb0334c5),
	.w4(32'hbb94d503),
	.w5(32'h3b096c08),
	.w6(32'h3be7f1d9),
	.w7(32'hbb37eca7),
	.w8(32'h3c6997a9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fbeae),
	.w1(32'h3bda4365),
	.w2(32'hbbd5ad39),
	.w3(32'hbc9c1fef),
	.w4(32'h3a1efdfa),
	.w5(32'hbc3b0766),
	.w6(32'hbb2069fd),
	.w7(32'hbc3e3c21),
	.w8(32'hbc89e3c6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4950c5),
	.w1(32'h3b9041b6),
	.w2(32'h3a24faa7),
	.w3(32'h3c91f4d8),
	.w4(32'h3c20e5ae),
	.w5(32'h3b25e2df),
	.w6(32'h3c8b4227),
	.w7(32'hbb9c3d90),
	.w8(32'h3ac9e137),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd5b68c),
	.w1(32'hbc816b5a),
	.w2(32'hbc4ac646),
	.w3(32'h3c9c2627),
	.w4(32'hbcc5ca8e),
	.w5(32'hbba29f61),
	.w6(32'h3ce33da7),
	.w7(32'hbc058219),
	.w8(32'h3cdb0b76),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5767a7),
	.w1(32'h3b8d5ac0),
	.w2(32'hba33abe2),
	.w3(32'hbbddfc39),
	.w4(32'hba49a142),
	.w5(32'hbc2fdc52),
	.w6(32'h3b03242c),
	.w7(32'h38aaeca9),
	.w8(32'hbbb22c08),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc06f72),
	.w1(32'hbc0f52c1),
	.w2(32'h3b6294ad),
	.w3(32'hbb3c2332),
	.w4(32'hbc81ee60),
	.w5(32'h3bd8eba7),
	.w6(32'h3c519ab6),
	.w7(32'hbb8abb7b),
	.w8(32'h3c0036b7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3116ca),
	.w1(32'h3aed7ee7),
	.w2(32'h3b8d39a1),
	.w3(32'h3b19362e),
	.w4(32'h3c05ce17),
	.w5(32'hbbbbaf5d),
	.w6(32'h3b2726ac),
	.w7(32'hbaf1b09f),
	.w8(32'hbc7be885),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf13d5b),
	.w1(32'hbccf9274),
	.w2(32'h3d2b01df),
	.w3(32'h3cd1b6ef),
	.w4(32'hbd03cf03),
	.w5(32'h3d3568b3),
	.w6(32'h3b4cd24c),
	.w7(32'hbc96081c),
	.w8(32'h3c4280f9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77550),
	.w1(32'h3c00fb3d),
	.w2(32'h3c0aa081),
	.w3(32'h3c3790a3),
	.w4(32'h3b8c44ca),
	.w5(32'h3b7ddd88),
	.w6(32'h3d053e20),
	.w7(32'hbb9fb6e7),
	.w8(32'h3c1c5d3b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ba231),
	.w1(32'hbcaf6b66),
	.w2(32'h3842076a),
	.w3(32'h39a03702),
	.w4(32'hbba2a214),
	.w5(32'h3c03abf9),
	.w6(32'hbc44b1fd),
	.w7(32'h3aed1efd),
	.w8(32'h3d282b55),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32b5a9),
	.w1(32'h3bb62156),
	.w2(32'hbb3db65b),
	.w3(32'hbc2c375d),
	.w4(32'h3cc8e1fa),
	.w5(32'hbad902a5),
	.w6(32'hbcb2ef44),
	.w7(32'h3c889dae),
	.w8(32'hbc02b8ca),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b574b4),
	.w1(32'hbc150f1e),
	.w2(32'h3c41f13d),
	.w3(32'h3c4d3ea6),
	.w4(32'h3ae63afb),
	.w5(32'h3bbe1285),
	.w6(32'h3b2edc33),
	.w7(32'hbba8fff5),
	.w8(32'hba43efd6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4f35e),
	.w1(32'hbb90ce71),
	.w2(32'h3c8a7162),
	.w3(32'hbb0df9c5),
	.w4(32'h3be04187),
	.w5(32'h3c9892d4),
	.w6(32'h39c38b0d),
	.w7(32'hbbbd80a7),
	.w8(32'h3c55ae2c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917fc5a),
	.w1(32'h3c0dd9e9),
	.w2(32'h3b22359a),
	.w3(32'h3bc81777),
	.w4(32'h3b51a505),
	.w5(32'h3ba2810d),
	.w6(32'h3bae77f0),
	.w7(32'h3bfc2f84),
	.w8(32'h3b873958),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c8fb7),
	.w1(32'h3bb93a03),
	.w2(32'h3c9e1ea2),
	.w3(32'hbc399f38),
	.w4(32'h3b03d9ae),
	.w5(32'h3cb52866),
	.w6(32'h3b602574),
	.w7(32'h3c10a320),
	.w8(32'h3c55e54c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c92c0),
	.w1(32'h3b9ccac7),
	.w2(32'h3d1ea879),
	.w3(32'h3c940415),
	.w4(32'h3c564c85),
	.w5(32'h3d06ad6e),
	.w6(32'h3be3823a),
	.w7(32'h3c86162a),
	.w8(32'h3cd1734d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a69c1),
	.w1(32'hbbf1ac9e),
	.w2(32'hb9a4ac64),
	.w3(32'hba7efbeb),
	.w4(32'hbb900a04),
	.w5(32'hbc9ee5d1),
	.w6(32'h3b9c86a9),
	.w7(32'hbbe42af0),
	.w8(32'hbcbc0328),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c173b11),
	.w1(32'hbc95ee17),
	.w2(32'h3c21d5d7),
	.w3(32'h3ca1e22f),
	.w4(32'hbc02f27a),
	.w5(32'h3b3dd86f),
	.w6(32'hbafd2e54),
	.w7(32'h3b9bf0af),
	.w8(32'hbadda713),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1728b8),
	.w1(32'h39c23f0f),
	.w2(32'h3d067eb8),
	.w3(32'h3c675811),
	.w4(32'hbb3c9b8e),
	.w5(32'h3cd64d9e),
	.w6(32'h3c24dc89),
	.w7(32'h3a6d8b6a),
	.w8(32'hba198517),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd8205),
	.w1(32'hbc6fb9c7),
	.w2(32'hbc800e7a),
	.w3(32'h3cebb97b),
	.w4(32'hbce8294e),
	.w5(32'hbc800d70),
	.w6(32'h3cd4fd29),
	.w7(32'hbd4d6308),
	.w8(32'hbd2db7cf),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d62a6),
	.w1(32'hbbd75023),
	.w2(32'hbd1a3435),
	.w3(32'h3c5f6b04),
	.w4(32'hbb00231a),
	.w5(32'hbd04220b),
	.w6(32'hbc9b0263),
	.w7(32'hbc9f60b8),
	.w8(32'hbce988d0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e6886),
	.w1(32'h3bc0b7ac),
	.w2(32'h3bae9f81),
	.w3(32'h3bab7297),
	.w4(32'h3b7741a3),
	.w5(32'h3c30639b),
	.w6(32'h3b981b27),
	.w7(32'hbb15b81e),
	.w8(32'h3c749dbb),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6dcadc),
	.w1(32'hbcd2d8c3),
	.w2(32'h3ca08fe1),
	.w3(32'hbcbf25b3),
	.w4(32'hbd2f8441),
	.w5(32'h3c90bf77),
	.w6(32'hbcfdff2a),
	.w7(32'hbcbfb478),
	.w8(32'h3d223288),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d9323),
	.w1(32'hb9b6856e),
	.w2(32'h3c3c1e8a),
	.w3(32'h3d181e76),
	.w4(32'h3ce83f0d),
	.w5(32'h3cac1fbc),
	.w6(32'h3bf0db3e),
	.w7(32'h3b9584ce),
	.w8(32'hbaf14c8e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c7a4c),
	.w1(32'hbb9c6c2b),
	.w2(32'hbc22a9ec),
	.w3(32'h3b7d3292),
	.w4(32'hbbd6973e),
	.w5(32'hbcac9266),
	.w6(32'h3b7e1554),
	.w7(32'hbc1df523),
	.w8(32'hbc46b414),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4299ca),
	.w1(32'hbc4bd41c),
	.w2(32'hba78d76a),
	.w3(32'hbbf90ee7),
	.w4(32'h3af45d2d),
	.w5(32'hbb038ad4),
	.w6(32'hbc8d161b),
	.w7(32'h3c1f880f),
	.w8(32'h3a4f1b8d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07ba0d),
	.w1(32'hb9c08162),
	.w2(32'hbad3e01f),
	.w3(32'hbc587ca9),
	.w4(32'hbc1a838c),
	.w5(32'h37cf74ac),
	.w6(32'hb9f9db15),
	.w7(32'hbb045e94),
	.w8(32'h3bfaefb3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c16c3),
	.w1(32'h3c435a68),
	.w2(32'h3a522d6e),
	.w3(32'h3b166f4b),
	.w4(32'h3b01fdba),
	.w5(32'h3b210342),
	.w6(32'h3b4c6268),
	.w7(32'h3b94b6f5),
	.w8(32'h3b66be64),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90edad),
	.w1(32'hbca22e5b),
	.w2(32'hbcae2716),
	.w3(32'hbc53e54d),
	.w4(32'hbcd44569),
	.w5(32'hbc9ea188),
	.w6(32'hbc034f36),
	.w7(32'hbce541ea),
	.w8(32'hbc1a20f1),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5de318),
	.w1(32'h3c1d78a0),
	.w2(32'hbbbfacb8),
	.w3(32'h39289d0c),
	.w4(32'hbb9a4ff7),
	.w5(32'h3ac14ebc),
	.w6(32'h3c2f7b5d),
	.w7(32'h391a4685),
	.w8(32'h3c79b32f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6de2b3),
	.w1(32'hbba3e702),
	.w2(32'h3bfc4e9f),
	.w3(32'h3b78d5e1),
	.w4(32'hbc2a40af),
	.w5(32'h3b48b3bb),
	.w6(32'h3c9ba9a3),
	.w7(32'hbbb050b8),
	.w8(32'hbb44d890),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba091276),
	.w1(32'h3b9afda4),
	.w2(32'hb9e79533),
	.w3(32'h3b8a9255),
	.w4(32'h3b4de43c),
	.w5(32'hbae0d8a6),
	.w6(32'h3a25e3a3),
	.w7(32'h3bd33216),
	.w8(32'h3bb71521),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c007202),
	.w1(32'hbc01a11b),
	.w2(32'h3aa747a6),
	.w3(32'hbb9682e8),
	.w4(32'hbca104fc),
	.w5(32'h3beb4549),
	.w6(32'hbc4515fd),
	.w7(32'hbca3951d),
	.w8(32'h3cb4e9e7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05d95c),
	.w1(32'h3c5ce704),
	.w2(32'hbc61d791),
	.w3(32'hbc22109d),
	.w4(32'h3c397798),
	.w5(32'hbcf81595),
	.w6(32'hbc1a47fc),
	.w7(32'hbb713e2f),
	.w8(32'hbcca527e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fad5),
	.w1(32'hbbca77ee),
	.w2(32'hbbb7cce5),
	.w3(32'h3c13c4a3),
	.w4(32'hbc4f538a),
	.w5(32'hb9373560),
	.w6(32'h3c19e5a2),
	.w7(32'hbb0fcb75),
	.w8(32'h3ba21284),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97d7f2),
	.w1(32'h3c38910d),
	.w2(32'h3bcf7cbc),
	.w3(32'h3cb80f52),
	.w4(32'h3c63e295),
	.w5(32'h3c578b55),
	.w6(32'h3bd34f99),
	.w7(32'h3ccd1a57),
	.w8(32'hbb960b98),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1245f),
	.w1(32'hba30f683),
	.w2(32'hbb49c627),
	.w3(32'hbc589f99),
	.w4(32'hbc836b9e),
	.w5(32'hbbaff551),
	.w6(32'h3b89e6a1),
	.w7(32'hbceb477e),
	.w8(32'hbbeb04b9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd5c34),
	.w1(32'hbbceb4c3),
	.w2(32'hbbf92034),
	.w3(32'h3bb5c2e2),
	.w4(32'hbbe4c1e9),
	.w5(32'hb9984c04),
	.w6(32'h3ba33a54),
	.w7(32'hbc22d5b7),
	.w8(32'hbc18edee),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf40f98),
	.w1(32'hbc491ad9),
	.w2(32'hbb0259df),
	.w3(32'h3c603489),
	.w4(32'hb7b01ea0),
	.w5(32'h3c44b5d4),
	.w6(32'h3ce1c4b3),
	.w7(32'h3c04fde9),
	.w8(32'h3a8776b9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0945c8),
	.w1(32'h3b3a294d),
	.w2(32'h3be7686f),
	.w3(32'h3c700413),
	.w4(32'hbb40a0b2),
	.w5(32'h3bd80074),
	.w6(32'h3cadb04d),
	.w7(32'hbaac4a0b),
	.w8(32'h3a7a9a25),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f12eb),
	.w1(32'h3c062f17),
	.w2(32'hbbe7d5c4),
	.w3(32'h3c4d18d5),
	.w4(32'hbb4b5755),
	.w5(32'hbb8a1028),
	.w6(32'h3ca25caa),
	.w7(32'hbb27d6ec),
	.w8(32'hbbe40c83),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d338774),
	.w1(32'hbc75aaf4),
	.w2(32'h3a830d09),
	.w3(32'h3d83779e),
	.w4(32'h3cb9f710),
	.w5(32'h3b4be1bc),
	.w6(32'h3d30d70f),
	.w7(32'h3d472e2f),
	.w8(32'h3b654c2b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91868f),
	.w1(32'h3b7c25cf),
	.w2(32'h3c5cfa42),
	.w3(32'hbb829440),
	.w4(32'h3aeda5e2),
	.w5(32'h3c166726),
	.w6(32'h3ba60d72),
	.w7(32'h3bb215bd),
	.w8(32'h3cb018e5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2b442),
	.w1(32'hbc16d723),
	.w2(32'h3c0a8c22),
	.w3(32'hbb4050cf),
	.w4(32'hbc960576),
	.w5(32'h397a7602),
	.w6(32'hbc35cd09),
	.w7(32'hbcbf7d7b),
	.w8(32'h3bafa0f2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29643e),
	.w1(32'h3bea0c52),
	.w2(32'hbb2302c8),
	.w3(32'hbbd535ed),
	.w4(32'h3a3886be),
	.w5(32'h3b410f45),
	.w6(32'h39a68fb6),
	.w7(32'h3b453f82),
	.w8(32'h3c4724a4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01d1dd),
	.w1(32'h3c59e36e),
	.w2(32'hbc149c3b),
	.w3(32'hbb20be4c),
	.w4(32'h3c14aec9),
	.w5(32'hbc50a9e9),
	.w6(32'hbbb89ffe),
	.w7(32'hb9b109c5),
	.w8(32'h3ad28382),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2f1a9),
	.w1(32'hbc1e0b43),
	.w2(32'hbc805042),
	.w3(32'h3b64de60),
	.w4(32'hbcaae11d),
	.w5(32'hbd1997b9),
	.w6(32'h3c1d08f6),
	.w7(32'hbcae074d),
	.w8(32'h3cf2af1d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cedc529),
	.w1(32'hbb852457),
	.w2(32'h3b7ccbf0),
	.w3(32'h3c8f482c),
	.w4(32'h3b39eb3a),
	.w5(32'h3c3ee285),
	.w6(32'h3c07edf7),
	.w7(32'h3c8ebcd1),
	.w8(32'h3cbc5b67),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fc803),
	.w1(32'h3aa506a7),
	.w2(32'h3c0c510b),
	.w3(32'h3cafa265),
	.w4(32'h39220975),
	.w5(32'h3bba283e),
	.w6(32'h3d633f29),
	.w7(32'hbc90f1e1),
	.w8(32'h3c2c9186),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6759c7),
	.w1(32'hbd164301),
	.w2(32'hbc20bd4e),
	.w3(32'h3c7cf7d9),
	.w4(32'hbd41c072),
	.w5(32'hbc187669),
	.w6(32'hbc71d6ab),
	.w7(32'hbd4270c1),
	.w8(32'hbbf088a4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36810b),
	.w1(32'hbbbbb4bd),
	.w2(32'h3ca2eec3),
	.w3(32'hbc22574e),
	.w4(32'hbbdc7e90),
	.w5(32'h3c5c785c),
	.w6(32'hbbf5b8c6),
	.w7(32'hbb664795),
	.w8(32'h3c1f39bf),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83ca09),
	.w1(32'h3b5009d1),
	.w2(32'h3c1853b1),
	.w3(32'hbc2533f7),
	.w4(32'hba98e596),
	.w5(32'h3b44cb76),
	.w6(32'h3a201930),
	.w7(32'h3bec2cbf),
	.w8(32'h3c5b20f9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdf17a1),
	.w1(32'hbc9b645f),
	.w2(32'hbda4452f),
	.w3(32'hb8555524),
	.w4(32'hbd735e34),
	.w5(32'hbd749f28),
	.w6(32'h3c480cd6),
	.w7(32'hbda76e42),
	.w8(32'hbc186006),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07fe2),
	.w1(32'hbce94550),
	.w2(32'h3c53b5b4),
	.w3(32'hbc8576b2),
	.w4(32'hbd362f2b),
	.w5(32'h3beaee9e),
	.w6(32'hbc8f0332),
	.w7(32'hbd03bbe0),
	.w8(32'h3cb402e0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1c96a),
	.w1(32'h3c00e8fa),
	.w2(32'hbcf45d09),
	.w3(32'h3c8757b1),
	.w4(32'hba58aa84),
	.w5(32'hbc7435ce),
	.w6(32'hbcaa60c4),
	.w7(32'hbcf3a06a),
	.w8(32'hbc6162f8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf495b5),
	.w1(32'hbc5bd4f8),
	.w2(32'h3b832e57),
	.w3(32'hbb312995),
	.w4(32'hbbb86dbc),
	.w5(32'h3c09a133),
	.w6(32'h3b4beeec),
	.w7(32'hbb8e688f),
	.w8(32'h3c6d2392),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15f812),
	.w1(32'hbbc45776),
	.w2(32'h3c0ad06c),
	.w3(32'h3c405a7a),
	.w4(32'h3c0b4a54),
	.w5(32'h3c929eec),
	.w6(32'h3c3f6f97),
	.w7(32'h3b67568c),
	.w8(32'h3c52b5a4),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb871aea),
	.w1(32'h3b07dfc1),
	.w2(32'hbcc20591),
	.w3(32'h3b4f1691),
	.w4(32'h3b363960),
	.w5(32'hbce42310),
	.w6(32'hba882ce8),
	.w7(32'h3b865cda),
	.w8(32'hbbc35358),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31f7b5),
	.w1(32'h3a886dcc),
	.w2(32'hbbdf447a),
	.w3(32'hbd0a32c8),
	.w4(32'hbcaa7e06),
	.w5(32'hbc8d930d),
	.w6(32'hbcc9c2e9),
	.w7(32'hbc9bd012),
	.w8(32'hbcad03cf),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c0ee2),
	.w1(32'hbc24c07e),
	.w2(32'hbb37dc03),
	.w3(32'hbbdd1241),
	.w4(32'hbc0738c9),
	.w5(32'hbc67923b),
	.w6(32'hbb7787be),
	.w7(32'hbb74a56a),
	.w8(32'h39e78699),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6053a),
	.w1(32'hbc6babfd),
	.w2(32'h3c17d306),
	.w3(32'h3a016a16),
	.w4(32'hbb1226fe),
	.w5(32'h3c5693a4),
	.w6(32'hbc8dd0f9),
	.w7(32'h3be05b4f),
	.w8(32'h3b37612a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6af20f),
	.w1(32'hbc69e0dc),
	.w2(32'hbc3bd1eb),
	.w3(32'hbc8a997b),
	.w4(32'hbcf90b5e),
	.w5(32'hbc6b8379),
	.w6(32'h3c7dd1f7),
	.w7(32'hbcbe3289),
	.w8(32'hbb2554aa),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba18eb0),
	.w1(32'hbb333e57),
	.w2(32'h3c2b73c1),
	.w3(32'hbbfe661c),
	.w4(32'hbbba26be),
	.w5(32'h3d19c1fb),
	.w6(32'hbb52f1e8),
	.w7(32'hbbfd935f),
	.w8(32'h3d27aff1),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac7e7a),
	.w1(32'h3baeb1c6),
	.w2(32'h3bcf04b5),
	.w3(32'h3c9ddfec),
	.w4(32'hbab4802f),
	.w5(32'h3c362bc8),
	.w6(32'h3cb35154),
	.w7(32'h3be40c3e),
	.w8(32'h3c6c9ea8),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96bb7b7),
	.w1(32'h3c3bb447),
	.w2(32'h3aa97ce3),
	.w3(32'h3a9a14af),
	.w4(32'h3a12ea1c),
	.w5(32'hbb700f0e),
	.w6(32'h3c821a89),
	.w7(32'h3bff1a29),
	.w8(32'h3b8a4d1d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba867c5),
	.w1(32'hbce3d968),
	.w2(32'hbcf550f9),
	.w3(32'h3c3f3c15),
	.w4(32'hbd11de4e),
	.w5(32'hbc8c5430),
	.w6(32'h3bc7dba3),
	.w7(32'hbd706aab),
	.w8(32'hba0f34f4),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1e990),
	.w1(32'hbc1d8c2d),
	.w2(32'hbaf02b2e),
	.w3(32'hbbb8fb97),
	.w4(32'hbc57e944),
	.w5(32'h3bd66ce2),
	.w6(32'hbc6880fa),
	.w7(32'hbc6be389),
	.w8(32'h3c9a275c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c1a32),
	.w1(32'hbb8e237a),
	.w2(32'h38a1f49a),
	.w3(32'hbb4662c8),
	.w4(32'hbb3d3913),
	.w5(32'hbadb2a10),
	.w6(32'h3ba0ccbf),
	.w7(32'h3b081465),
	.w8(32'hbc19442b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe9348),
	.w1(32'hbcba0628),
	.w2(32'hbb8e5ae1),
	.w3(32'hbb850127),
	.w4(32'hbca3062b),
	.w5(32'hbb9cfb8d),
	.w6(32'hbbcecf29),
	.w7(32'hbc3962ec),
	.w8(32'hb9f4b8b7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13900f),
	.w1(32'hbc14880d),
	.w2(32'hbc167cb9),
	.w3(32'hbade17fc),
	.w4(32'hbc4f759b),
	.w5(32'hbc058415),
	.w6(32'hbb7c96ad),
	.w7(32'hbbc924a8),
	.w8(32'hba372350),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388922be),
	.w1(32'h3bf2679a),
	.w2(32'h3b457a22),
	.w3(32'hbc44b4cf),
	.w4(32'hbb198763),
	.w5(32'hbbd16335),
	.w6(32'hbc1a92e0),
	.w7(32'hbc026812),
	.w8(32'hbbcbf2cb),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35a7e3),
	.w1(32'hbbb60841),
	.w2(32'h3c36dad8),
	.w3(32'h3cd71ef8),
	.w4(32'hb92c913c),
	.w5(32'h3be7b83d),
	.w6(32'h3c192754),
	.w7(32'h3bbc16b4),
	.w8(32'hba205f2e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c0170),
	.w1(32'h3a93526a),
	.w2(32'h3bd3b99b),
	.w3(32'h3c920975),
	.w4(32'hbbef2918),
	.w5(32'hbb124475),
	.w6(32'h3c784de6),
	.w7(32'hb828bd9a),
	.w8(32'hbba9f3d7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0aa4ca),
	.w1(32'hbc542789),
	.w2(32'hbbd8b33f),
	.w3(32'h3bb9e46c),
	.w4(32'hbc6d3af1),
	.w5(32'h3ad650db),
	.w6(32'hbb436e77),
	.w7(32'hbc23a6af),
	.w8(32'hb96b0f42),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b7291),
	.w1(32'hbcbe2425),
	.w2(32'h3d25b651),
	.w3(32'h3c8db14c),
	.w4(32'hbcc430d4),
	.w5(32'h3d297726),
	.w6(32'h3be1a1da),
	.w7(32'hbd0bdb1a),
	.w8(32'h3ce6f566),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e8479),
	.w1(32'hbbf5279a),
	.w2(32'h3c4952d3),
	.w3(32'h3b5f2fc2),
	.w4(32'hbbc74447),
	.w5(32'h3b89eb4b),
	.w6(32'h3b48b1a0),
	.w7(32'hbc7119d6),
	.w8(32'h3c6618aa),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fda4d),
	.w1(32'hbc304a05),
	.w2(32'h3c898e2a),
	.w3(32'hbb4e4f4d),
	.w4(32'hbcc9fcc4),
	.w5(32'h3b6d7871),
	.w6(32'hbc96e5c4),
	.w7(32'hbd04811f),
	.w8(32'h3ba2b047),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35ceec),
	.w1(32'h3b9bdae0),
	.w2(32'hbba7722c),
	.w3(32'hbc090ccb),
	.w4(32'hbc72bf93),
	.w5(32'hbb774c60),
	.w6(32'hba60afc9),
	.w7(32'hbc7655ad),
	.w8(32'h3b4c6e57),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5ea6e),
	.w1(32'h3baae7fc),
	.w2(32'h3bf7dbf1),
	.w3(32'hbc719fad),
	.w4(32'hba577fb0),
	.w5(32'hbbdff0ad),
	.w6(32'hbb888b35),
	.w7(32'h3ad48708),
	.w8(32'hbc05d98f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27cc44),
	.w1(32'h3bc96a2b),
	.w2(32'hbb620f69),
	.w3(32'h3b24b5c4),
	.w4(32'h3ab75624),
	.w5(32'hbb439358),
	.w6(32'hbbbf2df2),
	.w7(32'hbbd52eb9),
	.w8(32'h3b61c80b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad35fec),
	.w1(32'h39136620),
	.w2(32'hbb8c2249),
	.w3(32'hbc13603d),
	.w4(32'hbbd5e48b),
	.w5(32'h3bc5ac71),
	.w6(32'h395a7f13),
	.w7(32'hb8b970b9),
	.w8(32'hbc3152f1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc394cf5),
	.w1(32'hbb6e5d36),
	.w2(32'h3d16c3c4),
	.w3(32'h3a82c83f),
	.w4(32'hbc5182f1),
	.w5(32'h3d24540e),
	.w6(32'h3be2e8b6),
	.w7(32'hbc1c161f),
	.w8(32'h3d079d9c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc50b0),
	.w1(32'h3c14924e),
	.w2(32'hbbc8c401),
	.w3(32'h3af3b519),
	.w4(32'hbaa31b13),
	.w5(32'h3bb19630),
	.w6(32'h3ca6469a),
	.w7(32'h3aec9a1f),
	.w8(32'hbb83bfac),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb387c4),
	.w1(32'hbbedcae2),
	.w2(32'hbb4bcf2a),
	.w3(32'hbb966510),
	.w4(32'h3ae56f17),
	.w5(32'h3b148fc7),
	.w6(32'hbba46498),
	.w7(32'h3bb3715e),
	.w8(32'h3a20d926),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc412a),
	.w1(32'h3b33412b),
	.w2(32'h3a911af8),
	.w3(32'h3b9d6d5e),
	.w4(32'h3bf89672),
	.w5(32'h3a001c67),
	.w6(32'h3be907a2),
	.w7(32'h3b96fa26),
	.w8(32'hba0d8b24),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c17cf),
	.w1(32'hba181635),
	.w2(32'hba942b96),
	.w3(32'h3b44b3d8),
	.w4(32'h3aaa2985),
	.w5(32'hbc72f866),
	.w6(32'h3ab5bf2c),
	.w7(32'h3baf3f79),
	.w8(32'hbca16e88),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc22b69),
	.w1(32'hbcceccea),
	.w2(32'hbaf26566),
	.w3(32'h3cc17906),
	.w4(32'hbb13eca1),
	.w5(32'h3a4908d3),
	.w6(32'hbc137d65),
	.w7(32'h3c6c8d48),
	.w8(32'hb99e76e0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba50cc6),
	.w1(32'hbb74c2c4),
	.w2(32'hbbd7714b),
	.w3(32'h3b30963f),
	.w4(32'h3aa47025),
	.w5(32'hbbbad193),
	.w6(32'h3b461bfd),
	.w7(32'h3b535c64),
	.w8(32'hbb736382),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4af092),
	.w1(32'hbcb64123),
	.w2(32'h3d6731cb),
	.w3(32'h3cb8bc78),
	.w4(32'hbb802e23),
	.w5(32'h3d798b64),
	.w6(32'h3c3e694d),
	.w7(32'h3c86637f),
	.w8(32'h3d60c254),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc297411),
	.w1(32'hbbfed070),
	.w2(32'hbb26e6ce),
	.w3(32'hbbb2f5b9),
	.w4(32'hbc90d312),
	.w5(32'h3b0cb35f),
	.w6(32'hbb5b753a),
	.w7(32'hbbea26a1),
	.w8(32'h3b344594),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80a5e5),
	.w1(32'hbc353727),
	.w2(32'h3be49c3f),
	.w3(32'h3cd44207),
	.w4(32'hbc0edaff),
	.w5(32'h3be9c5e2),
	.w6(32'h3d0bd1e7),
	.w7(32'h3c8d600f),
	.w8(32'h3c6ab584),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule