module layer_10_featuremap_476(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ae904),
	.w1(32'hbb0622ca),
	.w2(32'h38e7b378),
	.w3(32'hb9debafc),
	.w4(32'hbb92f7e2),
	.w5(32'hbb1a3773),
	.w6(32'hbb3faa2f),
	.w7(32'h3b47c6db),
	.w8(32'h3b549b8e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b23b2b),
	.w1(32'h39e37090),
	.w2(32'h3a55349d),
	.w3(32'hba0021a6),
	.w4(32'hbb3f03e7),
	.w5(32'hbb9cbfbf),
	.w6(32'h3b85cd14),
	.w7(32'hb91503d1),
	.w8(32'hbb4da4b8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5d1c3),
	.w1(32'h3ad846df),
	.w2(32'h3a8221d8),
	.w3(32'h3a030837),
	.w4(32'hba80d128),
	.w5(32'hba03fc34),
	.w6(32'hbad15c39),
	.w7(32'h3a222943),
	.w8(32'hba4341af),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fc29f),
	.w1(32'h38ce5008),
	.w2(32'h3ad0db6f),
	.w3(32'hba8e63fc),
	.w4(32'hbb8bc955),
	.w5(32'hbaf41d64),
	.w6(32'hb90cd4c2),
	.w7(32'hbb5e2c27),
	.w8(32'h3b04e7f9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6b62f),
	.w1(32'hbaa4cc9c),
	.w2(32'hba9215b1),
	.w3(32'h3b9e5628),
	.w4(32'h3b34cd6e),
	.w5(32'hbac5364d),
	.w6(32'h3b9500b2),
	.w7(32'h3995489e),
	.w8(32'h3b03d20e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9fbbc),
	.w1(32'h39267b3a),
	.w2(32'h3990a006),
	.w3(32'hbb177679),
	.w4(32'h3ba83347),
	.w5(32'h3ae7cc6f),
	.w6(32'h3b61583b),
	.w7(32'hb94ac2c1),
	.w8(32'hbb425ee2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a44ed),
	.w1(32'h3a0a686e),
	.w2(32'hbb038f09),
	.w3(32'h3a7eab6c),
	.w4(32'hba0a2aac),
	.w5(32'hbb173b45),
	.w6(32'hbb3a89bc),
	.w7(32'hbb077789),
	.w8(32'h390d6d91),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6baae),
	.w1(32'hbb03d0d4),
	.w2(32'h3b078212),
	.w3(32'hbb720a9d),
	.w4(32'hbbbe0b17),
	.w5(32'hbb9b49fb),
	.w6(32'hbae0fba9),
	.w7(32'hba8217d2),
	.w8(32'hbb15be3a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27069e),
	.w1(32'hba1dbc2d),
	.w2(32'h3b03c6bb),
	.w3(32'hbbccca63),
	.w4(32'h3aa87716),
	.w5(32'h3b3d6860),
	.w6(32'hbbbf83ab),
	.w7(32'hb80172e2),
	.w8(32'hbb6975c1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e0bdf),
	.w1(32'hbb88b361),
	.w2(32'hbb18e510),
	.w3(32'h3bbc70c6),
	.w4(32'h3a52f415),
	.w5(32'h3b8c07b2),
	.w6(32'h3acdb849),
	.w7(32'hba65bc1e),
	.w8(32'h3ae88b68),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978a02),
	.w1(32'hbb533b11),
	.w2(32'hba8e2a5f),
	.w3(32'h3b52492c),
	.w4(32'h3c30be80),
	.w5(32'h3c801484),
	.w6(32'hba45f155),
	.w7(32'hbb68d0c4),
	.w8(32'hba6bfb9d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a1aff),
	.w1(32'hb9e92017),
	.w2(32'h398c77db),
	.w3(32'h3c081857),
	.w4(32'h3b426034),
	.w5(32'h3addac1e),
	.w6(32'h3a50a617),
	.w7(32'h3b8475c0),
	.w8(32'h390ba915),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83656a),
	.w1(32'hb9ae9792),
	.w2(32'h3ae649a1),
	.w3(32'hbac0ab94),
	.w4(32'hbb0f3054),
	.w5(32'hbacf387a),
	.w6(32'hba31500f),
	.w7(32'hb82f277a),
	.w8(32'h3a1b86f7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb754172),
	.w1(32'hba2f05d1),
	.w2(32'hb9105706),
	.w3(32'h3b2b3da5),
	.w4(32'h3bcc8d6d),
	.w5(32'h3b5dfaea),
	.w6(32'h3b0e6d08),
	.w7(32'h3b5a3470),
	.w8(32'h3c0c47fe),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd1385),
	.w1(32'hba68c7b0),
	.w2(32'hba1d99dc),
	.w3(32'h39891ea1),
	.w4(32'h3b94e67e),
	.w5(32'h3b626527),
	.w6(32'h3c1e5afd),
	.w7(32'h3987beee),
	.w8(32'hbb3f27e6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0980b6),
	.w1(32'hba8e73b6),
	.w2(32'hba833e16),
	.w3(32'h3a59704d),
	.w4(32'h3904b65b),
	.w5(32'h3ac651fa),
	.w6(32'hbb1b9fd1),
	.w7(32'h3b605198),
	.w8(32'h3b0cbf69),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07e476),
	.w1(32'h3b88012a),
	.w2(32'h3b3573b8),
	.w3(32'h3a81bf89),
	.w4(32'h3a45c89b),
	.w5(32'hb6c5b03d),
	.w6(32'h3a71b3ef),
	.w7(32'hbac901ef),
	.w8(32'hbb3e4327),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba636fba),
	.w1(32'h3b1a6ff3),
	.w2(32'h39eb99bf),
	.w3(32'hba0ecce9),
	.w4(32'hbb52a39a),
	.w5(32'hb98b2b78),
	.w6(32'hbb9a85f9),
	.w7(32'hbb1e4eae),
	.w8(32'hbb7b2b38),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af132b5),
	.w1(32'hbb20a575),
	.w2(32'hb94ae840),
	.w3(32'h39903d31),
	.w4(32'h3aa0ef48),
	.w5(32'hba7f9498),
	.w6(32'hbae90286),
	.w7(32'hba5e04ff),
	.w8(32'hbb96c0dc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0caa8e),
	.w1(32'h3a95f446),
	.w2(32'hbb9ba844),
	.w3(32'hb8af5edb),
	.w4(32'hba7949ec),
	.w5(32'h3ab9c2d4),
	.w6(32'hbacf74ac),
	.w7(32'hbacc3aff),
	.w8(32'hbac9adf4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e57dd),
	.w1(32'h3aff6948),
	.w2(32'hbb0d947e),
	.w3(32'h3b16b0c9),
	.w4(32'h3b8e40b8),
	.w5(32'h3a7c5212),
	.w6(32'hbaa5fb75),
	.w7(32'h3adef31b),
	.w8(32'hba185cf3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb81e0),
	.w1(32'hb94ef7ca),
	.w2(32'h3a3e1d88),
	.w3(32'hbaa2bd94),
	.w4(32'hbb34f88c),
	.w5(32'h39577ec1),
	.w6(32'h3793a422),
	.w7(32'hbadd1ccf),
	.w8(32'hbb753589),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d5876),
	.w1(32'h3b1c6f2e),
	.w2(32'h3b136d75),
	.w3(32'h3b5fd831),
	.w4(32'h3b84a170),
	.w5(32'h3bbb823a),
	.w6(32'h3ade05d0),
	.w7(32'h3adb1a94),
	.w8(32'h3955e4fe),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28ea56),
	.w1(32'h3abb4f60),
	.w2(32'hba506e6f),
	.w3(32'h3bbbad15),
	.w4(32'hb93b673a),
	.w5(32'hbb219698),
	.w6(32'hbb081b84),
	.w7(32'h39b7b4f7),
	.w8(32'hbb221a54),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfe395),
	.w1(32'h3a578101),
	.w2(32'h39be86c3),
	.w3(32'hb8f8b4cb),
	.w4(32'h3b8b7cb2),
	.w5(32'h3b3fa933),
	.w6(32'h3979323f),
	.w7(32'h3b0ddeb3),
	.w8(32'hbabbe675),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf2e69),
	.w1(32'h3b887f1f),
	.w2(32'h3af250bc),
	.w3(32'h3a8a4b7d),
	.w4(32'h3a8831df),
	.w5(32'hbaf33ec6),
	.w6(32'h3a2af686),
	.w7(32'hbbb0af6a),
	.w8(32'hbaeca679),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38040eb4),
	.w1(32'hba9e35d1),
	.w2(32'hbb4803d3),
	.w3(32'hbb85f549),
	.w4(32'hbabc98cb),
	.w5(32'hbb2cfcbf),
	.w6(32'hbb32b197),
	.w7(32'hbb21d3b9),
	.w8(32'hbb366996),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44077d),
	.w1(32'hb9dfff6b),
	.w2(32'hb99c86d3),
	.w3(32'hbb16d73d),
	.w4(32'h3a88b395),
	.w5(32'hba212445),
	.w6(32'hbb3a25d1),
	.w7(32'hbb1080e5),
	.w8(32'hbb32ab85),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993f2ce),
	.w1(32'hbb440b53),
	.w2(32'hbb6bbd6a),
	.w3(32'hbb0ddbfb),
	.w4(32'hb9901529),
	.w5(32'hbb4a0ee9),
	.w6(32'hbaec082a),
	.w7(32'hbabb8583),
	.w8(32'hbae0b568),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c8b10),
	.w1(32'h3ab627aa),
	.w2(32'hba547b7e),
	.w3(32'h3b69fb40),
	.w4(32'h3b7f01af),
	.w5(32'h39a434a4),
	.w6(32'h3aab3dd6),
	.w7(32'h39bd3e4e),
	.w8(32'hba19853b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0f66),
	.w1(32'hb8fa1eb1),
	.w2(32'hbaf81086),
	.w3(32'hb9998a96),
	.w4(32'h3ac88d08),
	.w5(32'h3b87bd53),
	.w6(32'hbb72ddf7),
	.w7(32'h3a3bb4d6),
	.w8(32'h39dddb6f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383faee4),
	.w1(32'hb74a884d),
	.w2(32'h3adc30ad),
	.w3(32'h3b24e1de),
	.w4(32'h3af5d300),
	.w5(32'hba0c41c9),
	.w6(32'hb953c783),
	.w7(32'hba858be2),
	.w8(32'h39abcd3d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab26571),
	.w1(32'h3ab2b514),
	.w2(32'h3a1f96cf),
	.w3(32'h3ae6ad58),
	.w4(32'hba8c151c),
	.w5(32'h384b7f2b),
	.w6(32'hb970072e),
	.w7(32'h3b6d9370),
	.w8(32'h3b8d0809),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeefd55),
	.w1(32'h39b8c178),
	.w2(32'h3a69ada1),
	.w3(32'hba9e2b4b),
	.w4(32'hbacebb11),
	.w5(32'hba348157),
	.w6(32'h39eb8821),
	.w7(32'hbb19b484),
	.w8(32'h3702e7d0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54a464),
	.w1(32'hbb2685d7),
	.w2(32'hbace40ec),
	.w3(32'hbb897c0e),
	.w4(32'hbbb1aef7),
	.w5(32'hbb8c50d5),
	.w6(32'hbb106f5b),
	.w7(32'h38ec6ea2),
	.w8(32'h3b35ead9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e811d),
	.w1(32'hb9b9252b),
	.w2(32'h389440b5),
	.w3(32'hbb8a6184),
	.w4(32'hba2d381e),
	.w5(32'h3acc2fac),
	.w6(32'h3b117fcc),
	.w7(32'h3a9d5ae6),
	.w8(32'h3b554c25),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66975f),
	.w1(32'hba487113),
	.w2(32'h3abac1b6),
	.w3(32'h3b5bdf5a),
	.w4(32'h3bce8258),
	.w5(32'h3bddb8ff),
	.w6(32'h3b92f7a1),
	.w7(32'hbaf802b1),
	.w8(32'h3990e718),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba269f6b),
	.w1(32'hbad337fa),
	.w2(32'h3aa2cde0),
	.w3(32'h3b145f32),
	.w4(32'hba852875),
	.w5(32'hbaebea53),
	.w6(32'h39fc9eb9),
	.w7(32'hbabcf7c2),
	.w8(32'hb8fd6a2a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381e4ca6),
	.w1(32'hbb8b0eab),
	.w2(32'hbb224d4f),
	.w3(32'h3a943cd8),
	.w4(32'h3bbe9c6b),
	.w5(32'h3adca4d5),
	.w6(32'hbb41b939),
	.w7(32'h3ab5a71f),
	.w8(32'hbb1121d8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc856),
	.w1(32'h3977ffca),
	.w2(32'h3b40f8d5),
	.w3(32'h3b1c8f66),
	.w4(32'hbb49757b),
	.w5(32'hbabf35df),
	.w6(32'h3a634ebe),
	.w7(32'hbb81cdaa),
	.w8(32'hbab973c7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a982f6d),
	.w1(32'hba54b06b),
	.w2(32'hb9339c5c),
	.w3(32'h3a3b41aa),
	.w4(32'hbb6f2271),
	.w5(32'hbbcea4d8),
	.w6(32'hbb23cb1b),
	.w7(32'h3b211240),
	.w8(32'h3b78543e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8583b8),
	.w1(32'hba90a87a),
	.w2(32'hba8241c8),
	.w3(32'hbbc48b29),
	.w4(32'h3b07f44c),
	.w5(32'hbafa907e),
	.w6(32'h3b20b913),
	.w7(32'hba923a75),
	.w8(32'hbba8e827),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a84e98),
	.w1(32'h39506a47),
	.w2(32'hba5899db),
	.w3(32'hbb767a28),
	.w4(32'hbb098793),
	.w5(32'hbb4f68c9),
	.w6(32'hbb1946d6),
	.w7(32'hbb1aa100),
	.w8(32'hbac52a54),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb05220),
	.w1(32'hb9d57f04),
	.w2(32'h3b3e2d9c),
	.w3(32'h3bb12b29),
	.w4(32'hb9354d17),
	.w5(32'h3ac548dc),
	.w6(32'h38ffbdc3),
	.w7(32'hba928029),
	.w8(32'hb7f38657),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07d434),
	.w1(32'h3a327731),
	.w2(32'hba8cf08e),
	.w3(32'h3ab8ee61),
	.w4(32'hba35d70e),
	.w5(32'hba849dbd),
	.w6(32'hba22bfeb),
	.w7(32'h3b113a2c),
	.w8(32'h3aa92178),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab55f66),
	.w1(32'hba739ab1),
	.w2(32'hbba4af4d),
	.w3(32'hbaa24924),
	.w4(32'h3aa607f5),
	.w5(32'h3aca6fbe),
	.w6(32'h3aa7d718),
	.w7(32'h3bbd343f),
	.w8(32'h3b77b81c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8459e6),
	.w1(32'hbaaf2feb),
	.w2(32'h3b0f7f27),
	.w3(32'h3b4a1125),
	.w4(32'h3c05c8ef),
	.w5(32'h3be50d41),
	.w6(32'h3b28acb8),
	.w7(32'h3aa85aaf),
	.w8(32'h39ed8935),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6705e),
	.w1(32'hba81a7ae),
	.w2(32'hba47093c),
	.w3(32'h3c0de201),
	.w4(32'hbb022b36),
	.w5(32'hbb05e4b0),
	.w6(32'h3b248cb6),
	.w7(32'hba62bd3f),
	.w8(32'hbac60ad1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0143c0),
	.w1(32'hbadfa59d),
	.w2(32'hbb5ae00b),
	.w3(32'h3b07efc4),
	.w4(32'h3b10473d),
	.w5(32'hb9f63952),
	.w6(32'h3b45aa13),
	.w7(32'h3ba14c34),
	.w8(32'h3b06004e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb400427),
	.w1(32'h39ee6b7c),
	.w2(32'hba42e641),
	.w3(32'hbb5a4dcf),
	.w4(32'h3b93f7d3),
	.w5(32'h3b6b19bb),
	.w6(32'hbaa53a3c),
	.w7(32'h3b344368),
	.w8(32'h3b142b87),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bb2fd),
	.w1(32'hbb06e126),
	.w2(32'hbaf20362),
	.w3(32'hbaf9c1c5),
	.w4(32'hb9d99661),
	.w5(32'hbb2df0e3),
	.w6(32'hb8dae5a7),
	.w7(32'h3b2fb95e),
	.w8(32'hb9ec57c3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1c2fc),
	.w1(32'hba66cbcb),
	.w2(32'hbae5f61b),
	.w3(32'hba2c9276),
	.w4(32'hb9dc8a53),
	.w5(32'h3a9145b7),
	.w6(32'h3b642d0d),
	.w7(32'hb9a67387),
	.w8(32'hbae5940f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a786b0),
	.w1(32'h378d6095),
	.w2(32'h3ab7a8e8),
	.w3(32'h3b3f66f3),
	.w4(32'hbb028353),
	.w5(32'hba2ba9de),
	.w6(32'h3ad38d83),
	.w7(32'h39608361),
	.w8(32'h3954df61),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b8796),
	.w1(32'h3983f6e1),
	.w2(32'hb9ed881e),
	.w3(32'hbb3f88dd),
	.w4(32'hbb7e03f6),
	.w5(32'hbadbe605),
	.w6(32'hbb2f8a7f),
	.w7(32'h3a8ef396),
	.w8(32'h3a88795f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa2a66),
	.w1(32'hba10904b),
	.w2(32'h3b155ecd),
	.w3(32'hbb3b820d),
	.w4(32'hbb51be22),
	.w5(32'hba1c476b),
	.w6(32'hbaed42b7),
	.w7(32'hbb63590b),
	.w8(32'hb9f72e39),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42cda5),
	.w1(32'h3b03c37b),
	.w2(32'hb9d7b5d3),
	.w3(32'h3885e22c),
	.w4(32'h3aa743db),
	.w5(32'hb9310424),
	.w6(32'hbb8679a5),
	.w7(32'h3abf9621),
	.w8(32'h392ff636),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aec31),
	.w1(32'hbaa2a5b3),
	.w2(32'hbaad537c),
	.w3(32'h3b368e04),
	.w4(32'h3a72b6ac),
	.w5(32'hbaf3243c),
	.w6(32'hba0f1657),
	.w7(32'hb9fa8187),
	.w8(32'hbac5ab06),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb987a27),
	.w1(32'h3ac60786),
	.w2(32'hb97fafff),
	.w3(32'hba93fe36),
	.w4(32'h3b762d06),
	.w5(32'h3acd53ad),
	.w6(32'h3a70f008),
	.w7(32'hbb2bb173),
	.w8(32'hba5e7964),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26ce3b),
	.w1(32'hbb626ad2),
	.w2(32'hbb4db7d4),
	.w3(32'h3b066ab5),
	.w4(32'hbbb7bfdf),
	.w5(32'hbbad2f33),
	.w6(32'hba1a12e7),
	.w7(32'hbb7b3d26),
	.w8(32'hbba49572),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7347c4),
	.w1(32'h3bb50063),
	.w2(32'h3ba4fdb5),
	.w3(32'hbb6bba19),
	.w4(32'h3b03999b),
	.w5(32'hba2c6252),
	.w6(32'hbb976979),
	.w7(32'h39ed45bc),
	.w8(32'hba417fe9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c2486),
	.w1(32'h3bdaf720),
	.w2(32'h3b96d9fe),
	.w3(32'h3ac6d41c),
	.w4(32'hb9e26795),
	.w5(32'h3af3d48b),
	.w6(32'hba728bce),
	.w7(32'hbb873220),
	.w8(32'hbb377281),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e748a),
	.w1(32'hbb95c1ee),
	.w2(32'hbb725d96),
	.w3(32'h3a5e5eb4),
	.w4(32'h3b8a56d2),
	.w5(32'h3ab82df9),
	.w6(32'hbb39e15a),
	.w7(32'hba68dfd4),
	.w8(32'hbb6cf759),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcb47e),
	.w1(32'h3a563169),
	.w2(32'hbb163dff),
	.w3(32'hba97ad0c),
	.w4(32'hbb6a1634),
	.w5(32'hbbc9108d),
	.w6(32'hbb19d661),
	.w7(32'hbb8bbf18),
	.w8(32'hbbb1090e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb779d8e),
	.w1(32'hb9ef8a6f),
	.w2(32'hbb26496a),
	.w3(32'h3ace16f8),
	.w4(32'h3a4faae0),
	.w5(32'hbac03c1c),
	.w6(32'hba9e394e),
	.w7(32'h3b355afc),
	.w8(32'h3b1a3596),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04c879),
	.w1(32'h3b116e07),
	.w2(32'h3ace7095),
	.w3(32'hbb5346ce),
	.w4(32'h3a07963a),
	.w5(32'h392e5555),
	.w6(32'h3b13726f),
	.w7(32'h38c5920d),
	.w8(32'hb839cebe),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa9092),
	.w1(32'hbb6737a7),
	.w2(32'hbb10092c),
	.w3(32'h3b2ee3fd),
	.w4(32'h3bb718df),
	.w5(32'hb934aa45),
	.w6(32'h3abda0ea),
	.w7(32'h3a97e764),
	.w8(32'hbb732bd5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87f5ab),
	.w1(32'h395dab21),
	.w2(32'hb9e20bf4),
	.w3(32'hbb12cdaf),
	.w4(32'hbb156169),
	.w5(32'hbacaa0c9),
	.w6(32'hbb8215dc),
	.w7(32'hb975cae3),
	.w8(32'hb9c9884c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e6de0),
	.w1(32'h3ba60f0c),
	.w2(32'h3b3d356f),
	.w3(32'h3ae05fbb),
	.w4(32'h3a3c0138),
	.w5(32'hbb7b1c39),
	.w6(32'h3ae0d620),
	.w7(32'h3a662553),
	.w8(32'hbbc05870),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9991513),
	.w1(32'h3a2d6216),
	.w2(32'h3a8e7f4b),
	.w3(32'hbba8c4d0),
	.w4(32'hb95d856d),
	.w5(32'hba92f15d),
	.w6(32'hbb4fba1b),
	.w7(32'hb8ad73fb),
	.w8(32'hbaa647d8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebaa79),
	.w1(32'hbb871729),
	.w2(32'hbbb20fa8),
	.w3(32'h3a5f2fd3),
	.w4(32'hbc154480),
	.w5(32'hbaeb71f4),
	.w6(32'hb9ecb0e8),
	.w7(32'hbbe0ec14),
	.w8(32'h3b9de93f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69896e),
	.w1(32'hbb704a0e),
	.w2(32'h3b560012),
	.w3(32'hbb90b913),
	.w4(32'h3bba9252),
	.w5(32'h3c45f77a),
	.w6(32'hbb8b30a5),
	.w7(32'hbb4b663f),
	.w8(32'h38a43e14),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394824e0),
	.w1(32'h3b824386),
	.w2(32'hbb90fead),
	.w3(32'hb9f3a818),
	.w4(32'hbaac37c6),
	.w5(32'h3c430545),
	.w6(32'hbb8cdfe8),
	.w7(32'hb98193a5),
	.w8(32'hbbefc580),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc082392),
	.w1(32'hbb39867f),
	.w2(32'h3afee84b),
	.w3(32'hbbe92168),
	.w4(32'h3af2f362),
	.w5(32'h3bfd1bb8),
	.w6(32'hbbce54b9),
	.w7(32'h3ab3fb3a),
	.w8(32'h3b1e049a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b980644),
	.w1(32'h3961f6ea),
	.w2(32'hb9b4c391),
	.w3(32'h3a0a1a8b),
	.w4(32'hbba2a11a),
	.w5(32'h3b92545b),
	.w6(32'hbb39eba8),
	.w7(32'hbb2c33a1),
	.w8(32'hbabba3a2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb891f4e8),
	.w1(32'h3b3fc1a8),
	.w2(32'hba6d5116),
	.w3(32'hbb367a3d),
	.w4(32'h3bafdb2e),
	.w5(32'h3b113e99),
	.w6(32'h3b2bb58c),
	.w7(32'h3bd8efc1),
	.w8(32'h3a919539),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd4783),
	.w1(32'h3b6cc6ab),
	.w2(32'h3b77fe96),
	.w3(32'h3b710364),
	.w4(32'hbbfb5d6c),
	.w5(32'hbbf739f2),
	.w6(32'h3aef2b47),
	.w7(32'hbbb466a7),
	.w8(32'hbba7ce71),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ff2df),
	.w1(32'hba3f3191),
	.w2(32'hba7a5c3d),
	.w3(32'hba6f6b59),
	.w4(32'hbb5ddf53),
	.w5(32'hbbf09db9),
	.w6(32'h3b882433),
	.w7(32'hbb1911bb),
	.w8(32'hbbcbae8e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2e7a9),
	.w1(32'h3a530596),
	.w2(32'hbb94a369),
	.w3(32'hbc1f771e),
	.w4(32'h39eaa8de),
	.w5(32'hbb9250f0),
	.w6(32'hbb99c7a1),
	.w7(32'h3b1aca4c),
	.w8(32'h38a4a33c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbb9ff),
	.w1(32'hbb2e9f8f),
	.w2(32'hbbb1c899),
	.w3(32'hbb980b11),
	.w4(32'hbb8e145e),
	.w5(32'hbbca1dd1),
	.w6(32'hbb5c67a7),
	.w7(32'hbb58fc10),
	.w8(32'hbb4c2ebf),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00cf4d),
	.w1(32'hba845751),
	.w2(32'h3b26d3fa),
	.w3(32'hbb16fbf5),
	.w4(32'h3b2d237f),
	.w5(32'h3b6a394d),
	.w6(32'h3a29608d),
	.w7(32'hbbb5cf2c),
	.w8(32'h3b14a375),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5040be),
	.w1(32'h3b9afc73),
	.w2(32'h3c57160c),
	.w3(32'h3be4957b),
	.w4(32'h3b92ba9f),
	.w5(32'h3bacdf1d),
	.w6(32'h3a8be1da),
	.w7(32'h3badfc61),
	.w8(32'h3b041ffb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bba10),
	.w1(32'hbb041780),
	.w2(32'h3be3cd73),
	.w3(32'h3c071132),
	.w4(32'h3b821466),
	.w5(32'h3c082386),
	.w6(32'h3ae8e344),
	.w7(32'h3b1d41db),
	.w8(32'hba808870),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6aeac),
	.w1(32'h3b9cf5c3),
	.w2(32'h3bc1ca48),
	.w3(32'hbb2d4e3b),
	.w4(32'h3bcea043),
	.w5(32'h3c7c5f5a),
	.w6(32'hbbf447d4),
	.w7(32'h3bed90c9),
	.w8(32'h3b0ff0fb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c167454),
	.w1(32'hbba5ed50),
	.w2(32'h3a30fa84),
	.w3(32'h3c028d3c),
	.w4(32'hba9b9f2f),
	.w5(32'h3ccff2ee),
	.w6(32'h3b03140c),
	.w7(32'h3bd48ef7),
	.w8(32'h3c7169da),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f6f07),
	.w1(32'h3729d9e9),
	.w2(32'hbbb59b5b),
	.w3(32'h3c8993de),
	.w4(32'hba6a8992),
	.w5(32'hbc171165),
	.w6(32'hbae14b0a),
	.w7(32'h3a1a2ac5),
	.w8(32'hbb094b11),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba08645),
	.w1(32'h3af4476e),
	.w2(32'h3b862b58),
	.w3(32'hbaf64af8),
	.w4(32'hbaba7772),
	.w5(32'h3c8b881d),
	.w6(32'hbb33d731),
	.w7(32'h3bc7be39),
	.w8(32'h3a490fb8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78e51f),
	.w1(32'h3b34d2b2),
	.w2(32'hbbad33d6),
	.w3(32'h3bb9d063),
	.w4(32'h3b1252d7),
	.w5(32'hbc35584f),
	.w6(32'h3c04dfec),
	.w7(32'h381fb969),
	.w8(32'hbb17eda4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba850e78),
	.w1(32'h3b3e6f6d),
	.w2(32'hbba4977d),
	.w3(32'hbbc6d60f),
	.w4(32'h3bb62a9d),
	.w5(32'h3b935483),
	.w6(32'hbb735803),
	.w7(32'h3bae42a7),
	.w8(32'h3b5b8a29),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b435276),
	.w1(32'hb81b20bd),
	.w2(32'hbbd78ac5),
	.w3(32'h39111c8c),
	.w4(32'hbb651899),
	.w5(32'hbbde1c60),
	.w6(32'hbb57fadd),
	.w7(32'hbba4bfbd),
	.w8(32'h3b9f16a4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb874a),
	.w1(32'h3a252a0a),
	.w2(32'hbb2a62b9),
	.w3(32'h3c312fa5),
	.w4(32'hba8bdee8),
	.w5(32'hbbf18161),
	.w6(32'h38b9257c),
	.w7(32'hbb36d42c),
	.w8(32'hbba242f4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e98b0),
	.w1(32'h3b45e9fe),
	.w2(32'hbb8b69bf),
	.w3(32'hb9e24541),
	.w4(32'hbb74aa24),
	.w5(32'hbbf876af),
	.w6(32'h3b40c2fb),
	.w7(32'hbbc564e4),
	.w8(32'hba1f43c6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb821d703),
	.w1(32'hbc16e860),
	.w2(32'hbc194731),
	.w3(32'h390c631d),
	.w4(32'h3c0042d6),
	.w5(32'h3bc768ae),
	.w6(32'hbb92bd07),
	.w7(32'hbaea8500),
	.w8(32'hbb0b233d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e4002),
	.w1(32'h3ae2c5cd),
	.w2(32'hbab9cb27),
	.w3(32'h3b557ebe),
	.w4(32'hbb0c9996),
	.w5(32'hbb581693),
	.w6(32'h3b043146),
	.w7(32'hbb2a0f38),
	.w8(32'h39bad723),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26a729),
	.w1(32'hbaf9b7b5),
	.w2(32'hbb0070c0),
	.w3(32'h3a182a3d),
	.w4(32'hbc174133),
	.w5(32'hbbcad4ca),
	.w6(32'h3bf459a0),
	.w7(32'hba954e1f),
	.w8(32'h3b277654),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02ff44),
	.w1(32'hbbb653a9),
	.w2(32'hbb500eb9),
	.w3(32'hbb74bd32),
	.w4(32'hb8ac5af8),
	.w5(32'h3bcc89f7),
	.w6(32'h3bae1db6),
	.w7(32'h3aaf5b2e),
	.w8(32'hbb9abc19),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7a08d),
	.w1(32'h3b2ab95e),
	.w2(32'h3ba95e50),
	.w3(32'h3c800dbe),
	.w4(32'h3b0c42bd),
	.w5(32'h3c9c1196),
	.w6(32'hbb381a22),
	.w7(32'h3b8e9dae),
	.w8(32'h3b4cf3b2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87e2b8),
	.w1(32'h3bec9c09),
	.w2(32'h3bcc5d8a),
	.w3(32'hba83ced0),
	.w4(32'h3b0a833f),
	.w5(32'h3c4c39a5),
	.w6(32'hbb1328bc),
	.w7(32'hba85282e),
	.w8(32'hbb86e93d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9834d6d),
	.w1(32'hbb82dbff),
	.w2(32'h3b0cb6c7),
	.w3(32'hbbbe33d7),
	.w4(32'hbbc1ef6a),
	.w5(32'hbb49fa1f),
	.w6(32'hbc183bd1),
	.w7(32'hb8a289be),
	.w8(32'h3b3a9537),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd77fd),
	.w1(32'hbb628d96),
	.w2(32'hbc1f5045),
	.w3(32'h3c0c8581),
	.w4(32'hbb8ce163),
	.w5(32'hbb5be839),
	.w6(32'h3be7600b),
	.w7(32'hbb55bcde),
	.w8(32'hba953e38),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819d5f),
	.w1(32'hb9fab2bd),
	.w2(32'hbba0954b),
	.w3(32'h3b29054c),
	.w4(32'h3b4ef7cb),
	.w5(32'hbb6b2c19),
	.w6(32'hbb766722),
	.w7(32'hba16981f),
	.w8(32'h3b057fe9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ab889),
	.w1(32'h3b1ad66a),
	.w2(32'h3aa8fb9b),
	.w3(32'h3baeac00),
	.w4(32'hbc073df3),
	.w5(32'hbb9a0b0f),
	.w6(32'h3b5237d9),
	.w7(32'hbafe0809),
	.w8(32'hbbafe8a2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08c7e1),
	.w1(32'h3b8e45e4),
	.w2(32'h3b6563f7),
	.w3(32'hbbd3aeba),
	.w4(32'h3b4707da),
	.w5(32'hbab0b20f),
	.w6(32'hbbb24b8b),
	.w7(32'hba8ece0d),
	.w8(32'hbb275a4a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b756c6),
	.w1(32'hbbb3636f),
	.w2(32'hbba4ef2d),
	.w3(32'h3a6fccfd),
	.w4(32'hbb02a2aa),
	.w5(32'h3d1f73fb),
	.w6(32'h3a84c337),
	.w7(32'h3bdb220e),
	.w8(32'hbb333f00),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a556bb4),
	.w1(32'hbb4bba7c),
	.w2(32'hbbe386c8),
	.w3(32'h3bebce22),
	.w4(32'hba423b32),
	.w5(32'hbc0e8160),
	.w6(32'hbc758645),
	.w7(32'h3b11997b),
	.w8(32'hbbb905ac),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12e5b7),
	.w1(32'h3bc18692),
	.w2(32'h3bbf8228),
	.w3(32'h3b2b2302),
	.w4(32'h3b61df32),
	.w5(32'h3ac9b950),
	.w6(32'h3a0c2cff),
	.w7(32'h3aec7981),
	.w8(32'hbb424eca),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac78da1),
	.w1(32'h3b604834),
	.w2(32'h3b536dea),
	.w3(32'hbb8e707a),
	.w4(32'h3b7dcbd4),
	.w5(32'h3bb6c547),
	.w6(32'h3b0e7efd),
	.w7(32'h3bdfe793),
	.w8(32'h3b82b1c1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2cb55),
	.w1(32'h3b876291),
	.w2(32'h3c2c594a),
	.w3(32'h3a69aa1f),
	.w4(32'h3c156097),
	.w5(32'h3bd23af7),
	.w6(32'hbafe23af),
	.w7(32'h3a57d7e8),
	.w8(32'hb9f4e3ed),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b566027),
	.w1(32'h3bf707c8),
	.w2(32'hbbd773d6),
	.w3(32'hbade1165),
	.w4(32'h3b7873c7),
	.w5(32'hbb897950),
	.w6(32'hbbb29803),
	.w7(32'hba168dea),
	.w8(32'hbb94a7b7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1673a),
	.w1(32'h3b3e60b0),
	.w2(32'h3ad2ae2e),
	.w3(32'hbbdce8cb),
	.w4(32'hbaaddaf5),
	.w5(32'hbb2e82fc),
	.w6(32'hbae32a00),
	.w7(32'h39dd2d45),
	.w8(32'hbbb2ea7b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3aeb81),
	.w1(32'h3b9e1127),
	.w2(32'h3bfe7a22),
	.w3(32'h3b00a7d2),
	.w4(32'h3b6cbb12),
	.w5(32'hbc6a2fff),
	.w6(32'h39e5c802),
	.w7(32'h3bbf61f6),
	.w8(32'h3b99b1cf),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50f5f3),
	.w1(32'hb8a101b4),
	.w2(32'h3b52b3f8),
	.w3(32'hbbe4965c),
	.w4(32'hba12643d),
	.w5(32'h39954e2a),
	.w6(32'h3b651a48),
	.w7(32'hbbe277ec),
	.w8(32'hbb660a1b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa45c32),
	.w1(32'h3ab805a0),
	.w2(32'h3b2183b9),
	.w3(32'h3b45c919),
	.w4(32'h3a8d9507),
	.w5(32'h3bdd8363),
	.w6(32'h3c0bf34e),
	.w7(32'h3bf22d8b),
	.w8(32'hbae4c052),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8115628),
	.w1(32'h3b098a1d),
	.w2(32'h3c8c2f9d),
	.w3(32'hba959ca3),
	.w4(32'h3c0a6ca1),
	.w5(32'h3ce97b8c),
	.w6(32'hbbccdcc3),
	.w7(32'h3bc4e8c3),
	.w8(32'h3c0c7e50),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62e333),
	.w1(32'h3c7f7613),
	.w2(32'h3c29688d),
	.w3(32'h3c4ea275),
	.w4(32'h3bc039a1),
	.w5(32'hbc3ca03a),
	.w6(32'h3b45332f),
	.w7(32'hbb8ff684),
	.w8(32'hbc3f8fae),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30889b),
	.w1(32'hbbeb0d90),
	.w2(32'hbc0c6c7c),
	.w3(32'hbc6ccd8a),
	.w4(32'hbc3e45ae),
	.w5(32'hba8c79bd),
	.w6(32'hbb368b0a),
	.w7(32'hbbc8ea6b),
	.w8(32'hbb940278),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2154db),
	.w1(32'h3ba1e4c1),
	.w2(32'h395518a6),
	.w3(32'hbb1a1023),
	.w4(32'h3bf443ae),
	.w5(32'hbbb2e7d0),
	.w6(32'h3b482c8d),
	.w7(32'hbac5200c),
	.w8(32'hbb5bcadf),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b1047),
	.w1(32'hb996dce2),
	.w2(32'h3c22dcd3),
	.w3(32'hbb76e2bc),
	.w4(32'h38cdc592),
	.w5(32'hbae0704d),
	.w6(32'h3ab2585e),
	.w7(32'hbae59621),
	.w8(32'h3c21e4fa),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ee736),
	.w1(32'h35dcb0e3),
	.w2(32'hbc44a40f),
	.w3(32'hbb43b8c9),
	.w4(32'hbc54b119),
	.w5(32'hbc8f0263),
	.w6(32'hbae89ed9),
	.w7(32'hbc4def6d),
	.w8(32'hbc1c2bc4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e2c19),
	.w1(32'h3adc1d5a),
	.w2(32'hb995858e),
	.w3(32'hbc28fcc2),
	.w4(32'hbb1f00d9),
	.w5(32'h3b28fbc4),
	.w6(32'h3bdde588),
	.w7(32'hbc177811),
	.w8(32'hbb4d5144),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfbf6e),
	.w1(32'hbb94012d),
	.w2(32'h3c32f41b),
	.w3(32'hbb3b9215),
	.w4(32'h3c0c351d),
	.w5(32'h3d0943c9),
	.w6(32'hbb836b4d),
	.w7(32'h3bad10dc),
	.w8(32'h3bca0f09),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02ef94),
	.w1(32'hba8b006e),
	.w2(32'hba3726ed),
	.w3(32'h3bcceb2e),
	.w4(32'h3a413d26),
	.w5(32'hbb4c92ae),
	.w6(32'hbbb1c3c6),
	.w7(32'hb9709f8d),
	.w8(32'hbb0d486d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f2121),
	.w1(32'h3b0f60da),
	.w2(32'hbc023a55),
	.w3(32'hba10a9b1),
	.w4(32'h3ab0e9d1),
	.w5(32'hbb9d26b1),
	.w6(32'h3a0ed713),
	.w7(32'h3b4905dd),
	.w8(32'hbb159a85),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3b615),
	.w1(32'hbb2c520d),
	.w2(32'h3c259187),
	.w3(32'hbb675fd7),
	.w4(32'h3c4be89a),
	.w5(32'h3d03c7e8),
	.w6(32'hbc25166d),
	.w7(32'h3b4e3198),
	.w8(32'hb9abd322),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99092e),
	.w1(32'hbb3ac2a3),
	.w2(32'h3c1ce042),
	.w3(32'h3a71d9cf),
	.w4(32'h3c1744ea),
	.w5(32'h3c58a6d2),
	.w6(32'hbc35fdde),
	.w7(32'h3c5055a7),
	.w8(32'h3b2612e9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3d080),
	.w1(32'h3c33aa19),
	.w2(32'hbaa36b61),
	.w3(32'h3b781ade),
	.w4(32'h3b2f45d8),
	.w5(32'hbc2a70c3),
	.w6(32'h3b093373),
	.w7(32'h3b057a95),
	.w8(32'hbb6e3090),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf23bdf),
	.w1(32'h39de7e20),
	.w2(32'hbb11e200),
	.w3(32'hbb97645f),
	.w4(32'hbb9a1b0a),
	.w5(32'h39aeb0d7),
	.w6(32'h398aea9e),
	.w7(32'hbbab830d),
	.w8(32'hbb7a5cfb),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf39a91),
	.w1(32'hbbd17b66),
	.w2(32'hbc57cee3),
	.w3(32'hbc1beceb),
	.w4(32'hbbf584aa),
	.w5(32'hbb7ed409),
	.w6(32'h3b6cb6dd),
	.w7(32'hbab85fd3),
	.w8(32'h3b7148ec),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb367715),
	.w1(32'hbb9bab07),
	.w2(32'hbc6102c3),
	.w3(32'h3bb68a61),
	.w4(32'hbbe9dfb4),
	.w5(32'h3ac1ca59),
	.w6(32'h3b2dedfa),
	.w7(32'hbb04b681),
	.w8(32'hbc4c79b9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe6723),
	.w1(32'h3a22cd1f),
	.w2(32'hbb020bed),
	.w3(32'hbc4658bc),
	.w4(32'hba559c98),
	.w5(32'hbb27b365),
	.w6(32'hbc465b7a),
	.w7(32'h3a1ac8d4),
	.w8(32'h392de170),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f944b),
	.w1(32'h3bb7f30c),
	.w2(32'h39469746),
	.w3(32'h3af2d782),
	.w4(32'h3bb3a8b0),
	.w5(32'h39cca294),
	.w6(32'h3b016d50),
	.w7(32'h3b7e0a87),
	.w8(32'h3b51d9c1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45d03b),
	.w1(32'hbba68659),
	.w2(32'h3bb25395),
	.w3(32'h3b219b89),
	.w4(32'hbc8ba268),
	.w5(32'hbc9c518c),
	.w6(32'h3b7c7c01),
	.w7(32'hbb93ac56),
	.w8(32'h3b1ab3d9),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e7678),
	.w1(32'h3ba25d39),
	.w2(32'h3b5b642c),
	.w3(32'hbc3927c3),
	.w4(32'hbb6f067d),
	.w5(32'h3b1f6ae6),
	.w6(32'hbab42b0f),
	.w7(32'hb9ac16c5),
	.w8(32'h3b75f2af),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5acfef),
	.w1(32'hba2ca8f0),
	.w2(32'h3b891825),
	.w3(32'hbbc90907),
	.w4(32'h397b9f8e),
	.w5(32'h3b855b3b),
	.w6(32'h3ba1e9de),
	.w7(32'h3b201bee),
	.w8(32'h39bf7f67),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3943732b),
	.w1(32'hba04ef9a),
	.w2(32'hbb1838eb),
	.w3(32'h3b15a248),
	.w4(32'hbb877bb8),
	.w5(32'hba9334da),
	.w6(32'h3a0aa5de),
	.w7(32'h3b17a9d8),
	.w8(32'h3b962748),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bc3a9),
	.w1(32'h3b68bdcf),
	.w2(32'h3b251926),
	.w3(32'h39b56353),
	.w4(32'h3a7ce159),
	.w5(32'h3c918134),
	.w6(32'hbb4634cf),
	.w7(32'h3bda11c3),
	.w8(32'h3bab3fa2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ba988),
	.w1(32'hbbff909a),
	.w2(32'hbb908dd5),
	.w3(32'h3b71588f),
	.w4(32'hbbdfd9b9),
	.w5(32'hbbdc5c4f),
	.w6(32'h3a0b5b45),
	.w7(32'hba3c4fb5),
	.w8(32'h3b21f70f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb724f14),
	.w1(32'h3a1b1de0),
	.w2(32'hbaf5421e),
	.w3(32'hbb97737b),
	.w4(32'h3af376b4),
	.w5(32'h3b340104),
	.w6(32'h3bcd28ae),
	.w7(32'h396d5dfc),
	.w8(32'hb8a6ac91),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8af8b),
	.w1(32'hba08cddc),
	.w2(32'hbb7153c0),
	.w3(32'hba586338),
	.w4(32'h3a03d424),
	.w5(32'h3b091cd5),
	.w6(32'h3b8e2491),
	.w7(32'h3bfac4a2),
	.w8(32'h3b750344),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b1853b),
	.w1(32'hba22f629),
	.w2(32'hb9eef4db),
	.w3(32'h3c005d73),
	.w4(32'h3b9ad115),
	.w5(32'hba8e6c70),
	.w6(32'h3b73d1c5),
	.w7(32'h3c0b9d0d),
	.w8(32'h3ba9e219),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c6e13),
	.w1(32'h3b96ac73),
	.w2(32'h3c28bae8),
	.w3(32'h3a1ce89c),
	.w4(32'h3bccccfc),
	.w5(32'h3ba75734),
	.w6(32'h3b2dc56e),
	.w7(32'h3ba73a62),
	.w8(32'hbb1098cf),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ee02b),
	.w1(32'h3c01fbc3),
	.w2(32'h3b5d9247),
	.w3(32'h39d58591),
	.w4(32'h3b83a387),
	.w5(32'h3c6f6425),
	.w6(32'hbbf21138),
	.w7(32'hbb193ead),
	.w8(32'hbb2da4c4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39744f2d),
	.w1(32'hbb91bb63),
	.w2(32'hbc016f32),
	.w3(32'hbb9d1f4e),
	.w4(32'hbb48dfd9),
	.w5(32'hbac466e4),
	.w6(32'h3b3cb966),
	.w7(32'h3bbe375c),
	.w8(32'hbb36c4c4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06b02a),
	.w1(32'h3ae61dcd),
	.w2(32'h3c149ae8),
	.w3(32'h3c10bfb2),
	.w4(32'h3b19df11),
	.w5(32'h3bca6b30),
	.w6(32'hbae63484),
	.w7(32'hba2609eb),
	.w8(32'h3ba90f54),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a444107),
	.w1(32'h3a5f8fcc),
	.w2(32'h3bee2f98),
	.w3(32'hbb55b654),
	.w4(32'h3c0e08a8),
	.w5(32'h3be26d72),
	.w6(32'hbb7c50a3),
	.w7(32'hb9cb5ace),
	.w8(32'hba9d0c30),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9916677),
	.w1(32'h3a8a49b1),
	.w2(32'h3b108f0d),
	.w3(32'h3aa3920e),
	.w4(32'h3abb6185),
	.w5(32'hb94dcaac),
	.w6(32'hbb871f2f),
	.w7(32'hbb92ee1f),
	.w8(32'hbb6e5157),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad48c8a),
	.w1(32'hbbd5faf4),
	.w2(32'hbbeb55b4),
	.w3(32'hbb0da8e6),
	.w4(32'hbc0dafb6),
	.w5(32'hbc07d894),
	.w6(32'hbb37508c),
	.w7(32'hbb762580),
	.w8(32'hb98836db),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe6414),
	.w1(32'h3b8b1510),
	.w2(32'h3b3c79e4),
	.w3(32'hbbc9acae),
	.w4(32'h3b62fa25),
	.w5(32'h3adabe45),
	.w6(32'h3c07bb54),
	.w7(32'hba9c4fe2),
	.w8(32'hbbb73c67),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc7601),
	.w1(32'h3a9d7b69),
	.w2(32'hba1ea6c0),
	.w3(32'hba34d2c1),
	.w4(32'h3ab64821),
	.w5(32'hbbadf571),
	.w6(32'hbb4ff737),
	.w7(32'h3bae7cd3),
	.w8(32'h3b6ac3f3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88c1dd),
	.w1(32'h3bf1c2ef),
	.w2(32'h3c04bec6),
	.w3(32'hbac31fff),
	.w4(32'h3b76c8d7),
	.w5(32'h3b24d806),
	.w6(32'h3b32966c),
	.w7(32'h3bda45bd),
	.w8(32'h3b92f6d9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a913d8d),
	.w1(32'h3abdf74a),
	.w2(32'h3afa45a1),
	.w3(32'hb9934ef8),
	.w4(32'hbb9872d4),
	.w5(32'hbb95bef6),
	.w6(32'hbb738d1a),
	.w7(32'hbc1625c2),
	.w8(32'h3b0f57f7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59b4e3),
	.w1(32'h3b38a1f6),
	.w2(32'hbc10db2b),
	.w3(32'h3a9320ad),
	.w4(32'hb99960dc),
	.w5(32'hba90f51c),
	.w6(32'h3afd3c8b),
	.w7(32'h398e66e9),
	.w8(32'hbc15a787),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02cdc8),
	.w1(32'h3bbc0935),
	.w2(32'h3bafeb7d),
	.w3(32'hbba7cb41),
	.w4(32'h3b3b0862),
	.w5(32'h3a879a32),
	.w6(32'hbb173617),
	.w7(32'hbaa48832),
	.w8(32'hbb94d67c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1eca2),
	.w1(32'h3866ccce),
	.w2(32'hbaf876b9),
	.w3(32'hbbb0cb24),
	.w4(32'h3bd64e72),
	.w5(32'h3b82a99e),
	.w6(32'hbb75cfa5),
	.w7(32'h3b8ddde1),
	.w8(32'h3c10e19f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b717641),
	.w1(32'hbc1d0f81),
	.w2(32'hbc0e69eb),
	.w3(32'h3a9cf62d),
	.w4(32'hbbe7c59d),
	.w5(32'hbc1ebdb6),
	.w6(32'hbb88b1ab),
	.w7(32'hbb9a21c9),
	.w8(32'hbba0bd80),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedade1),
	.w1(32'h3bc0613e),
	.w2(32'h3b8e8fc5),
	.w3(32'hbb05e110),
	.w4(32'h3b6281c1),
	.w5(32'h3c0617f7),
	.w6(32'h3b896238),
	.w7(32'h3980ec38),
	.w8(32'h3b6b7ab7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b6be9),
	.w1(32'h3af59c6e),
	.w2(32'hba742dde),
	.w3(32'h3bc3cdeb),
	.w4(32'h3bb0b858),
	.w5(32'h3c1a7cbe),
	.w6(32'h3c23da4b),
	.w7(32'h3bd9ce76),
	.w8(32'h3b893b07),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07032d),
	.w1(32'h3c108041),
	.w2(32'hbbeb31ea),
	.w3(32'h3babed20),
	.w4(32'h3b8410ad),
	.w5(32'hbb10867c),
	.w6(32'hbbd15380),
	.w7(32'h3ba87ffd),
	.w8(32'hbb9ec974),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe708c7),
	.w1(32'hbb1d1a11),
	.w2(32'h3b78709c),
	.w3(32'hbc0743a8),
	.w4(32'hba3c1d8b),
	.w5(32'h3b4b4ea9),
	.w6(32'h3c4445be),
	.w7(32'h3b4f6c12),
	.w8(32'h3b453dfa),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d1e1f),
	.w1(32'hbbc21431),
	.w2(32'hbbf0d862),
	.w3(32'h3bbbc58d),
	.w4(32'hbbbf144f),
	.w5(32'hbb44171d),
	.w6(32'hbb2703f2),
	.w7(32'hbac29c60),
	.w8(32'hbbb6b09a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8e2a5),
	.w1(32'h3af75e40),
	.w2(32'h3c7552d0),
	.w3(32'hbbe2b8e5),
	.w4(32'h3c077805),
	.w5(32'h3c8c6a3f),
	.w6(32'hbb0d3a1c),
	.w7(32'h3b6f59d9),
	.w8(32'h3c0fd17d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35060a),
	.w1(32'hba3083bf),
	.w2(32'hbb00c613),
	.w3(32'h3b5b63ac),
	.w4(32'hbbbe4f5f),
	.w5(32'hbb837625),
	.w6(32'hbb8167a9),
	.w7(32'h3a10688f),
	.w8(32'hbb56bfb7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ff887),
	.w1(32'hbb8aee71),
	.w2(32'hba2f2f54),
	.w3(32'hba0f7a86),
	.w4(32'h3b072787),
	.w5(32'h3c5a5def),
	.w6(32'hbb8558b9),
	.w7(32'h3bb151f2),
	.w8(32'h3ba9eb4b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9e7ab),
	.w1(32'h39d47b38),
	.w2(32'h3b255c95),
	.w3(32'h3bbe00f1),
	.w4(32'h3bc433cf),
	.w5(32'h3c3ba1b0),
	.w6(32'hbbee309e),
	.w7(32'h3c1f25d4),
	.w8(32'h3c15b538),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37cbc5),
	.w1(32'hbb10986c),
	.w2(32'hbc14b5d7),
	.w3(32'h3c01eacf),
	.w4(32'hbc0baf45),
	.w5(32'hbc2d71b1),
	.w6(32'h3bcb970b),
	.w7(32'hbc062c66),
	.w8(32'hbbc45148),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43aeb3),
	.w1(32'hbb3de8d1),
	.w2(32'hba82dbaf),
	.w3(32'hbbf97157),
	.w4(32'h38a8ef76),
	.w5(32'h3b639754),
	.w6(32'h3b359cf8),
	.w7(32'hbb03185a),
	.w8(32'h3b49928f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b375a84),
	.w1(32'hba8498a7),
	.w2(32'h3abe716b),
	.w3(32'h3bef9c87),
	.w4(32'hbb327ff1),
	.w5(32'h3b2fe4b0),
	.w6(32'h3aa3984c),
	.w7(32'hb9f88468),
	.w8(32'hbb4e386f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b979e6e),
	.w1(32'hba8522ac),
	.w2(32'hb742670f),
	.w3(32'hbad13ca6),
	.w4(32'hbb6e83ee),
	.w5(32'hbb4f9222),
	.w6(32'hbb4e3cff),
	.w7(32'hba93d29c),
	.w8(32'hbb2bc9d5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06186f),
	.w1(32'h3b257410),
	.w2(32'hbbb36019),
	.w3(32'hba87f277),
	.w4(32'hb9fb0dac),
	.w5(32'hbad491c4),
	.w6(32'hbc195150),
	.w7(32'h3a9d29a6),
	.w8(32'h3b505001),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a880579),
	.w1(32'hbc5c2c65),
	.w2(32'hbc820db0),
	.w3(32'h3af1f85f),
	.w4(32'hbc0656f5),
	.w5(32'h3be54255),
	.w6(32'h3a69913a),
	.w7(32'h3b1eb2b5),
	.w8(32'h3abfcff1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f6b87),
	.w1(32'hbb935159),
	.w2(32'hba42080e),
	.w3(32'h3bf7b843),
	.w4(32'hbb2918d3),
	.w5(32'h3c12b754),
	.w6(32'h3b30d226),
	.w7(32'hbbcbde15),
	.w8(32'h3a9c66e1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0360c2),
	.w1(32'h3aaa5c2a),
	.w2(32'hbaa24ed2),
	.w3(32'h3b826d64),
	.w4(32'hbb38d58e),
	.w5(32'h3a6f6c19),
	.w6(32'hbbb1ce10),
	.w7(32'hbbd68b1f),
	.w8(32'hbbb6ebb5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69394b),
	.w1(32'h3b63549e),
	.w2(32'h3b0f7cda),
	.w3(32'hbbd18fb2),
	.w4(32'h3bb2d0b0),
	.w5(32'h3b37ffd8),
	.w6(32'h3ba4e5dc),
	.w7(32'h3c01b271),
	.w8(32'h3c36006a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b68b7),
	.w1(32'hbb2195a4),
	.w2(32'h3b7a6792),
	.w3(32'h3bb1142c),
	.w4(32'h3b8e8c97),
	.w5(32'h3c52e6f4),
	.w6(32'h3b23cc0a),
	.w7(32'h3b0a2372),
	.w8(32'h39729bbf),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a61f7),
	.w1(32'hbafd4ccb),
	.w2(32'h3bd31376),
	.w3(32'h3a928556),
	.w4(32'h3c14a51b),
	.w5(32'h3bbeb89e),
	.w6(32'h3aa83a74),
	.w7(32'hbb1cb098),
	.w8(32'h3b00ddee),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c7b07),
	.w1(32'h3b89725c),
	.w2(32'hba989b5e),
	.w3(32'hbaced575),
	.w4(32'h3a9b92a3),
	.w5(32'h3b738837),
	.w6(32'hbb93dff2),
	.w7(32'hb8f511d3),
	.w8(32'hba960ef2),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7dbed),
	.w1(32'hbc0234c7),
	.w2(32'hbbb4ecb4),
	.w3(32'hbbb63e0a),
	.w4(32'hbbfa9844),
	.w5(32'h3b064d8c),
	.w6(32'hba0420dd),
	.w7(32'hbb2b3213),
	.w8(32'h3b5e9168),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5632ed),
	.w1(32'hbb96992a),
	.w2(32'hbc346ce6),
	.w3(32'h3b6416b7),
	.w4(32'hbb927340),
	.w5(32'hbc45c8cb),
	.w6(32'h3a90deff),
	.w7(32'hbb8de918),
	.w8(32'hbb8a2fb8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2cf95),
	.w1(32'h3a906076),
	.w2(32'h3c3aa359),
	.w3(32'hbaf52678),
	.w4(32'h3c439a76),
	.w5(32'h3c2cb320),
	.w6(32'hbb1e89fd),
	.w7(32'h3bf725d3),
	.w8(32'h3b8c21e2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb24f80),
	.w1(32'h3b88fd38),
	.w2(32'h38e3cac7),
	.w3(32'h3c1f3aa8),
	.w4(32'h3b520b58),
	.w5(32'h3b4ef74a),
	.w6(32'h3a9f3feb),
	.w7(32'h39942124),
	.w8(32'hbc2b7ab7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebe8c3),
	.w1(32'h3bef6619),
	.w2(32'h3b6f40b0),
	.w3(32'hbc0c6782),
	.w4(32'h3aa1d48a),
	.w5(32'h3b0466b2),
	.w6(32'hbbb537fa),
	.w7(32'hbb968f35),
	.w8(32'h3b543564),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba481df4),
	.w1(32'hbbf66e18),
	.w2(32'hbb4e67f8),
	.w3(32'hbaeed0b0),
	.w4(32'hbb2c3775),
	.w5(32'h3bb0396f),
	.w6(32'h3ac4a3dd),
	.w7(32'h3a13ab55),
	.w8(32'h3bcade9c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddc913),
	.w1(32'h3861b36b),
	.w2(32'h3bad204a),
	.w3(32'h3bc5f492),
	.w4(32'h3b0ec962),
	.w5(32'h3b84a769),
	.w6(32'h3bbecd32),
	.w7(32'h3b9c4cb6),
	.w8(32'h3bce3e84),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73f499),
	.w1(32'h3bab6aaa),
	.w2(32'hbbceb708),
	.w3(32'h3a076009),
	.w4(32'h3b9fd8f3),
	.w5(32'hbb5374b0),
	.w6(32'hb8d30695),
	.w7(32'h3a87e3e8),
	.w8(32'h3a95be29),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99b8eb),
	.w1(32'hbb20a877),
	.w2(32'hbbc41b75),
	.w3(32'hbad072bb),
	.w4(32'hbbca6599),
	.w5(32'hbc4f2ae3),
	.w6(32'h3b82407b),
	.w7(32'hbb908fc6),
	.w8(32'hbbeab947),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8093cb),
	.w1(32'h3a4566da),
	.w2(32'hba9e4081),
	.w3(32'hba32d4ae),
	.w4(32'h3ab0123b),
	.w5(32'hbaea7485),
	.w6(32'h3aadd2d5),
	.w7(32'hba9d1edf),
	.w8(32'hbc1fd306),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f8b0e),
	.w1(32'h38f01569),
	.w2(32'hbb853732),
	.w3(32'hbbb1402e),
	.w4(32'hbbc046ba),
	.w5(32'hbc130a6e),
	.w6(32'hbb8b528a),
	.w7(32'hbbd01aee),
	.w8(32'hbaa481eb),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6c192),
	.w1(32'h3ab4a2ef),
	.w2(32'hbc44608a),
	.w3(32'hbab26b22),
	.w4(32'hbbe9fd98),
	.w5(32'hbc6e3a1e),
	.w6(32'h3b40f157),
	.w7(32'hbb733d81),
	.w8(32'hbbc0c6c8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc285829),
	.w1(32'h3b2d01e5),
	.w2(32'hba7da9c8),
	.w3(32'hbc1796d0),
	.w4(32'h3be2fe1a),
	.w5(32'h3a973e1f),
	.w6(32'hba7864f4),
	.w7(32'h3b5948fb),
	.w8(32'h3aab1575),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82e019),
	.w1(32'h3b178ba3),
	.w2(32'hbc521eea),
	.w3(32'h3bb565e2),
	.w4(32'h3b435e75),
	.w5(32'hbbdb3498),
	.w6(32'hbab0e8a4),
	.w7(32'h3abe17d1),
	.w8(32'hbb8650d5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5f836),
	.w1(32'h3a1017da),
	.w2(32'h3c1cec7a),
	.w3(32'hbb18f80f),
	.w4(32'h3baf6bee),
	.w5(32'h3c086c82),
	.w6(32'h3b3f8299),
	.w7(32'h3ba5c29a),
	.w8(32'h3be57caa),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b353e),
	.w1(32'h3bdbaa20),
	.w2(32'hbbbcc747),
	.w3(32'h3b83b921),
	.w4(32'h3ba020b3),
	.w5(32'h3b82b677),
	.w6(32'hbaa6277e),
	.w7(32'h3b43b948),
	.w8(32'hbb23bc72),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe817f),
	.w1(32'hbaafac06),
	.w2(32'h3ad3990d),
	.w3(32'hbb54eff5),
	.w4(32'h3b2ef6a0),
	.w5(32'hbbee2f53),
	.w6(32'h3ae4e73b),
	.w7(32'hbb637860),
	.w8(32'hbc1b8fbe),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf553ae),
	.w1(32'h3b1d4145),
	.w2(32'h3ad548c3),
	.w3(32'hbc1a3f2e),
	.w4(32'h3b7af5f0),
	.w5(32'hbb265dda),
	.w6(32'hbc09e2bd),
	.w7(32'h3b05c673),
	.w8(32'hbb00164b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c83bb9),
	.w1(32'hbad6bb3f),
	.w2(32'hba8ae1f6),
	.w3(32'h3b41ac58),
	.w4(32'hbad12ffb),
	.w5(32'h3a67764d),
	.w6(32'h3b0bdf2b),
	.w7(32'hbb1c089c),
	.w8(32'h3ae73eb0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c0065),
	.w1(32'hba828989),
	.w2(32'hbba560f0),
	.w3(32'h3a775ac7),
	.w4(32'hbac71cb5),
	.w5(32'h3a29ecf0),
	.w6(32'h3805089e),
	.w7(32'h3b9b6f92),
	.w8(32'h3c1e0b2f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1b772),
	.w1(32'h3bc70651),
	.w2(32'hbbc5d6ab),
	.w3(32'h3b4efd81),
	.w4(32'h3bf79429),
	.w5(32'hbb890e41),
	.w6(32'h39a8130e),
	.w7(32'h3ab36442),
	.w8(32'h3a58cce6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad2ebc),
	.w1(32'h3b51e9a0),
	.w2(32'hba15921d),
	.w3(32'h3aee72cc),
	.w4(32'h3ae2d12f),
	.w5(32'h3c0f82c4),
	.w6(32'hb96fa2b4),
	.w7(32'h3bf14792),
	.w8(32'h3b350301),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37768fdb),
	.w1(32'hbaeb1486),
	.w2(32'hba518157),
	.w3(32'hbb5d2c09),
	.w4(32'h3970ebca),
	.w5(32'h3ab0e079),
	.w6(32'hba2821e1),
	.w7(32'hbb9878fe),
	.w8(32'hbb7f0b69),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf9fc9),
	.w1(32'hbaf9590b),
	.w2(32'h3b06ca75),
	.w3(32'h3a7b49f0),
	.w4(32'hb9a82c64),
	.w5(32'hbb33d7ff),
	.w6(32'hbaebf0dd),
	.w7(32'hba15cb17),
	.w8(32'h3b2b94dd),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a2d4b),
	.w1(32'h3b6dddd4),
	.w2(32'hbab5101e),
	.w3(32'hba4ab6ed),
	.w4(32'h3aa48125),
	.w5(32'hbb0c75c5),
	.w6(32'h3b2efec2),
	.w7(32'h3b075895),
	.w8(32'h3b899956),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ac9a7),
	.w1(32'hba8df505),
	.w2(32'hbb92390a),
	.w3(32'h3b7e033b),
	.w4(32'h3a809564),
	.w5(32'h3b0b0246),
	.w6(32'h3b8ade09),
	.w7(32'hbb8abd47),
	.w8(32'hbba46e09),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa59671),
	.w1(32'hbae2917f),
	.w2(32'hba94821b),
	.w3(32'hbb8792c9),
	.w4(32'h3a34cd9a),
	.w5(32'hb9faf587),
	.w6(32'hbad47f4c),
	.w7(32'h3a085aef),
	.w8(32'hbb07c478),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31b1ff),
	.w1(32'hbb0b8f0a),
	.w2(32'hb98b8c9e),
	.w3(32'hba32402d),
	.w4(32'hbb9c7e1c),
	.w5(32'hba490f27),
	.w6(32'hbb025215),
	.w7(32'h39ef767d),
	.w8(32'h3ae42b05),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04f744),
	.w1(32'hbb0001bb),
	.w2(32'hbb0795d5),
	.w3(32'hbb652861),
	.w4(32'hba83df18),
	.w5(32'hb935cf40),
	.w6(32'hb9c4e56b),
	.w7(32'hb8f4eb0d),
	.w8(32'h39adbcbe),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cde29),
	.w1(32'h3bc34f32),
	.w2(32'h3bc97302),
	.w3(32'hba7c3caf),
	.w4(32'h3a12b263),
	.w5(32'h3b506412),
	.w6(32'hb9bfbdf2),
	.w7(32'h38d8f755),
	.w8(32'hbae318f1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4e16a),
	.w1(32'hbb960a6b),
	.w2(32'hbba0b79d),
	.w3(32'h3b1fec0f),
	.w4(32'h3a6d0843),
	.w5(32'hbb6eb8ce),
	.w6(32'hba0bf24f),
	.w7(32'h3af18ef0),
	.w8(32'h3b34e2d3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af914),
	.w1(32'hbb89a37b),
	.w2(32'hbacf9952),
	.w3(32'hb8293d93),
	.w4(32'hb7b522ec),
	.w5(32'hba8cd284),
	.w6(32'h3b01ae58),
	.w7(32'h3b4f5ef6),
	.w8(32'h3ba750d1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16c42e),
	.w1(32'h3be9c795),
	.w2(32'h3ba48545),
	.w3(32'h3aa3cbfa),
	.w4(32'hbaef2fc2),
	.w5(32'h3a889e75),
	.w6(32'h3b044d25),
	.w7(32'h3a92f0ef),
	.w8(32'hba003b91),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a3824),
	.w1(32'h3b65adeb),
	.w2(32'h3a59ce7f),
	.w3(32'hbb394069),
	.w4(32'h3badbccf),
	.w5(32'h3b08eb97),
	.w6(32'hba7733c2),
	.w7(32'h3b2d1cd9),
	.w8(32'h3a0c4a1e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70b18a),
	.w1(32'hbb2c5dfe),
	.w2(32'hbb914f9e),
	.w3(32'h3b6a3072),
	.w4(32'hbb051e1f),
	.w5(32'hbb4a324d),
	.w6(32'hba35f108),
	.w7(32'hbb29c9b2),
	.w8(32'hbb4d8ba9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2c194),
	.w1(32'h3b9aa306),
	.w2(32'h3ac123bc),
	.w3(32'hbaf3e7e9),
	.w4(32'hbb05d790),
	.w5(32'hbaf4c706),
	.w6(32'hbb02e1cf),
	.w7(32'hba639eef),
	.w8(32'h3ac60a01),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d2bb3),
	.w1(32'hbb3ac05b),
	.w2(32'h3b0ffd14),
	.w3(32'h3b2a16db),
	.w4(32'hba47e8e1),
	.w5(32'hba60e440),
	.w6(32'h399705d0),
	.w7(32'hbb03ace2),
	.w8(32'hbadc86fe),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cc6d3),
	.w1(32'hb9298bae),
	.w2(32'hba4c05ac),
	.w3(32'h3a313111),
	.w4(32'hba553ea7),
	.w5(32'h3bfe4c09),
	.w6(32'hb9b53a92),
	.w7(32'h3aee2ac2),
	.w8(32'h3a2d3bf3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a157b),
	.w1(32'hba73e1fa),
	.w2(32'h3906532f),
	.w3(32'hbb94eb4a),
	.w4(32'hba492081),
	.w5(32'hbb46cabf),
	.w6(32'h3acaa49b),
	.w7(32'h3aafd04a),
	.w8(32'hbbb6dd50),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21526c),
	.w1(32'hbac9dfe8),
	.w2(32'h3b451570),
	.w3(32'h39c1fad2),
	.w4(32'h3aedde55),
	.w5(32'hba9c4f91),
	.w6(32'h39bf3c4d),
	.w7(32'h3ba010d9),
	.w8(32'h3bc3bab0),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fffda),
	.w1(32'hbb1be3bc),
	.w2(32'h3ab4341a),
	.w3(32'h3b423d6b),
	.w4(32'h3ba48b55),
	.w5(32'hbb3d7219),
	.w6(32'h3b7905fc),
	.w7(32'h3b650f91),
	.w8(32'h3a009ebc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9942d9),
	.w1(32'hbaa4482d),
	.w2(32'hbb107e48),
	.w3(32'hbb36b4c1),
	.w4(32'hbb273341),
	.w5(32'hba1555e7),
	.w6(32'hb8cf91d0),
	.w7(32'hbb30f7cb),
	.w8(32'hbac80ed4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0539f),
	.w1(32'h3b1d7c72),
	.w2(32'h392c1fa7),
	.w3(32'h39179bfd),
	.w4(32'h3b074c15),
	.w5(32'hbb28cb90),
	.w6(32'hbba29862),
	.w7(32'hbb73f5da),
	.w8(32'h3b592f37),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa21c1e),
	.w1(32'hbb49d144),
	.w2(32'hbafed0b2),
	.w3(32'hb91938ec),
	.w4(32'hbad2e8eb),
	.w5(32'hbb0e5c13),
	.w6(32'h3a575c15),
	.w7(32'hba81155a),
	.w8(32'hba73d84e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7a147),
	.w1(32'h3b51aa9c),
	.w2(32'h3b5fead6),
	.w3(32'hbb045d43),
	.w4(32'h3bf97e1b),
	.w5(32'h3b307da0),
	.w6(32'h3a7c9cdf),
	.w7(32'hbb01ab0d),
	.w8(32'hbb118d8b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b675467),
	.w1(32'h3af9ba1f),
	.w2(32'hbb39071b),
	.w3(32'h3a68004c),
	.w4(32'hbaa9d948),
	.w5(32'hbb823abf),
	.w6(32'hbb4ac7a2),
	.w7(32'hbb905082),
	.w8(32'hbb91044c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba409330),
	.w1(32'hbb00878a),
	.w2(32'hb979c31f),
	.w3(32'h3ad86cd4),
	.w4(32'h3b10befe),
	.w5(32'hbb242e74),
	.w6(32'hbb86a68a),
	.w7(32'hbb33e270),
	.w8(32'hbb9ae7df),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9572344),
	.w1(32'h3bc0baa6),
	.w2(32'h3bcd6111),
	.w3(32'h373f4afa),
	.w4(32'h3b8c28bd),
	.w5(32'h3b9655a9),
	.w6(32'hbad485d7),
	.w7(32'h3aa47102),
	.w8(32'h3aeaccbd),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b0ba7),
	.w1(32'hba82d5b3),
	.w2(32'h3bc6c915),
	.w3(32'hbb453fdf),
	.w4(32'h3ac14901),
	.w5(32'h3c4b5a39),
	.w6(32'hbb7c02be),
	.w7(32'h3a5fdc70),
	.w8(32'hbbe84928),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e152a),
	.w1(32'hbae5bb29),
	.w2(32'h3bd13891),
	.w3(32'hbb422aa2),
	.w4(32'hbaa197c1),
	.w5(32'h3c2291ff),
	.w6(32'h3a240027),
	.w7(32'hba6d6064),
	.w8(32'hbb1919cb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fb0a2),
	.w1(32'h3babd924),
	.w2(32'h3b5c27d8),
	.w3(32'hb9839d05),
	.w4(32'h3a1fbe76),
	.w5(32'hba66412c),
	.w6(32'hb989d0c6),
	.w7(32'h3afe379f),
	.w8(32'h3af4d24b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb0b61),
	.w1(32'hba026af7),
	.w2(32'hba244a65),
	.w3(32'h3b22cb9b),
	.w4(32'h3a8b943d),
	.w5(32'h3a68b43b),
	.w6(32'h3a224b8b),
	.w7(32'hbaf87a61),
	.w8(32'h3a6bdeae),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab60b0),
	.w1(32'h3a6eada1),
	.w2(32'hba646cef),
	.w3(32'hb95808fa),
	.w4(32'hba3b6305),
	.w5(32'hbaee98ad),
	.w6(32'hbaebcf93),
	.w7(32'hb9f570b2),
	.w8(32'h3b68f9cf),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92a16b),
	.w1(32'hba3d2665),
	.w2(32'h3b6ff6b2),
	.w3(32'h3a9a18da),
	.w4(32'h3a97d143),
	.w5(32'h3aa8f9cd),
	.w6(32'hbb4cf294),
	.w7(32'hba1fe88a),
	.w8(32'hba7c3a4f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b095d40),
	.w1(32'h3b023431),
	.w2(32'h3b79c92f),
	.w3(32'h3a5f3738),
	.w4(32'hbad079cb),
	.w5(32'h3c2988a5),
	.w6(32'hba607b7b),
	.w7(32'hbb0f8fd2),
	.w8(32'hbb643c63),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd590e),
	.w1(32'hba09fc62),
	.w2(32'hbaa7dddc),
	.w3(32'hba42aece),
	.w4(32'hbb897b2e),
	.w5(32'hbbaa92c1),
	.w6(32'h3bbf6ed8),
	.w7(32'h3b704f8e),
	.w8(32'h3b89ac9e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e7fb4),
	.w1(32'h3a198e34),
	.w2(32'h3b7214b2),
	.w3(32'hbb013bc4),
	.w4(32'h3a9145c1),
	.w5(32'h3b2cc43b),
	.w6(32'hb9cb4e4b),
	.w7(32'hba1b80d1),
	.w8(32'h3b13cc11),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2b55d),
	.w1(32'h3bc2d120),
	.w2(32'h3aeb8061),
	.w3(32'hbb63f5d1),
	.w4(32'hbb13e7ad),
	.w5(32'hbaeb1dde),
	.w6(32'h3b9df253),
	.w7(32'hba81ab69),
	.w8(32'h3b613a1c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4c337),
	.w1(32'hbb3b5d04),
	.w2(32'hbb603599),
	.w3(32'h3b4b4706),
	.w4(32'hb9087261),
	.w5(32'hbb48576d),
	.w6(32'h3b5447df),
	.w7(32'hbaa40899),
	.w8(32'hba8b1c38),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f00bb),
	.w1(32'hba82e740),
	.w2(32'hba6bd8e0),
	.w3(32'h39c42329),
	.w4(32'h38996ee7),
	.w5(32'hbb29cc69),
	.w6(32'hba59a88d),
	.w7(32'hbaa8f927),
	.w8(32'hbaa1a640),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb8469),
	.w1(32'hba09b64c),
	.w2(32'hbb7b57ff),
	.w3(32'hba178379),
	.w4(32'h3b5ab7fc),
	.w5(32'h3bad6908),
	.w6(32'h3a731e0d),
	.w7(32'h3a847253),
	.w8(32'h3a33b044),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ed546),
	.w1(32'h3b8464fb),
	.w2(32'hbb11dedd),
	.w3(32'h3a826d18),
	.w4(32'hbb4e5219),
	.w5(32'hba5af596),
	.w6(32'h3b1ecec5),
	.w7(32'hbba411db),
	.w8(32'h3b43f34f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ad061),
	.w1(32'h3be1d109),
	.w2(32'h3c06a1a4),
	.w3(32'hbab2c6a1),
	.w4(32'hbae442b2),
	.w5(32'h3b59cefd),
	.w6(32'h3aeadb10),
	.w7(32'hbb324008),
	.w8(32'h3a94fdd4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f57173),
	.w1(32'h3b269802),
	.w2(32'hb767e685),
	.w3(32'h3b212b2e),
	.w4(32'h3b808092),
	.w5(32'h3b28027c),
	.w6(32'h3b28ce46),
	.w7(32'hba8d2b59),
	.w8(32'hba6b6c1b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb299fba),
	.w1(32'hba42b573),
	.w2(32'h3a7deaa0),
	.w3(32'h3b0ff289),
	.w4(32'hbaa1b404),
	.w5(32'h3b50518f),
	.w6(32'h3afe7a52),
	.w7(32'hbb1d8df2),
	.w8(32'h3a6f1768),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb00b0),
	.w1(32'hb966116f),
	.w2(32'h3b17a831),
	.w3(32'h39e27862),
	.w4(32'h3a834192),
	.w5(32'h3bbf329a),
	.w6(32'hb9a7a7a6),
	.w7(32'hbae9a2e0),
	.w8(32'hbbbe9b49),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39292a),
	.w1(32'h3b2e794c),
	.w2(32'h3b03304d),
	.w3(32'hbaaf0b26),
	.w4(32'hbbbe8efa),
	.w5(32'h3b655d0e),
	.w6(32'hb9a26312),
	.w7(32'hbad3251e),
	.w8(32'hbbeb9b49),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83185f),
	.w1(32'hb85b9824),
	.w2(32'hba6b8e62),
	.w3(32'h3b3d2e82),
	.w4(32'h39933051),
	.w5(32'hbb33d104),
	.w6(32'hbba6f2f1),
	.w7(32'h3a0d6e79),
	.w8(32'hbb2a506c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f848f),
	.w1(32'hba7e516f),
	.w2(32'hbaa129c0),
	.w3(32'hba187e80),
	.w4(32'hb92e22ac),
	.w5(32'hb9b4a620),
	.w6(32'hbaa46bfc),
	.w7(32'hb9e554fb),
	.w8(32'hba8f1e52),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b6ea8f),
	.w1(32'h3b5acff9),
	.w2(32'h3b323501),
	.w3(32'h38a522c1),
	.w4(32'h39e33df9),
	.w5(32'h3aab4eb0),
	.w6(32'hbaa4e1b2),
	.w7(32'h3afc2895),
	.w8(32'hba79c0b3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81ea0a),
	.w1(32'h394ca1ab),
	.w2(32'hbb96d235),
	.w3(32'h39d343e8),
	.w4(32'h3aa987d5),
	.w5(32'hbb27ae79),
	.w6(32'h3b45626d),
	.w7(32'hbb5a9a8c),
	.w8(32'hbaef3002),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b445),
	.w1(32'hbb4472c2),
	.w2(32'hba7e44ee),
	.w3(32'h38ddc34b),
	.w4(32'h3af7a087),
	.w5(32'hbb96dd11),
	.w6(32'hbb5ed9c8),
	.w7(32'h3b4b54d1),
	.w8(32'hb67591f9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2c3b0),
	.w1(32'h3ac7653d),
	.w2(32'hbb5bba80),
	.w3(32'hbb214f61),
	.w4(32'h39fb2ef0),
	.w5(32'h3a430be9),
	.w6(32'h3a58a54b),
	.w7(32'h3b059c51),
	.w8(32'hbb55129c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afffc8a),
	.w1(32'h3b14d8df),
	.w2(32'hba83260f),
	.w3(32'h3a7b3f38),
	.w4(32'h38a740c9),
	.w5(32'h39b73dd6),
	.w6(32'hbb899e42),
	.w7(32'hbac6fe9c),
	.w8(32'hbbace3c2),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0055ee),
	.w1(32'hbb853c6b),
	.w2(32'hba213995),
	.w3(32'h3ab66bd5),
	.w4(32'h3a1e5575),
	.w5(32'hba8a1041),
	.w6(32'hbb5d30c3),
	.w7(32'hbada5874),
	.w8(32'h386b7398),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7b63b),
	.w1(32'hb9eb0630),
	.w2(32'h3b09d012),
	.w3(32'hbac255c0),
	.w4(32'hba90440a),
	.w5(32'h3ae3bb22),
	.w6(32'hbb6a45d9),
	.w7(32'h3a266b2e),
	.w8(32'hb8c12edd),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81eeb6),
	.w1(32'hbaa5691a),
	.w2(32'h39e31248),
	.w3(32'hbabbaa76),
	.w4(32'hbb4a0bff),
	.w5(32'h3bdbdc16),
	.w6(32'h3a25a6a8),
	.w7(32'hbb1220e6),
	.w8(32'hbb192d23),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ae5ac),
	.w1(32'h3a8bc0c0),
	.w2(32'hbba59f3a),
	.w3(32'h3ade7f11),
	.w4(32'h396c0d52),
	.w5(32'hba500bb5),
	.w6(32'h3ad3af03),
	.w7(32'hba53f4eb),
	.w8(32'h3b053f37),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb058326),
	.w1(32'hba22c144),
	.w2(32'hbb8da742),
	.w3(32'hbabc65e3),
	.w4(32'hbb87cf5f),
	.w5(32'hbb752265),
	.w6(32'h3abc8f10),
	.w7(32'hbafa0593),
	.w8(32'hbac15071),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb498ae6),
	.w1(32'hbb77621b),
	.w2(32'h3abcf195),
	.w3(32'h383b9a93),
	.w4(32'hbbcd5ef5),
	.w5(32'hbbb9d977),
	.w6(32'hba5aca5d),
	.w7(32'hbb0c7107),
	.w8(32'h39b9c5e5),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f205a),
	.w1(32'h39ccfc2b),
	.w2(32'h3a86d93f),
	.w3(32'hbbb3cca7),
	.w4(32'hbae02780),
	.w5(32'h3aec3dbd),
	.w6(32'hba3d08ce),
	.w7(32'hbb1d3d52),
	.w8(32'hbb1a7381),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule