module layer_8_featuremap_151(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b252395),
	.w1(32'hbc514208),
	.w2(32'hbd3a67ff),
	.w3(32'h3bf16da9),
	.w4(32'h3bb41dad),
	.w5(32'hbbe51a16),
	.w6(32'h3c0908b0),
	.w7(32'hbcb0a8fd),
	.w8(32'hbc99c7fb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b85fb4),
	.w1(32'hbb7a0e59),
	.w2(32'hbc861d04),
	.w3(32'hbb61d3b1),
	.w4(32'hbbd2e9b2),
	.w5(32'h3c9d1ec0),
	.w6(32'hbb9705cd),
	.w7(32'h3c96e5a2),
	.w8(32'h3d139b38),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd871e25),
	.w1(32'hbd25c214),
	.w2(32'hbc7fe56b),
	.w3(32'h3c8448fe),
	.w4(32'hbc1b5f9a),
	.w5(32'hbb70a710),
	.w6(32'h3c99e86d),
	.w7(32'hbbb08db6),
	.w8(32'h3bb1ba24),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85b0b0),
	.w1(32'hbb925e53),
	.w2(32'hbc5fd6b0),
	.w3(32'hb9f4710e),
	.w4(32'hbad23e16),
	.w5(32'h3b696c37),
	.w6(32'hbc042619),
	.w7(32'hbc8773a4),
	.w8(32'hbc6e03cc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98af9e),
	.w1(32'h3a866d40),
	.w2(32'hbac836e7),
	.w3(32'hbb03bc18),
	.w4(32'hbc0d42ac),
	.w5(32'h3a5dad33),
	.w6(32'hbc067628),
	.w7(32'hbc84dfde),
	.w8(32'hbcda7660),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c733844),
	.w1(32'hbc3eab0e),
	.w2(32'h3c17f3dc),
	.w3(32'hbc24035c),
	.w4(32'hbb31fab0),
	.w5(32'h3c9484eb),
	.w6(32'hbce3fe7d),
	.w7(32'h3c1217d5),
	.w8(32'h3cb33308),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc602c99),
	.w1(32'hbb8af3f7),
	.w2(32'h3be006a8),
	.w3(32'hbb5a825e),
	.w4(32'hbc162edf),
	.w5(32'h3bf29084),
	.w6(32'h3cd9fbfc),
	.w7(32'h3b37b461),
	.w8(32'hbc4688df),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d047099),
	.w1(32'hbbedc34e),
	.w2(32'h3c8918d4),
	.w3(32'h3c823d98),
	.w4(32'hbb271191),
	.w5(32'hba8a97b6),
	.w6(32'hbc62a2b7),
	.w7(32'hbcb000b2),
	.w8(32'hbcb75652),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95f41c),
	.w1(32'hbbfeba5e),
	.w2(32'h3b55b39e),
	.w3(32'hba50d55d),
	.w4(32'hbcb8d4c4),
	.w5(32'hbcb52867),
	.w6(32'h3cb2e4e4),
	.w7(32'hbc1caa69),
	.w8(32'hbbc682ef),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb6b22),
	.w1(32'hb977357c),
	.w2(32'hbc8235ea),
	.w3(32'hbca285fc),
	.w4(32'hbc7a0ca4),
	.w5(32'hbc6f465d),
	.w6(32'h3b8393fe),
	.w7(32'hbc483a6b),
	.w8(32'hbb51edc1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfbb6e3),
	.w1(32'h3c7e12c3),
	.w2(32'h3c7f7fdb),
	.w3(32'h3b51db54),
	.w4(32'hbb4e7aba),
	.w5(32'h3baa4ce1),
	.w6(32'h3bf7b0bf),
	.w7(32'hbc754a8b),
	.w8(32'hbd10af63),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d75c25d),
	.w1(32'h3d1bda3a),
	.w2(32'h3c900b65),
	.w3(32'h3b982254),
	.w4(32'hbc4876c4),
	.w5(32'hbbbea98d),
	.w6(32'hbbbe9666),
	.w7(32'hbcaa0043),
	.w8(32'hbbf2d518),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b0a5e),
	.w1(32'hbc2119ee),
	.w2(32'hbb989e76),
	.w3(32'hbc2f4091),
	.w4(32'hbbb1cf47),
	.w5(32'hbc0945ce),
	.w6(32'h3c9f9d6e),
	.w7(32'h3c6bdcaf),
	.w8(32'h3c55ef67),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad81628),
	.w1(32'hba4e5ffe),
	.w2(32'h3a9c3694),
	.w3(32'hbadb1a6c),
	.w4(32'h3b1b9d0b),
	.w5(32'hbaf21c5b),
	.w6(32'h3b630fdd),
	.w7(32'h3b3e1231),
	.w8(32'hbb4b2dfc),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f5609),
	.w1(32'hbb61183f),
	.w2(32'h3680ae9a),
	.w3(32'h3a79a010),
	.w4(32'h3a836bbc),
	.w5(32'h39d07489),
	.w6(32'hb9cdd030),
	.w7(32'h399a870c),
	.w8(32'hb9e22967),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ace7e),
	.w1(32'hbb050d10),
	.w2(32'h3ae75195),
	.w3(32'h3b0135e9),
	.w4(32'hbb44a766),
	.w5(32'hb6cb7741),
	.w6(32'h37a62063),
	.w7(32'h3b8a5726),
	.w8(32'h3b34783b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53019f),
	.w1(32'h3ab6d261),
	.w2(32'hbc48b158),
	.w3(32'h3aba6676),
	.w4(32'h3b479fd8),
	.w5(32'hba938698),
	.w6(32'h3ba06005),
	.w7(32'h3c153f7b),
	.w8(32'h3ba958e4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba30f46),
	.w1(32'hbbc3fc83),
	.w2(32'hbb96f331),
	.w3(32'h3b68ddf5),
	.w4(32'hbb0599d2),
	.w5(32'hbc726134),
	.w6(32'h3b326702),
	.w7(32'hbb591aec),
	.w8(32'hbb2840c9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d86785c),
	.w1(32'h3d402b04),
	.w2(32'hbb0b1b02),
	.w3(32'h3c6175bc),
	.w4(32'h3bd8ce3b),
	.w5(32'hbcd13c76),
	.w6(32'hbbe0fd5d),
	.w7(32'hbcb8d240),
	.w8(32'hbd5963f4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d5011),
	.w1(32'h3c018f4d),
	.w2(32'hbb886358),
	.w3(32'h3b2a6138),
	.w4(32'h3a63805b),
	.w5(32'h3b5de6b8),
	.w6(32'hb85ddce3),
	.w7(32'hbb92308e),
	.w8(32'hbbe76ff2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca765f),
	.w1(32'hbb8f8393),
	.w2(32'h3c6b1c8c),
	.w3(32'hbc37f234),
	.w4(32'hbbb2bc35),
	.w5(32'h3c81e86c),
	.w6(32'hbc899f0f),
	.w7(32'h3ca1a387),
	.w8(32'h3cb94d1b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac0e4a),
	.w1(32'hbc1a9a2e),
	.w2(32'hbc22cea0),
	.w3(32'h3ab3ab2f),
	.w4(32'hb921ff57),
	.w5(32'hbb538d40),
	.w6(32'h3c80fb0d),
	.w7(32'h3a49f8ac),
	.w8(32'hbb0b1dc3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d0b0e),
	.w1(32'h3cd1ac99),
	.w2(32'hbc891cf9),
	.w3(32'h3c787673),
	.w4(32'hbac8e684),
	.w5(32'hbce9411d),
	.w6(32'h3be98ee1),
	.w7(32'hbc4dc96b),
	.w8(32'hbd3283e8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb34fd9),
	.w1(32'hbc20fd93),
	.w2(32'hbbe45f57),
	.w3(32'hba97dcf1),
	.w4(32'h38fb4a47),
	.w5(32'hbb4ebd76),
	.w6(32'hbab91940),
	.w7(32'h3b8d995b),
	.w8(32'h3b7fb481),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28fab0),
	.w1(32'hbac3c5c4),
	.w2(32'h3b98a4fb),
	.w3(32'hbacf8e6f),
	.w4(32'h3c2f9465),
	.w5(32'h3c9d42eb),
	.w6(32'h3a89c737),
	.w7(32'h3bda5acb),
	.w8(32'h3cb26966),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d27b30a),
	.w1(32'h3ce6fed6),
	.w2(32'hbb7999a0),
	.w3(32'h3c9802a8),
	.w4(32'h3c29e1a6),
	.w5(32'h3b951cfa),
	.w6(32'h3bf32c6d),
	.w7(32'hbb9bafc9),
	.w8(32'h3a51e632),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba831883),
	.w1(32'h3b1933dc),
	.w2(32'h3b227456),
	.w3(32'h3ab68f6c),
	.w4(32'hba2c80f3),
	.w5(32'hbbce5c47),
	.w6(32'h3ba0276f),
	.w7(32'h3ab8ea41),
	.w8(32'h39fead49),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1b84d7),
	.w1(32'h3cac0a60),
	.w2(32'h3c637c56),
	.w3(32'hbd51aab7),
	.w4(32'hbd3853b4),
	.w5(32'h3d0db6d7),
	.w6(32'h3d1008c0),
	.w7(32'h3cda13c8),
	.w8(32'hbc99ceec),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50a736),
	.w1(32'h3c05c3a0),
	.w2(32'h3b218050),
	.w3(32'h3c303ef6),
	.w4(32'hba52a664),
	.w5(32'hbc2cc656),
	.w6(32'h3c13cf10),
	.w7(32'hbc4a5c2d),
	.w8(32'hbc8a3de6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0b4c6),
	.w1(32'hbb5e7e5c),
	.w2(32'h3b936044),
	.w3(32'hbb56b164),
	.w4(32'h3bbd432d),
	.w5(32'h3b1b7fc2),
	.w6(32'hbbce7793),
	.w7(32'h3c09b6e5),
	.w8(32'h3c5d7b27),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c74af),
	.w1(32'hbc6486c3),
	.w2(32'hb994d393),
	.w3(32'h3ae05cfd),
	.w4(32'h3b4399c6),
	.w5(32'h3b33329a),
	.w6(32'h3c76515c),
	.w7(32'h3b3cc960),
	.w8(32'h3abefb86),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe8062),
	.w1(32'hb98f4388),
	.w2(32'hbb872c99),
	.w3(32'h3a0c3b51),
	.w4(32'hbb7a49cc),
	.w5(32'h3a94b66c),
	.w6(32'h3abab423),
	.w7(32'h3bad4429),
	.w8(32'h3c3b8c75),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19d423),
	.w1(32'hbbbcc585),
	.w2(32'hb9cf3695),
	.w3(32'hbbb45f17),
	.w4(32'hb80c7849),
	.w5(32'h3b757553),
	.w6(32'h3ba44add),
	.w7(32'hbc415b79),
	.w8(32'hbbef3baa),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacb9fd),
	.w1(32'h3bf90747),
	.w2(32'h3ad6bafe),
	.w3(32'h3b6962f4),
	.w4(32'hbc02cf20),
	.w5(32'hbc1b3350),
	.w6(32'hbc149446),
	.w7(32'hba3b4519),
	.w8(32'h3a79fabb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e91cc),
	.w1(32'hbbaf816d),
	.w2(32'hbaee0f8a),
	.w3(32'hbc5a0865),
	.w4(32'hb9cb1185),
	.w5(32'h3b1b4007),
	.w6(32'h3c04a9fd),
	.w7(32'h3bcc8fe9),
	.w8(32'h3bbca3d3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9155c),
	.w1(32'h3c2466d7),
	.w2(32'hba79ce9b),
	.w3(32'h3c4416f5),
	.w4(32'hbb8b0c5e),
	.w5(32'hbc3909bf),
	.w6(32'h3c01603e),
	.w7(32'hbc25c6c7),
	.w8(32'hbca8585f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc368ba1),
	.w1(32'hbc1dded1),
	.w2(32'hbb6164a0),
	.w3(32'hbc639d21),
	.w4(32'h391d41b1),
	.w5(32'h38eb6537),
	.w6(32'hbc912b38),
	.w7(32'hbc13cb35),
	.w8(32'hbc2617ed),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb06d2),
	.w1(32'hbbb5605b),
	.w2(32'hbba86e20),
	.w3(32'h3b27d5c1),
	.w4(32'hbb64fb14),
	.w5(32'h3c556a46),
	.w6(32'hbc4ae9f6),
	.w7(32'hbc1db97a),
	.w8(32'h3bb08df1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ce994),
	.w1(32'h3c80e10a),
	.w2(32'hbb50b082),
	.w3(32'h3bb8a789),
	.w4(32'h3b1f0445),
	.w5(32'h3aaddeb9),
	.w6(32'h3c225b8e),
	.w7(32'h3c3e8210),
	.w8(32'h3c885961),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cd867),
	.w1(32'h3b917984),
	.w2(32'h3adc5032),
	.w3(32'h3b20c8cf),
	.w4(32'h3c8ad262),
	.w5(32'h3c8d4697),
	.w6(32'h3c8438c2),
	.w7(32'h3cd0e619),
	.w8(32'h3d1732ea),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2dfcb1),
	.w1(32'h3d1b7be4),
	.w2(32'h3c821f0d),
	.w3(32'h3d114921),
	.w4(32'h3b92a9f3),
	.w5(32'h3a349eae),
	.w6(32'h3d2ee6ec),
	.w7(32'hbb36f1de),
	.w8(32'h3b88a5a2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c2f1e),
	.w1(32'hba963bfb),
	.w2(32'hbc050b09),
	.w3(32'hbaa62202),
	.w4(32'h3ae58f3e),
	.w5(32'h3bded590),
	.w6(32'hba5c0e5e),
	.w7(32'h3bd8357f),
	.w8(32'hbb19061a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e5349),
	.w1(32'hbc1cff41),
	.w2(32'h3c31eabd),
	.w3(32'h3bbdf12d),
	.w4(32'h3ba57c4f),
	.w5(32'hb9fb3f81),
	.w6(32'h3b0a9f2a),
	.w7(32'h3c48f917),
	.w8(32'h3c19ce58),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c348cfd),
	.w1(32'h3c21049b),
	.w2(32'h3b3d8a91),
	.w3(32'h3be648b4),
	.w4(32'h3b9c1963),
	.w5(32'hbaa27304),
	.w6(32'h3c501c99),
	.w7(32'h3c2c27e0),
	.w8(32'h39d94c8c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b375f),
	.w1(32'h3c972a12),
	.w2(32'hbb8a320e),
	.w3(32'h3b838e66),
	.w4(32'h3a9759b2),
	.w5(32'hbca1e132),
	.w6(32'hbbbf3a5a),
	.w7(32'hbc7e8c1d),
	.w8(32'hbcf25eae),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cb11b),
	.w1(32'h3abfc553),
	.w2(32'hbc263728),
	.w3(32'hbbc4e835),
	.w4(32'hbaf5f3cc),
	.w5(32'hbc810c60),
	.w6(32'hbb88b91e),
	.w7(32'h390f4ece),
	.w8(32'hbc2ed6db),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399546e2),
	.w1(32'h3bf0eff1),
	.w2(32'hbbaf5031),
	.w3(32'hbc173141),
	.w4(32'h3bf6c642),
	.w5(32'h3b0abc98),
	.w6(32'hbb6f619c),
	.w7(32'h3c23dbcb),
	.w8(32'h3c3075b9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c524f),
	.w1(32'h3c8f1a6b),
	.w2(32'hbc18766c),
	.w3(32'h38d2f031),
	.w4(32'h3c34f7f9),
	.w5(32'hbc221713),
	.w6(32'h3bf40930),
	.w7(32'hbc3a1161),
	.w8(32'hbcc727aa),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdc907),
	.w1(32'h3b87c28f),
	.w2(32'hba82f737),
	.w3(32'hbc170212),
	.w4(32'hbb838b22),
	.w5(32'hba5694bb),
	.w6(32'hbc0fddd0),
	.w7(32'hbb1c18c0),
	.w8(32'hbb1691f0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b416d),
	.w1(32'h3c03eafc),
	.w2(32'hbb0555c0),
	.w3(32'h3c12725a),
	.w4(32'hbb43103b),
	.w5(32'hbc1fff1c),
	.w6(32'hbb897d96),
	.w7(32'hbc15b775),
	.w8(32'hbc07c20f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bb964),
	.w1(32'hbbdb7006),
	.w2(32'h3aa39296),
	.w3(32'hbcc88c2b),
	.w4(32'hbcd6aaf2),
	.w5(32'hbc026fdf),
	.w6(32'hbca0e6f9),
	.w7(32'hbcd17af5),
	.w8(32'hbc4c6ea3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb30c8),
	.w1(32'h3ca92356),
	.w2(32'h3a24853b),
	.w3(32'h3cb63aff),
	.w4(32'h3d01f214),
	.w5(32'h3b587097),
	.w6(32'hbc933eca),
	.w7(32'hbc1f41e0),
	.w8(32'hbc9b7ae4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6f8da),
	.w1(32'h3b19ccd7),
	.w2(32'hbb4f2180),
	.w3(32'h3c505fe3),
	.w4(32'h3bf9e6d3),
	.w5(32'h3b0c027c),
	.w6(32'h3c194753),
	.w7(32'h3b09a94e),
	.w8(32'hbb2af5bc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c0bf3),
	.w1(32'h3c40df13),
	.w2(32'hbad8ba2c),
	.w3(32'h3bd2a906),
	.w4(32'h3a732b94),
	.w5(32'hbc84440a),
	.w6(32'h3c6b0f04),
	.w7(32'h3bfb1f65),
	.w8(32'hbc0acf7e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b5407),
	.w1(32'hba88cb06),
	.w2(32'h3b9dd9ba),
	.w3(32'hba13bed3),
	.w4(32'h3bd044c9),
	.w5(32'h3b28cc1c),
	.w6(32'hbab34b76),
	.w7(32'h3a4ef3c1),
	.w8(32'h3c018887),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7f81c),
	.w1(32'h3d129f92),
	.w2(32'hb99000d4),
	.w3(32'hbb9224db),
	.w4(32'hbaa6b31a),
	.w5(32'hbca859bc),
	.w6(32'h3ce2845a),
	.w7(32'hbb4f6cb2),
	.w8(32'hbcebbcf2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3e76f),
	.w1(32'hbbc0d59d),
	.w2(32'hbc04f378),
	.w3(32'hbbc9cf55),
	.w4(32'h3ad50566),
	.w5(32'h3b02c183),
	.w6(32'hbabaa8f9),
	.w7(32'h3ca59686),
	.w8(32'h3c848586),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc10408),
	.w1(32'h3a910fca),
	.w2(32'h3b787b0f),
	.w3(32'h3ca28b6f),
	.w4(32'h3bd01283),
	.w5(32'hbaf0908b),
	.w6(32'h3c3b1839),
	.w7(32'h3c259c88),
	.w8(32'h3a257cee),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9916f),
	.w1(32'h3bb16ac2),
	.w2(32'h3b1f8027),
	.w3(32'h3bcbc9e0),
	.w4(32'h3c2c6e10),
	.w5(32'hbafbddb6),
	.w6(32'h3c41f41e),
	.w7(32'h3c4213be),
	.w8(32'hbbc61595),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f2789),
	.w1(32'h3a9cc6fc),
	.w2(32'h3b2920de),
	.w3(32'h3a658743),
	.w4(32'hbb594df4),
	.w5(32'hbb66f8c6),
	.w6(32'h3a9c9f50),
	.w7(32'h3b805e38),
	.w8(32'h3be0a74f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0740f1),
	.w1(32'h3c19f9c1),
	.w2(32'hbb8895d0),
	.w3(32'h3b38f329),
	.w4(32'hbc3ada08),
	.w5(32'hbc19f67b),
	.w6(32'h3bfe32c2),
	.w7(32'h381de4f8),
	.w8(32'hbb064b64),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe48453),
	.w1(32'hbbe94177),
	.w2(32'h3a887bca),
	.w3(32'hba1fd1f6),
	.w4(32'hba753fd1),
	.w5(32'hbb8f9154),
	.w6(32'h3c29fe89),
	.w7(32'hbc09090e),
	.w8(32'hbc438b6f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8afafa),
	.w1(32'h3c97d4f4),
	.w2(32'h3c6fe2f3),
	.w3(32'h3c5c2d31),
	.w4(32'hbb2b1485),
	.w5(32'hbb3ac6d0),
	.w6(32'hbc0afa61),
	.w7(32'hbc2302b4),
	.w8(32'hbc6680bd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa17e8),
	.w1(32'hbbbb76db),
	.w2(32'hbbdb8faa),
	.w3(32'hbaf84ef0),
	.w4(32'hbb6ade65),
	.w5(32'hbb379ee6),
	.w6(32'h3b45e8bf),
	.w7(32'h3c89d8b9),
	.w8(32'h3cc78787),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfef34f),
	.w1(32'hbba10110),
	.w2(32'h3be57704),
	.w3(32'hbbb81ddb),
	.w4(32'h394a9dfa),
	.w5(32'h3b7b701e),
	.w6(32'h3c96b700),
	.w7(32'h3c0f6871),
	.w8(32'h3c43c613),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c337cf7),
	.w1(32'h3c0c2311),
	.w2(32'hbb86a496),
	.w3(32'h3bcbc779),
	.w4(32'h3b1444e9),
	.w5(32'h3be93788),
	.w6(32'h3c637a24),
	.w7(32'hbbdbbb64),
	.w8(32'hbab47056),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c156784),
	.w1(32'h3ac31d08),
	.w2(32'hbabb1e3b),
	.w3(32'h3b044ed5),
	.w4(32'hbaa00b53),
	.w5(32'h3ba13e05),
	.w6(32'hbb98eb3d),
	.w7(32'hbafb6185),
	.w8(32'h3bba7883),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7242e2),
	.w1(32'h3bdc7450),
	.w2(32'h3aef6c06),
	.w3(32'hbbd224d8),
	.w4(32'hbbd9844e),
	.w5(32'hbb69c4d8),
	.w6(32'h3bde1e1d),
	.w7(32'hbbebb129),
	.w8(32'hbb379bef),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e7c2c),
	.w1(32'hbbad5475),
	.w2(32'h3ba3a3e3),
	.w3(32'hbb01a740),
	.w4(32'hbb3d089e),
	.w5(32'hbbef6c80),
	.w6(32'hbb039184),
	.w7(32'hbb94dad0),
	.w8(32'hbbf326de),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9b4da),
	.w1(32'h3ca78df8),
	.w2(32'h3c651339),
	.w3(32'hbbf5ec7b),
	.w4(32'h3c30205e),
	.w5(32'h3c5bb7e7),
	.w6(32'h3b02cbec),
	.w7(32'hbb6c45d3),
	.w8(32'hbcd46a00),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac974ce),
	.w1(32'hbb83664e),
	.w2(32'h3a796ddc),
	.w3(32'hbaacfb78),
	.w4(32'hbc2a731b),
	.w5(32'hbba3d0ec),
	.w6(32'hbb3e65d7),
	.w7(32'hbb992547),
	.w8(32'hbbf9a0e7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0795f),
	.w1(32'hbbbf8282),
	.w2(32'h3bdd4b92),
	.w3(32'hbb43e35d),
	.w4(32'h3b724aa8),
	.w5(32'h3a03ca30),
	.w6(32'hbbabd1bf),
	.w7(32'h3c40b4c8),
	.w8(32'h3c4c9e68),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e5627),
	.w1(32'h3b8737d3),
	.w2(32'hbbda94e4),
	.w3(32'hbb889ead),
	.w4(32'hb9e1bbfe),
	.w5(32'hb9691180),
	.w6(32'h3b8c654a),
	.w7(32'hbc2c32b1),
	.w8(32'hbc234a43),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba985d68),
	.w1(32'hbb31b525),
	.w2(32'h3bbec62d),
	.w3(32'hbb3c6096),
	.w4(32'hbcacc5ee),
	.w5(32'hbca2163c),
	.w6(32'hbc06c485),
	.w7(32'h3ad22cf3),
	.w8(32'hbbc73fd1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb41cbc),
	.w1(32'h3b88a6f4),
	.w2(32'hba337cd3),
	.w3(32'h397571de),
	.w4(32'h3b97051b),
	.w5(32'h3ba7ac8f),
	.w6(32'hbb364096),
	.w7(32'hb8b4c1f4),
	.w8(32'h3b24aba6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cb382),
	.w1(32'h3bc46ce9),
	.w2(32'h39934f93),
	.w3(32'hbaa7cc15),
	.w4(32'h3a3a15fc),
	.w5(32'hbbc788e0),
	.w6(32'h3b82a5a8),
	.w7(32'hbb139bc4),
	.w8(32'hbbbe20c2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03f90f),
	.w1(32'hbbb1170f),
	.w2(32'hb8963449),
	.w3(32'h3a419d44),
	.w4(32'hb7970e8a),
	.w5(32'hb8c8faa9),
	.w6(32'h3a874f94),
	.w7(32'hb88754c9),
	.w8(32'hb8e03500),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9fd77d),
	.w1(32'h3c877ef2),
	.w2(32'h3b5e9aea),
	.w3(32'h3bedfbaa),
	.w4(32'h3bb165b1),
	.w5(32'hb9c96668),
	.w6(32'h3b337810),
	.w7(32'hbc154bdd),
	.w8(32'hbc6f08f7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafd137),
	.w1(32'h3bbfdc5e),
	.w2(32'hbbe3125d),
	.w3(32'h3b605eba),
	.w4(32'hbb3d2a5d),
	.w5(32'hbc4c89db),
	.w6(32'h3baaa521),
	.w7(32'hbb08bf93),
	.w8(32'hbc2f6d2b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b47b5),
	.w1(32'hba5c35e6),
	.w2(32'hba351d3f),
	.w3(32'hbaa7a85e),
	.w4(32'hba80e95f),
	.w5(32'hba86b9f3),
	.w6(32'hba28ca41),
	.w7(32'hb86f3bf8),
	.w8(32'hb9d0a4cb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8949761),
	.w1(32'hb929f7af),
	.w2(32'hb9fdcf5e),
	.w3(32'hb8271e52),
	.w4(32'hb8e98f5d),
	.w5(32'hb9dd4144),
	.w6(32'hb909f516),
	.w7(32'hb9014cad),
	.w8(32'hb9ae075c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83aed9),
	.w1(32'hbb92be78),
	.w2(32'h3a9b0ef7),
	.w3(32'h38834682),
	.w4(32'h3a3d14bb),
	.w5(32'h3b9ae7c9),
	.w6(32'h3b70cff3),
	.w7(32'h3bc5ce06),
	.w8(32'h3bacfb22),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41ccc6),
	.w1(32'h3c66809b),
	.w2(32'h3b804dc1),
	.w3(32'h3b9ad6d0),
	.w4(32'h3bc11ba2),
	.w5(32'hb98d7dfc),
	.w6(32'hbad2ba73),
	.w7(32'hbc13f4c6),
	.w8(32'hbc40e378),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1177cd),
	.w1(32'h3ceda036),
	.w2(32'h3cffed49),
	.w3(32'h3ca205d7),
	.w4(32'h3b8eb0e8),
	.w5(32'h3c4d3e66),
	.w6(32'h3b57084f),
	.w7(32'hbc441d83),
	.w8(32'h3ba4a581),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce5e8bd),
	.w1(32'h3ccdb1ed),
	.w2(32'hb9aa3221),
	.w3(32'h3c097f89),
	.w4(32'h3bc1a432),
	.w5(32'hbc128016),
	.w6(32'hbb0f9a36),
	.w7(32'hbc8c2334),
	.w8(32'hbcde0c08),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7553e),
	.w1(32'h3b3cf58c),
	.w2(32'hb857ef28),
	.w3(32'h3bc20e6d),
	.w4(32'h3bb8fffb),
	.w5(32'h3b62691e),
	.w6(32'hbb37659e),
	.w7(32'hba92929f),
	.w8(32'hbac31dc1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e60b66),
	.w1(32'h391f30ad),
	.w2(32'hb90834a1),
	.w3(32'h38cd724f),
	.w4(32'hb7cb97bd),
	.w5(32'hb99f2721),
	.w6(32'h38158a26),
	.w7(32'h386e6431),
	.w8(32'h3810df58),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e33cb3),
	.w1(32'h38eb139b),
	.w2(32'hb6aa0289),
	.w3(32'h38ef570b),
	.w4(32'h38dd152f),
	.w5(32'hb7bc7bb8),
	.w6(32'h386a9891),
	.w7(32'h38527384),
	.w8(32'hb7c8a16a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389820b5),
	.w1(32'h3894eec7),
	.w2(32'h38ecb9bb),
	.w3(32'h391c5735),
	.w4(32'h38dc1125),
	.w5(32'hb6ad313b),
	.w6(32'h3955405e),
	.w7(32'h3991b9c1),
	.w8(32'h3919ce94),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d62e4d),
	.w1(32'h3b1edbf4),
	.w2(32'h3b2d7aa1),
	.w3(32'h3a8d00aa),
	.w4(32'h3b5a7e03),
	.w5(32'h3ab03761),
	.w6(32'h3a939c6f),
	.w7(32'h3b3d9f94),
	.w8(32'h394afa7b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7d40f),
	.w1(32'h3b50bffa),
	.w2(32'h3a8eb5bc),
	.w3(32'h3b7f8a3d),
	.w4(32'h3b8748a9),
	.w5(32'h3b93eeff),
	.w6(32'h3b8d545c),
	.w7(32'h3b9d8561),
	.w8(32'h3b958160),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab4a65),
	.w1(32'hba00e932),
	.w2(32'h3aeee93e),
	.w3(32'hbab57d5b),
	.w4(32'hba7c1d6c),
	.w5(32'h3a2a342e),
	.w6(32'hb9e1b7c7),
	.w7(32'h3a3715f5),
	.w8(32'h3af45a6d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45f63a),
	.w1(32'hbb959095),
	.w2(32'h3a312b0b),
	.w3(32'hba319ede),
	.w4(32'h3ac92665),
	.w5(32'h3b827fc4),
	.w6(32'h3b63135f),
	.w7(32'h3bce9029),
	.w8(32'h3bce7a3b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd19281),
	.w1(32'h3bb54829),
	.w2(32'h3af19a07),
	.w3(32'h3b73be10),
	.w4(32'h3ac77c65),
	.w5(32'hbb44db08),
	.w6(32'h39443251),
	.w7(32'hbb360d2f),
	.w8(32'hbba18dc2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8939e55),
	.w1(32'hbb13f0cc),
	.w2(32'hbb69e5c2),
	.w3(32'hbb095675),
	.w4(32'hbb981f2a),
	.w5(32'hbb95e985),
	.w6(32'h3affc51c),
	.w7(32'hb9e17e93),
	.w8(32'hb93d57d4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1aee1),
	.w1(32'h3bff4d11),
	.w2(32'h3bb54035),
	.w3(32'h3ae49a9b),
	.w4(32'h3ba89704),
	.w5(32'h3ac3abff),
	.w6(32'h3b74e577),
	.w7(32'h3b9c6dba),
	.w8(32'hbb04a4a4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f5642),
	.w1(32'h3b90c824),
	.w2(32'hbb8030cb),
	.w3(32'h39e59d3a),
	.w4(32'hbaf7c3ba),
	.w5(32'hbc1aff37),
	.w6(32'hbc092ef8),
	.w7(32'hbc043937),
	.w8(32'hbc1cda9a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3813be07),
	.w1(32'h38c2084b),
	.w2(32'hb8954222),
	.w3(32'h37e59036),
	.w4(32'h38b640dd),
	.w5(32'hb8d5a421),
	.w6(32'h38beb2fa),
	.w7(32'h39341dcf),
	.w8(32'hb825f50e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d53300),
	.w1(32'hb9426ab7),
	.w2(32'hb90ac5f8),
	.w3(32'hb919c5e2),
	.w4(32'h38fb21f0),
	.w5(32'h390e0406),
	.w6(32'hb8a1baaa),
	.w7(32'h38fa71d8),
	.w8(32'hb7cea453),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959d1f1),
	.w1(32'hb9382e59),
	.w2(32'hb8c4dbde),
	.w3(32'hb8cdc41f),
	.w4(32'h36a97853),
	.w5(32'h384f2e44),
	.w6(32'hb64079dc),
	.w7(32'h38d037f5),
	.w8(32'h388c55df),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3941c0cb),
	.w1(32'h391aeca5),
	.w2(32'h39f71e1b),
	.w3(32'h3a0bbd3f),
	.w4(32'h3a68240d),
	.w5(32'h3a60a5cd),
	.w6(32'h3940bef8),
	.w7(32'h3a0ac1ed),
	.w8(32'h3a330b7d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab24793),
	.w1(32'hba978825),
	.w2(32'h38524e33),
	.w3(32'hb9f3b848),
	.w4(32'hb9ebd632),
	.w5(32'h3a71d6f7),
	.w6(32'h3b0dad4b),
	.w7(32'h3ac13ce8),
	.w8(32'h39860ae3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46d5af),
	.w1(32'hba04fcd7),
	.w2(32'h3a293b3d),
	.w3(32'hbb17e93e),
	.w4(32'hbafddd06),
	.w5(32'hba18433e),
	.w6(32'hbafdd0be),
	.w7(32'hbaf45f81),
	.w8(32'hba8f98de),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab60c3e),
	.w1(32'hbc3a0b9c),
	.w2(32'hbc00a65f),
	.w3(32'hbb4216c4),
	.w4(32'hbb94e07b),
	.w5(32'hb9e7c2d7),
	.w6(32'hbab76566),
	.w7(32'h3afa4173),
	.w8(32'h3bd2ba68),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf2255),
	.w1(32'hbba3da26),
	.w2(32'hbb29205e),
	.w3(32'hbb6f3304),
	.w4(32'hbb373c87),
	.w5(32'hba3fd9e2),
	.w6(32'h39508f7b),
	.w7(32'h3ac8733a),
	.w8(32'h3b103851),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05cd6d),
	.w1(32'h3c42bb4c),
	.w2(32'hbafcef56),
	.w3(32'h3b62cb02),
	.w4(32'h3bd52875),
	.w5(32'hbb17cfa1),
	.w6(32'h3a9c97ca),
	.w7(32'hbb8cb385),
	.w8(32'hbc7d8eaf),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b46dc),
	.w1(32'h3b6d62f0),
	.w2(32'h3a15f023),
	.w3(32'h3a533c28),
	.w4(32'h3b12893e),
	.w5(32'h39cc1dfb),
	.w6(32'hb88dc058),
	.w7(32'h3954bed7),
	.w8(32'hba691db5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb961c28),
	.w1(32'hbb85590b),
	.w2(32'hbb1216e2),
	.w3(32'hbb150349),
	.w4(32'h39be9473),
	.w5(32'h3a8aec1b),
	.w6(32'h3aa8006b),
	.w7(32'h3b78919a),
	.w8(32'h3b679d32),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa65ed),
	.w1(32'hbb0a30e0),
	.w2(32'h3aae1c18),
	.w3(32'h3a338b98),
	.w4(32'h398bf169),
	.w5(32'h3b22c52f),
	.w6(32'h3b30f9bf),
	.w7(32'h3b48e28a),
	.w8(32'h3b808a1f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878853),
	.w1(32'hb99d7b85),
	.w2(32'hbb726501),
	.w3(32'hbb60281a),
	.w4(32'hbb94e2d3),
	.w5(32'hbbc91115),
	.w6(32'hb9b9c17d),
	.w7(32'h35ca670e),
	.w8(32'hbb916495),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bfc4a),
	.w1(32'h3b819bf7),
	.w2(32'h3b82dab0),
	.w3(32'hbb080fcc),
	.w4(32'hbb8ac5f1),
	.w5(32'hba8434bf),
	.w6(32'h3b4679d7),
	.w7(32'h3ac6f553),
	.w8(32'h3b6f0584),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf86eb),
	.w1(32'h3b840196),
	.w2(32'h3b86c497),
	.w3(32'hba4f37a1),
	.w4(32'hba837838),
	.w5(32'h3b28cae7),
	.w6(32'h3a2753b2),
	.w7(32'h3abe9c05),
	.w8(32'h3b4a8b8c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ffee7),
	.w1(32'hbc4763e9),
	.w2(32'hbbfeb5ce),
	.w3(32'hbbbf20cc),
	.w4(32'hbbe14c1e),
	.w5(32'hbb4531ce),
	.w6(32'h3adf6f92),
	.w7(32'h39e9526a),
	.w8(32'h3b1ec1bd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68077d),
	.w1(32'h3a0cb198),
	.w2(32'h3862c50f),
	.w3(32'h3a6ee1de),
	.w4(32'h3a20e3ae),
	.w5(32'h39a8a422),
	.w6(32'h3997e36f),
	.w7(32'h3a0381e3),
	.w8(32'h3a19a218),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d928f),
	.w1(32'h3b0daa81),
	.w2(32'h396f40b0),
	.w3(32'h3b5423bb),
	.w4(32'h3b437870),
	.w5(32'h39ef5ba5),
	.w6(32'h3ac8f957),
	.w7(32'h3aa719cf),
	.w8(32'hba191e27),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac629fe),
	.w1(32'hba9dd440),
	.w2(32'hb983ef34),
	.w3(32'hbb8085ae),
	.w4(32'hbb4fb306),
	.w5(32'hbb0977ba),
	.w6(32'hbb8fdbcb),
	.w7(32'hbb253e0d),
	.w8(32'hbaf3a935),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46031e),
	.w1(32'hbadcd3ef),
	.w2(32'h3a16a392),
	.w3(32'hba550a21),
	.w4(32'h3ac33d05),
	.w5(32'h3b00bb58),
	.w6(32'h3b564e51),
	.w7(32'h3bafd334),
	.w8(32'h3b81a511),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0440a),
	.w1(32'h3c1a1080),
	.w2(32'h3b8d81f6),
	.w3(32'h3b943846),
	.w4(32'h3b6301ce),
	.w5(32'h3a0bb632),
	.w6(32'h3b2f22eb),
	.w7(32'hbb96b4a8),
	.w8(32'hbbd6f07b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ae660),
	.w1(32'hb87b74dc),
	.w2(32'hb79704e3),
	.w3(32'hb7e74e09),
	.w4(32'hb7678000),
	.w5(32'hb69ada44),
	.w6(32'hb737a0d3),
	.w7(32'h3771d8aa),
	.w8(32'h35f80aa2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a15a62),
	.w1(32'h39377f27),
	.w2(32'hba5aed7b),
	.w3(32'hb9618ba5),
	.w4(32'hba330035),
	.w5(32'hbaf2c49d),
	.w6(32'hb80fbbb4),
	.w7(32'hba5c58a1),
	.w8(32'hbabad3d3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b06b0),
	.w1(32'hbb8680f9),
	.w2(32'hbbb61254),
	.w3(32'h3b1b8024),
	.w4(32'hba11acda),
	.w5(32'hbb99c5cc),
	.w6(32'h3c065c2b),
	.w7(32'h3c3cf36d),
	.w8(32'h3b94353d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41fd4e),
	.w1(32'h3b5d149d),
	.w2(32'h3aeb8293),
	.w3(32'h3b3a3603),
	.w4(32'hbb8f3739),
	.w5(32'hbb5354ce),
	.w6(32'h3b512ecb),
	.w7(32'h3a559d90),
	.w8(32'h3acb8e23),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaccf55),
	.w1(32'h3a3e0e34),
	.w2(32'h3aa53c1b),
	.w3(32'h3af4eb44),
	.w4(32'h3ac5d97f),
	.w5(32'h3acd25d5),
	.w6(32'h3b07bf1f),
	.w7(32'h3b40b6a1),
	.w8(32'h3b1f7256),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11bceb),
	.w1(32'hbb82fa88),
	.w2(32'h3a1794c8),
	.w3(32'hb9c093ae),
	.w4(32'hbab8de13),
	.w5(32'h3afa8d5b),
	.w6(32'h3ad82c56),
	.w7(32'h3a745238),
	.w8(32'h3b84def7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb619332),
	.w1(32'hbb88c48d),
	.w2(32'hbb03601d),
	.w3(32'hbb875f6c),
	.w4(32'hbb97f754),
	.w5(32'hbb155d05),
	.w6(32'hbb9e0682),
	.w7(32'hbb8d1def),
	.w8(32'hbb28b3be),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8070a),
	.w1(32'h3ade8cf0),
	.w2(32'h3b7c6363),
	.w3(32'hbb524961),
	.w4(32'h3b63beee),
	.w5(32'h3a8bd3e4),
	.w6(32'h3b067890),
	.w7(32'h3abc2267),
	.w8(32'hbb20e6fe),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada67e1),
	.w1(32'hba9d3885),
	.w2(32'hbb8059c5),
	.w3(32'hbb2742ed),
	.w4(32'hbbe0b598),
	.w5(32'hbbddc82f),
	.w6(32'hba8b3ab9),
	.w7(32'hbb4eaca9),
	.w8(32'hba85d2b3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb878718),
	.w1(32'h3b85d3da),
	.w2(32'h3b43c1e8),
	.w3(32'hb8afeb31),
	.w4(32'h3bcb66c1),
	.w5(32'h3ac93eec),
	.w6(32'h3b854230),
	.w7(32'h3b90f88e),
	.w8(32'hbb290e52),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule