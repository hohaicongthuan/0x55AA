module layer_10_featuremap_260(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9714e7),
	.w1(32'hbba86a2b),
	.w2(32'hba7f45d0),
	.w3(32'hbb967ecd),
	.w4(32'h3bbda984),
	.w5(32'hbb2eab14),
	.w6(32'hbbf93d73),
	.w7(32'h3a82d690),
	.w8(32'hbb95c62d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fa0fc),
	.w1(32'h3b7497da),
	.w2(32'hbbea6384),
	.w3(32'hbab91aeb),
	.w4(32'hba30c32a),
	.w5(32'hbb75cd97),
	.w6(32'h3a70c95f),
	.w7(32'hbb5f7e0a),
	.w8(32'hbbff659d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b762f41),
	.w1(32'h3bdf9b35),
	.w2(32'h3b968783),
	.w3(32'h3b13a13a),
	.w4(32'hb9c8a978),
	.w5(32'h37e75994),
	.w6(32'hb926785d),
	.w7(32'hbaa57ca6),
	.w8(32'h3a368c4b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268a69),
	.w1(32'hbb8b4d3a),
	.w2(32'hbb1b3b9f),
	.w3(32'hbafa02cc),
	.w4(32'hba31a624),
	.w5(32'h3a68b40e),
	.w6(32'hbab8b6c6),
	.w7(32'h39bf20ff),
	.w8(32'hbb92c5e5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9aad4),
	.w1(32'hbbc7e4ad),
	.w2(32'hb9da5556),
	.w3(32'h3b28fa21),
	.w4(32'h3be35c14),
	.w5(32'h3a569b1b),
	.w6(32'hbb14c9e3),
	.w7(32'h3a762e63),
	.w8(32'hba81dfd3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c5694),
	.w1(32'hbba8a751),
	.w2(32'hbb5ca9d0),
	.w3(32'h3b1e2cf1),
	.w4(32'h3b6c40ab),
	.w5(32'h3bb51e17),
	.w6(32'hbae3f6f0),
	.w7(32'hb99d7d16),
	.w8(32'h3a8d5054),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b282c2f),
	.w1(32'hbbcda2c5),
	.w2(32'hbbd8c212),
	.w3(32'h3b44ac6f),
	.w4(32'hbaeace3e),
	.w5(32'hbb1e3f09),
	.w6(32'hba337c67),
	.w7(32'hbb2c1bba),
	.w8(32'h3b2daec0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b06298),
	.w1(32'hbb7c41b2),
	.w2(32'hba588ac3),
	.w3(32'hbc28e675),
	.w4(32'hbc0e5392),
	.w5(32'h39a35430),
	.w6(32'hbc342bdc),
	.w7(32'hbb309998),
	.w8(32'hbb4e05a9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7fea5),
	.w1(32'hbb26c4b8),
	.w2(32'hbb97ba17),
	.w3(32'h3a013883),
	.w4(32'h3a2a910d),
	.w5(32'hbb35b6f5),
	.w6(32'hbb7a16a6),
	.w7(32'hbb910c04),
	.w8(32'hbb9b7340),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50aaf2),
	.w1(32'hbc4c7cd8),
	.w2(32'hbc8c337d),
	.w3(32'hbbfe8dd8),
	.w4(32'hb9171f7a),
	.w5(32'hbbe348f0),
	.w6(32'hbc4f477f),
	.w7(32'hbb9df897),
	.w8(32'hbc1ae8e0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d01ab),
	.w1(32'hbbeec2c2),
	.w2(32'hbb4c93ba),
	.w3(32'hbb664de1),
	.w4(32'h3aebebec),
	.w5(32'h3b7d5d23),
	.w6(32'hbbb413e3),
	.w7(32'hbb13f246),
	.w8(32'hbc0c0e5c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b151206),
	.w1(32'h3c14a023),
	.w2(32'h3bb6aac3),
	.w3(32'h3ae54fc6),
	.w4(32'h3b0fd45a),
	.w5(32'hbc3830a9),
	.w6(32'hbb90e45e),
	.w7(32'hbb749972),
	.w8(32'hbc2b63c3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc867754),
	.w1(32'hbc3bc210),
	.w2(32'hbc6d7e9e),
	.w3(32'hbc3685e9),
	.w4(32'hbc057ff8),
	.w5(32'hbc33f909),
	.w6(32'hbbb55ff5),
	.w7(32'hbbe5df56),
	.w8(32'hbc5ac818),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1787ad),
	.w1(32'hbb68f10c),
	.w2(32'hbb5783b0),
	.w3(32'hbaeb799a),
	.w4(32'hbaf245a7),
	.w5(32'h3a5ac05f),
	.w6(32'hbab27811),
	.w7(32'hba17f528),
	.w8(32'h39e8baa9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cb6f9),
	.w1(32'hb92ebac8),
	.w2(32'h382b07cc),
	.w3(32'hbac8e8c0),
	.w4(32'h3b7d6786),
	.w5(32'hbb51e326),
	.w6(32'hbbcbd87d),
	.w7(32'h3b7144a8),
	.w8(32'hbb9c2b48),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e1c2d),
	.w1(32'hbc04362a),
	.w2(32'hbc2feaf0),
	.w3(32'hbc0ac78c),
	.w4(32'hba9d39f2),
	.w5(32'h3a250354),
	.w6(32'hbc327370),
	.w7(32'hbbe17ccd),
	.w8(32'hbbc888ef),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dc5bd),
	.w1(32'h3be36831),
	.w2(32'h3af64dd6),
	.w3(32'h3ad561bc),
	.w4(32'h3b08aad1),
	.w5(32'hbae59ef6),
	.w6(32'hbaeb5e7b),
	.w7(32'h394100e7),
	.w8(32'h3b11bae6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d55d4),
	.w1(32'hbbc546ab),
	.w2(32'hbc217be9),
	.w3(32'hbbcd2343),
	.w4(32'hbbc111e3),
	.w5(32'hbc31679e),
	.w6(32'hbb9c5815),
	.w7(32'hbaef8c7a),
	.w8(32'h3a150500),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f38b),
	.w1(32'hbbab098b),
	.w2(32'hbbc902cd),
	.w3(32'hbbcd22f9),
	.w4(32'hbba82913),
	.w5(32'hbc388cff),
	.w6(32'h3ba03cb6),
	.w7(32'h3baff688),
	.w8(32'hbc6cd34f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d3bd4),
	.w1(32'hbaf08ee0),
	.w2(32'hbb0b7dc0),
	.w3(32'hb9525bec),
	.w4(32'hbb40913a),
	.w5(32'hbb940a21),
	.w6(32'hba02ba2f),
	.w7(32'hbb646b10),
	.w8(32'hbb2aa6b3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cc293),
	.w1(32'hbaf34ec6),
	.w2(32'hbb73ad00),
	.w3(32'hbabba9ed),
	.w4(32'hbb37d2d2),
	.w5(32'h3b5f3438),
	.w6(32'hb9b7d4e6),
	.w7(32'hbb3f765b),
	.w8(32'h3b086302),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f47b7),
	.w1(32'h369a297e),
	.w2(32'h3b0cb17e),
	.w3(32'h3b9f0a90),
	.w4(32'h3c04c401),
	.w5(32'hbb4e2e5b),
	.w6(32'h392b1b90),
	.w7(32'h3c148086),
	.w8(32'hbc01512a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc146a20),
	.w1(32'h3a817697),
	.w2(32'hbc06c8eb),
	.w3(32'hbba8df87),
	.w4(32'h3ab1ff6c),
	.w5(32'hbc3ecb55),
	.w6(32'hbc47783a),
	.w7(32'hbbc758c1),
	.w8(32'hbcaf3bdb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f4dfe),
	.w1(32'hbb6615f3),
	.w2(32'hbca40e49),
	.w3(32'hbbbbdc40),
	.w4(32'hbbbc7754),
	.w5(32'hbbe95003),
	.w6(32'hbb8b3d72),
	.w7(32'hbc22e700),
	.w8(32'hbc03bb42),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8efd6a),
	.w1(32'hbbf24ac8),
	.w2(32'hbc8447ba),
	.w3(32'hbbbd6e16),
	.w4(32'hbab9f9f4),
	.w5(32'h3a695675),
	.w6(32'hbbe7b491),
	.w7(32'hbbc98bcc),
	.w8(32'hbc19a8b6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a277f),
	.w1(32'hbb148495),
	.w2(32'h3b7ffef1),
	.w3(32'h3a1a3a90),
	.w4(32'h3b6139da),
	.w5(32'h393fb17f),
	.w6(32'hbaf87f36),
	.w7(32'h3b99b6b7),
	.w8(32'hbb077ee0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9802a9),
	.w1(32'h3b0e02d7),
	.w2(32'h3bfebf44),
	.w3(32'h3b98fac8),
	.w4(32'h3b976d65),
	.w5(32'hba6de284),
	.w6(32'h3a85a8c5),
	.w7(32'h3b594691),
	.w8(32'h39e8ffdc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f21a3),
	.w1(32'h38bf515d),
	.w2(32'hbbee1f74),
	.w3(32'h3aa771f8),
	.w4(32'h3c233cef),
	.w5(32'hbab5d772),
	.w6(32'hbb1c5f5f),
	.w7(32'h3b29d9d2),
	.w8(32'hbb3cb77a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f1042),
	.w1(32'h3b677885),
	.w2(32'h3aa4c47a),
	.w3(32'h3a95c865),
	.w4(32'hbaeade35),
	.w5(32'hbb312a35),
	.w6(32'h3b0facaa),
	.w7(32'hb858a73d),
	.w8(32'hbb955d71),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8e8d7),
	.w1(32'hb8702a17),
	.w2(32'hbbc73a11),
	.w3(32'hbbd9cdd6),
	.w4(32'hbb591c37),
	.w5(32'hbc1786d0),
	.w6(32'hbc19be53),
	.w7(32'hbb69286c),
	.w8(32'hbc08d27e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc011712),
	.w1(32'hbbef6d91),
	.w2(32'h3a99861a),
	.w3(32'hbb9d9338),
	.w4(32'hbba6de08),
	.w5(32'hbb3b5e47),
	.w6(32'hbb889026),
	.w7(32'hbbdcdc3f),
	.w8(32'hbbe52f0c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc92bb7),
	.w1(32'h3c22aa2d),
	.w2(32'h3ab67f77),
	.w3(32'hba43b181),
	.w4(32'h3bb29e54),
	.w5(32'h3ab965bb),
	.w6(32'hbb9376db),
	.w7(32'hbaa83ffe),
	.w8(32'h3bcdb92a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d013b),
	.w1(32'hbba7e440),
	.w2(32'h3a163c9a),
	.w3(32'hbad82c00),
	.w4(32'h3bd8d272),
	.w5(32'hbbbee9ad),
	.w6(32'hbaf021ba),
	.w7(32'h3bbec2f1),
	.w8(32'hbbe6cbee),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc240a9e),
	.w1(32'hbb88e4e0),
	.w2(32'hbb86b726),
	.w3(32'hbb8a3e0f),
	.w4(32'hbb23c654),
	.w5(32'h3b1aa80b),
	.w6(32'hbbd582a8),
	.w7(32'h376c5bba),
	.w8(32'hba13e834),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fecb1),
	.w1(32'hbb019d75),
	.w2(32'h3aae796c),
	.w3(32'hb6c0c158),
	.w4(32'hbb945501),
	.w5(32'hbc02baf5),
	.w6(32'h3ba86804),
	.w7(32'h3a3c6157),
	.w8(32'hbb2acd22),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb511b03),
	.w1(32'hbb4a0b7d),
	.w2(32'hbbf2a708),
	.w3(32'hb99c1738),
	.w4(32'hbb9035d0),
	.w5(32'h3b400534),
	.w6(32'hba390c60),
	.w7(32'hbb5ab02a),
	.w8(32'hba13f783),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd0bc0),
	.w1(32'hbb22e5eb),
	.w2(32'hbbf19ef7),
	.w3(32'h3b92907c),
	.w4(32'h3b5435c0),
	.w5(32'h39211f2a),
	.w6(32'h3b9ad257),
	.w7(32'h3c36786e),
	.w8(32'hbbf8a720),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc027b29),
	.w1(32'h3b70c54f),
	.w2(32'h3b17f672),
	.w3(32'hbb481a43),
	.w4(32'h3c92920d),
	.w5(32'h3acbe0df),
	.w6(32'hbc132e38),
	.w7(32'h3c0f142d),
	.w8(32'hbbeec069),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70e677),
	.w1(32'h3c3da49b),
	.w2(32'hbc0f5179),
	.w3(32'hbb40b523),
	.w4(32'h3c4bb674),
	.w5(32'hbc02aa9b),
	.w6(32'hbc65f5f8),
	.w7(32'h38c9646b),
	.w8(32'hbc603104),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8c6b5),
	.w1(32'hb9c519ae),
	.w2(32'hbb0cd235),
	.w3(32'h3b18d6ac),
	.w4(32'h3ba4c5d2),
	.w5(32'hbaf41e8b),
	.w6(32'h3a8ba5e2),
	.w7(32'h3bb9151c),
	.w8(32'hbb996d69),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb961c6c),
	.w1(32'hbb1c1a1a),
	.w2(32'hbaf8069c),
	.w3(32'hbb8b6b7e),
	.w4(32'hbb8c3285),
	.w5(32'h3b4d87f8),
	.w6(32'hbb368df2),
	.w7(32'hbb5dfc3b),
	.w8(32'hbb8bcd3a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00cf50),
	.w1(32'hbb31b213),
	.w2(32'h3b877c5c),
	.w3(32'h3b8393e0),
	.w4(32'h3befa021),
	.w5(32'hba6f7679),
	.w6(32'hba9e426a),
	.w7(32'h3b18abd8),
	.w8(32'h3c2865ac),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa39e9a),
	.w1(32'hbc368174),
	.w2(32'hbc214bad),
	.w3(32'hbc476d3e),
	.w4(32'hbbc0ab14),
	.w5(32'hbac8cab7),
	.w6(32'hbaec5161),
	.w7(32'hbb62ca1a),
	.w8(32'hbab5e831),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91d5c2),
	.w1(32'h3b02927b),
	.w2(32'hbba0d104),
	.w3(32'hbbba2ebd),
	.w4(32'hbaf8b60b),
	.w5(32'hbaca739c),
	.w6(32'hbc5ef8f9),
	.w7(32'hbc0b9d25),
	.w8(32'hbc1a6db3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6d887),
	.w1(32'hbbe1be8b),
	.w2(32'hbbcc1fa2),
	.w3(32'hba914ba6),
	.w4(32'h3c5c7dac),
	.w5(32'h3a546b13),
	.w6(32'hbc6022aa),
	.w7(32'h3b76df53),
	.w8(32'hbc030e56),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a8b69),
	.w1(32'hbb89aaf5),
	.w2(32'hbc7d6f58),
	.w3(32'h3bc06b79),
	.w4(32'h3bd942e9),
	.w5(32'hbc1679f1),
	.w6(32'hbb587f52),
	.w7(32'hbb28db61),
	.w8(32'hbc7b2d0b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2e66),
	.w1(32'h3b5b3263),
	.w2(32'hba1f3fb7),
	.w3(32'hbb8f53d4),
	.w4(32'h3af990be),
	.w5(32'hbb992431),
	.w6(32'hbbb247f9),
	.w7(32'h3a406166),
	.w8(32'hbbd93ed4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb97eb2),
	.w1(32'hbc5cb596),
	.w2(32'hbc6db8a5),
	.w3(32'hbba73803),
	.w4(32'hbc49406e),
	.w5(32'hbc94b187),
	.w6(32'hbc04f936),
	.w7(32'hbc39b213),
	.w8(32'hbc88cab7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79661b),
	.w1(32'hbb0a172f),
	.w2(32'hbb85ea62),
	.w3(32'hba813375),
	.w4(32'hbb9421dd),
	.w5(32'h3b63bcac),
	.w6(32'h396c4793),
	.w7(32'hbb3f4704),
	.w8(32'hbaa3c85b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff2ecf),
	.w1(32'hbb999d09),
	.w2(32'h3b30901c),
	.w3(32'h3b8db73e),
	.w4(32'h3bcdf552),
	.w5(32'hbb8e6f47),
	.w6(32'hbb19a7bb),
	.w7(32'h3be5a817),
	.w8(32'hba826291),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46ab81),
	.w1(32'h39da7b6e),
	.w2(32'hbbda45fc),
	.w3(32'h3b86180d),
	.w4(32'hbb63059a),
	.w5(32'hbb00d55b),
	.w6(32'h3bbfe411),
	.w7(32'hbbea8071),
	.w8(32'h3b199a04),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa31c9),
	.w1(32'h3a70075e),
	.w2(32'h3ad80912),
	.w3(32'hbbc09065),
	.w4(32'hb9e42216),
	.w5(32'hbb760c26),
	.w6(32'h3b72a2a8),
	.w7(32'h3ac4ef36),
	.w8(32'hbb58161f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8d1cf),
	.w1(32'hbb28d713),
	.w2(32'hbb813c17),
	.w3(32'hbaca0310),
	.w4(32'h3b685342),
	.w5(32'hbbbee05a),
	.w6(32'hbad1ddd3),
	.w7(32'hb95a2663),
	.w8(32'hbc0ca8c5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a502a),
	.w1(32'hbb60374c),
	.w2(32'hbc10d3a5),
	.w3(32'h3a54c757),
	.w4(32'hbbf43300),
	.w5(32'hbc337635),
	.w6(32'hbb007f25),
	.w7(32'hbb7e84e5),
	.w8(32'hbc49e4c9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60da72),
	.w1(32'hbb73064b),
	.w2(32'hbba030ec),
	.w3(32'hba245af8),
	.w4(32'hb89bd380),
	.w5(32'h3a329003),
	.w6(32'hbac882fd),
	.w7(32'hbabcf77e),
	.w8(32'hbb282a41),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2badfd),
	.w1(32'h393f9adf),
	.w2(32'hb9a9e82d),
	.w3(32'hbb360388),
	.w4(32'hbb092bc3),
	.w5(32'hbb728b5d),
	.w6(32'h3b535770),
	.w7(32'h39fe1805),
	.w8(32'hbb9a4367),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8edde0),
	.w1(32'hbb304f01),
	.w2(32'hbb0a5790),
	.w3(32'hbb3a59c8),
	.w4(32'hbb936ee4),
	.w5(32'hbbb16eee),
	.w6(32'hb9d319f8),
	.w7(32'hb965d0c9),
	.w8(32'hbbd6f38d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12f65e),
	.w1(32'hbb326470),
	.w2(32'h3acb3dcc),
	.w3(32'hbb8b8bcd),
	.w4(32'hb99ebfd3),
	.w5(32'h3b9822be),
	.w6(32'hbb83b2e8),
	.w7(32'hb93fd0ad),
	.w8(32'hbaa214a2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63f086),
	.w1(32'hbaf3a756),
	.w2(32'h3b452285),
	.w3(32'h3bc83101),
	.w4(32'h3c257876),
	.w5(32'h3be3547f),
	.w6(32'hbb6d8bb5),
	.w7(32'h3bd5f86d),
	.w8(32'h3bd7e056),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a4d88),
	.w1(32'h398ace66),
	.w2(32'h3c024be7),
	.w3(32'h3c27657d),
	.w4(32'h3bae8abe),
	.w5(32'hbb2cb48c),
	.w6(32'h3c0daab3),
	.w7(32'h3c17133c),
	.w8(32'hbbab6bf5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd887d5),
	.w1(32'hbba75374),
	.w2(32'hbbc08967),
	.w3(32'hbc03a7f0),
	.w4(32'hbb60358b),
	.w5(32'hbbcaaf43),
	.w6(32'hbc55d40a),
	.w7(32'hbb578f60),
	.w8(32'hbc00803e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0df2ef),
	.w1(32'hbb6bdec4),
	.w2(32'hbb096924),
	.w3(32'hbbbc2e3d),
	.w4(32'hbb2467a4),
	.w5(32'h3b1eadcc),
	.w6(32'hbb9ecc77),
	.w7(32'hb95b7862),
	.w8(32'h3bbbcd56),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc55e40),
	.w1(32'hbb8eb4fd),
	.w2(32'hbb4a133d),
	.w3(32'h3bbf68e7),
	.w4(32'h3b910065),
	.w5(32'hb9f9c630),
	.w6(32'h3c2acaa9),
	.w7(32'h3b8f58bb),
	.w8(32'hbb93fe25),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb254521),
	.w1(32'h3a8cb369),
	.w2(32'h3b337179),
	.w3(32'hbb032063),
	.w4(32'hbaf660b0),
	.w5(32'hbb0c8c6c),
	.w6(32'hb9d6639c),
	.w7(32'h3a76d2df),
	.w8(32'hbb735479),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8b3aa),
	.w1(32'h3b1a87b8),
	.w2(32'hbaab0220),
	.w3(32'h38856acc),
	.w4(32'hbb1966ef),
	.w5(32'h376e463b),
	.w6(32'h3b2def62),
	.w7(32'hb9704227),
	.w8(32'h3a180b66),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8cdab),
	.w1(32'hbbee2118),
	.w2(32'hbbc72693),
	.w3(32'h3a596c22),
	.w4(32'h3abbd9f8),
	.w5(32'hba07d7fd),
	.w6(32'h3b64388e),
	.w7(32'hba7984cb),
	.w8(32'h3a4061d8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb596375),
	.w1(32'hbbcbbaea),
	.w2(32'hbb57ded7),
	.w3(32'hbbe9d5e8),
	.w4(32'hbc0f13ac),
	.w5(32'hbb8fad09),
	.w6(32'hbb858510),
	.w7(32'hbb04739a),
	.w8(32'hbb070580),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fbef6),
	.w1(32'h3b0fe9f3),
	.w2(32'hbc1f16a1),
	.w3(32'hbb59a529),
	.w4(32'hbb453224),
	.w5(32'hbc398f70),
	.w6(32'hbc12ee52),
	.w7(32'hbbb8fffe),
	.w8(32'hbc1e0a5f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd02e23),
	.w1(32'hbb4440d5),
	.w2(32'hbc0973ed),
	.w3(32'hbb46a2b1),
	.w4(32'h3bb6eccc),
	.w5(32'hbb9bac3c),
	.w6(32'hbc5f2b75),
	.w7(32'hbab8e60e),
	.w8(32'hbbe54d57),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b5c37),
	.w1(32'hbb379fd1),
	.w2(32'hbcbc7bb6),
	.w3(32'hbb7bea44),
	.w4(32'h3bf0d38e),
	.w5(32'hbb536edc),
	.w6(32'hbc71f86a),
	.w7(32'hbb8e4e56),
	.w8(32'hbc014269),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e14169),
	.w1(32'hbb92ead3),
	.w2(32'hbab5586d),
	.w3(32'h38a91fd6),
	.w4(32'h3b3e9870),
	.w5(32'hba664efb),
	.w6(32'h3b164f31),
	.w7(32'h3b7802a6),
	.w8(32'h3896936a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b511ec2),
	.w1(32'h3bc29228),
	.w2(32'hbb380c26),
	.w3(32'hb9fbfa4d),
	.w4(32'h3a3c5717),
	.w5(32'h3b9e8212),
	.w6(32'h38cc3d9b),
	.w7(32'hbb4ce17c),
	.w8(32'hb9b47b42),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8f63f),
	.w1(32'hb9c5b44f),
	.w2(32'hba514bbd),
	.w3(32'h3b7ba99c),
	.w4(32'h3b320b36),
	.w5(32'hbb5f2d87),
	.w6(32'hbb0d4d4d),
	.w7(32'hbae67227),
	.w8(32'hbab3b318),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb862f8b),
	.w1(32'hbb2212a5),
	.w2(32'hbbaa55a1),
	.w3(32'hbb3732f2),
	.w4(32'hbb2483e6),
	.w5(32'hbb925a7d),
	.w6(32'h39e18811),
	.w7(32'hb91e735f),
	.w8(32'hbb84d830),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39468040),
	.w1(32'h3aab0e82),
	.w2(32'h3ba9dc37),
	.w3(32'h3ae08ff3),
	.w4(32'hbb5ca297),
	.w5(32'hbc0cda77),
	.w6(32'h384d6258),
	.w7(32'hbb356605),
	.w8(32'hbb526c31),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e5fd4),
	.w1(32'hbb4b0f34),
	.w2(32'hbc0c5c65),
	.w3(32'hbbff3f07),
	.w4(32'hbc100e80),
	.w5(32'hbb417024),
	.w6(32'h39b855d5),
	.w7(32'hbb8a347e),
	.w8(32'hbb0b2f0f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc816535),
	.w1(32'hbb9b2381),
	.w2(32'hbbb1cb76),
	.w3(32'hbc40cd26),
	.w4(32'hbaad1ff9),
	.w5(32'hbb5e9f90),
	.w6(32'hbc0ff95e),
	.w7(32'hbb50fdf8),
	.w8(32'hbc36d81c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a1554),
	.w1(32'hbbe4e080),
	.w2(32'hbbfdd08d),
	.w3(32'hbbdaa380),
	.w4(32'h3b056f58),
	.w5(32'hbc256d62),
	.w6(32'hbc2e3584),
	.w7(32'hbb9790fb),
	.w8(32'hbc0989d8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb782aa1),
	.w1(32'hbab75a7f),
	.w2(32'hbbf0b588),
	.w3(32'hbbf8c6e8),
	.w4(32'hbba8ac42),
	.w5(32'hbb91cb63),
	.w6(32'hbb93a3b9),
	.w7(32'hbbad5f2d),
	.w8(32'hbb835c0b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7ca9e),
	.w1(32'hbb159f5b),
	.w2(32'hbbb06083),
	.w3(32'hb9a48e9c),
	.w4(32'hbb39fe56),
	.w5(32'hbc3de362),
	.w6(32'h3aae2cad),
	.w7(32'hbb0a82ef),
	.w8(32'hbbaa7a87),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba994206),
	.w1(32'hbb75937c),
	.w2(32'hbbfc41a8),
	.w3(32'hbc1bd171),
	.w4(32'hbc0ae258),
	.w5(32'hbb88693a),
	.w6(32'hbbbf7e57),
	.w7(32'hbbc326be),
	.w8(32'h3aee3538),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2596),
	.w1(32'hbbb99724),
	.w2(32'hbc0ad915),
	.w3(32'hbba43202),
	.w4(32'hbbb3ec0c),
	.w5(32'hbbd285d1),
	.w6(32'hbb1b962f),
	.w7(32'hbb6856d0),
	.w8(32'hbc0aa63b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81b600),
	.w1(32'hbb1d0445),
	.w2(32'hba4f25bb),
	.w3(32'hbb0ccbc2),
	.w4(32'hba880692),
	.w5(32'h3968bfe8),
	.w6(32'hbb5c932d),
	.w7(32'hbb47b02c),
	.w8(32'hba3f6c3d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51887e),
	.w1(32'h3bb63cfe),
	.w2(32'h3a81db07),
	.w3(32'h3bb9d497),
	.w4(32'hbb18fd4b),
	.w5(32'hbb052776),
	.w6(32'h3bb038d3),
	.w7(32'hbb0d7a01),
	.w8(32'hbb79be24),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e770d6),
	.w1(32'hba4dfaff),
	.w2(32'hbb10f00f),
	.w3(32'hba6e5de0),
	.w4(32'h3a83a612),
	.w5(32'hbb995366),
	.w6(32'hb996d75d),
	.w7(32'hbace11d5),
	.w8(32'hbb7fa643),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba70904),
	.w1(32'h3aa3dec0),
	.w2(32'hbb726a87),
	.w3(32'h3ac93c68),
	.w4(32'hbb065ca5),
	.w5(32'h3ada4fb0),
	.w6(32'h3b3889fd),
	.w7(32'h3a86ea52),
	.w8(32'hbbabf037),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba738b74),
	.w1(32'h3c2cb298),
	.w2(32'h3a7f9c6e),
	.w3(32'h3c1ffd07),
	.w4(32'h3b6fd15b),
	.w5(32'hba3c317d),
	.w6(32'h3acf9a07),
	.w7(32'h3ab32c04),
	.w8(32'h3829fcf4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43efda),
	.w1(32'hbb599944),
	.w2(32'hb7526ac4),
	.w3(32'hb8e79b6a),
	.w4(32'h3b590d86),
	.w5(32'h3bc957f6),
	.w6(32'h3b93ee6f),
	.w7(32'h3ba8b84b),
	.w8(32'h3b5f84ee),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7da7b7),
	.w1(32'hbab47f29),
	.w2(32'hbb0405d4),
	.w3(32'h3b4fd652),
	.w4(32'h3b984b4d),
	.w5(32'hbc10a6b4),
	.w6(32'hba8be25a),
	.w7(32'h3b6f427f),
	.w8(32'hbc2549ea),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8657d5),
	.w1(32'hbc26f0a0),
	.w2(32'hbbf3bc88),
	.w3(32'hbc5b6bf8),
	.w4(32'hba9b4370),
	.w5(32'hbbcce4c7),
	.w6(32'hbc9a67b2),
	.w7(32'hbba0b96c),
	.w8(32'hbc1df642),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e0800),
	.w1(32'h3b17e087),
	.w2(32'hbbfe7b29),
	.w3(32'hbac20594),
	.w4(32'hb8cb89a2),
	.w5(32'hba206d49),
	.w6(32'hbb13552e),
	.w7(32'hbab0fbf0),
	.w8(32'h3a21afa2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba6d25),
	.w1(32'hbae9a9f9),
	.w2(32'hbb924776),
	.w3(32'hbc155c33),
	.w4(32'h3ab97393),
	.w5(32'h3b079912),
	.w6(32'hbb845a1d),
	.w7(32'hbb09924e),
	.w8(32'hbb49ef02),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2441e4),
	.w1(32'h3c59ab00),
	.w2(32'h3be5615a),
	.w3(32'h3b0e2054),
	.w4(32'h3c656479),
	.w5(32'hbbcba790),
	.w6(32'hbc077542),
	.w7(32'h3bff06f8),
	.w8(32'h3b87bcd6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0352ae),
	.w1(32'h3c2905bd),
	.w2(32'h3b37e8ba),
	.w3(32'hbb72c7e3),
	.w4(32'h3ab66089),
	.w5(32'hbb926903),
	.w6(32'h3b6442d9),
	.w7(32'h3b73b1d6),
	.w8(32'hbc04ba6c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf74637),
	.w1(32'hbba553ec),
	.w2(32'hbb635610),
	.w3(32'hbb1fb446),
	.w4(32'h3c4e0594),
	.w5(32'h3c373584),
	.w6(32'hbb2ab6e2),
	.w7(32'h3ba01cd9),
	.w8(32'h3b0cfc5c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91dd94),
	.w1(32'h3ba27bea),
	.w2(32'h3b13bdc5),
	.w3(32'h37a9f912),
	.w4(32'h3c5862e5),
	.w5(32'hbc1a778b),
	.w6(32'hbc2d8de9),
	.w7(32'h3b8dc47e),
	.w8(32'hbc0269d5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbf6e3),
	.w1(32'hba65158b),
	.w2(32'hbba30355),
	.w3(32'hbb97d914),
	.w4(32'hbba55600),
	.w5(32'h3b47845f),
	.w6(32'h3b7f2074),
	.w7(32'hbb1aad6a),
	.w8(32'h3c14ee7c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29bb47),
	.w1(32'hbc1d0d6a),
	.w2(32'hbc59cb1c),
	.w3(32'hbb714cfa),
	.w4(32'h3b80022e),
	.w5(32'hbc11884a),
	.w6(32'hbbbd5cef),
	.w7(32'hba723b58),
	.w8(32'hbc578b26),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4853ce),
	.w1(32'hb971c9a1),
	.w2(32'hbb9cc269),
	.w3(32'h3a689cb9),
	.w4(32'h3b3cd4ec),
	.w5(32'hb903c9ae),
	.w6(32'h3a9fea69),
	.w7(32'h3af7c52d),
	.w8(32'hbb626cfc),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cbae9),
	.w1(32'hbb5d065e),
	.w2(32'hbc319c23),
	.w3(32'hbabf585d),
	.w4(32'h3b76ecac),
	.w5(32'hbc25ca23),
	.w6(32'hbbbb23ed),
	.w7(32'h3a6f598b),
	.w8(32'hbc638cdf),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9a00f),
	.w1(32'h3c4dd13b),
	.w2(32'h39ab4798),
	.w3(32'h3c1229c5),
	.w4(32'h3c8f1a63),
	.w5(32'h39f79d93),
	.w6(32'h3bc65bea),
	.w7(32'h3c6f56c5),
	.w8(32'hbb5d27f0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc049d68),
	.w1(32'hbbc606ad),
	.w2(32'hbc3b9bf6),
	.w3(32'hbb9a2e89),
	.w4(32'h38d2543f),
	.w5(32'hbbd57394),
	.w6(32'hbbdff3f0),
	.w7(32'hbb0b7db5),
	.w8(32'hbc1de16d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acccd1c),
	.w1(32'hba805388),
	.w2(32'hbb633fbf),
	.w3(32'h3b1fb110),
	.w4(32'h3a7cd667),
	.w5(32'hbbd3daa6),
	.w6(32'h3bd6f7b5),
	.w7(32'h3b64a293),
	.w8(32'hbc037482),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695f80),
	.w1(32'hbae7efe5),
	.w2(32'h39346973),
	.w3(32'hba8e7524),
	.w4(32'hba377b68),
	.w5(32'hba8f8934),
	.w6(32'h38dfe4a8),
	.w7(32'h39e381a2),
	.w8(32'h3990f239),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5551ae),
	.w1(32'hbbd180fc),
	.w2(32'hbc419da6),
	.w3(32'hbbdb61c3),
	.w4(32'hb9c2ac67),
	.w5(32'hbc1a918f),
	.w6(32'hbb9298c9),
	.w7(32'h3a5b7a1e),
	.w8(32'hbbe2bf79),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb608d7f),
	.w1(32'hbb565a6b),
	.w2(32'hbbe4928a),
	.w3(32'hbb4c56bb),
	.w4(32'hbb92230c),
	.w5(32'hbb951771),
	.w6(32'hbae56ede),
	.w7(32'hbbb50be9),
	.w8(32'hbb48c121),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e3105),
	.w1(32'h3b2fe66c),
	.w2(32'h3b219c03),
	.w3(32'hba789f25),
	.w4(32'h3acbccc7),
	.w5(32'hb9bcfa91),
	.w6(32'h38dfb0b4),
	.w7(32'h3b26b861),
	.w8(32'hba3e81bc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1092b9),
	.w1(32'hbb25e683),
	.w2(32'hbae56eea),
	.w3(32'hbae24d08),
	.w4(32'hb979a602),
	.w5(32'hbb7a2bb2),
	.w6(32'hbb7025d4),
	.w7(32'hbae3953c),
	.w8(32'hbba16f93),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3de6d),
	.w1(32'hbc10fd4f),
	.w2(32'hbc05efcc),
	.w3(32'hbba61d4c),
	.w4(32'hbb9247cd),
	.w5(32'hbba86358),
	.w6(32'hbc142141),
	.w7(32'hbc0647ed),
	.w8(32'hbc1dcb2c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eea80),
	.w1(32'hbb395731),
	.w2(32'hbbc00fdc),
	.w3(32'hbb1e4e5a),
	.w4(32'h3b193093),
	.w5(32'hbb1631da),
	.w6(32'hbb4c9654),
	.w7(32'h3aee5bd8),
	.w8(32'hbaec317c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398019ca),
	.w1(32'hba046394),
	.w2(32'hbb717c58),
	.w3(32'hba158eb0),
	.w4(32'h3b0f8d9f),
	.w5(32'hbb442412),
	.w6(32'hbaf2e333),
	.w7(32'h38d4973b),
	.w8(32'hbbc82ce3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca9ee8),
	.w1(32'hbaa02c99),
	.w2(32'hbb67f032),
	.w3(32'hbb01d28c),
	.w4(32'hb9d6f5e7),
	.w5(32'h39ac08e0),
	.w6(32'hbb292890),
	.w7(32'hbad42e0c),
	.w8(32'hbae6bc40),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09d79f),
	.w1(32'h3a896bd5),
	.w2(32'hbb0d6771),
	.w3(32'hba0e571b),
	.w4(32'h3b2edc37),
	.w5(32'hbae9e70d),
	.w6(32'hbb67ae40),
	.w7(32'hb822925c),
	.w8(32'hbb9cfbef),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb903179),
	.w1(32'hbb4fcb1b),
	.w2(32'hbbb99a8a),
	.w3(32'hbb584684),
	.w4(32'hba2c2249),
	.w5(32'hbb556b46),
	.w6(32'hbb2ee1c7),
	.w7(32'hb947e78a),
	.w8(32'hbb856456),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55ece0),
	.w1(32'hba193bd1),
	.w2(32'hbabfcac2),
	.w3(32'hbb0adb1e),
	.w4(32'h39e22c8d),
	.w5(32'hba41e168),
	.w6(32'hbb820585),
	.w7(32'hba5e3ba5),
	.w8(32'hbb2dc867),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37802f3a),
	.w1(32'h399e065e),
	.w2(32'h3a563e32),
	.w3(32'hb8ae2c78),
	.w4(32'h39eb1ba4),
	.w5(32'h3b4beda3),
	.w6(32'h38c3f652),
	.w7(32'h3a418061),
	.w8(32'h3b4d80b2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c9eac),
	.w1(32'h3b20636b),
	.w2(32'h3ab527fc),
	.w3(32'h3b442c87),
	.w4(32'h3b04c41c),
	.w5(32'h3a9690df),
	.w6(32'h3b40da71),
	.w7(32'h3aebbaad),
	.w8(32'h3a1fa21d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c77b9c),
	.w1(32'hb9c52c8f),
	.w2(32'h3ab10650),
	.w3(32'h39daa527),
	.w4(32'h3ad23e9b),
	.w5(32'hbb2d9f2f),
	.w6(32'h37f5f29c),
	.w7(32'h3b14ad0f),
	.w8(32'hbb2a206d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb090dc6),
	.w1(32'hbb221ecf),
	.w2(32'hb9210df4),
	.w3(32'hbb5bd950),
	.w4(32'hba6fa5f8),
	.w5(32'hbb886a64),
	.w6(32'hbb4a6d15),
	.w7(32'hba2b6d41),
	.w8(32'hbbb94cb6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0037c9),
	.w1(32'hbb8b691a),
	.w2(32'hbbbf6281),
	.w3(32'hbbf0f457),
	.w4(32'h39a4d4a7),
	.w5(32'h3a2c1a95),
	.w6(32'hbc55eaf3),
	.w7(32'hbb96e335),
	.w8(32'hba5d459b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf4e8b),
	.w1(32'hb72a225b),
	.w2(32'hba7ee478),
	.w3(32'h398e49ed),
	.w4(32'h3a1f8a75),
	.w5(32'hba330aab),
	.w6(32'h3980ed98),
	.w7(32'h3a0bbd22),
	.w8(32'hb9bba7ce),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e66fb3),
	.w1(32'hbb001260),
	.w2(32'hbb55ba21),
	.w3(32'h3a96d167),
	.w4(32'hba99522b),
	.w5(32'hbb590f39),
	.w6(32'h3a721d0e),
	.w7(32'hb9221e6e),
	.w8(32'hbb60aa2b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd59244),
	.w1(32'hbb605130),
	.w2(32'hbb948fea),
	.w3(32'hbbb9c151),
	.w4(32'h3a69b2f6),
	.w5(32'hbb392511),
	.w6(32'hbc08a098),
	.w7(32'hbb16a805),
	.w8(32'hbc07e87c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bbd91),
	.w1(32'hb9a00ff6),
	.w2(32'h38dc184d),
	.w3(32'h39c4a46d),
	.w4(32'hb9f5877e),
	.w5(32'h3a344cf2),
	.w6(32'h39f7abb5),
	.w7(32'h3a3c3ffa),
	.w8(32'h38fb26a1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09ab20),
	.w1(32'h371caff6),
	.w2(32'hb7b95b98),
	.w3(32'h399a9f0f),
	.w4(32'h3a98521a),
	.w5(32'hba194aa8),
	.w6(32'h388dcd7c),
	.w7(32'h3987168f),
	.w8(32'hba82ec7d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f001fc),
	.w1(32'hb946049a),
	.w2(32'hb9b10634),
	.w3(32'hba137f73),
	.w4(32'hba46ee6c),
	.w5(32'h3a665a99),
	.w6(32'hba1683bc),
	.w7(32'hb995efb2),
	.w8(32'h3a15532c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0ebd6),
	.w1(32'hba2b1632),
	.w2(32'hbad7a1ca),
	.w3(32'h3a92fff6),
	.w4(32'h39aea1b1),
	.w5(32'h39f51350),
	.w6(32'h3a98b645),
	.w7(32'hb9bf7990),
	.w8(32'hbae85407),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60f539),
	.w1(32'hbb0269d6),
	.w2(32'hba38bd27),
	.w3(32'h3ad469b2),
	.w4(32'hbb25fc80),
	.w5(32'hbba7a1b8),
	.w6(32'hb9956b0b),
	.w7(32'hbaf25d09),
	.w8(32'hbb80f193),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb878546),
	.w1(32'hbb828c98),
	.w2(32'hbbf4aa29),
	.w3(32'hbb4d5522),
	.w4(32'hbaca39a9),
	.w5(32'hbb935006),
	.w6(32'hbb173076),
	.w7(32'hbace3335),
	.w8(32'hbb8df763),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc1c19),
	.w1(32'h39b89ce2),
	.w2(32'h3a87d7eb),
	.w3(32'hb715d94e),
	.w4(32'h398a580a),
	.w5(32'hb9acbeaa),
	.w6(32'h3a626c26),
	.w7(32'h3aa1583d),
	.w8(32'hbaa1365e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eb3ce),
	.w1(32'hbaf23ff2),
	.w2(32'hbb1d64b4),
	.w3(32'hbb65aebf),
	.w4(32'hbb33d099),
	.w5(32'hba90d81e),
	.w6(32'hbbde3809),
	.w7(32'hbb6f1b0e),
	.w8(32'hbb5854f6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3700e18d),
	.w1(32'h38f6dd38),
	.w2(32'hbad0f603),
	.w3(32'hba22d0e4),
	.w4(32'h396141d3),
	.w5(32'hbb849bab),
	.w6(32'hbabb8b19),
	.w7(32'hba015e29),
	.w8(32'hbb6f6350),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88906c),
	.w1(32'hbad2be89),
	.w2(32'hbb3e662d),
	.w3(32'hbb9e67d1),
	.w4(32'hbafcafae),
	.w5(32'h3a1106d8),
	.w6(32'hbb97fff7),
	.w7(32'hbb2fc541),
	.w8(32'hba9f7899),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad95f3f),
	.w1(32'hba9b864a),
	.w2(32'hbb856e8d),
	.w3(32'hbaa9a3d3),
	.w4(32'h3b283309),
	.w5(32'h3b33e7b0),
	.w6(32'hbb3449c0),
	.w7(32'h3a33705c),
	.w8(32'h3aa1b812),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a324ed8),
	.w1(32'hbae54180),
	.w2(32'hbbf8a917),
	.w3(32'hba32a21e),
	.w4(32'hbb16cf71),
	.w5(32'hbbc70797),
	.w6(32'h3a728601),
	.w7(32'hbb0e7e67),
	.w8(32'hbbdfa612),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1182e4),
	.w1(32'hbae56eaa),
	.w2(32'hbb045120),
	.w3(32'hbac82f5b),
	.w4(32'h3aeea522),
	.w5(32'h3ac92a90),
	.w6(32'hbaf00338),
	.w7(32'hb80d62bb),
	.w8(32'hbb214336),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d1340),
	.w1(32'hbaf599ee),
	.w2(32'hbb5842ee),
	.w3(32'h3b3b56f6),
	.w4(32'h3b56c863),
	.w5(32'h3a60d186),
	.w6(32'h3b3f3997),
	.w7(32'h3af3f8bf),
	.w8(32'hbb04057a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fe36a),
	.w1(32'hbb0072cd),
	.w2(32'hbb498c05),
	.w3(32'hbaa649bc),
	.w4(32'h38e17334),
	.w5(32'hbb0771f6),
	.w6(32'hbb008960),
	.w7(32'hba3043f8),
	.w8(32'hbb677b67),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eebb0),
	.w1(32'hba6ed4b0),
	.w2(32'hbae932b5),
	.w3(32'hbae962aa),
	.w4(32'h3b16aef8),
	.w5(32'h3a8e7e31),
	.w6(32'hbb7e1fdd),
	.w7(32'hb966ca4b),
	.w8(32'hbad22158),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8aed1),
	.w1(32'hba8e0e2f),
	.w2(32'hbb91e4cc),
	.w3(32'hbb0d873b),
	.w4(32'hbad9651c),
	.w5(32'hbbb92cbb),
	.w6(32'hbaad61c4),
	.w7(32'hb8e6541f),
	.w8(32'hbbd7ca58),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85438c),
	.w1(32'hbb403347),
	.w2(32'hbba89ad9),
	.w3(32'hbb734a8f),
	.w4(32'hbb4dd09f),
	.w5(32'hbaa28133),
	.w6(32'hbb8babc7),
	.w7(32'hbb6aa31b),
	.w8(32'hbb2691a0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f085f),
	.w1(32'h3b195d27),
	.w2(32'hbb6185c3),
	.w3(32'hbb8ad0da),
	.w4(32'h3b53265f),
	.w5(32'hbaec79b6),
	.w6(32'hbb7f3fc6),
	.w7(32'h3b0a5aad),
	.w8(32'hbbd34fbc),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe369b),
	.w1(32'h3b810b6c),
	.w2(32'h3a170202),
	.w3(32'h3b2ca2f7),
	.w4(32'h3b930c4b),
	.w5(32'h3a94e314),
	.w6(32'h3a9e5a0d),
	.w7(32'h3b25ae14),
	.w8(32'hbabea4d6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c89639),
	.w1(32'hb921f980),
	.w2(32'hb8578779),
	.w3(32'hb9ac4da8),
	.w4(32'h39204e3b),
	.w5(32'h3ac653e9),
	.w6(32'hb90734c8),
	.w7(32'hba25474e),
	.w8(32'h39e33bf0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57dade),
	.w1(32'hba1f1d53),
	.w2(32'hba02cd4d),
	.w3(32'h39e7ca96),
	.w4(32'hb9811cf4),
	.w5(32'hba9ddc92),
	.w6(32'hba4174f4),
	.w7(32'hba0108e0),
	.w8(32'hba3c266d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae47b00),
	.w1(32'hba656563),
	.w2(32'hba959ddf),
	.w3(32'hbb22daa5),
	.w4(32'h378bd3b7),
	.w5(32'hb97762f4),
	.w6(32'hbb27f264),
	.w7(32'hba7b6006),
	.w8(32'hba702ebc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb483bd2),
	.w1(32'hba06a493),
	.w2(32'hbb57b75b),
	.w3(32'h3aacc118),
	.w4(32'h3bd0a66d),
	.w5(32'h3abd859d),
	.w6(32'hb931e920),
	.w7(32'h3b9821e3),
	.w8(32'hbb1f4e2e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f2f53),
	.w1(32'hbb2e1b9f),
	.w2(32'hbb8d48f1),
	.w3(32'hbc1db2cc),
	.w4(32'hb9461879),
	.w5(32'hbb865156),
	.w6(32'hbc35570e),
	.w7(32'hbb819371),
	.w8(32'hbbfc7990),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fd1cf),
	.w1(32'h3a1be0be),
	.w2(32'h381c2538),
	.w3(32'h3a0f2cc4),
	.w4(32'hb97caa1b),
	.w5(32'h3b44b868),
	.w6(32'h3a959a94),
	.w7(32'hb9dbea4f),
	.w8(32'h3b2aa567),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d0fa),
	.w1(32'hba9fd953),
	.w2(32'hbbbec6f9),
	.w3(32'hbb0bbf4e),
	.w4(32'h3a7ddc63),
	.w5(32'hbba66f82),
	.w6(32'hbb542c4d),
	.w7(32'hbaedc8f4),
	.w8(32'hbbc2c3ea),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11c8f5),
	.w1(32'hbaf52e5a),
	.w2(32'hbb79fcd5),
	.w3(32'hb9d80e4e),
	.w4(32'h3a857668),
	.w5(32'hbb16a1b9),
	.w6(32'hbaa33647),
	.w7(32'hba102b86),
	.w8(32'hbb90fd11),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87e379),
	.w1(32'hbc0a9436),
	.w2(32'hbc3c9127),
	.w3(32'hbb949469),
	.w4(32'hbbee7ce2),
	.w5(32'hbbfbb73e),
	.w6(32'hbb16dd3d),
	.w7(32'hbbb144aa),
	.w8(32'hbbcf3143),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af33e64),
	.w1(32'h3b4a0f21),
	.w2(32'hbbd04a6a),
	.w3(32'hba046a88),
	.w4(32'h3b90c5ba),
	.w5(32'hbb517c0a),
	.w6(32'hbb2eea90),
	.w7(32'h3b967674),
	.w8(32'hbb1ba794),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa3dba),
	.w1(32'h3b4670c1),
	.w2(32'h3aac6424),
	.w3(32'h3b883e8a),
	.w4(32'h3bad388b),
	.w5(32'h3b563b3a),
	.w6(32'h3b15ad32),
	.w7(32'h3b188a64),
	.w8(32'h387b3f94),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18d756),
	.w1(32'h3a07a859),
	.w2(32'h3a39a0db),
	.w3(32'h3b062238),
	.w4(32'h3a0fedfe),
	.w5(32'h37f4259b),
	.w6(32'h3ab6d912),
	.w7(32'h3a264fd2),
	.w8(32'hb9c2dc6f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf34b9),
	.w1(32'hbb2bbe81),
	.w2(32'hbb388e75),
	.w3(32'hbb929e96),
	.w4(32'h3a2333be),
	.w5(32'hbb192c0e),
	.w6(32'hbbd3572a),
	.w7(32'hba8f401c),
	.w8(32'hbb8a7d04),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d82c80),
	.w1(32'h3bc96298),
	.w2(32'h3b3bc4f0),
	.w3(32'h3ba1fa1f),
	.w4(32'h3c5aa209),
	.w5(32'h3b397f18),
	.w6(32'h3ba6cb16),
	.w7(32'h3c21e9e2),
	.w8(32'hbb0d8218),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2884a),
	.w1(32'h3b304be6),
	.w2(32'hba7115aa),
	.w3(32'hbac333a7),
	.w4(32'h3b7e674d),
	.w5(32'h3939b698),
	.w6(32'hbb728d8d),
	.w7(32'h3adebac4),
	.w8(32'hba71dcae),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2899ab),
	.w1(32'hbb08cb55),
	.w2(32'hbaec1423),
	.w3(32'hbb4331ac),
	.w4(32'hbb0efbe8),
	.w5(32'hba8fa435),
	.w6(32'hba88529d),
	.w7(32'hba7f3065),
	.w8(32'hba374941),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40a204),
	.w1(32'hb9347402),
	.w2(32'hbad7f215),
	.w3(32'hba4c6cde),
	.w4(32'hba20d0c1),
	.w5(32'h3af40395),
	.w6(32'h37ba5304),
	.w7(32'hb9b5fc6a),
	.w8(32'h3a8a6dff),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacab620),
	.w1(32'hba31faa0),
	.w2(32'hbb6e4446),
	.w3(32'h3b1a06bd),
	.w4(32'h3ac337de),
	.w5(32'hbbd49139),
	.w6(32'h3a90b0dc),
	.w7(32'hba84064d),
	.w8(32'hbbc5b247),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944e205),
	.w1(32'hba0a8762),
	.w2(32'hba265002),
	.w3(32'hba752bd6),
	.w4(32'hb706b89d),
	.w5(32'h3ab0dbd8),
	.w6(32'hba0a9bcb),
	.w7(32'h39dc314d),
	.w8(32'h3a209184),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd09bf),
	.w1(32'hba509e38),
	.w2(32'hbb05c9f9),
	.w3(32'hba26eeff),
	.w4(32'h38ecc042),
	.w5(32'hba882782),
	.w6(32'hba80506e),
	.w7(32'h3a4250e3),
	.w8(32'h39b1e547),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a873d5),
	.w1(32'h3aa12258),
	.w2(32'hb9424487),
	.w3(32'h3ab2d4dd),
	.w4(32'h3a514bd0),
	.w5(32'h3a074755),
	.w6(32'h3a8d3ac6),
	.w7(32'h3a4f3783),
	.w8(32'h3a4eb353),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae5c1),
	.w1(32'hb8a4d44b),
	.w2(32'hbb8cb865),
	.w3(32'hbb89e3da),
	.w4(32'h3a4c5ed2),
	.w5(32'hbb0c0f0d),
	.w6(32'hbc00c53d),
	.w7(32'hb91c9279),
	.w8(32'hbb30b26d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14afe3),
	.w1(32'h3aa64c12),
	.w2(32'h3a018d84),
	.w3(32'h3b2ecaa6),
	.w4(32'h3ad42832),
	.w5(32'hb981a6eb),
	.w6(32'h3ad7b360),
	.w7(32'h3a2ea36a),
	.w8(32'h39cec745),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f73e1),
	.w1(32'hba2208bf),
	.w2(32'hb9e0b867),
	.w3(32'hb793d6a3),
	.w4(32'hb96320c6),
	.w5(32'hb9ebc873),
	.w6(32'h3857dbef),
	.w7(32'h3a3f8505),
	.w8(32'h3a4e4f44),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bbcd1),
	.w1(32'h3ae24fca),
	.w2(32'hba3ec87a),
	.w3(32'h3b9bd038),
	.w4(32'h3bb45465),
	.w5(32'hb81ad9ca),
	.w6(32'h3ba42ae8),
	.w7(32'h3b9634fd),
	.w8(32'hbb00c7fb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5f3c5),
	.w1(32'hba9cef54),
	.w2(32'hbbca6eba),
	.w3(32'hbbb686eb),
	.w4(32'hbb03747d),
	.w5(32'hbc056e6b),
	.w6(32'hbbe26185),
	.w7(32'hba5cb954),
	.w8(32'hbc076b89),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80dfcc),
	.w1(32'h3add3e92),
	.w2(32'hba9405a2),
	.w3(32'hba07c078),
	.w4(32'h3ad85b9d),
	.w5(32'hba161e70),
	.w6(32'hbb352869),
	.w7(32'hb9d286fa),
	.w8(32'hbadb1625),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ca331),
	.w1(32'hbb289b75),
	.w2(32'hbbab32ad),
	.w3(32'hbb834e1b),
	.w4(32'hb9e5a942),
	.w5(32'h3959b5ef),
	.w6(32'hbbd7f32d),
	.w7(32'hbb3041a3),
	.w8(32'hbb5b320b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b495b56),
	.w1(32'h39db6629),
	.w2(32'hb6c9e30c),
	.w3(32'h37d6cd0d),
	.w4(32'h3b091aee),
	.w5(32'hb9ba1db4),
	.w6(32'hba311a74),
	.w7(32'h3ab7d915),
	.w8(32'hbab2ba18),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc497f98),
	.w1(32'hbb9d65f6),
	.w2(32'hbc867875),
	.w3(32'hbbb5665d),
	.w4(32'h3b8a4387),
	.w5(32'hbc2cc52b),
	.w6(32'hbc06fe8a),
	.w7(32'hba8422d7),
	.w8(32'hbc5c1506),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf37f61),
	.w1(32'hbb45394b),
	.w2(32'hbc0cc48c),
	.w3(32'hbbae09a7),
	.w4(32'h3a46c8dc),
	.w5(32'hbb33d092),
	.w6(32'hbbf7b9cb),
	.w7(32'hbadffd81),
	.w8(32'hbbc37893),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd002fb),
	.w1(32'hbb83c057),
	.w2(32'hbbd9aedc),
	.w3(32'hbbb36958),
	.w4(32'hba7176b7),
	.w5(32'hbb43ea3a),
	.w6(32'hbbbd0c1d),
	.w7(32'hbab14c62),
	.w8(32'hbb558f37),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bd7b9),
	.w1(32'h3abd6a1f),
	.w2(32'h3a572527),
	.w3(32'h3b077a37),
	.w4(32'h3aba9032),
	.w5(32'hb8c2fcbd),
	.w6(32'h3b18a9b1),
	.w7(32'h3aa40f6b),
	.w8(32'h398aa10a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb142c75),
	.w1(32'hbad65a5f),
	.w2(32'hbb8207c4),
	.w3(32'hba637f9d),
	.w4(32'hba1c4048),
	.w5(32'h3b291509),
	.w6(32'h3a2280d1),
	.w7(32'h39472e4d),
	.w8(32'h3b2090f7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3259d5),
	.w1(32'h3ada43b1),
	.w2(32'h3a650d7c),
	.w3(32'h3b2a1fa3),
	.w4(32'h3abc4e2b),
	.w5(32'hbac8604e),
	.w6(32'h3b2b6206),
	.w7(32'h3a586873),
	.w8(32'hba386b17),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08f15b),
	.w1(32'hbb0ec870),
	.w2(32'hbb32877f),
	.w3(32'hbb59b001),
	.w4(32'hbaa19584),
	.w5(32'hba1c482f),
	.w6(32'hbb7e85f4),
	.w7(32'hbb1e184f),
	.w8(32'hbae02089),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39165faf),
	.w1(32'h3ab6558f),
	.w2(32'h3a8f87fe),
	.w3(32'hba8d263f),
	.w4(32'h3a945c7f),
	.w5(32'hb909ce23),
	.w6(32'hba279be2),
	.w7(32'h3aee12b0),
	.w8(32'hba9e57f5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4bc62),
	.w1(32'hbb7e85a1),
	.w2(32'hbc088541),
	.w3(32'hbb8d8091),
	.w4(32'hb998d6df),
	.w5(32'hbba54114),
	.w6(32'hbbb7df61),
	.w7(32'hbb583722),
	.w8(32'hbbd7f73c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de0ae0),
	.w1(32'hb972325c),
	.w2(32'hb8f966d2),
	.w3(32'h39aa0ba1),
	.w4(32'h39fe48cc),
	.w5(32'h3a2913c1),
	.w6(32'h39c215e9),
	.w7(32'hb8791ea0),
	.w8(32'h3a2b8b10),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7db9cc7),
	.w1(32'h3a3bd0ff),
	.w2(32'h39b3c184),
	.w3(32'h3885911b),
	.w4(32'h39507a33),
	.w5(32'hba330ab7),
	.w6(32'h3ac71655),
	.w7(32'h39a45ae4),
	.w8(32'hba2cd954),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34b880),
	.w1(32'hb98a24de),
	.w2(32'hb95521fe),
	.w3(32'hbab668b8),
	.w4(32'h3a69b74c),
	.w5(32'h3866e43a),
	.w6(32'hbb323076),
	.w7(32'hba1fd0fc),
	.w8(32'hbab2b6c5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2b539),
	.w1(32'hbb33bef9),
	.w2(32'hbb8968c5),
	.w3(32'hb9ffd02f),
	.w4(32'hbad63b2e),
	.w5(32'hbb395f31),
	.w6(32'hbb0dbe44),
	.w7(32'hbb9e1952),
	.w8(32'hbbcc8503),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f6b84),
	.w1(32'hba9f6859),
	.w2(32'hba845d3b),
	.w3(32'hbb38b5d5),
	.w4(32'hb8c07aec),
	.w5(32'h3b0788b4),
	.w6(32'hba8c2ab9),
	.w7(32'h3b2fd7a3),
	.w8(32'h3abd65d9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13b474),
	.w1(32'h3b1b14fe),
	.w2(32'h39b4fa39),
	.w3(32'h3b1ce13f),
	.w4(32'h3aac08be),
	.w5(32'hbaca2f63),
	.w6(32'h3b2bbe8d),
	.w7(32'h3a6a3e92),
	.w8(32'hbb741709),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac4bcd),
	.w1(32'hbc81adda),
	.w2(32'hbcc5e722),
	.w3(32'hbc98e64f),
	.w4(32'hbc135503),
	.w5(32'hbc679a89),
	.w6(32'hbc59eb65),
	.w7(32'hbc0c5d88),
	.w8(32'hbbe1cc8f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a7571),
	.w1(32'h3b27d62e),
	.w2(32'hbb8e386d),
	.w3(32'hbb51d0af),
	.w4(32'h3c103425),
	.w5(32'h3b1afe09),
	.w6(32'h3b197ce2),
	.w7(32'h3c2709ad),
	.w8(32'h3a086874),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af01617),
	.w1(32'hba0950d4),
	.w2(32'hbaa6a067),
	.w3(32'h3a1f56b0),
	.w4(32'hb9a285a8),
	.w5(32'hbae4f740),
	.w6(32'h3a3b9c8a),
	.w7(32'hb928382c),
	.w8(32'hbada7142),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bf39d),
	.w1(32'hba2c402c),
	.w2(32'hb8c5f684),
	.w3(32'hba3084a7),
	.w4(32'hba44345f),
	.w5(32'h3a0f165b),
	.w6(32'hb8d2d31b),
	.w7(32'hb82b0c9d),
	.w8(32'h3a41cd40),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86e130a),
	.w1(32'h39fa970e),
	.w2(32'h3a3580df),
	.w3(32'h3a60de1e),
	.w4(32'h395c579b),
	.w5(32'h3a08bb4a),
	.w6(32'h3b16d0a8),
	.w7(32'h3a9b972a),
	.w8(32'h38e7e07c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2490a),
	.w1(32'h3a1881a1),
	.w2(32'h390df710),
	.w3(32'h3a2d03a3),
	.w4(32'h3a1e5464),
	.w5(32'h39bee72b),
	.w6(32'h3ab77772),
	.w7(32'h390629a5),
	.w8(32'h3a4ddb2d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b4cd),
	.w1(32'hba1d02be),
	.w2(32'hbaeb15ce),
	.w3(32'h3ab9ba0d),
	.w4(32'hba5b394d),
	.w5(32'hba11b7ab),
	.w6(32'h3b08966d),
	.w7(32'h38251ec9),
	.w8(32'hba2688b8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04980f),
	.w1(32'h3b01cec4),
	.w2(32'hbac89b21),
	.w3(32'h3b003564),
	.w4(32'h3b7cc022),
	.w5(32'h3aa7da30),
	.w6(32'h3903a428),
	.w7(32'h3b2668a6),
	.w8(32'hbb8992c0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05eceb),
	.w1(32'hbb95b238),
	.w2(32'hbc07bc61),
	.w3(32'hbbf3e8ca),
	.w4(32'h39cb6b1b),
	.w5(32'hbb372304),
	.w6(32'hbc2d1bbd),
	.w7(32'hbb483a83),
	.w8(32'hbbbb9bb8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd1a26),
	.w1(32'h3aba264a),
	.w2(32'h39e0778f),
	.w3(32'hb8ddd6fa),
	.w4(32'h3a73b125),
	.w5(32'h3afd6ba4),
	.w6(32'h392f6e23),
	.w7(32'hba194f0f),
	.w8(32'h3a007c5d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fc0b1),
	.w1(32'hbbdd5e68),
	.w2(32'hbc3f2824),
	.w3(32'hb8eb1d19),
	.w4(32'hbb3266db),
	.w5(32'hbc067f25),
	.w6(32'hbbb85901),
	.w7(32'hbbcb2840),
	.w8(32'hbc2db813),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38eff8),
	.w1(32'hbb5dbad6),
	.w2(32'hbb4d9b0b),
	.w3(32'hbb00d1a5),
	.w4(32'hbb3af9cc),
	.w5(32'hbb50d2a4),
	.w6(32'hbb9cc6fc),
	.w7(32'hbb977f37),
	.w8(32'hbb1c8cf1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a1d48),
	.w1(32'hb7c09190),
	.w2(32'hb921d302),
	.w3(32'hba1fdfeb),
	.w4(32'hba805c0d),
	.w5(32'h3a2b1fc2),
	.w6(32'h3a1f8088),
	.w7(32'h38ad965e),
	.w8(32'h3ad590cd),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85b7e1),
	.w1(32'hbac5d4da),
	.w2(32'hba79c989),
	.w3(32'hbaa98184),
	.w4(32'hbaa0b91f),
	.w5(32'hba5da09c),
	.w6(32'hb9a9f4dd),
	.w7(32'h399e5bd8),
	.w8(32'hba3f8eb8),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df236f),
	.w1(32'hba5bb91a),
	.w2(32'hba2269f5),
	.w3(32'hba5f579e),
	.w4(32'hbab4c068),
	.w5(32'h3b19aa63),
	.w6(32'hba7e3221),
	.w7(32'hba0ddc79),
	.w8(32'h3af6422c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34dd35),
	.w1(32'hb9aac07d),
	.w2(32'hba6502f5),
	.w3(32'hbabf1132),
	.w4(32'h3b0ee2de),
	.w5(32'hbb72414a),
	.w6(32'hbb8035a6),
	.w7(32'hbabb3be1),
	.w8(32'hbbcc325d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd59405),
	.w1(32'h3bda6918),
	.w2(32'hbae61dfd),
	.w3(32'hba006733),
	.w4(32'h3c2980a9),
	.w5(32'h3a494343),
	.w6(32'hbb4248d1),
	.w7(32'h3bebac93),
	.w8(32'hbaca3d8f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164807),
	.w1(32'hba38d2d3),
	.w2(32'hbbd3107d),
	.w3(32'hba99b980),
	.w4(32'h3b17e2e2),
	.w5(32'hbb44b7b1),
	.w6(32'hbb569b87),
	.w7(32'hba1161dc),
	.w8(32'hbbd6b3d5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a71cd5),
	.w1(32'h3b0366a0),
	.w2(32'h3b0144b1),
	.w3(32'hb8367435),
	.w4(32'h3b186179),
	.w5(32'hbb6a8f47),
	.w6(32'hbacfba18),
	.w7(32'h3a72e6a3),
	.w8(32'hbb63243d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb39ef),
	.w1(32'hbb7e2178),
	.w2(32'hbc0d6a35),
	.w3(32'hbb91ba40),
	.w4(32'h3aaf4abf),
	.w5(32'hbb254a73),
	.w6(32'hbbcf9189),
	.w7(32'hbb15ef53),
	.w8(32'hbbdbf2a7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c9d90),
	.w1(32'hbb66b451),
	.w2(32'hbb9d5533),
	.w3(32'hbb8c8d4f),
	.w4(32'hba95c94a),
	.w5(32'hbbb0d4d8),
	.w6(32'hbb966d21),
	.w7(32'hbabbc3db),
	.w8(32'hbbc49944),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc917d9d),
	.w1(32'hbc197169),
	.w2(32'hbc35cfa6),
	.w3(32'hbc81d1fb),
	.w4(32'hbbc54e03),
	.w5(32'hbbad9306),
	.w6(32'hbc8f4c08),
	.w7(32'hbc191674),
	.w8(32'hbc0623c6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3011cc),
	.w1(32'hbae1fb59),
	.w2(32'hbac8f16b),
	.w3(32'hbac0463c),
	.w4(32'hbac9ba68),
	.w5(32'hba94c13c),
	.w6(32'hbad1481d),
	.w7(32'hbab5d2e4),
	.w8(32'h39215f95),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b3dd5),
	.w1(32'h3a18e05a),
	.w2(32'h3975cc2c),
	.w3(32'hb97f7ea3),
	.w4(32'hba0557d6),
	.w5(32'h3a954282),
	.w6(32'h3a38b401),
	.w7(32'hb9a2076a),
	.w8(32'h3a2d15e7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5086e),
	.w1(32'h3a4a3c33),
	.w2(32'hbbc838f0),
	.w3(32'hbaa5eda9),
	.w4(32'h3aa3b903),
	.w5(32'hbbd15c84),
	.w6(32'hbba02f43),
	.w7(32'hbb07f3e5),
	.w8(32'hbc0591b4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafa3d4),
	.w1(32'h390279bd),
	.w2(32'hbbcc3a8e),
	.w3(32'hbb43d3e4),
	.w4(32'h39c37ef0),
	.w5(32'hbbcd74d7),
	.w6(32'hbbd2be0d),
	.w7(32'hbae6c56c),
	.w8(32'hbbb0bc0f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd3a3d),
	.w1(32'hbba13ddc),
	.w2(32'hbc1a1994),
	.w3(32'hbb7d6285),
	.w4(32'h3ac762f0),
	.w5(32'hbb8608f8),
	.w6(32'hbbde892d),
	.w7(32'hbad85db0),
	.w8(32'hbbfe7b79),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d03e4),
	.w1(32'hbb040054),
	.w2(32'hb9f08ef4),
	.w3(32'hbb79442f),
	.w4(32'hbb803b46),
	.w5(32'hbb35b7a9),
	.w6(32'hb6823fdd),
	.w7(32'hb9ba76fb),
	.w8(32'hbb329308),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93deaba),
	.w1(32'hba07c3db),
	.w2(32'hba027fb7),
	.w3(32'hbaca8494),
	.w4(32'hbabb4e37),
	.w5(32'h3afe9647),
	.w6(32'hba8e7c87),
	.w7(32'hba605f8d),
	.w8(32'h3ae1dd47),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a407494),
	.w1(32'hb84fd672),
	.w2(32'h390285c2),
	.w3(32'h3903effd),
	.w4(32'h39862cad),
	.w5(32'h3a11f52c),
	.w6(32'hb890e8e2),
	.w7(32'hba128908),
	.w8(32'hb9384624),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1b5e8),
	.w1(32'hb902eac4),
	.w2(32'hbb939714),
	.w3(32'hba151ded),
	.w4(32'hbb8f844a),
	.w5(32'hbc02ebbe),
	.w6(32'h39299a20),
	.w7(32'h38852f54),
	.w8(32'hbba42722),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73b25d),
	.w1(32'hbba52fc8),
	.w2(32'hbc21504f),
	.w3(32'hbc19b1c8),
	.w4(32'hbb892c0e),
	.w5(32'hbc01cf04),
	.w6(32'hbc242103),
	.w7(32'hbba269d3),
	.w8(32'hbc0cd6ed),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b32c3c),
	.w1(32'hbb3aff6c),
	.w2(32'hbb80a930),
	.w3(32'h3abbc299),
	.w4(32'hb67001b6),
	.w5(32'hbbf1f06b),
	.w6(32'h3aecce0e),
	.w7(32'h39e7c53a),
	.w8(32'hbc05e59d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee999e),
	.w1(32'h3b30d533),
	.w2(32'hbad11eaa),
	.w3(32'hba778952),
	.w4(32'h3b680b3e),
	.w5(32'h3a3c36be),
	.w6(32'hbb8ae8a8),
	.w7(32'h3a4e4ef2),
	.w8(32'hbafa0c0f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af6e8),
	.w1(32'hbb893330),
	.w2(32'hbbc9ea42),
	.w3(32'hbc088d5e),
	.w4(32'h3ac47824),
	.w5(32'hbb2d253c),
	.w6(32'hbc09650f),
	.w7(32'hba0b0d2c),
	.w8(32'hbbc5872b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46bb0d),
	.w1(32'hb8e7a8ed),
	.w2(32'hb904d119),
	.w3(32'h399453d9),
	.w4(32'hb829ca12),
	.w5(32'h38a76c35),
	.w6(32'h37be06f6),
	.w7(32'hba24ccc4),
	.w8(32'h3998d627),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af856f3),
	.w1(32'h3b11294d),
	.w2(32'h3a8d1d13),
	.w3(32'hbb06e7f1),
	.w4(32'hbab5746c),
	.w5(32'hbb58b97e),
	.w6(32'hba9ea316),
	.w7(32'hba86bea9),
	.w8(32'hbb2c77a7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf986d3),
	.w1(32'hba6ca3c0),
	.w2(32'h38e9967e),
	.w3(32'hbaf79d3f),
	.w4(32'hbaab27b4),
	.w5(32'hba68f58a),
	.w6(32'hbab221d9),
	.w7(32'hba6c0c18),
	.w8(32'hba68642d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cb7cf),
	.w1(32'h3960e51d),
	.w2(32'hb9a79a69),
	.w3(32'h3a5ee272),
	.w4(32'h384cdaea),
	.w5(32'h3b727d36),
	.w6(32'h3a86a436),
	.w7(32'hbab932e2),
	.w8(32'h3ba29f28),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59198),
	.w1(32'hbad6bf51),
	.w2(32'h39a759f4),
	.w3(32'hb9bce42f),
	.w4(32'h39fcfcb4),
	.w5(32'hbae9119e),
	.w6(32'h3924966b),
	.w7(32'h3a5aef5f),
	.w8(32'hbb8a791b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13f8dc),
	.w1(32'hbc254fc1),
	.w2(32'hbba87e47),
	.w3(32'hbbc1374c),
	.w4(32'hba8fcd27),
	.w5(32'hbc003018),
	.w6(32'hbbf25d50),
	.w7(32'hbb011b35),
	.w8(32'hbc1ece7f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae8ba5),
	.w1(32'h3b1bc9a0),
	.w2(32'hbb3a6986),
	.w3(32'h398cf053),
	.w4(32'hbaf3e7e7),
	.w5(32'h3b24d4a0),
	.w6(32'hbb6bc2ea),
	.w7(32'hbb3965cd),
	.w8(32'hbbcc7849),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01d6a9),
	.w1(32'hbb50d8f2),
	.w2(32'h3addd1e8),
	.w3(32'hbb42d701),
	.w4(32'hbb22320a),
	.w5(32'h3bd3e69d),
	.w6(32'hba288b0d),
	.w7(32'h39d1906b),
	.w8(32'h3b895d3f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf79d6),
	.w1(32'hbbf4c4b0),
	.w2(32'hbc1104e4),
	.w3(32'hbba0a9f3),
	.w4(32'hbbd07d64),
	.w5(32'hbc28c301),
	.w6(32'hbb299ab1),
	.w7(32'hbb9533e4),
	.w8(32'hbc6e0a76),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe82a48),
	.w1(32'hbb2bc728),
	.w2(32'hbaca898f),
	.w3(32'hbb514dae),
	.w4(32'hbabd8feb),
	.w5(32'hb737b3c3),
	.w6(32'hbb6dcdb1),
	.w7(32'hbb02dbce),
	.w8(32'hbbc3c523),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d2efb3),
	.w1(32'hbb230cb7),
	.w2(32'hbbc219a7),
	.w3(32'hba5d4459),
	.w4(32'hbb862722),
	.w5(32'h39de882f),
	.w6(32'hbbb60106),
	.w7(32'hbba0c8d6),
	.w8(32'hbaef628d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe12c55),
	.w1(32'hbbde632b),
	.w2(32'hbbd501c8),
	.w3(32'hbaa967f3),
	.w4(32'hbb839ea0),
	.w5(32'hbaffe4a0),
	.w6(32'hbb1f0ce7),
	.w7(32'hbba9999c),
	.w8(32'hbb3d90df),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38a8f2),
	.w1(32'hbb83f62d),
	.w2(32'hbbb2b483),
	.w3(32'hba09da63),
	.w4(32'hbb15fe1d),
	.w5(32'h3a0393dd),
	.w6(32'h3babaa44),
	.w7(32'hbb37886e),
	.w8(32'h3b0db67e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87bdf1),
	.w1(32'h3b94dab1),
	.w2(32'h3ba4ec7a),
	.w3(32'h3bb46cd6),
	.w4(32'h3ac64b5e),
	.w5(32'h3b687453),
	.w6(32'h3bd281d0),
	.w7(32'h3b614ae2),
	.w8(32'h3bb6964e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a1c82),
	.w1(32'h3a661adc),
	.w2(32'h3b845e46),
	.w3(32'h3ad4ec65),
	.w4(32'h3b91a609),
	.w5(32'hbb2c9b72),
	.w6(32'h3a885b59),
	.w7(32'h3b12fc7e),
	.w8(32'h3b9b60d2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd016e2),
	.w1(32'h3ba45ddb),
	.w2(32'h3a6ee2c3),
	.w3(32'h3bcc7747),
	.w4(32'h3ae52040),
	.w5(32'hbc0f6d85),
	.w6(32'h3c5068ab),
	.w7(32'h3a8d92d1),
	.w8(32'hbbbe3e43),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eb747),
	.w1(32'hbbad3f93),
	.w2(32'hbbcd6c7a),
	.w3(32'hbba68b23),
	.w4(32'hbaadf8ee),
	.w5(32'h3b388a50),
	.w6(32'h3a5c2bb8),
	.w7(32'hbbc17b34),
	.w8(32'hbb2bc282),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51edce),
	.w1(32'hbc23c0b9),
	.w2(32'hbc1668da),
	.w3(32'hbb84859f),
	.w4(32'hbbb6a350),
	.w5(32'hbbc6971a),
	.w6(32'hbbd0948b),
	.w7(32'hbc166fbf),
	.w8(32'hbba406bb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b8e68),
	.w1(32'h3b2b59ef),
	.w2(32'hbbb69282),
	.w3(32'hbb3a11cf),
	.w4(32'h3a77b4f3),
	.w5(32'h3adbcc5b),
	.w6(32'h3be92aa0),
	.w7(32'hba8a4bfc),
	.w8(32'h3b6b7c6b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7bcf5),
	.w1(32'hbba0c474),
	.w2(32'hbbb969f5),
	.w3(32'hbbb157e5),
	.w4(32'hbbbe85a1),
	.w5(32'hbb83e13c),
	.w6(32'hbc0a9155),
	.w7(32'hbb9e6c3a),
	.w8(32'hbbafb40c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b013397),
	.w1(32'h39fccae6),
	.w2(32'hbb130180),
	.w3(32'h3a12138f),
	.w4(32'h3b38d70a),
	.w5(32'h3b5a7def),
	.w6(32'hbb2c012c),
	.w7(32'hbaa8aac4),
	.w8(32'hbb887521),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae232fa),
	.w1(32'hb9fcbf7b),
	.w2(32'h39c481d3),
	.w3(32'h3b063930),
	.w4(32'hbaa0bb38),
	.w5(32'h3c16765e),
	.w6(32'h3bb9b73d),
	.w7(32'hbb6c59da),
	.w8(32'h3c001a79),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c267db0),
	.w1(32'h3a62e652),
	.w2(32'h3b83daf8),
	.w3(32'hbb0f8c77),
	.w4(32'hbb9a6de9),
	.w5(32'hbb0ac853),
	.w6(32'hbbb3d54a),
	.w7(32'hba719d0c),
	.w8(32'hbb7870a2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba89b1f),
	.w1(32'hbb50c7df),
	.w2(32'h3b499f6c),
	.w3(32'hbb98d450),
	.w4(32'h3abd6d29),
	.w5(32'h3c159011),
	.w6(32'hbaa3857d),
	.w7(32'h3ae12f4a),
	.w8(32'h3b9ffe6b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aa66e),
	.w1(32'hbc23d707),
	.w2(32'hbc59d607),
	.w3(32'hbb0ee6c6),
	.w4(32'h3a5faab4),
	.w5(32'hbad6edae),
	.w6(32'hbb6b53b5),
	.w7(32'hbadfbee3),
	.w8(32'hbb3e0d80),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e5dbe),
	.w1(32'hba7acc06),
	.w2(32'hba32a61b),
	.w3(32'hbb8aa326),
	.w4(32'hbb165cc2),
	.w5(32'h3b07deaf),
	.w6(32'hba8a481b),
	.w7(32'h3a987ca3),
	.w8(32'hbac9ed3f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba438a7),
	.w1(32'h3b54a681),
	.w2(32'hb93e99f2),
	.w3(32'h3a5f7a01),
	.w4(32'h3a94bb60),
	.w5(32'hbc893f03),
	.w6(32'h3a77c831),
	.w7(32'hbb02d8f7),
	.w8(32'hbc8031c4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c51e2),
	.w1(32'h3be40293),
	.w2(32'hbbc32e3c),
	.w3(32'hbbf4efa7),
	.w4(32'h3aaf61b8),
	.w5(32'hbbe85d84),
	.w6(32'h3c25629e),
	.w7(32'h3afede7a),
	.w8(32'h3b620681),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80978b),
	.w1(32'hbafc578a),
	.w2(32'hbc06a444),
	.w3(32'h399c1ed6),
	.w4(32'h3c0f79d5),
	.w5(32'hbc02f22b),
	.w6(32'h3c5c4afc),
	.w7(32'hbb56f0d0),
	.w8(32'hbc72d1eb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc16bb6),
	.w1(32'h3ba75c03),
	.w2(32'hbbd1c74f),
	.w3(32'h3b2105b1),
	.w4(32'hbbcd3f81),
	.w5(32'hbbc15c6d),
	.w6(32'h3bd7dd6d),
	.w7(32'hbb8e8fac),
	.w8(32'hbb36f4cd),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf6cf2),
	.w1(32'hbbd67a84),
	.w2(32'hbbc658f6),
	.w3(32'hbb470eb9),
	.w4(32'h3b0db397),
	.w5(32'h3ad24a5d),
	.w6(32'h3b004b2c),
	.w7(32'hbb1318e4),
	.w8(32'hb9f8c332),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850571),
	.w1(32'hbbe5431c),
	.w2(32'hbbda9cdc),
	.w3(32'h3ade2f8d),
	.w4(32'hba6545b4),
	.w5(32'hbb219881),
	.w6(32'hbb40e3fb),
	.w7(32'hba30bb91),
	.w8(32'hbae1d37e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad337c3),
	.w1(32'h389d8e20),
	.w2(32'h3b085903),
	.w3(32'hb9664102),
	.w4(32'hb9b1d401),
	.w5(32'hb4e7103d),
	.w6(32'hbacce8ee),
	.w7(32'hba1206ec),
	.w8(32'hbada855d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb14a7),
	.w1(32'h3bd330c6),
	.w2(32'h3bbe76ae),
	.w3(32'h3bad5b45),
	.w4(32'h3b9bfc89),
	.w5(32'h3b7eb81a),
	.w6(32'hbbb417bb),
	.w7(32'h3aa25f86),
	.w8(32'h39d84bbc),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule