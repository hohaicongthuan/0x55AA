module layer_8_featuremap_23(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b8901),
	.w1(32'h39fdab84),
	.w2(32'h3aadf40b),
	.w3(32'hb8ede1f8),
	.w4(32'h3a5164c2),
	.w5(32'h3ad84a99),
	.w6(32'h3b5c839c),
	.w7(32'h3b385863),
	.w8(32'h3b4e0c2b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01a69c),
	.w1(32'hb9669e86),
	.w2(32'hbaa111c3),
	.w3(32'hbab3b3a9),
	.w4(32'hb9ab481b),
	.w5(32'hbab35353),
	.w6(32'h39bc7e3e),
	.w7(32'hba16371d),
	.w8(32'hba8b7c09),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91ecfb),
	.w1(32'hba7209d6),
	.w2(32'h3a1409fa),
	.w3(32'hbb59740c),
	.w4(32'hbac3e2e3),
	.w5(32'hbac471b9),
	.w6(32'hbbb7509b),
	.w7(32'hbb9a8632),
	.w8(32'hbb69b25e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f9c7f),
	.w1(32'h3ab4c842),
	.w2(32'h3b32178c),
	.w3(32'h39baa245),
	.w4(32'h3a436243),
	.w5(32'h3ae4e166),
	.w6(32'hba2ac24c),
	.w7(32'h38ce3ecc),
	.w8(32'h3860aa25),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff1dea),
	.w1(32'hbbb4e61c),
	.w2(32'hba98650f),
	.w3(32'hbb26498c),
	.w4(32'hbb8262bf),
	.w5(32'hbac11d23),
	.w6(32'h3aecc922),
	.w7(32'h3938a61a),
	.w8(32'h3bd8aa30),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b2079),
	.w1(32'h3bc5ccf0),
	.w2(32'h3bdf36b5),
	.w3(32'h3b153c1c),
	.w4(32'h3b492fe6),
	.w5(32'h3b97002a),
	.w6(32'h3a8da498),
	.w7(32'h3b64f0cd),
	.w8(32'hbaf9e436),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15f9a9),
	.w1(32'h39faf071),
	.w2(32'h38ef6b4e),
	.w3(32'hba8d40df),
	.w4(32'hb9a36347),
	.w5(32'hb88299ff),
	.w6(32'h398002a2),
	.w7(32'hb963961d),
	.w8(32'hba35b3b2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabca976),
	.w1(32'hbaab0080),
	.w2(32'h38bf641f),
	.w3(32'hbb9d80c3),
	.w4(32'hbbb3fdd2),
	.w5(32'hbb428307),
	.w6(32'hba8ac11a),
	.w7(32'hba9336ce),
	.w8(32'h399efdd7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e79d2),
	.w1(32'hbafb5c3b),
	.w2(32'h3a02e9ab),
	.w3(32'hbb39bdb8),
	.w4(32'hbb2c9e20),
	.w5(32'h3af8b695),
	.w6(32'hbabaac12),
	.w7(32'hbaea16a0),
	.w8(32'h3b01b852),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c02272),
	.w1(32'h3b0732da),
	.w2(32'h3afb37a5),
	.w3(32'h39f0d750),
	.w4(32'h3b041f4e),
	.w5(32'h3b172b0b),
	.w6(32'hb67263e8),
	.w7(32'hb9976281),
	.w8(32'h3b0beba1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f5c7d),
	.w1(32'hbbd7fd53),
	.w2(32'hbbc064a9),
	.w3(32'hbb71a943),
	.w4(32'hbbc859f4),
	.w5(32'hbb6daf65),
	.w6(32'h3a3df457),
	.w7(32'hba3c336d),
	.w8(32'hbabb5074),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba629eb9),
	.w1(32'h37f1572e),
	.w2(32'hba093dbb),
	.w3(32'hbaeaecfa),
	.w4(32'hba08858a),
	.w5(32'h39dce445),
	.w6(32'h3968fab8),
	.w7(32'h3a071f9a),
	.w8(32'h3aac7056),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fb091),
	.w1(32'h3a73ee11),
	.w2(32'h3a7b9cdd),
	.w3(32'hba8a58da),
	.w4(32'h39d4ec51),
	.w5(32'h3a98c317),
	.w6(32'hbb02f1f8),
	.w7(32'hbb0bbd18),
	.w8(32'h3ba16067),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4ef42),
	.w1(32'h3b73958b),
	.w2(32'h3ba36378),
	.w3(32'h3b853374),
	.w4(32'h3b3f0b93),
	.w5(32'h3b901dc3),
	.w6(32'h3ba33bd5),
	.w7(32'h3bb60ec5),
	.w8(32'h3b3bb445),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ae377),
	.w1(32'h3b12f2cd),
	.w2(32'h3b1dfbf4),
	.w3(32'h3b092e1c),
	.w4(32'h3afa11fb),
	.w5(32'h3b119be4),
	.w6(32'h3b31588e),
	.w7(32'h3b4a029c),
	.w8(32'hb91e9291),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa59222),
	.w1(32'hb9c95b98),
	.w2(32'hba51c8a5),
	.w3(32'hbac141e0),
	.w4(32'hba4a5f69),
	.w5(32'hba224f02),
	.w6(32'hb9da5432),
	.w7(32'hba5c0464),
	.w8(32'hb8fd6e92),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b2a85),
	.w1(32'h3a153948),
	.w2(32'hb9eabab2),
	.w3(32'hba84236f),
	.w4(32'hba80ab49),
	.w5(32'hba21de9f),
	.w6(32'h3a14d59e),
	.w7(32'hba165fd6),
	.w8(32'hbabb45b9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85aaac),
	.w1(32'hbb692a87),
	.w2(32'hbab6d596),
	.w3(32'hbb8a25a1),
	.w4(32'hbba347b2),
	.w5(32'hbb44831b),
	.w6(32'hbb88e0f4),
	.w7(32'hbba51985),
	.w8(32'hbb43cb90),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc975924),
	.w1(32'hbcbd970c),
	.w2(32'hbc4e828e),
	.w3(32'hbc63827b),
	.w4(32'hbc5865a5),
	.w5(32'hbc0b69ae),
	.w6(32'h38d83786),
	.w7(32'hbb04c014),
	.w8(32'hbb52d948),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6a75e),
	.w1(32'hbc3f0689),
	.w2(32'hbbf03fc1),
	.w3(32'hbbf4f8a8),
	.w4(32'hbc3d8242),
	.w5(32'hbc137b19),
	.w6(32'h391afe11),
	.w7(32'hbb318700),
	.w8(32'hbb839b44),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb691b7b),
	.w1(32'hbb2c825f),
	.w2(32'hbb9dcc9a),
	.w3(32'hbb41893a),
	.w4(32'hbb545c83),
	.w5(32'hbb548101),
	.w6(32'hbad731f3),
	.w7(32'hbb643917),
	.w8(32'h3a624250),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6a41c),
	.w1(32'h3b5fa4b8),
	.w2(32'h3b376370),
	.w3(32'hb9c6fbe4),
	.w4(32'h3b45707e),
	.w5(32'h3b3fde81),
	.w6(32'hbb211f28),
	.w7(32'hb9833800),
	.w8(32'hbb9bec40),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55ea96),
	.w1(32'hbc7b4c15),
	.w2(32'hbc166a4f),
	.w3(32'hbbd01646),
	.w4(32'hbc7ac879),
	.w5(32'hbc06d02a),
	.w6(32'h3b78ac1e),
	.w7(32'hb9dce932),
	.w8(32'h3bdeb846),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394534ff),
	.w1(32'hbb452a8b),
	.w2(32'hbb57a171),
	.w3(32'hbb52aa6a),
	.w4(32'hbbbbc84c),
	.w5(32'hbba2e9bb),
	.w6(32'hb89ce209),
	.w7(32'hbb471cc9),
	.w8(32'hbb843883),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50792d),
	.w1(32'hbb59acc9),
	.w2(32'hbb559246),
	.w3(32'hbafdec92),
	.w4(32'hbb587f13),
	.w5(32'hbb82cb00),
	.w6(32'hbb7aaaac),
	.w7(32'hbb3bd7d9),
	.w8(32'hbb27cbad),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31672a),
	.w1(32'hbc309662),
	.w2(32'hbc0089cd),
	.w3(32'hbab36162),
	.w4(32'hbbd87c1e),
	.w5(32'hbbb77225),
	.w6(32'h3bd108ba),
	.w7(32'hb922510e),
	.w8(32'h3ab41795),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dadbc5),
	.w1(32'hba76e213),
	.w2(32'hba63a2e0),
	.w3(32'hb9a6a680),
	.w4(32'hba864b98),
	.w5(32'hba5144f7),
	.w6(32'hba77af4b),
	.w7(32'hba514c8c),
	.w8(32'h399ec246),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce308a1),
	.w1(32'hbd1acbdf),
	.w2(32'hbd480064),
	.w3(32'hbd4274e6),
	.w4(32'hbd419ba7),
	.w5(32'hbcdd2903),
	.w6(32'hbc57c9a8),
	.w7(32'h3d14ff0e),
	.w8(32'h3cd9b4ba),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3a60f),
	.w1(32'hbb68e8df),
	.w2(32'hbb15f85c),
	.w3(32'hbb91a35f),
	.w4(32'hbadd6d78),
	.w5(32'h392ad192),
	.w6(32'h3aba481f),
	.w7(32'h3a95408c),
	.w8(32'h3aa9013d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8042d6),
	.w1(32'hb9885419),
	.w2(32'hb8f8654e),
	.w3(32'hba8a126f),
	.w4(32'hb9af5a92),
	.w5(32'hb9bcda51),
	.w6(32'hbaa5cd9e),
	.w7(32'hba653085),
	.w8(32'hbb519ca9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05cf0f),
	.w1(32'h3b837988),
	.w2(32'h3b6f18c5),
	.w3(32'h3b7d87ce),
	.w4(32'h3bb8d20a),
	.w5(32'h3b53e6d8),
	.w6(32'h39e75d5b),
	.w7(32'h3b3c19c5),
	.w8(32'hbaa9a073),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80e842),
	.w1(32'hbbb4e113),
	.w2(32'hbb983fb8),
	.w3(32'hbb52fd4d),
	.w4(32'hbb8330f3),
	.w5(32'hbb7d3182),
	.w6(32'hbb18001e),
	.w7(32'hbb559209),
	.w8(32'hb9bd0a5f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09a142),
	.w1(32'h385de22f),
	.w2(32'hba11fd1d),
	.w3(32'hba3ef7e3),
	.w4(32'hba837205),
	.w5(32'hba29d7f5),
	.w6(32'hba42c0a0),
	.w7(32'hb9e6e867),
	.w8(32'hba8a3d15),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9c00b),
	.w1(32'hb89550f4),
	.w2(32'h3987872d),
	.w3(32'hba15992f),
	.w4(32'h3a4c6720),
	.w5(32'h372c7309),
	.w6(32'hba3f9721),
	.w7(32'h3a5eb3cc),
	.w8(32'h3bb93132),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc048e0),
	.w1(32'h3b73bce9),
	.w2(32'h3b531e49),
	.w3(32'h3b8c3c80),
	.w4(32'h3ae859dc),
	.w5(32'h3a25e7e2),
	.w6(32'h3b82b8ad),
	.w7(32'h3b4449d7),
	.w8(32'hbbab4b4d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba359c97),
	.w1(32'hbba9b08b),
	.w2(32'hbbc18eff),
	.w3(32'hb920e516),
	.w4(32'hbb669254),
	.w5(32'hbb63a917),
	.w6(32'h3baa1f37),
	.w7(32'h3a4e9825),
	.w8(32'hbb85e8b8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a868e),
	.w1(32'hbb5573c9),
	.w2(32'hbb29bb86),
	.w3(32'hbb879ed4),
	.w4(32'hbb875f5c),
	.w5(32'hbb5a0e00),
	.w6(32'hbb6c8348),
	.w7(32'hbb410ccd),
	.w8(32'hb9d0d40c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bd012),
	.w1(32'hb9bc9554),
	.w2(32'hb9e26043),
	.w3(32'h39c479c6),
	.w4(32'h3b1d2713),
	.w5(32'h3b3a72c2),
	.w6(32'h3af4a6d0),
	.w7(32'h3b5abce8),
	.w8(32'h3c11c3af),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96421f),
	.w1(32'h3b861d75),
	.w2(32'h3b94eaf7),
	.w3(32'h3b663b13),
	.w4(32'h3b41f099),
	.w5(32'h3b6d9b93),
	.w6(32'h3b9aa156),
	.w7(32'h3ba5706b),
	.w8(32'hbaecb93e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f60fe1),
	.w1(32'hba00afeb),
	.w2(32'hbaaa4883),
	.w3(32'hbb0f66a2),
	.w4(32'hbb20a46f),
	.w5(32'hbb34cd3c),
	.w6(32'hbb0feb58),
	.w7(32'hbb3861d0),
	.w8(32'hba1a74c8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabca6d1),
	.w1(32'hbb951797),
	.w2(32'hbbbcb54f),
	.w3(32'h3aa10d22),
	.w4(32'hbae6457d),
	.w5(32'hbb7665a3),
	.w6(32'h3ab36399),
	.w7(32'hbb07a109),
	.w8(32'hbb8765f2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3305bb),
	.w1(32'hbb1e40ce),
	.w2(32'h3998e61f),
	.w3(32'hbb35dc00),
	.w4(32'hbb4b6f8c),
	.w5(32'hbac59793),
	.w6(32'hbb2e3185),
	.w7(32'hba6b731c),
	.w8(32'hbc0f5942),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18f64b),
	.w1(32'hbb55c617),
	.w2(32'h3b45dc0c),
	.w3(32'hbbdeedb2),
	.w4(32'hb90c8cbf),
	.w5(32'hbb12a6af),
	.w6(32'h3b3bcf05),
	.w7(32'hb9b9fa42),
	.w8(32'hb9ba21b6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9818cfd),
	.w1(32'hbb124160),
	.w2(32'hba8bf41f),
	.w3(32'hbad84a0f),
	.w4(32'hbaaceb34),
	.w5(32'hbac7a59f),
	.w6(32'h3abd4330),
	.w7(32'h3ac0ab52),
	.w8(32'h3a501fe7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b0939),
	.w1(32'hbb9a5be0),
	.w2(32'h399ed409),
	.w3(32'hbba36c5b),
	.w4(32'hbb4f9f34),
	.w5(32'hb9b7d197),
	.w6(32'h3b2bcad0),
	.w7(32'h3bc5c6f0),
	.w8(32'h3ba4c033),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933678a),
	.w1(32'hba961f8f),
	.w2(32'hba44657c),
	.w3(32'h3a2aaaa1),
	.w4(32'hb98e7355),
	.w5(32'hb664ac14),
	.w6(32'hb8e40b04),
	.w7(32'h3b478746),
	.w8(32'hbc1ffb05),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a1185),
	.w1(32'h39dcd91b),
	.w2(32'hbc018d96),
	.w3(32'hbb219a82),
	.w4(32'h3b7b742c),
	.w5(32'h3a877235),
	.w6(32'hbb9cbc63),
	.w7(32'h3aa76ac0),
	.w8(32'hba97cd52),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8bd76),
	.w1(32'hbc30c131),
	.w2(32'hbb4bb94a),
	.w3(32'hbc02c802),
	.w4(32'hbc0da08e),
	.w5(32'hbae2c90d),
	.w6(32'hbb68b335),
	.w7(32'hbb6a4f0e),
	.w8(32'h3a736e64),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f591e),
	.w1(32'hb982f12a),
	.w2(32'h3af13476),
	.w3(32'hba8460ec),
	.w4(32'hba32296e),
	.w5(32'h3ac9b1c2),
	.w6(32'hbaaa9887),
	.w7(32'hb9b5a027),
	.w8(32'hb9ef874b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb314f26),
	.w1(32'hbb2dfe46),
	.w2(32'h3a177a7e),
	.w3(32'hbaca17b6),
	.w4(32'h39b38e25),
	.w5(32'h3b645cf8),
	.w6(32'hb9214eff),
	.w7(32'h3b78e8e0),
	.w8(32'h3b2aa6eb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79c6ef),
	.w1(32'h36b07a71),
	.w2(32'h3a35c431),
	.w3(32'hbb3fc47c),
	.w4(32'h3aa0d609),
	.w5(32'h3ae8ba59),
	.w6(32'hbb367488),
	.w7(32'h3ad7d217),
	.w8(32'h3b063882),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34bdd0),
	.w1(32'hbc78888b),
	.w2(32'hbc0a2f32),
	.w3(32'hbc9fe3a7),
	.w4(32'hbcb4eb49),
	.w5(32'hbc8e9cc0),
	.w6(32'hbbdf8a81),
	.w7(32'hbbb1377a),
	.w8(32'hbbe181d2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e340c1),
	.w1(32'hbbd3f623),
	.w2(32'hbc3c4726),
	.w3(32'hbc370a0d),
	.w4(32'hbc38f3fd),
	.w5(32'hbc1dfc9b),
	.w6(32'hba9a341d),
	.w7(32'hbbba4a81),
	.w8(32'h3b569f21),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3a911),
	.w1(32'hbb687df8),
	.w2(32'hbac5f864),
	.w3(32'hbae01c99),
	.w4(32'hbb65b134),
	.w5(32'hb9d6a759),
	.w6(32'hba9988d8),
	.w7(32'hbab4680b),
	.w8(32'hb8fa43dc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04a348),
	.w1(32'hbb1cc9d3),
	.w2(32'hbc1bd8e5),
	.w3(32'hba268b93),
	.w4(32'h3b4cbf59),
	.w5(32'hbb88f6ea),
	.w6(32'h3b2b5930),
	.w7(32'hbbe67116),
	.w8(32'hbb976281),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc212232),
	.w1(32'hbc32eb6a),
	.w2(32'hbc5377c0),
	.w3(32'hbc4c8996),
	.w4(32'hbc20eb4a),
	.w5(32'hbbda7c12),
	.w6(32'hbb6d9df7),
	.w7(32'h3b5e057b),
	.w8(32'h3bed365c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c2540),
	.w1(32'h3b6ab0d6),
	.w2(32'h3a4c6d66),
	.w3(32'hbafd9e12),
	.w4(32'hbab057dd),
	.w5(32'h3ab566b4),
	.w6(32'h3b3d327d),
	.w7(32'h3b57b95a),
	.w8(32'h3b89151c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab93286),
	.w1(32'hbb396f98),
	.w2(32'hbaa25fdd),
	.w3(32'h3b131694),
	.w4(32'hbaa6cafc),
	.w5(32'hbb919c30),
	.w6(32'h3b555664),
	.w7(32'hbb307e61),
	.w8(32'h3adcae49),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31ecae),
	.w1(32'hbb6e3457),
	.w2(32'h39595fef),
	.w3(32'hbbb983fa),
	.w4(32'hbb8a9564),
	.w5(32'hb9b19549),
	.w6(32'hbaa16313),
	.w7(32'h3b4b9dba),
	.w8(32'hbb75cbdc),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb772493),
	.w1(32'hbb503078),
	.w2(32'hbb827940),
	.w3(32'hbb81c5d6),
	.w4(32'hbba3952a),
	.w5(32'hbb96293b),
	.w6(32'hbb3b1ba1),
	.w7(32'hbbda2c64),
	.w8(32'h3a0c2ec8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc245c51),
	.w1(32'h39fac736),
	.w2(32'h3b062abf),
	.w3(32'h3b0d3b3e),
	.w4(32'h3ba1a604),
	.w5(32'hbb2945c8),
	.w6(32'hbb57d06e),
	.w7(32'hbb312357),
	.w8(32'hbb1f791f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a93ae8),
	.w1(32'hbb8865cc),
	.w2(32'hbb230e3d),
	.w3(32'h3921cf46),
	.w4(32'hba2c001e),
	.w5(32'h3a5918b6),
	.w6(32'hbb976086),
	.w7(32'hba9d9c46),
	.w8(32'h39b2eeb2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc7146),
	.w1(32'hbb98dcc4),
	.w2(32'hbb78a2f4),
	.w3(32'hbb43dd8a),
	.w4(32'hbbab49d0),
	.w5(32'hbb9ef040),
	.w6(32'h399ea4cf),
	.w7(32'h3b12c019),
	.w8(32'h3a9e2bcd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb630d10),
	.w1(32'hbc10508c),
	.w2(32'hbbdf43c1),
	.w3(32'hbb8104c6),
	.w4(32'hbb83c93b),
	.w5(32'hbc21c873),
	.w6(32'h392e6d43),
	.w7(32'hbbdf9365),
	.w8(32'hbbaefa9e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19a8ea),
	.w1(32'hb976c714),
	.w2(32'h3ac5c9fe),
	.w3(32'h3a2b8cb0),
	.w4(32'hba98e7f9),
	.w5(32'hba1fa730),
	.w6(32'h3aca547c),
	.w7(32'hb9918eb9),
	.w8(32'hb8ab875d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c4768),
	.w1(32'hbb080836),
	.w2(32'hbae78fed),
	.w3(32'hbac8b277),
	.w4(32'hbb41fdb7),
	.w5(32'hbb52fee8),
	.w6(32'h39af7c7a),
	.w7(32'hba64fdbc),
	.w8(32'hbadb9584),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c2de),
	.w1(32'hbbbf8e0c),
	.w2(32'hbb86bc99),
	.w3(32'hbb97b7ee),
	.w4(32'hbbbcdb48),
	.w5(32'hbbaf5437),
	.w6(32'hbb8ec221),
	.w7(32'hbb6e3d4c),
	.w8(32'hbba3b516),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a7935),
	.w1(32'h3a51b054),
	.w2(32'h39e1f702),
	.w3(32'hbb2c7e8b),
	.w4(32'h3afa830a),
	.w5(32'h3a8e8c71),
	.w6(32'hba8f8f0b),
	.w7(32'hbab366da),
	.w8(32'h3b19bc4f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a950e4d),
	.w1(32'h39a23235),
	.w2(32'h3ab8899c),
	.w3(32'h392f2d80),
	.w4(32'h39a1ef5f),
	.w5(32'h3abf4bc3),
	.w6(32'hb9243a5e),
	.w7(32'h3ad0fd8f),
	.w8(32'h3b8c10db),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf1ec5),
	.w1(32'hbc2db0e9),
	.w2(32'hbc01cb0c),
	.w3(32'hbc0a6184),
	.w4(32'hbc2b2f56),
	.w5(32'hbbec6a72),
	.w6(32'h3b86a79a),
	.w7(32'h3be5faf2),
	.w8(32'h3a423f51),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a227cac),
	.w1(32'h3926bd76),
	.w2(32'h3a91719a),
	.w3(32'hba01b3f1),
	.w4(32'hb9278404),
	.w5(32'h36f61cc1),
	.w6(32'hb9ae96cb),
	.w7(32'h3aa35838),
	.w8(32'h3ae35169),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8922962),
	.w1(32'hbb6db121),
	.w2(32'hbae9749f),
	.w3(32'hbb9dbb55),
	.w4(32'hbbab81bb),
	.w5(32'hbae0c624),
	.w6(32'hbae5858a),
	.w7(32'hba20f6da),
	.w8(32'h3a961819),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb966547f),
	.w1(32'hb9fa5ed2),
	.w2(32'h39e6ccd9),
	.w3(32'hbaec5bba),
	.w4(32'hbaece4bc),
	.w5(32'hba665120),
	.w6(32'hbb03a666),
	.w7(32'h35489c50),
	.w8(32'hbaae1711),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedfbbc),
	.w1(32'hba52d2ea),
	.w2(32'hbc36aa96),
	.w3(32'hbb37443a),
	.w4(32'hba08522e),
	.w5(32'h3a775fb0),
	.w6(32'hbbb21576),
	.w7(32'hbc078aaa),
	.w8(32'hb9e371d0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01a11c),
	.w1(32'hba5e5c39),
	.w2(32'hb9d047ad),
	.w3(32'hbacbce55),
	.w4(32'hbb03494d),
	.w5(32'hbb17dc20),
	.w6(32'hbadd1d56),
	.w7(32'hbab7f920),
	.w8(32'hb9202228),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa9438),
	.w1(32'hbb3bdb62),
	.w2(32'hb99b7168),
	.w3(32'hbad6592b),
	.w4(32'hba70e21b),
	.w5(32'h3a0f53c5),
	.w6(32'h3aeeaec2),
	.w7(32'h3b4043b7),
	.w8(32'h3ad9726e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc624f),
	.w1(32'hba7cbd9c),
	.w2(32'hb96eab11),
	.w3(32'hbaaaed4f),
	.w4(32'hbac44c38),
	.w5(32'hba915c62),
	.w6(32'hba99c9a2),
	.w7(32'hb92ce36f),
	.w8(32'h3b63c901),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d9e9d),
	.w1(32'hbbf79d3d),
	.w2(32'hbb52c558),
	.w3(32'hbba6781d),
	.w4(32'hbbaf44d2),
	.w5(32'hbb73330c),
	.w6(32'h3bcbf84a),
	.w7(32'h3c0c7cc1),
	.w8(32'h3b41b9ed),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7a462),
	.w1(32'hbb2c3ef9),
	.w2(32'hbb325933),
	.w3(32'hb9bfac0b),
	.w4(32'hba970cde),
	.w5(32'hbb25a9c2),
	.w6(32'h3acf68b7),
	.w7(32'h3b8c457e),
	.w8(32'h39ff4703),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905d2be),
	.w1(32'h38afb34b),
	.w2(32'hba99ef78),
	.w3(32'hba679dc8),
	.w4(32'hba198f05),
	.w5(32'hb9994cdd),
	.w6(32'hb9893832),
	.w7(32'hbad5e26f),
	.w8(32'h3a868449),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d956f),
	.w1(32'h3b248fb0),
	.w2(32'hba781fad),
	.w3(32'hbb2b21e8),
	.w4(32'h3ba73152),
	.w5(32'hbab6d924),
	.w6(32'h3bd63dac),
	.w7(32'h3bb36517),
	.w8(32'hba52b072),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6116b5),
	.w1(32'hbb549abf),
	.w2(32'hba818ecc),
	.w3(32'hbb3f27d3),
	.w4(32'hbabd3d5f),
	.w5(32'h39f29f85),
	.w6(32'hbb5f5a06),
	.w7(32'hb94e2a7c),
	.w8(32'h3aa6f25b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981275b),
	.w1(32'hbbc18d99),
	.w2(32'hbbac3058),
	.w3(32'hbb8076ee),
	.w4(32'hbbd904a7),
	.w5(32'hbb995a85),
	.w6(32'h3afebc82),
	.w7(32'h3aa79c0c),
	.w8(32'h3aba7c17),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e1221),
	.w1(32'hbc402a59),
	.w2(32'hbc40caba),
	.w3(32'hbc05c283),
	.w4(32'hbc06f69a),
	.w5(32'hbbb5959d),
	.w6(32'hbb5c322c),
	.w7(32'hbbb19de9),
	.w8(32'hba16aec2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb599419),
	.w1(32'hbc3941fc),
	.w2(32'hbba38ac9),
	.w3(32'hbbe4be6d),
	.w4(32'hbc305c6e),
	.w5(32'hbb6a71a1),
	.w6(32'h3b99b1de),
	.w7(32'h3b3800c0),
	.w8(32'h3bce2566),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53cc81),
	.w1(32'hbb226ae8),
	.w2(32'hbb0e8556),
	.w3(32'hbb06b3c3),
	.w4(32'hbbc228b7),
	.w5(32'hbbaec8fa),
	.w6(32'h3abce1ef),
	.w7(32'hb99d108d),
	.w8(32'h3ae34f9d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5ebd5),
	.w1(32'h3a18b554),
	.w2(32'h3b753594),
	.w3(32'h3b04b21c),
	.w4(32'h3a9af45c),
	.w5(32'h3b9b4409),
	.w6(32'h3ae4f6b2),
	.w7(32'h3aaf062c),
	.w8(32'h394f6506),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39914f31),
	.w1(32'hbaf2d987),
	.w2(32'h3a5b9b07),
	.w3(32'hb6d6a21b),
	.w4(32'h3aa90b21),
	.w5(32'h3aebc00f),
	.w6(32'hba94eca0),
	.w7(32'h3a332d98),
	.w8(32'hbba93669),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb56a7a),
	.w1(32'hbb4b7944),
	.w2(32'hbb8813db),
	.w3(32'hbb50a3ad),
	.w4(32'hbb71155a),
	.w5(32'hbb5f99f6),
	.w6(32'hbb45e011),
	.w7(32'hbbc555fa),
	.w8(32'h3a22d4f2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6453ff),
	.w1(32'hba8c2271),
	.w2(32'h3a965037),
	.w3(32'h3af46415),
	.w4(32'hbb5079f6),
	.w5(32'h3ad0d343),
	.w6(32'h3b7e269c),
	.w7(32'h3a66d13e),
	.w8(32'h3a5bfc11),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c3412),
	.w1(32'hba4b454d),
	.w2(32'h3b1b2258),
	.w3(32'hbaaa7d4b),
	.w4(32'hbac21ee6),
	.w5(32'h3b0ca07d),
	.w6(32'hba98767b),
	.w7(32'h3a3e3260),
	.w8(32'hbaa5ddab),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a858d1e),
	.w1(32'hba0dc223),
	.w2(32'hb9581361),
	.w3(32'h3a4c78c2),
	.w4(32'hbaa89c9c),
	.w5(32'hba537bc9),
	.w6(32'hba3dfcbd),
	.w7(32'hba1de5c5),
	.w8(32'hbbacbdf1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc241e36),
	.w1(32'hbb8983ed),
	.w2(32'hbaf8a5d8),
	.w3(32'hbbac3c59),
	.w4(32'hb85471ae),
	.w5(32'hbb01a80c),
	.w6(32'h3aa993a6),
	.w7(32'hbb44e07f),
	.w8(32'h3aa4601b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4edeec),
	.w1(32'hbb89f48d),
	.w2(32'hbb2add21),
	.w3(32'hbbc32390),
	.w4(32'hbbb99cff),
	.w5(32'hbb92c83d),
	.w6(32'hbb8d758b),
	.w7(32'hbb7ea62a),
	.w8(32'hba1ec423),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e396c),
	.w1(32'hbbc85e50),
	.w2(32'hbc184732),
	.w3(32'hba01fb11),
	.w4(32'h39b4dbbe),
	.w5(32'h3982ffe1),
	.w6(32'h3ab74cee),
	.w7(32'hbb0866ab),
	.w8(32'hbb1fc39c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ef7f0),
	.w1(32'h3b700901),
	.w2(32'h3b866fe5),
	.w3(32'h3b3fef72),
	.w4(32'hb98253ac),
	.w5(32'h3abc0a84),
	.w6(32'h3bb46f3f),
	.w7(32'h3b760b77),
	.w8(32'h3c0d68ee),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef54a5),
	.w1(32'hbbbd1eef),
	.w2(32'hbaa456f0),
	.w3(32'hbbb2d51d),
	.w4(32'hbba84b7a),
	.w5(32'h3a8a1d63),
	.w6(32'h3c2629f5),
	.w7(32'h3b995e9c),
	.w8(32'h3bc071c5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4ce3),
	.w1(32'hba872a5c),
	.w2(32'hbae6f46d),
	.w3(32'h39c654e3),
	.w4(32'h3a56a2e6),
	.w5(32'h3939ec9b),
	.w6(32'h3ad4da80),
	.w7(32'hbae77dc9),
	.w8(32'h3b4b6e9e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9674972),
	.w1(32'hba0c2498),
	.w2(32'h3aa8b77f),
	.w3(32'hbaac6c17),
	.w4(32'h39886b88),
	.w5(32'hb943e956),
	.w6(32'h3b3f077c),
	.w7(32'h3bd7e90b),
	.w8(32'hb82c6792),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c378a),
	.w1(32'hba7e6e57),
	.w2(32'hb953af5d),
	.w3(32'hba2a7ff1),
	.w4(32'h39b80a44),
	.w5(32'h399d2d47),
	.w6(32'hba0a932f),
	.w7(32'h3a4a28ed),
	.w8(32'hbae5963e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ba199),
	.w1(32'hbaf97a24),
	.w2(32'hbb7f8b77),
	.w3(32'hbac1e1e6),
	.w4(32'hbb0cb324),
	.w5(32'hbba306ba),
	.w6(32'hb99f890f),
	.w7(32'hbbb0b088),
	.w8(32'hba2b42da),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9d9bf),
	.w1(32'hbb573829),
	.w2(32'hbb14c708),
	.w3(32'hbb1cfdb8),
	.w4(32'hbb35ce84),
	.w5(32'hbb2859df),
	.w6(32'h38b71c26),
	.w7(32'h3a60eeb6),
	.w8(32'h3b5c742d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2177f),
	.w1(32'hbaddf0bb),
	.w2(32'h3965277d),
	.w3(32'h3a9d1429),
	.w4(32'h3aa9aa27),
	.w5(32'h3ac46036),
	.w6(32'h3ae3d2e3),
	.w7(32'h3c004da9),
	.w8(32'h39dc96d2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d823e),
	.w1(32'hb9db1dfd),
	.w2(32'h3a32be43),
	.w3(32'hbb337eb2),
	.w4(32'hbaa953e5),
	.w5(32'hba9171c9),
	.w6(32'hbb6ef3e3),
	.w7(32'hbb416c42),
	.w8(32'hb8497d0e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f52a5),
	.w1(32'h39922d39),
	.w2(32'h3a2cf747),
	.w3(32'h38a072d4),
	.w4(32'hb9165b95),
	.w5(32'h398e2d47),
	.w6(32'hba8d68d9),
	.w7(32'hbaa7e6eb),
	.w8(32'hba9eacea),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dd4e3),
	.w1(32'hbc0a219f),
	.w2(32'hbba92004),
	.w3(32'hbbdd893b),
	.w4(32'hbc290bc0),
	.w5(32'hbbb4c167),
	.w6(32'hb9e285d4),
	.w7(32'hbb22bb0f),
	.w8(32'hbaaf3691),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef8db7),
	.w1(32'hbb176b2c),
	.w2(32'hbaa42db6),
	.w3(32'hbb554cd5),
	.w4(32'hbb938c03),
	.w5(32'h39428fdb),
	.w6(32'h3b164be7),
	.w7(32'hbb1b2fba),
	.w8(32'h399388c3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b698f2),
	.w1(32'hbae2a083),
	.w2(32'hbaaadcdf),
	.w3(32'hbb6419ac),
	.w4(32'hbb5e261c),
	.w5(32'hbb4f8fd7),
	.w6(32'hbb156435),
	.w7(32'hbb56a499),
	.w8(32'hbac4aaa0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab77855),
	.w1(32'h3b4fb049),
	.w2(32'h3b0ea440),
	.w3(32'h3a8fce62),
	.w4(32'h3b24e9db),
	.w5(32'h3b16ae50),
	.w6(32'h37e1661f),
	.w7(32'h3b200280),
	.w8(32'h3b4c7ded),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf1bf3),
	.w1(32'hbbf5c1f4),
	.w2(32'hbb451712),
	.w3(32'hbb724031),
	.w4(32'hbb8a406c),
	.w5(32'hb8d22177),
	.w6(32'h3a8fd83c),
	.w7(32'h38c5442f),
	.w8(32'hbb5e259f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ab42),
	.w1(32'hb7f93db3),
	.w2(32'hbb1653e5),
	.w3(32'hba29b052),
	.w4(32'h3b88423a),
	.w5(32'h3ac9a4c0),
	.w6(32'h3aab9891),
	.w7(32'h3b1b09e5),
	.w8(32'h3a64ad13),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdab5e5),
	.w1(32'hbbbeaaff),
	.w2(32'hbbb948e4),
	.w3(32'hbbb06722),
	.w4(32'hbb4356d7),
	.w5(32'hbb4fdc9b),
	.w6(32'hbb4423de),
	.w7(32'hbb322bb6),
	.w8(32'hbb834ec6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cec33),
	.w1(32'h3acbbb79),
	.w2(32'h3b1cb386),
	.w3(32'h3af889b1),
	.w4(32'h3b13379f),
	.w5(32'h3b072435),
	.w6(32'hbb28b610),
	.w7(32'hbac78c91),
	.w8(32'hb9fd1e1a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b52a6),
	.w1(32'hba691638),
	.w2(32'h39719071),
	.w3(32'h380a5ff4),
	.w4(32'hba41a75a),
	.w5(32'h35e2b772),
	.w6(32'h3a18805a),
	.w7(32'h3a3f42de),
	.w8(32'h39accc36),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38864b59),
	.w1(32'hb9cb191e),
	.w2(32'hb7e9eb9c),
	.w3(32'hb9adb3ff),
	.w4(32'hba3f4f5d),
	.w5(32'hb9a9498b),
	.w6(32'hb88ae1dd),
	.w7(32'h37be4560),
	.w8(32'h3a7e2314),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a623cf6),
	.w1(32'h38d7b74f),
	.w2(32'hb9b6f38f),
	.w3(32'h3a0a8e1a),
	.w4(32'h39dfcb49),
	.w5(32'hb92cb151),
	.w6(32'h3b20698d),
	.w7(32'h3b1c53b0),
	.w8(32'h390cabf7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdeeb9),
	.w1(32'hbae40da4),
	.w2(32'hbbef74df),
	.w3(32'h3b07df3e),
	.w4(32'h3a0106e4),
	.w5(32'hbb17fad3),
	.w6(32'hbb187aff),
	.w7(32'hbaf847bb),
	.w8(32'h3a5b254d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad505ed),
	.w1(32'hbab12f51),
	.w2(32'h38614b19),
	.w3(32'hb9d00266),
	.w4(32'h3a29151c),
	.w5(32'h3ac5e63d),
	.w6(32'hbb11c0a1),
	.w7(32'hba17fbc9),
	.w8(32'hbb1a7024),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e2e95),
	.w1(32'hbb9958fd),
	.w2(32'hbb94a108),
	.w3(32'hbb89c7c5),
	.w4(32'hbab3dfe8),
	.w5(32'h3b02a8d0),
	.w6(32'hbb8d5423),
	.w7(32'hbb9b96d2),
	.w8(32'h39620a28),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa19628),
	.w1(32'hba7f4252),
	.w2(32'hbb0a5852),
	.w3(32'hbac372a5),
	.w4(32'hbb1b581a),
	.w5(32'hbb61aa7d),
	.w6(32'hbb100511),
	.w7(32'hba550723),
	.w8(32'hbae7a8be),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a746733),
	.w1(32'h38395f2a),
	.w2(32'hba62c910),
	.w3(32'hbb5c1f97),
	.w4(32'hbb866579),
	.w5(32'hbb8dd3f2),
	.w6(32'hbb1a5be9),
	.w7(32'h39755d37),
	.w8(32'h3a05de75),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b3adc),
	.w1(32'hbb9bb525),
	.w2(32'hbc142746),
	.w3(32'h3aa9b967),
	.w4(32'hbb01fd73),
	.w5(32'hba6dcdfd),
	.w6(32'h3b6c6db3),
	.w7(32'hb9a47aca),
	.w8(32'hbb783beb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17c474),
	.w1(32'hba076746),
	.w2(32'hb720ef48),
	.w3(32'hb9b4cd80),
	.w4(32'h3a43663c),
	.w5(32'h3a391a05),
	.w6(32'hb97ce0f1),
	.w7(32'hb979c9f3),
	.w8(32'h370777f0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40db48),
	.w1(32'h3b94cf1b),
	.w2(32'h3b8743c8),
	.w3(32'h3b182246),
	.w4(32'h3b093f90),
	.w5(32'h3b1c41be),
	.w6(32'h3a8411f7),
	.w7(32'h3a41544c),
	.w8(32'hb9d021e9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf549fa),
	.w1(32'hbb597ab2),
	.w2(32'hbb22d4e9),
	.w3(32'hbb0d2e02),
	.w4(32'h3bad66e2),
	.w5(32'h3b650012),
	.w6(32'hbb43ddc7),
	.w7(32'hbb2568d0),
	.w8(32'hb8837236),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb148df2),
	.w1(32'hbb61176c),
	.w2(32'hba56eba5),
	.w3(32'hbaf9da0a),
	.w4(32'hba846817),
	.w5(32'h3a4e3c77),
	.w6(32'hbae498eb),
	.w7(32'hb9d35d90),
	.w8(32'h3b0719de),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a437bdb),
	.w1(32'h393a7912),
	.w2(32'h39dbce7b),
	.w3(32'h3abf85e6),
	.w4(32'h3af6374c),
	.w5(32'h39cc2eb8),
	.w6(32'h3b13a0c3),
	.w7(32'h3b228980),
	.w8(32'hb7f9c806),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b645aee),
	.w1(32'h3c2e7ce2),
	.w2(32'h3bbdf89d),
	.w3(32'hbabc4804),
	.w4(32'h3a9799d4),
	.w5(32'h3a456dab),
	.w6(32'hbadaf0cb),
	.w7(32'hb990c71f),
	.w8(32'h378de62b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule