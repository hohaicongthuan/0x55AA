module layer_10_featuremap_507(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf6be4),
	.w1(32'hbcc00436),
	.w2(32'hbb2f7632),
	.w3(32'h3bcc5769),
	.w4(32'hbc02bfec),
	.w5(32'h3cfe16cc),
	.w6(32'h3abce111),
	.w7(32'hbc0535c4),
	.w8(32'hbb88f074),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe41e6),
	.w1(32'h3b4f66e3),
	.w2(32'h3c11bd26),
	.w3(32'h3ac26fcb),
	.w4(32'hbcfe2ea0),
	.w5(32'hbc39cfc6),
	.w6(32'hbbbedc5b),
	.w7(32'hbbac093f),
	.w8(32'hba38ca57),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b33d4),
	.w1(32'hbbbb78ed),
	.w2(32'hbca36bc6),
	.w3(32'hb9c6998f),
	.w4(32'h3cde0351),
	.w5(32'h3bf9b309),
	.w6(32'hbc0886c2),
	.w7(32'hbc1c0a14),
	.w8(32'hbc9c3bd8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11d34a),
	.w1(32'h3b0bc356),
	.w2(32'hbbfc0a1b),
	.w3(32'h3b24372e),
	.w4(32'hbbd85760),
	.w5(32'hbcbe22c0),
	.w6(32'h3c671272),
	.w7(32'h3a62b601),
	.w8(32'hbc39d420),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b0010),
	.w1(32'h39668730),
	.w2(32'hbaedd0c8),
	.w3(32'h3c076d6e),
	.w4(32'h3be50580),
	.w5(32'h3ad85022),
	.w6(32'h3ae727c4),
	.w7(32'h3c010390),
	.w8(32'h3b424e2a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6eee9e),
	.w1(32'h3c3c4769),
	.w2(32'hbc7e36dc),
	.w3(32'hbcb19885),
	.w4(32'h3c1cbbcd),
	.w5(32'h3ba86910),
	.w6(32'h3ba44b48),
	.w7(32'hbc286d88),
	.w8(32'hbc5d7f9c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8241bb),
	.w1(32'h3c21e100),
	.w2(32'h3bea56c3),
	.w3(32'h3c1c8a23),
	.w4(32'hbbafab9c),
	.w5(32'hbb434113),
	.w6(32'hbbcaae08),
	.w7(32'h3d4934dc),
	.w8(32'hb9c0014c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e0539),
	.w1(32'h3c65017a),
	.w2(32'h3b95d146),
	.w3(32'hbca89147),
	.w4(32'hbb6136ab),
	.w5(32'hbc56c8e5),
	.w6(32'hbc4efe9a),
	.w7(32'hbc7e255b),
	.w8(32'hbce4513f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb365311),
	.w1(32'h3c6b89e3),
	.w2(32'h3c228820),
	.w3(32'h3bad90cc),
	.w4(32'h3bfbf1fa),
	.w5(32'h3bea9480),
	.w6(32'hbc07c11e),
	.w7(32'hbc300a31),
	.w8(32'h3bfb25fd),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63f683),
	.w1(32'h3c933f13),
	.w2(32'h3cc40c4b),
	.w3(32'h3c2ba20d),
	.w4(32'hbbb1b31d),
	.w5(32'h3c2b7837),
	.w6(32'hbbaad265),
	.w7(32'h3b7d7a61),
	.w8(32'hbc857352),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56d539),
	.w1(32'h3bbf0818),
	.w2(32'hbc47921c),
	.w3(32'hb9d46dcd),
	.w4(32'h3bf524f4),
	.w5(32'hbb99a28a),
	.w6(32'h3c935e9b),
	.w7(32'hbc7bd370),
	.w8(32'h3b50d432),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c21d9),
	.w1(32'hbbe0c57d),
	.w2(32'hba76a3ba),
	.w3(32'h3b4ba91b),
	.w4(32'h3be146da),
	.w5(32'hbbc43bba),
	.w6(32'hbc7ae330),
	.w7(32'h3861904b),
	.w8(32'h3c039ccd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6aa7b),
	.w1(32'hbc345b4d),
	.w2(32'h3c48541a),
	.w3(32'hbc520f43),
	.w4(32'hbc214951),
	.w5(32'hb98eb4ca),
	.w6(32'h3c9043d8),
	.w7(32'hbbfb1e3b),
	.w8(32'hbbe7e609),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ce05d),
	.w1(32'hbc3fa44f),
	.w2(32'hb9e58c84),
	.w3(32'h3b2d71a0),
	.w4(32'hbc5075b4),
	.w5(32'hbc50544f),
	.w6(32'hbc1c9ffc),
	.w7(32'h3c3945a8),
	.w8(32'h3c301403),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47a777),
	.w1(32'h3c7d8e26),
	.w2(32'h3c5cb1eb),
	.w3(32'h3c5af2bc),
	.w4(32'hbb6c3d2d),
	.w5(32'hbbc7ae86),
	.w6(32'h3c0c12e3),
	.w7(32'hb9982c2c),
	.w8(32'h3c6180a3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5c4e1),
	.w1(32'hbc3b34d4),
	.w2(32'h3cadac11),
	.w3(32'hbc0335a3),
	.w4(32'hbb1822e9),
	.w5(32'h3b0a8264),
	.w6(32'hbbf9bb17),
	.w7(32'hbc3bd488),
	.w8(32'h3a38b570),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2138b0),
	.w1(32'h39c80dfd),
	.w2(32'hbbb28699),
	.w3(32'h3b94bcc6),
	.w4(32'h3a23119f),
	.w5(32'h3be96eaf),
	.w6(32'hbbdcde9c),
	.w7(32'hbc965b9f),
	.w8(32'hb95cf1f9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2394dc),
	.w1(32'hbb299009),
	.w2(32'hbc3062c7),
	.w3(32'hbd1573d5),
	.w4(32'hbcd2c5e1),
	.w5(32'hbc97083d),
	.w6(32'hbc211235),
	.w7(32'hbcd3059f),
	.w8(32'hbd0e8ded),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b067b),
	.w1(32'h3b180f45),
	.w2(32'hbc61719b),
	.w3(32'hbc1b83b0),
	.w4(32'hbc43f636),
	.w5(32'hbc6dbf8c),
	.w6(32'hbbcefe1b),
	.w7(32'hbc147297),
	.w8(32'hbcbfca11),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3826af),
	.w1(32'h3b84d1fc),
	.w2(32'hbb0a23a9),
	.w3(32'hbb79d1b0),
	.w4(32'hbbce5a6a),
	.w5(32'h3be3f845),
	.w6(32'h3a966d5f),
	.w7(32'h3aac5075),
	.w8(32'h3b18f75d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b251d03),
	.w1(32'hbba2b59b),
	.w2(32'h3b996be9),
	.w3(32'hbc49a251),
	.w4(32'h3ba69d83),
	.w5(32'hbc77d3ce),
	.w6(32'h3c014312),
	.w7(32'hb9ff940b),
	.w8(32'h3bad84d1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72e7cd),
	.w1(32'hba530991),
	.w2(32'hbc300609),
	.w3(32'h3c091b09),
	.w4(32'hbbac2b0f),
	.w5(32'h3b15d642),
	.w6(32'h3c82b520),
	.w7(32'h3ba27577),
	.w8(32'h3c30837f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fa8b7),
	.w1(32'hbca27147),
	.w2(32'hbc65ef3e),
	.w3(32'hbd1b5b65),
	.w4(32'hbca7aff5),
	.w5(32'hbc562680),
	.w6(32'hbcb85fb0),
	.w7(32'hbc9ab626),
	.w8(32'hbcfde8a9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4420f),
	.w1(32'hbb26d04d),
	.w2(32'h3c4db139),
	.w3(32'h3b789f4a),
	.w4(32'hba38939d),
	.w5(32'hbb6db28f),
	.w6(32'h3ba97fdf),
	.w7(32'h3c10476a),
	.w8(32'h3b97e694),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdba950),
	.w1(32'h3c28191f),
	.w2(32'h3c75e08c),
	.w3(32'h3b5471cd),
	.w4(32'h3b20d0f2),
	.w5(32'h3c17745e),
	.w6(32'h3c23495e),
	.w7(32'h39428cff),
	.w8(32'h3ba23ef9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69279f),
	.w1(32'hbcb6c907),
	.w2(32'h3b9690ec),
	.w3(32'hbbd170e4),
	.w4(32'h3c5ece77),
	.w5(32'hbcd95b2b),
	.w6(32'h3c6a5c7d),
	.w7(32'h3a3c6178),
	.w8(32'hbc41499a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd127a20),
	.w1(32'h3bd407ab),
	.w2(32'hbb4882a6),
	.w3(32'hbc075845),
	.w4(32'hbc0cc614),
	.w5(32'h3b81e7c9),
	.w6(32'hbc86d8fa),
	.w7(32'hbb2eb222),
	.w8(32'hbc071f65),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e7f29),
	.w1(32'hbac885f8),
	.w2(32'h3a57fd27),
	.w3(32'h3cd50e60),
	.w4(32'hbca27a98),
	.w5(32'h3bb2896d),
	.w6(32'h3d739669),
	.w7(32'h3a9d73d5),
	.w8(32'hbaae5f31),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa74118),
	.w1(32'hbc984c9c),
	.w2(32'h3a2f344c),
	.w3(32'h3be868fc),
	.w4(32'h3cc89b1c),
	.w5(32'hbce8c3de),
	.w6(32'hbaacb45c),
	.w7(32'hbc66acf2),
	.w8(32'h3af5bf87),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67c24e),
	.w1(32'h3c899c70),
	.w2(32'h3a576d56),
	.w3(32'h3c8def3a),
	.w4(32'h3b92a9a4),
	.w5(32'h3d0963c5),
	.w6(32'h3c1b9673),
	.w7(32'hbc08d786),
	.w8(32'h3d00547c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2607d),
	.w1(32'hbc7345f5),
	.w2(32'hbba65f94),
	.w3(32'hbb621472),
	.w4(32'h3c2960ba),
	.w5(32'h3bbb96cc),
	.w6(32'hbc3d3f6e),
	.w7(32'h3bc9bfa2),
	.w8(32'hbc391200),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9f2c0),
	.w1(32'hbbd02717),
	.w2(32'hbbe23b35),
	.w3(32'hb9c18964),
	.w4(32'h3c1a7fc9),
	.w5(32'hbb22efa8),
	.w6(32'h3cd8b65e),
	.w7(32'hbb2d41cc),
	.w8(32'hbb99a65f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936566),
	.w1(32'hbc83b683),
	.w2(32'h3cce2e28),
	.w3(32'hbbbf60e4),
	.w4(32'h3caaeb7a),
	.w5(32'hba85580a),
	.w6(32'hbc0754c8),
	.w7(32'h3a881eff),
	.w8(32'h3bb8def4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e8b70),
	.w1(32'hbb789a3c),
	.w2(32'hbb1fa8c7),
	.w3(32'h3d09c0d9),
	.w4(32'hbc156e52),
	.w5(32'h3c97bb02),
	.w6(32'h3aeee82b),
	.w7(32'h3d8d06c5),
	.w8(32'hb997b6f2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69971f),
	.w1(32'h3c6034da),
	.w2(32'hbca71df0),
	.w3(32'hbc805949),
	.w4(32'hbc1d7f3e),
	.w5(32'h3b7c1050),
	.w6(32'hbc65ad69),
	.w7(32'h3bf07238),
	.w8(32'h39fb705c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bbeb5),
	.w1(32'hbad210f4),
	.w2(32'hbc710263),
	.w3(32'hbba7df9b),
	.w4(32'h3afe39dc),
	.w5(32'h3b08b73f),
	.w6(32'h3991ac66),
	.w7(32'hbb9c6885),
	.w8(32'hbbb45405),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be35597),
	.w1(32'h3bd0e46a),
	.w2(32'h3b6c7528),
	.w3(32'hb996c712),
	.w4(32'h3ba2027b),
	.w5(32'h3b74ba97),
	.w6(32'hbc12f444),
	.w7(32'h3c089ab4),
	.w8(32'hbcdda1b3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd91ef4),
	.w1(32'h3c539518),
	.w2(32'h3baf3c0c),
	.w3(32'h3c2db622),
	.w4(32'h3c50b56d),
	.w5(32'h3b997a5f),
	.w6(32'hbb4231c6),
	.w7(32'h3bf7e306),
	.w8(32'hbb0ae601),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c583347),
	.w1(32'hbc1ea763),
	.w2(32'hbae0e922),
	.w3(32'h3c96ff6e),
	.w4(32'h3b6fc3f1),
	.w5(32'hba6c4751),
	.w6(32'h3c336401),
	.w7(32'h3c5d8ba3),
	.w8(32'h3a0c8101),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78dc26),
	.w1(32'h3c209ecc),
	.w2(32'hbbfe70ae),
	.w3(32'h3ba0347a),
	.w4(32'h3b553e78),
	.w5(32'h3bdbe855),
	.w6(32'h3a369ac6),
	.w7(32'h3b9a6274),
	.w8(32'hbc714531),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e73d8f),
	.w1(32'hbc6d5f36),
	.w2(32'hba9bef05),
	.w3(32'hbb29545f),
	.w4(32'hbb0c698a),
	.w5(32'h3cb73831),
	.w6(32'h3b3eb2a3),
	.w7(32'h3c96de19),
	.w8(32'h3c01a06b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98420fd),
	.w1(32'hb9191c80),
	.w2(32'hbb5dc0d5),
	.w3(32'hbc1398df),
	.w4(32'h3ade6c99),
	.w5(32'h3b3e4f79),
	.w6(32'hbc1aad77),
	.w7(32'h3c0ab849),
	.w8(32'h3bc24696),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0737b7),
	.w1(32'hbbb17904),
	.w2(32'hb9f9cabd),
	.w3(32'h3c1309a3),
	.w4(32'hbbcf5c84),
	.w5(32'h3cb0801f),
	.w6(32'hbbcd0a8d),
	.w7(32'hbc794962),
	.w8(32'hbbcee358),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2a551),
	.w1(32'hbb64f448),
	.w2(32'hbc16e26d),
	.w3(32'h3b8949e7),
	.w4(32'hbaaa4811),
	.w5(32'h3b7e2d87),
	.w6(32'h3d11e4f5),
	.w7(32'hbb88e0d5),
	.w8(32'hba81cc37),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e03ee),
	.w1(32'h3bfbfaac),
	.w2(32'hbbbcd559),
	.w3(32'h381008f0),
	.w4(32'h3c0f1f15),
	.w5(32'h3bc83256),
	.w6(32'h3b1e8aa2),
	.w7(32'h3c485f25),
	.w8(32'h3c1c19d9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cbaa9),
	.w1(32'h3aa49ad4),
	.w2(32'h3cdb0daa),
	.w3(32'h3b8049c4),
	.w4(32'h3c29b3be),
	.w5(32'h3caadce4),
	.w6(32'h3b90d9f2),
	.w7(32'hba72d9c2),
	.w8(32'hbc195c66),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdda585),
	.w1(32'hbb05aa4c),
	.w2(32'h3a686d0e),
	.w3(32'hb8acf2f4),
	.w4(32'h3b7a8c07),
	.w5(32'h39bdd401),
	.w6(32'h3b15b1fb),
	.w7(32'hba76af3a),
	.w8(32'hba814acb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c9ebf),
	.w1(32'hbc008a71),
	.w2(32'hbc9e2eb5),
	.w3(32'hbca3b21b),
	.w4(32'hbcb8aa7e),
	.w5(32'hbcafa666),
	.w6(32'hbce389dd),
	.w7(32'hbcd9b0eb),
	.w8(32'hbc8fd217),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb837a45),
	.w1(32'hbb9ee1c7),
	.w2(32'hb8e2327b),
	.w3(32'h3c03a76e),
	.w4(32'h3c3e7bf5),
	.w5(32'h3ca50a03),
	.w6(32'h3c40a71d),
	.w7(32'h3b6038f0),
	.w8(32'hbbe45d5c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91b1dc),
	.w1(32'h3be09c71),
	.w2(32'h3b87e4af),
	.w3(32'h3bb03047),
	.w4(32'hbba5fa6b),
	.w5(32'h3c08681f),
	.w6(32'h3b8b870f),
	.w7(32'h3a8399b2),
	.w8(32'hbb94080f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0931fa),
	.w1(32'h3b65b9f0),
	.w2(32'h3b516870),
	.w3(32'hbb9f9d42),
	.w4(32'h3cc5499d),
	.w5(32'h3bbbf07f),
	.w6(32'h3ade1750),
	.w7(32'hbb8cd452),
	.w8(32'h3b94d79d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64e89e),
	.w1(32'hbb1f6b19),
	.w2(32'hbcacb376),
	.w3(32'h3b4471e0),
	.w4(32'h3b9dfbef),
	.w5(32'h39b8d70c),
	.w6(32'hbc14e7c8),
	.w7(32'hbca15e98),
	.w8(32'h3c9e3bb5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd57489),
	.w1(32'hbbe12703),
	.w2(32'hbc151739),
	.w3(32'hb945ae1a),
	.w4(32'h3be41c42),
	.w5(32'hba0a73b1),
	.w6(32'hbd082a91),
	.w7(32'hbca7b11f),
	.w8(32'hbbe0dfd5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf0615),
	.w1(32'hbbaae754),
	.w2(32'hbac32873),
	.w3(32'hbc9759d2),
	.w4(32'hbcdbee74),
	.w5(32'h3c463f67),
	.w6(32'hbc968092),
	.w7(32'hbcda9152),
	.w8(32'hbc2c0731),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc138efe),
	.w1(32'hbc8da0c4),
	.w2(32'hb8ff3d64),
	.w3(32'h3b191f50),
	.w4(32'hbcf916a1),
	.w5(32'hbc67cf4f),
	.w6(32'h3bec1d65),
	.w7(32'hbbcce8ef),
	.w8(32'hbb234474),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18d103),
	.w1(32'h3b13ae82),
	.w2(32'hb6b55c51),
	.w3(32'hbbc0969e),
	.w4(32'h3b9a6212),
	.w5(32'hbb12f2b7),
	.w6(32'h3c66ba70),
	.w7(32'hbc96017c),
	.w8(32'h3b9c92a9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847bcf),
	.w1(32'hbb732639),
	.w2(32'h3c6d1d69),
	.w3(32'h3ab7814d),
	.w4(32'hbc109ecc),
	.w5(32'hbc1d035e),
	.w6(32'h3ad9ccf8),
	.w7(32'h3c9e431c),
	.w8(32'h3cc60fac),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07e359),
	.w1(32'hbbc010fc),
	.w2(32'h3b89b462),
	.w3(32'h3ac01f19),
	.w4(32'h3c2676e4),
	.w5(32'hbaaf6b85),
	.w6(32'h3b16e080),
	.w7(32'hbc2048ea),
	.w8(32'hba897a8a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a7b04),
	.w1(32'hbc108940),
	.w2(32'h3a7ff8eb),
	.w3(32'hbc5bc0c2),
	.w4(32'h3c8f313e),
	.w5(32'hb9e4b42e),
	.w6(32'hbc1e1a83),
	.w7(32'hbbb270f8),
	.w8(32'hbbc23e72),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e9370),
	.w1(32'hbbd3714e),
	.w2(32'h3b2da33c),
	.w3(32'h3a0bd8f5),
	.w4(32'h3c585c5f),
	.w5(32'hbbd302ba),
	.w6(32'h3bd4b5c9),
	.w7(32'hbc653478),
	.w8(32'hbb9cf474),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f35b),
	.w1(32'hbc326938),
	.w2(32'hbc81de7e),
	.w3(32'hbcb9de0b),
	.w4(32'hbc47c581),
	.w5(32'hbc4b6449),
	.w6(32'hbb892f2d),
	.w7(32'h3b671600),
	.w8(32'hbc843efa),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75a431),
	.w1(32'hbcc252ad),
	.w2(32'hbb9a5536),
	.w3(32'hbc46cea7),
	.w4(32'hbb3a9e00),
	.w5(32'hbc0a3781),
	.w6(32'h3b3be0cb),
	.w7(32'hbc5efe5d),
	.w8(32'hbc3f0a17),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaabef2),
	.w1(32'hbc10270f),
	.w2(32'h3cbe0a6f),
	.w3(32'hbb7eaff3),
	.w4(32'hba8615a0),
	.w5(32'hbc8e2ba6),
	.w6(32'h3b6964de),
	.w7(32'hbbc23035),
	.w8(32'hbbd2f7b9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07d74a),
	.w1(32'hbb8d4f79),
	.w2(32'hbaee6499),
	.w3(32'hbb410641),
	.w4(32'h3827e6be),
	.w5(32'h3ba0369a),
	.w6(32'hba31600b),
	.w7(32'h3bb98bda),
	.w8(32'hbb91ef5f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c68d7),
	.w1(32'hbc19e693),
	.w2(32'hbb90ef4b),
	.w3(32'h3c56a5ce),
	.w4(32'hbb8ab7a2),
	.w5(32'h3c10f4cc),
	.w6(32'hbb4ed4de),
	.w7(32'h3d03cc57),
	.w8(32'h3ad2f0e8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93f8cc),
	.w1(32'h3c18373c),
	.w2(32'hbaff5aa6),
	.w3(32'hbc46263e),
	.w4(32'hbbb43119),
	.w5(32'hbafd7cd0),
	.w6(32'h3c285ec9),
	.w7(32'hbb88f570),
	.w8(32'h3be43165),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30eb33),
	.w1(32'h3b21c0d1),
	.w2(32'h3bee48c8),
	.w3(32'hbc69e058),
	.w4(32'h3c7638b1),
	.w5(32'h3b489568),
	.w6(32'hbbba6e13),
	.w7(32'hbcc83aa4),
	.w8(32'hbc420c19),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cca2515),
	.w1(32'h3c482027),
	.w2(32'h3c37a39e),
	.w3(32'hbc0ed1d9),
	.w4(32'h3c7e055c),
	.w5(32'hbbebd41d),
	.w6(32'hbbaab5af),
	.w7(32'hbb09d143),
	.w8(32'h3c4b35fa),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cb1fa),
	.w1(32'h3a1c2ff3),
	.w2(32'hbc4432c1),
	.w3(32'hbc650d5d),
	.w4(32'hbc1fa9b1),
	.w5(32'hbc7c7ed1),
	.w6(32'hbc72d811),
	.w7(32'hbc76455d),
	.w8(32'hbd483d1e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f0d88),
	.w1(32'h3c316ce9),
	.w2(32'h3c32542a),
	.w3(32'h3b6c0b24),
	.w4(32'h3aa31f21),
	.w5(32'h3c9418d9),
	.w6(32'h3c8066d4),
	.w7(32'h3caa9b74),
	.w8(32'h3cdfc1d2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8357ef),
	.w1(32'h3bd2b7f3),
	.w2(32'hb9fb92c7),
	.w3(32'hbc75e898),
	.w4(32'h3ba3a322),
	.w5(32'h3c8916d9),
	.w6(32'h3c07c4a8),
	.w7(32'hbc8ad774),
	.w8(32'hbbb834cd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c891f49),
	.w1(32'hb9d41ea2),
	.w2(32'hbc0e2ef3),
	.w3(32'hb9f2214f),
	.w4(32'h3bbb9acf),
	.w5(32'h3c338269),
	.w6(32'h3d2989b5),
	.w7(32'h39ff6ca1),
	.w8(32'h3c307d79),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0b25d),
	.w1(32'hbbc66d12),
	.w2(32'h3a11657d),
	.w3(32'h3acbd507),
	.w4(32'hbc5fc436),
	.w5(32'h3bd9f026),
	.w6(32'h3b9d1a67),
	.w7(32'h3b6ad37a),
	.w8(32'h3c0725cd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad65877),
	.w1(32'hbb3f65d9),
	.w2(32'h3bfc0a05),
	.w3(32'h3ba58b99),
	.w4(32'h3b56a5fb),
	.w5(32'hbc36a872),
	.w6(32'hbbb9a65c),
	.w7(32'hbc41829b),
	.w8(32'hbc734d2f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b246d49),
	.w1(32'h3a7457e9),
	.w2(32'h3a863629),
	.w3(32'h3c94ff88),
	.w4(32'h3b776b48),
	.w5(32'h3bada7eb),
	.w6(32'hbad5fdc8),
	.w7(32'h3bc47d2e),
	.w8(32'h3bbc957f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21d0b5),
	.w1(32'hbc054a31),
	.w2(32'hbc535138),
	.w3(32'hbc406f8a),
	.w4(32'hbc0ffa1a),
	.w5(32'h3ba29a01),
	.w6(32'hbc77e64f),
	.w7(32'hbbb4215d),
	.w8(32'hbc446dd1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc712759),
	.w1(32'h3c53af3c),
	.w2(32'hbcb0830d),
	.w3(32'hbcc93d4e),
	.w4(32'hbc830fe2),
	.w5(32'hbcd1ffb9),
	.w6(32'hbc8b8b08),
	.w7(32'hbccd4f88),
	.w8(32'hbc39512e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a058d34),
	.w1(32'h3c80c6ab),
	.w2(32'hbc74c174),
	.w3(32'h3cc7c203),
	.w4(32'h3c4db098),
	.w5(32'h3b35f5df),
	.w6(32'h350030a4),
	.w7(32'hbb5b3a39),
	.w8(32'h3c680865),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9193916),
	.w1(32'h3b0019d9),
	.w2(32'h3c133133),
	.w3(32'hbbd7a597),
	.w4(32'hbb4c6f37),
	.w5(32'h3c1e91f0),
	.w6(32'hbb35a557),
	.w7(32'hbbd61de1),
	.w8(32'hbaf8e434),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb848835),
	.w1(32'hbbc6b161),
	.w2(32'hbbc6256d),
	.w3(32'hbb81fd52),
	.w4(32'hbba100f3),
	.w5(32'hbc0497e4),
	.w6(32'h3c48afa3),
	.w7(32'h38c7d4dd),
	.w8(32'h3a16f10b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71abf9),
	.w1(32'hbc2643b5),
	.w2(32'hbbbfe00b),
	.w3(32'hbaeab6c2),
	.w4(32'hbc6e52b0),
	.w5(32'hbbbcfa5c),
	.w6(32'h3cdfc383),
	.w7(32'hb9102563),
	.w8(32'hbc0ba769),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78244e),
	.w1(32'hbc512b6d),
	.w2(32'h3b8c3302),
	.w3(32'hbbe9ddb6),
	.w4(32'hbae165d1),
	.w5(32'hbcac44c7),
	.w6(32'hbcc647bb),
	.w7(32'h3b75938d),
	.w8(32'h3ab645ea),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc874471),
	.w1(32'hbc41c77b),
	.w2(32'hbbe08a26),
	.w3(32'h3be25503),
	.w4(32'hbb81689e),
	.w5(32'hbba582c0),
	.w6(32'h3b0fd2f4),
	.w7(32'h3d6728dd),
	.w8(32'hbb94bc63),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c400bdd),
	.w1(32'hbc0fba6d),
	.w2(32'hba36a916),
	.w3(32'h3c68cced),
	.w4(32'hbb6ce59b),
	.w5(32'h3ac5f8a5),
	.w6(32'hbb512570),
	.w7(32'hbb9d1635),
	.w8(32'hbaaaf6a5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf732cf),
	.w1(32'hbb72f6eb),
	.w2(32'h3af810fd),
	.w3(32'hbae01682),
	.w4(32'hbc2b1849),
	.w5(32'h3c2e5a54),
	.w6(32'h3ac58e40),
	.w7(32'h3c86ab36),
	.w8(32'hbb9ffc53),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85e52f),
	.w1(32'h3c0cef20),
	.w2(32'h3abe319c),
	.w3(32'hbb18cde9),
	.w4(32'h3a399df2),
	.w5(32'h3ba29267),
	.w6(32'h3bfe7de8),
	.w7(32'h3bf9731c),
	.w8(32'h3b5e1348),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01e1b5),
	.w1(32'h3b22dcf3),
	.w2(32'h3c5f98af),
	.w3(32'h3b15a0ee),
	.w4(32'h3ba96183),
	.w5(32'h3c07a4d0),
	.w6(32'hb9b1b350),
	.w7(32'h3c05d863),
	.w8(32'h3ba0932d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef3840),
	.w1(32'hbc851ca0),
	.w2(32'hbb5bff52),
	.w3(32'hbbd31986),
	.w4(32'hbae84ac7),
	.w5(32'h3b84b58b),
	.w6(32'h3c12ca16),
	.w7(32'hbc4eed93),
	.w8(32'hbbaaf5ae),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6ff69),
	.w1(32'hbc830607),
	.w2(32'hbc6206f2),
	.w3(32'hbc8b1b9c),
	.w4(32'h3be1d007),
	.w5(32'h3d1c8762),
	.w6(32'h3c1b1a54),
	.w7(32'hbb823278),
	.w8(32'hbc3fe8e4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2f020),
	.w1(32'hbbb19c27),
	.w2(32'hbc50ac70),
	.w3(32'hbc78169f),
	.w4(32'hbc778e37),
	.w5(32'hbce533c7),
	.w6(32'hbd12a2cc),
	.w7(32'hbd3fc93a),
	.w8(32'hbc1de1e0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021d2a),
	.w1(32'h3c1acfb0),
	.w2(32'h3c67bacb),
	.w3(32'h3ba5464d),
	.w4(32'hbb624876),
	.w5(32'hbac32115),
	.w6(32'h3b1d2db4),
	.w7(32'h3b91e6ab),
	.w8(32'hbcdbfb1b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ac491),
	.w1(32'h3b6b2adc),
	.w2(32'h3c016d96),
	.w3(32'hbc8ea40e),
	.w4(32'hbb80502f),
	.w5(32'h3c16bfd3),
	.w6(32'hbb63c16c),
	.w7(32'h3ca2453e),
	.w8(32'h3be390ea),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb052a13),
	.w1(32'h3c717382),
	.w2(32'h3c36c75d),
	.w3(32'h3bc95f97),
	.w4(32'h3c51a753),
	.w5(32'hbbcb3599),
	.w6(32'h391989b7),
	.w7(32'h3c480e2c),
	.w8(32'h3adbd616),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15bd09),
	.w1(32'hbc42aeda),
	.w2(32'h3ac4dc03),
	.w3(32'hbc29de2b),
	.w4(32'hbc8345da),
	.w5(32'h3b541d71),
	.w6(32'hb9d610c7),
	.w7(32'hba033a51),
	.w8(32'hbbf99776),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0843ac),
	.w1(32'h3b878b5f),
	.w2(32'h3c9f923a),
	.w3(32'h3c10439b),
	.w4(32'hbb050223),
	.w5(32'h3c9661a7),
	.w6(32'hbc4b4da3),
	.w7(32'hbbcbb4cf),
	.w8(32'h3b16b16e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd867eb),
	.w1(32'hbb101267),
	.w2(32'h3ca450b8),
	.w3(32'h3b638687),
	.w4(32'h3b7a1d49),
	.w5(32'h3c21d1e5),
	.w6(32'hbb1d0347),
	.w7(32'hb9e3a13a),
	.w8(32'h3c769ddf),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fb85d),
	.w1(32'hb9f15418),
	.w2(32'h3c3bc1a6),
	.w3(32'hbbf6c234),
	.w4(32'hbc2b3720),
	.w5(32'hbc0769f1),
	.w6(32'hbb1901f8),
	.w7(32'hbc0e8353),
	.w8(32'h3791bb46),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae76682),
	.w1(32'h3c2967d9),
	.w2(32'h3c915cf1),
	.w3(32'h3aba34eb),
	.w4(32'hbbce8d32),
	.w5(32'hba9f2e27),
	.w6(32'hbc2f3f20),
	.w7(32'h3c8ce690),
	.w8(32'hbc69ff39),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfab5cf),
	.w1(32'hbb8e09c6),
	.w2(32'h3bc0afeb),
	.w3(32'h3c881a20),
	.w4(32'hbae7011c),
	.w5(32'h3c07daf2),
	.w6(32'h3bea9c80),
	.w7(32'h3b9c0feb),
	.w8(32'hba476d4c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ca953),
	.w1(32'hbc221a4e),
	.w2(32'hbcb18e12),
	.w3(32'hbd05b0a1),
	.w4(32'hbc726d26),
	.w5(32'hbc1ae2db),
	.w6(32'hbcb1a3a7),
	.w7(32'h3a8a5399),
	.w8(32'hbbeeb74d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a515246),
	.w1(32'hbc0f2cc7),
	.w2(32'h3b88d9d1),
	.w3(32'h3cb4907a),
	.w4(32'h3c13c00c),
	.w5(32'h3c519334),
	.w6(32'h3d0b9d7a),
	.w7(32'hb91492d5),
	.w8(32'h3bdb12ec),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc025b83),
	.w1(32'h3c7b7e8d),
	.w2(32'h3ca7da64),
	.w3(32'h3c69face),
	.w4(32'h3c8157c8),
	.w5(32'h3ca09128),
	.w6(32'h3c67dcb0),
	.w7(32'h3b9849cc),
	.w8(32'h3c523e27),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd153dd),
	.w1(32'hbbaf5659),
	.w2(32'h3bda2e8c),
	.w3(32'hbc184083),
	.w4(32'hbbcc2803),
	.w5(32'hbd0023a4),
	.w6(32'hbc10c380),
	.w7(32'hbbb4c745),
	.w8(32'hbc48c56c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f1085),
	.w1(32'h390a00a9),
	.w2(32'hbc58e1cc),
	.w3(32'hba42453e),
	.w4(32'hbaef7b85),
	.w5(32'hb9389d68),
	.w6(32'hba987358),
	.w7(32'h3c69fc5c),
	.w8(32'h3c3c6e1d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc318ba),
	.w1(32'hbc8b3846),
	.w2(32'hbcafe900),
	.w3(32'hbd1d0d46),
	.w4(32'hbcca749d),
	.w5(32'hbb4541ef),
	.w6(32'hbcf918b7),
	.w7(32'hbcb54785),
	.w8(32'hbca176af),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5963ee),
	.w1(32'hbbc83335),
	.w2(32'hba3a24a5),
	.w3(32'h3c9b3cd5),
	.w4(32'h3bfd56be),
	.w5(32'hbc382a9c),
	.w6(32'h3b7c804d),
	.w7(32'h3bc2654c),
	.w8(32'h3aa29ddc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba78c4b),
	.w1(32'hbc448ab0),
	.w2(32'hbc289e03),
	.w3(32'h3c0aa74b),
	.w4(32'h3abd7a18),
	.w5(32'hbbd266d7),
	.w6(32'hbbd1f814),
	.w7(32'hba29dd70),
	.w8(32'h3b3f6bfe),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985533b),
	.w1(32'hbb2a10da),
	.w2(32'h3bf2bcce),
	.w3(32'hbba5986b),
	.w4(32'hba25989b),
	.w5(32'hbbca22df),
	.w6(32'hbaf7b3ae),
	.w7(32'h3acdce1e),
	.w8(32'h3cab55b1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30dc9b),
	.w1(32'h3b492fda),
	.w2(32'h3be815f1),
	.w3(32'h3bc174ee),
	.w4(32'h3c3bf3e6),
	.w5(32'h3c913b80),
	.w6(32'h3c646b4c),
	.w7(32'hba91a6d4),
	.w8(32'hbc4ed176),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec4326),
	.w1(32'h3bbb2795),
	.w2(32'hbb76b168),
	.w3(32'h3c673cb8),
	.w4(32'h3c14aea0),
	.w5(32'h3ba09661),
	.w6(32'h3bc34451),
	.w7(32'h3be7a1f1),
	.w8(32'h3be096da),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c8337),
	.w1(32'hbc2947b0),
	.w2(32'hbb4f1f3f),
	.w3(32'h3c93f7d7),
	.w4(32'h3d069e80),
	.w5(32'hbbb48e39),
	.w6(32'h3ab61d81),
	.w7(32'hbae9cb76),
	.w8(32'hbbfb8185),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2bbf7),
	.w1(32'h3c05a377),
	.w2(32'h3c586860),
	.w3(32'h3b4ad775),
	.w4(32'hbadc2903),
	.w5(32'h3b2c1e9f),
	.w6(32'hbb8368af),
	.w7(32'h3b226b21),
	.w8(32'hba31fc92),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aa434),
	.w1(32'h3c3c82fa),
	.w2(32'hbb435b2a),
	.w3(32'h3b5142d0),
	.w4(32'hbc9e2470),
	.w5(32'hbce5fc99),
	.w6(32'hbc902a03),
	.w7(32'hbb4a45c7),
	.w8(32'h3a9de570),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ee5b7),
	.w1(32'h3b4e7f19),
	.w2(32'hbc5bfe32),
	.w3(32'h3b0665d0),
	.w4(32'hbc06138e),
	.w5(32'h3aa0ac70),
	.w6(32'hbbc73ea6),
	.w7(32'hbb2be042),
	.w8(32'hb887871a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24321c),
	.w1(32'hbc0f9c3b),
	.w2(32'hba40b2b8),
	.w3(32'hbd007940),
	.w4(32'hba13b6c6),
	.w5(32'h3c050f26),
	.w6(32'h3c79a368),
	.w7(32'h3c98011e),
	.w8(32'h3c051b5c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba32559),
	.w1(32'hbb437908),
	.w2(32'h3c8a1ad6),
	.w3(32'h3a43648f),
	.w4(32'hbc31e1a5),
	.w5(32'h3afc2849),
	.w6(32'hbab924a3),
	.w7(32'hbc1c64c1),
	.w8(32'h3b53a9f1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2bdfe),
	.w1(32'hbc942fc1),
	.w2(32'hba6fbb4c),
	.w3(32'h3a831e75),
	.w4(32'h3bd7e704),
	.w5(32'h38985ed5),
	.w6(32'h3c064857),
	.w7(32'h3d1ec565),
	.w8(32'hbc0a9b52),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c703c84),
	.w1(32'hbba9c485),
	.w2(32'hbc992297),
	.w3(32'h3b4a075e),
	.w4(32'hbae37e5e),
	.w5(32'h3c8046bf),
	.w6(32'hbbaf82a2),
	.w7(32'hbb08b1e2),
	.w8(32'h3ace95f4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8651d4),
	.w1(32'h3ba3db31),
	.w2(32'h3bf79f25),
	.w3(32'h3a2d1276),
	.w4(32'hbb1191d3),
	.w5(32'hbbdf1d44),
	.w6(32'hbb2ba60a),
	.w7(32'h39feb932),
	.w8(32'hbc408047),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f0145),
	.w1(32'hbad71f66),
	.w2(32'h3922f23a),
	.w3(32'h3c19de40),
	.w4(32'h3beec0a5),
	.w5(32'h3adbef1a),
	.w6(32'h3af24b73),
	.w7(32'h3b09ece7),
	.w8(32'h3c1cff38),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0b052),
	.w1(32'h3d27045e),
	.w2(32'hbb1d4afe),
	.w3(32'h3b804152),
	.w4(32'hbb5dc57c),
	.w5(32'hbc0ad22a),
	.w6(32'hbb632ea1),
	.w7(32'h3b63e470),
	.w8(32'hbbcd9933),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfb8aa0),
	.w1(32'h3bc3efa3),
	.w2(32'h3bd01abb),
	.w3(32'h3b9a9726),
	.w4(32'hbb9f2434),
	.w5(32'hbbbb0dfe),
	.w6(32'hbbc02c5b),
	.w7(32'hbc042834),
	.w8(32'hbaac4141),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f9449),
	.w1(32'hbb1095e3),
	.w2(32'h3c4ce5ba),
	.w3(32'h3bceafc5),
	.w4(32'h3acb9e35),
	.w5(32'h3c2411c1),
	.w6(32'h3cda36ed),
	.w7(32'hbb92c9cf),
	.w8(32'h3bf0f9a6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba09a58),
	.w1(32'hbb261a67),
	.w2(32'hbbbc2d06),
	.w3(32'hba61950b),
	.w4(32'h3c999fff),
	.w5(32'h3acd2102),
	.w6(32'h3bb437e8),
	.w7(32'hbc65bffa),
	.w8(32'hbc0047b4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5759de),
	.w1(32'hbbdeac95),
	.w2(32'hbca3dca1),
	.w3(32'hbb480ff2),
	.w4(32'hbc8ba538),
	.w5(32'hba96d846),
	.w6(32'hbbaf40fb),
	.w7(32'h3ae708c1),
	.w8(32'h3cb9198b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b16ed),
	.w1(32'h39a61393),
	.w2(32'h3c435348),
	.w3(32'hbc6ab148),
	.w4(32'hbac8253f),
	.w5(32'hbb445baf),
	.w6(32'hbb80a9e6),
	.w7(32'hba807525),
	.w8(32'hb9c8a3a1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95df23),
	.w1(32'h3c39af73),
	.w2(32'hbb6a0964),
	.w3(32'hbb35774e),
	.w4(32'hb816172e),
	.w5(32'hbc367553),
	.w6(32'hbbe35b2c),
	.w7(32'h3b0057e4),
	.w8(32'hbb9021c2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44a4bb),
	.w1(32'h3b6813a5),
	.w2(32'hbc1c6802),
	.w3(32'h3af08bec),
	.w4(32'h3c80058f),
	.w5(32'h3b78f7a5),
	.w6(32'hbbbf54e0),
	.w7(32'h3c0c0b79),
	.w8(32'hbc4e26fa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86fab4),
	.w1(32'h3bd328e0),
	.w2(32'h3c076bb5),
	.w3(32'h3bb2da18),
	.w4(32'h3bb54ac1),
	.w5(32'h3c657155),
	.w6(32'h3b8ff13f),
	.w7(32'h3bdb35db),
	.w8(32'hbad48286),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3bc79),
	.w1(32'hbba27c60),
	.w2(32'hbbd18413),
	.w3(32'hbb4b4ddf),
	.w4(32'h3b77bc96),
	.w5(32'hbb34b786),
	.w6(32'h3b4223e7),
	.w7(32'hbbe03fb1),
	.w8(32'h3b58b992),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d5739),
	.w1(32'hbc3baa1e),
	.w2(32'hbba1e413),
	.w3(32'hbc25868b),
	.w4(32'h3b8977fc),
	.w5(32'hbbd2d333),
	.w6(32'hbad9bbd5),
	.w7(32'h39cc6036),
	.w8(32'hbc28de50),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64a905),
	.w1(32'hb9c05c34),
	.w2(32'hbbc87851),
	.w3(32'h39b2b771),
	.w4(32'hbbcf140e),
	.w5(32'h3b2605a2),
	.w6(32'h3c6f5d60),
	.w7(32'hba84cdf2),
	.w8(32'h3c9bf132),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17676f),
	.w1(32'h3bd85d85),
	.w2(32'hbc4bae29),
	.w3(32'hbbff00ff),
	.w4(32'h3c3ad96e),
	.w5(32'h3b5feb2f),
	.w6(32'hbc5bd5ec),
	.w7(32'hbb4760f0),
	.w8(32'h3aacb06e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66387e),
	.w1(32'hbbbd4acb),
	.w2(32'h3c020557),
	.w3(32'hbc388e38),
	.w4(32'h3b1ab707),
	.w5(32'hbc8d251a),
	.w6(32'h39bb7656),
	.w7(32'h3b7a7031),
	.w8(32'hbb8c3745),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c8cac),
	.w1(32'hbbfb61b5),
	.w2(32'hbb6e100b),
	.w3(32'hbc9d6282),
	.w4(32'hbc8472fd),
	.w5(32'hbc4e0877),
	.w6(32'hbbc6b222),
	.w7(32'hbc97dd23),
	.w8(32'hbc5cc661),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d67f9),
	.w1(32'h3b9c31de),
	.w2(32'h3c039548),
	.w3(32'h3b33958c),
	.w4(32'hbbe40c4c),
	.w5(32'h3c0d4912),
	.w6(32'h3a4744fc),
	.w7(32'hbb9b8742),
	.w8(32'hba81351e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2ab8b),
	.w1(32'h3bb81646),
	.w2(32'hbc0b6ce5),
	.w3(32'h3b3cfd67),
	.w4(32'h3bc9f26d),
	.w5(32'h3a8ba2c7),
	.w6(32'hb9988d7a),
	.w7(32'h3ba00111),
	.w8(32'h3ce01576),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce0448),
	.w1(32'hbc3530fe),
	.w2(32'hbc801a42),
	.w3(32'hbb9400d1),
	.w4(32'hbc949426),
	.w5(32'hbc518817),
	.w6(32'hbc8e971e),
	.w7(32'hbcf6e636),
	.w8(32'hbc6cacf1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d5e44),
	.w1(32'h3afb8a09),
	.w2(32'h3be152b7),
	.w3(32'hba9917a3),
	.w4(32'h3b3bf9fb),
	.w5(32'h3b173f20),
	.w6(32'hbb23c13a),
	.w7(32'hb9831abe),
	.w8(32'hbc16220e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015dcc),
	.w1(32'h3ac95036),
	.w2(32'hbb3c8169),
	.w3(32'hbbfabbf7),
	.w4(32'h3b8b537b),
	.w5(32'hbba872ca),
	.w6(32'h3b4c946e),
	.w7(32'hbce4ebf6),
	.w8(32'hbad21a4f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58f596),
	.w1(32'h3c77b11c),
	.w2(32'h3c1011c4),
	.w3(32'h3a08e4ad),
	.w4(32'h3b8eebc8),
	.w5(32'h3c01b9c8),
	.w6(32'hbabf5310),
	.w7(32'h3c7bbb72),
	.w8(32'hbc1953f2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3360ba),
	.w1(32'h3aca7ea1),
	.w2(32'h3c024cf5),
	.w3(32'h3bce44a6),
	.w4(32'hbca650a8),
	.w5(32'h3c700978),
	.w6(32'h3bea17a5),
	.w7(32'h3c659217),
	.w8(32'h3b86dc4b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d12f2),
	.w1(32'hbb7fc890),
	.w2(32'hbb5cd47f),
	.w3(32'h3b891472),
	.w4(32'hbc00cc49),
	.w5(32'hbb85879d),
	.w6(32'hbb4b4cb9),
	.w7(32'h3b5f307b),
	.w8(32'hbc0518aa),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92e79e),
	.w1(32'h3c245d66),
	.w2(32'h3bdd0cbe),
	.w3(32'h3b94afb1),
	.w4(32'hbc02194e),
	.w5(32'h3c0d54b2),
	.w6(32'hbb1a8265),
	.w7(32'h3c7c6c7b),
	.w8(32'hbbacb54c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83bd18),
	.w1(32'h3bcde5b3),
	.w2(32'h3b1e9f35),
	.w3(32'hb9565786),
	.w4(32'h3bcf7932),
	.w5(32'hb9960b97),
	.w6(32'h3b17dd63),
	.w7(32'h3ba3c982),
	.w8(32'hbbdfa316),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd99b36),
	.w1(32'hbc6851ca),
	.w2(32'hbcdb0de0),
	.w3(32'hbbb66342),
	.w4(32'h3c6d57e2),
	.w5(32'hbbcd5f86),
	.w6(32'hbc0ad040),
	.w7(32'h3b363007),
	.w8(32'hbaabf035),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c468dc3),
	.w1(32'hbb980038),
	.w2(32'hbc8c92ca),
	.w3(32'h3a103f06),
	.w4(32'h3cb82bd4),
	.w5(32'h3b3c3e84),
	.w6(32'h3b837155),
	.w7(32'h3c9bd7c1),
	.w8(32'hbbeb7591),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900b2ab),
	.w1(32'h3bbaa5f4),
	.w2(32'h3aecdf0e),
	.w3(32'hbb0d7f58),
	.w4(32'h3bbe2d7c),
	.w5(32'h3c28ebf4),
	.w6(32'hb9823c29),
	.w7(32'hb92f4fac),
	.w8(32'hbacaaebf),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aece8c6),
	.w1(32'hbc4e6f99),
	.w2(32'h3b80ad73),
	.w3(32'hba92c37c),
	.w4(32'h3bd3eeb8),
	.w5(32'hbc3c3c69),
	.w6(32'hbb8aebb1),
	.w7(32'hbc20b288),
	.w8(32'hbc931eaf),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bc347),
	.w1(32'h3c0a00fd),
	.w2(32'h398e0118),
	.w3(32'h3ba5e323),
	.w4(32'hbc6691f2),
	.w5(32'h3c046054),
	.w6(32'hbb4fec84),
	.w7(32'hbb152837),
	.w8(32'h3c1cdaae),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f9505),
	.w1(32'h3c1ff1af),
	.w2(32'h3c2687fc),
	.w3(32'h3ccea9d2),
	.w4(32'hbbda61b4),
	.w5(32'h3cc50819),
	.w6(32'h3be3e33f),
	.w7(32'hbb77a03a),
	.w8(32'hba2d42c9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb362f04),
	.w1(32'h3a279e9d),
	.w2(32'hbb1c4c1b),
	.w3(32'hbb8ed7b8),
	.w4(32'h3c298c55),
	.w5(32'hbb99fa9d),
	.w6(32'hbbd54909),
	.w7(32'hbb5565cf),
	.w8(32'h3b0d1cd7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07cf1e),
	.w1(32'hbc0ab8d6),
	.w2(32'h3c0f5a8e),
	.w3(32'h3bd4da1c),
	.w4(32'h3bd28c36),
	.w5(32'hbb0c3bbb),
	.w6(32'h3c5ef0a8),
	.w7(32'hbb414e4f),
	.w8(32'h3c08831d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a9ec7),
	.w1(32'hbc004899),
	.w2(32'hbba07db3),
	.w3(32'hbc4bbb49),
	.w4(32'hbb25fd5a),
	.w5(32'hba1cc86c),
	.w6(32'h3b5ce564),
	.w7(32'hbaf73c67),
	.w8(32'hb94e8283),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45e7b2),
	.w1(32'hbbbf6544),
	.w2(32'hbbf7b7dd),
	.w3(32'h3c244285),
	.w4(32'h3be5b592),
	.w5(32'h3afca580),
	.w6(32'h3b3e817f),
	.w7(32'h3c3371b6),
	.w8(32'h3c8f7a38),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94a76b),
	.w1(32'hbaa61636),
	.w2(32'h3b1f5418),
	.w3(32'hbc5c1f3c),
	.w4(32'h3cae27ad),
	.w5(32'h3c113b26),
	.w6(32'h3b396e4b),
	.w7(32'h3be429c1),
	.w8(32'h3c2fd5cd),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc541631),
	.w1(32'h3b4b9dab),
	.w2(32'hbb1760ad),
	.w3(32'hbbac9af5),
	.w4(32'h3b9d2466),
	.w5(32'h3b298c59),
	.w6(32'h3c7af058),
	.w7(32'hbbd2f4ef),
	.w8(32'hbb86a6fc),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b0f37),
	.w1(32'h3ab3d93d),
	.w2(32'hb99a44d2),
	.w3(32'hba975a0e),
	.w4(32'h3c57068c),
	.w5(32'h3b78081b),
	.w6(32'h3c3bfc98),
	.w7(32'hbb5b883e),
	.w8(32'h3a94f4a7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96ce89),
	.w1(32'hbc139ff9),
	.w2(32'hbaca97ba),
	.w3(32'hbc1f6cfc),
	.w4(32'h3b26a4a4),
	.w5(32'hbae082bb),
	.w6(32'hbbcb2bdf),
	.w7(32'hbbac5793),
	.w8(32'h3bfe662e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43647f),
	.w1(32'h3a9c3ecd),
	.w2(32'h3a33b688),
	.w3(32'hbb5b7ead),
	.w4(32'hbae6f136),
	.w5(32'hbc7355e5),
	.w6(32'h3c1bfffd),
	.w7(32'h3b89c6dc),
	.w8(32'hbb02eddb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c116224),
	.w1(32'h3a421f72),
	.w2(32'h3c63a993),
	.w3(32'hbc44fd5a),
	.w4(32'h392fa740),
	.w5(32'h3c8cff29),
	.w6(32'hbaaafb5a),
	.w7(32'hbbc59f95),
	.w8(32'h3a235efe),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2eaf3),
	.w1(32'h3b4919dc),
	.w2(32'hbbf4c9c5),
	.w3(32'h3b27e61a),
	.w4(32'hbb9928bf),
	.w5(32'hbc54d5ae),
	.w6(32'h3bad4212),
	.w7(32'hbb2e7f5c),
	.w8(32'h3a3b5250),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd22da8),
	.w1(32'h3b776e5e),
	.w2(32'hb9834ce3),
	.w3(32'hbbdf85c2),
	.w4(32'h3b3b4011),
	.w5(32'h38feb6cc),
	.w6(32'h3c1f6446),
	.w7(32'h3ba1f0f3),
	.w8(32'hbb383184),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64eb7a),
	.w1(32'h3bb0acbc),
	.w2(32'h3aea8d44),
	.w3(32'hbb8596b3),
	.w4(32'hbc047160),
	.w5(32'h3a6513ce),
	.w6(32'h3b18733b),
	.w7(32'hbd05a9dd),
	.w8(32'hbb46aa24),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f99b92),
	.w1(32'hba5e3591),
	.w2(32'h3b0c084e),
	.w3(32'hbada299c),
	.w4(32'h3b9185e7),
	.w5(32'hbc3ce095),
	.w6(32'h3bb263ff),
	.w7(32'hbb0d373f),
	.w8(32'hbc22c313),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5a159),
	.w1(32'h39d86a14),
	.w2(32'hbc8eaeb5),
	.w3(32'hba76d516),
	.w4(32'hbb3c082c),
	.w5(32'h3c4dca52),
	.w6(32'hbc573cb2),
	.w7(32'h3ac74e91),
	.w8(32'h3b71006f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb4ea6),
	.w1(32'h3b9db09e),
	.w2(32'hbc0d67b9),
	.w3(32'hba9f7ce0),
	.w4(32'hbbb08c88),
	.w5(32'hbbd80cb4),
	.w6(32'hbbaafccc),
	.w7(32'h3c388015),
	.w8(32'hbba2ea7a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc798ae0),
	.w1(32'hbc2dc085),
	.w2(32'hbaaa05f3),
	.w3(32'hbc473366),
	.w4(32'hbc087b5b),
	.w5(32'h3c202d00),
	.w6(32'h3a3bb385),
	.w7(32'h3b7daaf3),
	.w8(32'hbbd174e6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ca650),
	.w1(32'hb9faa426),
	.w2(32'h3bf07ed2),
	.w3(32'h3af1debc),
	.w4(32'h3ab18355),
	.w5(32'h3aa0c0d7),
	.w6(32'hbc4babbe),
	.w7(32'hbbafd6e1),
	.w8(32'hbd100012),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eaf06),
	.w1(32'hbc071856),
	.w2(32'h3bdf0bb8),
	.w3(32'h3bb1d545),
	.w4(32'h3bf878f9),
	.w5(32'hbadf0dc2),
	.w6(32'hbb276a63),
	.w7(32'h3b740ed3),
	.w8(32'hbc81523a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9238423),
	.w1(32'hbc11f007),
	.w2(32'h3bf5652f),
	.w3(32'h3c66db0a),
	.w4(32'hbc723a45),
	.w5(32'h3b0dadad),
	.w6(32'h3c3e2f88),
	.w7(32'h3bccb058),
	.w8(32'h3bdc670a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e106e),
	.w1(32'hbc547052),
	.w2(32'hbc19cc48),
	.w3(32'hbc406e0e),
	.w4(32'hbc4b6f6b),
	.w5(32'hbc19aac2),
	.w6(32'h3c3c3e58),
	.w7(32'hbbf27921),
	.w8(32'hbc636c37),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf566aa),
	.w1(32'hbc064c58),
	.w2(32'hbc0d8acd),
	.w3(32'h3b5099df),
	.w4(32'h3ca746aa),
	.w5(32'hbc576942),
	.w6(32'h3bfaf27f),
	.w7(32'h3c46e67a),
	.w8(32'hbc14c9c7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a5321),
	.w1(32'hbaeb33e1),
	.w2(32'h3c43cc8e),
	.w3(32'hbb17baf3),
	.w4(32'hbbb54022),
	.w5(32'h3cc57395),
	.w6(32'h3b3dab6a),
	.w7(32'hbbd68fb2),
	.w8(32'hbbb84e81),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71163c),
	.w1(32'h3b1c88d2),
	.w2(32'h3c067437),
	.w3(32'h3c8a0ba6),
	.w4(32'h3c11b1ae),
	.w5(32'h3aff35e5),
	.w6(32'hbb4e756e),
	.w7(32'h3b8308e4),
	.w8(32'hbaf6a9f4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81a7f3),
	.w1(32'hbb5c3553),
	.w2(32'h3c398a13),
	.w3(32'hbac9a01c),
	.w4(32'h39bec7ec),
	.w5(32'h3b32113b),
	.w6(32'h3aee8f35),
	.w7(32'h3984824c),
	.w8(32'h3c21e9e5),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba91c42),
	.w1(32'hbba0c803),
	.w2(32'h3c68f0dc),
	.w3(32'h3a4980ba),
	.w4(32'h3c663c3e),
	.w5(32'hbc5ff92f),
	.w6(32'hbad6dd4a),
	.w7(32'hbbf6985a),
	.w8(32'hbc0bc517),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dbfb2),
	.w1(32'h3c2d2f4b),
	.w2(32'h3c0845b4),
	.w3(32'hbb64a159),
	.w4(32'hbb486b50),
	.w5(32'hbce23e33),
	.w6(32'hba8a5634),
	.w7(32'hbc1169f5),
	.w8(32'hbb49c0bd),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012b4f),
	.w1(32'h3c127158),
	.w2(32'hbb820c03),
	.w3(32'h3c11180b),
	.w4(32'h3aef6625),
	.w5(32'hbbd6eb8f),
	.w6(32'hbbf92556),
	.w7(32'h3c49c8fd),
	.w8(32'hbbea5644),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25b0c9),
	.w1(32'hbbfbaa5c),
	.w2(32'h39ba28b7),
	.w3(32'h3cba3c86),
	.w4(32'h3c50c107),
	.w5(32'hbc9283b1),
	.w6(32'hbaa93a8f),
	.w7(32'hb880472d),
	.w8(32'h3a404932),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc161e39),
	.w1(32'h3c21e875),
	.w2(32'hb88830da),
	.w3(32'hbba18a02),
	.w4(32'hb9db23bc),
	.w5(32'hbbb29a07),
	.w6(32'hb82d92c2),
	.w7(32'hbba6ed7a),
	.w8(32'h3bae3d48),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26a443),
	.w1(32'h3a017027),
	.w2(32'hbb99a87b),
	.w3(32'h3aaa38bc),
	.w4(32'h3bd886ef),
	.w5(32'hbbc9b99f),
	.w6(32'hbbaca3c7),
	.w7(32'h39502a8f),
	.w8(32'hbbe64e10),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83616a),
	.w1(32'h3a2909be),
	.w2(32'hbb25f03a),
	.w3(32'hbc0b2383),
	.w4(32'h3a0f11ff),
	.w5(32'hbba65d7f),
	.w6(32'h38e65ae3),
	.w7(32'h3c9834c5),
	.w8(32'hbb80feac),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6f483),
	.w1(32'hbb86aaf8),
	.w2(32'h3acae596),
	.w3(32'h3b0c36a6),
	.w4(32'hb988d1a8),
	.w5(32'h391b3468),
	.w6(32'hbc702b6d),
	.w7(32'hbbedf737),
	.w8(32'h3c9f7172),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93afcf),
	.w1(32'hba5c0dcf),
	.w2(32'hbc1f49fd),
	.w3(32'h3b6f1663),
	.w4(32'hbc2b3cc6),
	.w5(32'hbaeddf80),
	.w6(32'hbb6498bf),
	.w7(32'h3a0f78da),
	.w8(32'hbcaef78c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b949358),
	.w1(32'h3a30538e),
	.w2(32'h3c89f736),
	.w3(32'h3b7975a6),
	.w4(32'hbc08eaec),
	.w5(32'hbb653586),
	.w6(32'h3bcb638a),
	.w7(32'h39950987),
	.w8(32'h3c218b9d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4848f5),
	.w1(32'h3b42553a),
	.w2(32'h3c18c56e),
	.w3(32'hbb7b0b21),
	.w4(32'h3c215981),
	.w5(32'hbc207c06),
	.w6(32'hbbcee299),
	.w7(32'hbc2a730c),
	.w8(32'h3bf35b51),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51befa),
	.w1(32'hbc0441ba),
	.w2(32'hbbb8bb29),
	.w3(32'hbb630c7e),
	.w4(32'h3b87e93e),
	.w5(32'h3cb1b8a7),
	.w6(32'hbb00735b),
	.w7(32'h3b9c2164),
	.w8(32'h3a4310f5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f6d6a),
	.w1(32'h3c9a02a6),
	.w2(32'h3c1b55f0),
	.w3(32'h3c5c7a77),
	.w4(32'h3c8b15ae),
	.w5(32'hbb805b39),
	.w6(32'hbb4eb23f),
	.w7(32'h3c22025d),
	.w8(32'hbb8fa791),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b763881),
	.w1(32'hbbb5ac42),
	.w2(32'h3964fe98),
	.w3(32'h3c706cec),
	.w4(32'hbcffc3a7),
	.w5(32'hbc82800a),
	.w6(32'h3bf28968),
	.w7(32'hbbbb25f1),
	.w8(32'h3c8c50d1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd5faf),
	.w1(32'hbc624add),
	.w2(32'hbb8c7f68),
	.w3(32'hbbdf1b6e),
	.w4(32'hbc107709),
	.w5(32'hbb95b51b),
	.w6(32'h3b902afc),
	.w7(32'h3c59b62a),
	.w8(32'hba7f4206),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa123a),
	.w1(32'h39fb590b),
	.w2(32'hbc2e942e),
	.w3(32'h3bc27bce),
	.w4(32'hbc26eb8f),
	.w5(32'h3c799f5e),
	.w6(32'hbab6f287),
	.w7(32'hbc0e8181),
	.w8(32'h3b3e314f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d965b0),
	.w1(32'hba96db04),
	.w2(32'hbbe217a5),
	.w3(32'hbc0afe06),
	.w4(32'h3bb4d08a),
	.w5(32'hbb30925d),
	.w6(32'h39a06807),
	.w7(32'hbb773ea2),
	.w8(32'h3b3ad5d9),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1e630),
	.w1(32'h3c101f4f),
	.w2(32'hbb29a8bd),
	.w3(32'hba15dc9a),
	.w4(32'h3ba7f1b3),
	.w5(32'hba56c7b0),
	.w6(32'h3c1840bb),
	.w7(32'h3c8671fe),
	.w8(32'hbc63314b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25b653),
	.w1(32'hbb166749),
	.w2(32'hb9614bef),
	.w3(32'hbc576b1f),
	.w4(32'hbb15c2fd),
	.w5(32'hbc08b68f),
	.w6(32'hbc01ebe9),
	.w7(32'h3a198153),
	.w8(32'h3b5ac448),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb618ed),
	.w1(32'h3b72a127),
	.w2(32'h3c4d1bff),
	.w3(32'hbcbb1938),
	.w4(32'h3be917d2),
	.w5(32'h3c17c72b),
	.w6(32'hbaa818af),
	.w7(32'h3bea237f),
	.w8(32'h3caae7f3),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a8f99),
	.w1(32'hbb51bdf9),
	.w2(32'hbbc9f82e),
	.w3(32'h3a17e499),
	.w4(32'h3c4478a3),
	.w5(32'hbc989890),
	.w6(32'hbb7aad31),
	.w7(32'h3bdfb0c1),
	.w8(32'hba4195ae),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc156dea),
	.w1(32'hbbbead43),
	.w2(32'h3cd67d8b),
	.w3(32'h3b87d9dd),
	.w4(32'h3bae28f9),
	.w5(32'hbc30d421),
	.w6(32'h3a9a76b8),
	.w7(32'hbc4641a0),
	.w8(32'hbcbca615),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddf1d3),
	.w1(32'h3c79d893),
	.w2(32'hbc8cc5f2),
	.w3(32'hbb808ae5),
	.w4(32'h3b8e9148),
	.w5(32'hbc2054bb),
	.w6(32'h3a826c89),
	.w7(32'h3bd9cd6e),
	.w8(32'hbb7f1c07),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c518ead),
	.w1(32'h3b3aaedd),
	.w2(32'hbc3b912a),
	.w3(32'hbc70b0c6),
	.w4(32'hbd537955),
	.w5(32'h3b9eb6c7),
	.w6(32'h3bccaae8),
	.w7(32'hbc562b48),
	.w8(32'h3cdea6a3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c3ce7),
	.w1(32'hbbcd5f36),
	.w2(32'hbc01a7c0),
	.w3(32'hbb8cba3e),
	.w4(32'h3b991236),
	.w5(32'hbc4f7408),
	.w6(32'h3c6da1e9),
	.w7(32'h398d41b4),
	.w8(32'hbc922aa7),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98364e),
	.w1(32'h3c7551a8),
	.w2(32'hbc4f2cda),
	.w3(32'hbc26a292),
	.w4(32'hbbc4ba53),
	.w5(32'hbad36dcd),
	.w6(32'hbbcd01e8),
	.w7(32'hbc3482d9),
	.w8(32'h3cb006c0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce59458),
	.w1(32'h3b89be27),
	.w2(32'hbaac9ce0),
	.w3(32'hbb828543),
	.w4(32'h3c673ddd),
	.w5(32'hbbdfc82f),
	.w6(32'hbad585d5),
	.w7(32'hbb86e0b6),
	.w8(32'h3bae303a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb982e),
	.w1(32'h3c38f0f3),
	.w2(32'h3c24ffde),
	.w3(32'h3b713e7c),
	.w4(32'hbb9ecf92),
	.w5(32'hbc1d0b7d),
	.w6(32'hbc106b5f),
	.w7(32'hbb201130),
	.w8(32'h3c34959a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84f26f),
	.w1(32'h3c167a91),
	.w2(32'hba2346cf),
	.w3(32'h3beb0737),
	.w4(32'h3bc68762),
	.w5(32'hbc4ada57),
	.w6(32'hbc28219e),
	.w7(32'h3b9be9bf),
	.w8(32'h3bfd4898),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc122d05),
	.w1(32'hbc66bf67),
	.w2(32'hbbe17d34),
	.w3(32'hbb4c7580),
	.w4(32'h3b706f19),
	.w5(32'hbbdc8f0e),
	.w6(32'h3bdb1a9e),
	.w7(32'hbc0879cb),
	.w8(32'h3c3a570a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39826cb5),
	.w1(32'h3c54a020),
	.w2(32'h3ce14439),
	.w3(32'hbc89d9c0),
	.w4(32'h3d05a7ee),
	.w5(32'h3c04fae3),
	.w6(32'h3c07e6a0),
	.w7(32'h3b4e556a),
	.w8(32'h3bdf4cba),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c896e38),
	.w1(32'h3c8b46ec),
	.w2(32'hbbb91a96),
	.w3(32'hb90d6825),
	.w4(32'h3a17584c),
	.w5(32'h3b5bbcf8),
	.w6(32'hbcbb3ed3),
	.w7(32'hbc5d4c33),
	.w8(32'h3b757ddd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5900f8),
	.w1(32'h3c969463),
	.w2(32'h3c41d023),
	.w3(32'h3ba37a7f),
	.w4(32'h3c90f6b1),
	.w5(32'h3c899852),
	.w6(32'h3c2b69db),
	.w7(32'hbbefbf0c),
	.w8(32'h3a94c34f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeb843),
	.w1(32'h3be07654),
	.w2(32'hbc62193a),
	.w3(32'hbc88e223),
	.w4(32'hbb9bb743),
	.w5(32'hbc84e768),
	.w6(32'h3b8aad5c),
	.w7(32'hbaaf1951),
	.w8(32'h3b36437c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a46bf1),
	.w1(32'hbbfe51c0),
	.w2(32'h391b156f),
	.w3(32'h3b9f26f3),
	.w4(32'hbc2aae41),
	.w5(32'h392ca403),
	.w6(32'h3ba0bdf5),
	.w7(32'hbbcf19b5),
	.w8(32'hbb06d811),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd88de1),
	.w1(32'h3b5d163d),
	.w2(32'hbcbb6a7a),
	.w3(32'h3cc7aa48),
	.w4(32'hbc3b9ead),
	.w5(32'hbcbae112),
	.w6(32'hbbfcad06),
	.w7(32'hbbfbc9d8),
	.w8(32'h3cac066d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc410df4),
	.w1(32'h3c18b579),
	.w2(32'h3c28f712),
	.w3(32'hbc3a2f4a),
	.w4(32'h3bffde40),
	.w5(32'hbaab7db9),
	.w6(32'hbbfd4e8e),
	.w7(32'hbac7a5af),
	.w8(32'hbbd79fae),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6241a6),
	.w1(32'h3c683eff),
	.w2(32'h3ce08225),
	.w3(32'hbb6032a0),
	.w4(32'h3bec8113),
	.w5(32'hbc2c3dd4),
	.w6(32'hbb9f34d9),
	.w7(32'h3b96b3b8),
	.w8(32'h3c5cd5ab),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaac0db),
	.w1(32'hbc9d92be),
	.w2(32'hbc5cef02),
	.w3(32'hbbff56fa),
	.w4(32'hbb5e031c),
	.w5(32'h3c9909af),
	.w6(32'h37ee182e),
	.w7(32'hbbca6207),
	.w8(32'hbbe50fb1),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb92d5),
	.w1(32'hbc37cf23),
	.w2(32'h3b24d7da),
	.w3(32'hbc91166c),
	.w4(32'hb9262c33),
	.w5(32'hbbab5a97),
	.w6(32'hbc152125),
	.w7(32'h39307375),
	.w8(32'h3c18726c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9df3d7),
	.w1(32'h3b0195b1),
	.w2(32'hbb50cc23),
	.w3(32'h3b8b3cbb),
	.w4(32'hbb5da1a2),
	.w5(32'hba1c5c3a),
	.w6(32'hbbd27e05),
	.w7(32'hbb61cb32),
	.w8(32'h3c22ba06),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb497b6b),
	.w1(32'h3b93fff3),
	.w2(32'h3b255e3b),
	.w3(32'h3c05c96c),
	.w4(32'h3b6f24bc),
	.w5(32'hbc4b6720),
	.w6(32'h3bdb4c1f),
	.w7(32'hbc4b51fb),
	.w8(32'h3af9b745),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca54ae6),
	.w1(32'hbae01546),
	.w2(32'hbc815d81),
	.w3(32'hbc730a56),
	.w4(32'hbc431c15),
	.w5(32'h3c809a0a),
	.w6(32'hbc1be52c),
	.w7(32'hbcbf872c),
	.w8(32'hbc939e88),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb225df4),
	.w1(32'hbc1fdc1c),
	.w2(32'hbbc1bfbd),
	.w3(32'hbc276913),
	.w4(32'h3bd41c9b),
	.w5(32'hb94f602f),
	.w6(32'hbc979d5f),
	.w7(32'hbb6385bb),
	.w8(32'h3c42f236),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3f1f8),
	.w1(32'h3be1bcff),
	.w2(32'h3b935ca4),
	.w3(32'hbaf72288),
	.w4(32'h3c398ceb),
	.w5(32'hbc1da578),
	.w6(32'h3be3ebb6),
	.w7(32'hbb45fe0a),
	.w8(32'hbbba7e10),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c072de1),
	.w1(32'h3c801b73),
	.w2(32'h3c32f1ad),
	.w3(32'h3bc405f5),
	.w4(32'h3bfc8db2),
	.w5(32'h3c04f936),
	.w6(32'h3b800581),
	.w7(32'hb9b1ad04),
	.w8(32'h3b3ecfad),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca9c0a6),
	.w1(32'hbbf73f2d),
	.w2(32'hbb90a13e),
	.w3(32'hbbc81b8a),
	.w4(32'h3bbcdb9e),
	.w5(32'hbb077c92),
	.w6(32'hbba6f534),
	.w7(32'hbc9d1d96),
	.w8(32'hbc474054),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72888f),
	.w1(32'h3b76b4c0),
	.w2(32'hbcb557de),
	.w3(32'hbcd43e4b),
	.w4(32'h3a828925),
	.w5(32'h3b7e4e3b),
	.w6(32'h3a80d913),
	.w7(32'hbbf06467),
	.w8(32'h3a205406),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f2a01),
	.w1(32'hbb96aa58),
	.w2(32'hbb1d437d),
	.w3(32'h3b8acfe8),
	.w4(32'hba85c963),
	.w5(32'h3bac21f4),
	.w6(32'hbb019f50),
	.w7(32'hbc8f05a6),
	.w8(32'hbc44d75a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae459c),
	.w1(32'h3c4116f1),
	.w2(32'hbaa2fed3),
	.w3(32'hbd0b4f8a),
	.w4(32'hbbe8c68c),
	.w5(32'hbc7ef764),
	.w6(32'hbc78a4ee),
	.w7(32'hbc8a51d6),
	.w8(32'hbbbdaa2e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cbb6d),
	.w1(32'hbb3c692a),
	.w2(32'hbc5913f5),
	.w3(32'hbc1226cf),
	.w4(32'h3c873aea),
	.w5(32'hbba8982b),
	.w6(32'hbcc7cc2c),
	.w7(32'hbae61578),
	.w8(32'h3bb4f23f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0fa2c),
	.w1(32'h3ad516a2),
	.w2(32'h3c841937),
	.w3(32'hbae47e4c),
	.w4(32'h3cca8e64),
	.w5(32'hbbaabafa),
	.w6(32'hbc30e667),
	.w7(32'hbc69abca),
	.w8(32'hbbad3744),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c019bf2),
	.w1(32'h3cc55e3f),
	.w2(32'h3ce8ca22),
	.w3(32'hbc987502),
	.w4(32'h3b8242ee),
	.w5(32'h3c014b25),
	.w6(32'hba3f9110),
	.w7(32'h3b49570a),
	.w8(32'hbb72d8ff),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389fd887),
	.w1(32'hbcae005c),
	.w2(32'hbc2dfde5),
	.w3(32'h3c433446),
	.w4(32'hbc2d16da),
	.w5(32'h3b7fb050),
	.w6(32'hb9d9ddd3),
	.w7(32'hbc1f2dfa),
	.w8(32'hbb7aea1a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2d38a),
	.w1(32'hbcacae85),
	.w2(32'hbbeb944b),
	.w3(32'hbd193ec1),
	.w4(32'hbc8bafd2),
	.w5(32'hbcc7edab),
	.w6(32'hbce7d52d),
	.w7(32'hbc41c3bf),
	.w8(32'hbb3234f1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19ba2c),
	.w1(32'hbc23fac3),
	.w2(32'hbb385bf8),
	.w3(32'h3ca55a93),
	.w4(32'h3b54fda3),
	.w5(32'hbb699a93),
	.w6(32'hbc08621a),
	.w7(32'hbb748adf),
	.w8(32'hbbba3803),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c598b46),
	.w1(32'h3aa1da78),
	.w2(32'hbc8b6da4),
	.w3(32'hbc2f56e1),
	.w4(32'h3bb3b084),
	.w5(32'h3be873d1),
	.w6(32'hbc1ac592),
	.w7(32'h3c3cefb3),
	.w8(32'hbabdcd1a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88cb28),
	.w1(32'h3bbfc69c),
	.w2(32'h3aaba8b5),
	.w3(32'hbc68f4d5),
	.w4(32'hbc0b9491),
	.w5(32'hbb97eb03),
	.w6(32'h3c068f5b),
	.w7(32'h3c8451b3),
	.w8(32'hbb9cf067),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc790517),
	.w1(32'h3b5cf11e),
	.w2(32'hbbb0b76e),
	.w3(32'h3bb6757f),
	.w4(32'hbbb7cb6d),
	.w5(32'hbae756a5),
	.w6(32'h3be46d0a),
	.w7(32'h3c77822d),
	.w8(32'h3d3e1ee9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c2085),
	.w1(32'h3c1b49ee),
	.w2(32'hbc1cbb6d),
	.w3(32'h3c0ca44c),
	.w4(32'h3ce52a5b),
	.w5(32'hba8f5989),
	.w6(32'hbbbfd963),
	.w7(32'h3bce2c2b),
	.w8(32'hbaea8bb3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb813e),
	.w1(32'hbc2921f2),
	.w2(32'hbbdbcd4c),
	.w3(32'h3a89a3ee),
	.w4(32'hbc24442b),
	.w5(32'hbc7e7627),
	.w6(32'h3ca284da),
	.w7(32'hbad10f75),
	.w8(32'h3c380bc0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c822cac),
	.w1(32'h3bca2e52),
	.w2(32'h3a0db6bf),
	.w3(32'h3898a2b9),
	.w4(32'hbc39e84a),
	.w5(32'hbc5d5b88),
	.w6(32'h3b8c7884),
	.w7(32'hbb54a497),
	.w8(32'hb9a11841),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f2d0f),
	.w1(32'h3af913e4),
	.w2(32'hbb59e66f),
	.w3(32'hbbc5b7d6),
	.w4(32'hbcab2b28),
	.w5(32'hbbae35e5),
	.w6(32'hbbc4c368),
	.w7(32'h39fe8405),
	.w8(32'hba90ab97),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b246af2),
	.w1(32'h3aaa85e3),
	.w2(32'hbb4ecf5a),
	.w3(32'h3b1e25ee),
	.w4(32'h3954800d),
	.w5(32'h3c1bf53d),
	.w6(32'hbc033a32),
	.w7(32'h3c6d64c3),
	.w8(32'hb9ebdf53),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3871e2),
	.w1(32'hbb7567dd),
	.w2(32'h3c19fed2),
	.w3(32'hbc81f6d7),
	.w4(32'hbba1e5bb),
	.w5(32'h3c3b95a8),
	.w6(32'hbb8fa0e4),
	.w7(32'hbb8f1743),
	.w8(32'h3a1d4118),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ebb8f),
	.w1(32'h3d1b5d59),
	.w2(32'h3cd2ecbf),
	.w3(32'h3a0b3e1e),
	.w4(32'h3bdc1572),
	.w5(32'hbbc40e10),
	.w6(32'h3d2bd8d2),
	.w7(32'h3c42311d),
	.w8(32'h3a9d4369),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc699ea6),
	.w1(32'h3c3cf8a1),
	.w2(32'hba8390b4),
	.w3(32'h3c2445c3),
	.w4(32'h3b7c63ad),
	.w5(32'hbcb5e8b0),
	.w6(32'hbc94554e),
	.w7(32'h3c1047e5),
	.w8(32'hbc74450b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf88ccb),
	.w1(32'hbc04610a),
	.w2(32'hbbb8e4fd),
	.w3(32'hbc1571c5),
	.w4(32'h3b815ba2),
	.w5(32'hbc399138),
	.w6(32'h39d28fd9),
	.w7(32'hbb973140),
	.w8(32'hbabf2f09),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bbd74),
	.w1(32'h3b21a0e4),
	.w2(32'h3ba50772),
	.w3(32'h3b20d65d),
	.w4(32'h3a5b7a5b),
	.w5(32'hbc615987),
	.w6(32'h3c42c8ab),
	.w7(32'h3b185c56),
	.w8(32'h3aa10023),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9eca96),
	.w1(32'h3a2d9f17),
	.w2(32'hbbf15ce2),
	.w3(32'hbba780f1),
	.w4(32'hbc203d1e),
	.w5(32'hbbacee70),
	.w6(32'hbb3e42fd),
	.w7(32'hbb4400b1),
	.w8(32'h3aa7f4b3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef8da3),
	.w1(32'hbc1448cd),
	.w2(32'hbc4b68b0),
	.w3(32'hbcd7490a),
	.w4(32'hbbf84de8),
	.w5(32'hbc9ced07),
	.w6(32'hbbfd6163),
	.w7(32'hbc3838c2),
	.w8(32'hbb469018),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c895c),
	.w1(32'hbb8ff8d2),
	.w2(32'hbc2e25ab),
	.w3(32'hbba9e46c),
	.w4(32'h3b9e0bb0),
	.w5(32'h3aa9bb17),
	.w6(32'hbcb99792),
	.w7(32'hb8920612),
	.w8(32'h3cb8f95f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0e2f9),
	.w1(32'hbbd808fc),
	.w2(32'h3b00bbc6),
	.w3(32'hbb39d631),
	.w4(32'h3ba95027),
	.w5(32'hbb475cf8),
	.w6(32'hbbe2f585),
	.w7(32'hbc55e640),
	.w8(32'hbb660264),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82e779),
	.w1(32'hbb133e1e),
	.w2(32'h3c79b122),
	.w3(32'hba0f4d94),
	.w4(32'hbc06e42d),
	.w5(32'h3b379948),
	.w6(32'h3b8c4c0e),
	.w7(32'hbbe76a80),
	.w8(32'hbbb544bb),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb90ff),
	.w1(32'hbba38a69),
	.w2(32'hbbad8d3b),
	.w3(32'h3b8f5b27),
	.w4(32'h3b9581e2),
	.w5(32'hbc1be9f1),
	.w6(32'hbb07dc03),
	.w7(32'hbc90b8fb),
	.w8(32'hbb80b211),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc738f85),
	.w1(32'hbb993b15),
	.w2(32'h3c2dc826),
	.w3(32'hbc129924),
	.w4(32'hbb2680e3),
	.w5(32'hbc1f80f6),
	.w6(32'hbc872088),
	.w7(32'hbc243823),
	.w8(32'h3b038f42),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fdc11),
	.w1(32'h3ae62a1e),
	.w2(32'hbb8a6aba),
	.w3(32'hbb801e64),
	.w4(32'h3c86b697),
	.w5(32'hbb62631c),
	.w6(32'h3b9067dd),
	.w7(32'hbaefb8c7),
	.w8(32'h3a274700),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30ec3b),
	.w1(32'hbb525435),
	.w2(32'hbca509dd),
	.w3(32'hbb189340),
	.w4(32'hbc3c4c50),
	.w5(32'hbc36b73f),
	.w6(32'hbc08fde8),
	.w7(32'hbc1bf2a8),
	.w8(32'hbbc1479f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb866e408),
	.w1(32'h3ab7036c),
	.w2(32'h3bb1990a),
	.w3(32'h3cd4ce05),
	.w4(32'h3a38ca87),
	.w5(32'h3bbe3639),
	.w6(32'h3a6c9f3f),
	.w7(32'h3d067364),
	.w8(32'h3aa65e15),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4adb01),
	.w1(32'hbada2a11),
	.w2(32'h3c3b1b2a),
	.w3(32'hba875c27),
	.w4(32'h3b186d6c),
	.w5(32'hbc409186),
	.w6(32'hbca60f63),
	.w7(32'hbbd13c42),
	.w8(32'hbbc9f0df),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule