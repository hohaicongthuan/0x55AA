module layer_6_featuremap_17(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7665b),
	.w1(32'h3c032179),
	.w2(32'hbdf12dc5),
	.w3(32'hbd2c2bae),
	.w4(32'h3c6f73c4),
	.w5(32'h3d224342),
	.w6(32'hbb5cc7b8),
	.w7(32'h3d2fea1b),
	.w8(32'hbd7254af),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e0e455a),
	.w1(32'h3c4dede2),
	.w2(32'hbba5dc95),
	.w3(32'hbd4f81a1),
	.w4(32'h3c46b764),
	.w5(32'hbb40911d),
	.w6(32'h3c81910b),
	.w7(32'h3c13e3f0),
	.w8(32'h3c969078),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb37d54),
	.w1(32'h3c492e0a),
	.w2(32'hbcd6d881),
	.w3(32'h3b612ca6),
	.w4(32'h3cd316b5),
	.w5(32'hbc41be5f),
	.w6(32'h3c1762f3),
	.w7(32'hbc4266ad),
	.w8(32'h3c9e7ead),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9357a1),
	.w1(32'h3d56a000),
	.w2(32'hbd9f04e0),
	.w3(32'hbc40d9d0),
	.w4(32'hbd6e926d),
	.w5(32'h3da70925),
	.w6(32'h3bab1bea),
	.w7(32'hbbc7aaa1),
	.w8(32'hbbc59810),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d195918),
	.w1(32'hbb5ba193),
	.w2(32'hbb88b08f),
	.w3(32'hbd11eb1b),
	.w4(32'hbc1bf635),
	.w5(32'hb9b455a0),
	.w6(32'h3af4ec33),
	.w7(32'hb97d6b9c),
	.w8(32'hbb25545a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb477ec9),
	.w1(32'hbb1b6c2f),
	.w2(32'h3cdb260e),
	.w3(32'hba09ddf3),
	.w4(32'hbcaee826),
	.w5(32'hbc6a8e77),
	.w6(32'h3a5e1374),
	.w7(32'hbd2655ba),
	.w8(32'h3bd0f45f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd04edd3),
	.w1(32'h3b0029b5),
	.w2(32'hbb4b7b21),
	.w3(32'hbba63071),
	.w4(32'h3bd43b9b),
	.w5(32'h3bc101d8),
	.w6(32'h3bf6d149),
	.w7(32'h3b346977),
	.w8(32'h3c12c887),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7be4f8),
	.w1(32'hbc9a3b71),
	.w2(32'hbca7a25c),
	.w3(32'h3c7151f7),
	.w4(32'hbc00b3f2),
	.w5(32'hbb6f8916),
	.w6(32'h3b53fdc1),
	.w7(32'h3c8b0c32),
	.w8(32'hbcb4397b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd73c10),
	.w1(32'hbac16689),
	.w2(32'hbc110005),
	.w3(32'h3cfa562b),
	.w4(32'h3c236615),
	.w5(32'hbb976b76),
	.w6(32'h3bb8e540),
	.w7(32'hbb8b8cc5),
	.w8(32'h3a153b20),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb898531),
	.w1(32'h3b447901),
	.w2(32'h3a8c8259),
	.w3(32'h3c5fed00),
	.w4(32'h3bb60b9a),
	.w5(32'h3bfafea5),
	.w6(32'h3bebeec4),
	.w7(32'h3bfb508d),
	.w8(32'h3b3b2f0e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c9fee),
	.w1(32'h3b736592),
	.w2(32'h38426e6f),
	.w3(32'h3b92e04f),
	.w4(32'h3ce7b625),
	.w5(32'hbc1163f3),
	.w6(32'h3c3871a6),
	.w7(32'hbbce1a27),
	.w8(32'h3cb71c3a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f6dfa),
	.w1(32'hbc187762),
	.w2(32'hbb8b370f),
	.w3(32'hbb2b5c5c),
	.w4(32'hbc2433e0),
	.w5(32'h3b17b1c4),
	.w6(32'hbae943ac),
	.w7(32'h3c82a564),
	.w8(32'hbb8d57bd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd05d32),
	.w1(32'h3c9af669),
	.w2(32'h3d59e9ed),
	.w3(32'h3b7455b8),
	.w4(32'hbac4e706),
	.w5(32'h3c93b63a),
	.w6(32'hbd4216f8),
	.w7(32'h3aff48ef),
	.w8(32'h3b57957a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8edd85),
	.w1(32'hbb0c865e),
	.w2(32'h3b8d309c),
	.w3(32'hbd33881c),
	.w4(32'hbbf3b27d),
	.w5(32'hbc9c5557),
	.w6(32'hbb754ebc),
	.w7(32'hbc7ba632),
	.w8(32'hbbe95cf7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cca8f),
	.w1(32'hbcf1cf37),
	.w2(32'hbd290b1d),
	.w3(32'h3b1a31b3),
	.w4(32'h3d112140),
	.w5(32'hbc8d0152),
	.w6(32'h3c786e66),
	.w7(32'h3cbd5d90),
	.w8(32'hbd4119bd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2dd6a8),
	.w1(32'hbbe5b01c),
	.w2(32'hbc1027f3),
	.w3(32'hbc34ce59),
	.w4(32'h3cd3056c),
	.w5(32'hbd892bfd),
	.w6(32'hbb8dc739),
	.w7(32'hbc9760d4),
	.w8(32'h3c4bdd75),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fe77f),
	.w1(32'hbdb855f1),
	.w2(32'h3e5de0e3),
	.w3(32'h3af8f426),
	.w4(32'h3d3689c9),
	.w5(32'hbd36bbf0),
	.w6(32'h3d4f84a7),
	.w7(32'hbd996302),
	.w8(32'hbc0ae181),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd062224),
	.w1(32'hbd0af7b8),
	.w2(32'hbb4e367e),
	.w3(32'hbcb2f898),
	.w4(32'h3cb10001),
	.w5(32'hbb78dc23),
	.w6(32'hbbac0cdb),
	.w7(32'h3be69dab),
	.w8(32'hbc5103dc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c4b73),
	.w1(32'h3c1445d2),
	.w2(32'hbaa9cbe2),
	.w3(32'hbcf32008),
	.w4(32'h3b6ff1e8),
	.w5(32'h3bbc1906),
	.w6(32'h3baae24f),
	.w7(32'h3be7b755),
	.w8(32'hba874c32),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b8a7a),
	.w1(32'hbd9266d3),
	.w2(32'h3dad065f),
	.w3(32'h3beb7793),
	.w4(32'h3d916a79),
	.w5(32'hbdbf3004),
	.w6(32'hbc3f0a99),
	.w7(32'h3b979e4c),
	.w8(32'h3c170121),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7370d2),
	.w1(32'hbccfcd0f),
	.w2(32'h3caa080d),
	.w3(32'h3d0a0e4c),
	.w4(32'h3c543186),
	.w5(32'hbd019002),
	.w6(32'hbc1ae62c),
	.w7(32'hbaec7abd),
	.w8(32'hbd0e7a08),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bf10c),
	.w1(32'h3a99ed2e),
	.w2(32'h3bbd5ca0),
	.w3(32'hbc252c42),
	.w4(32'hbac3754d),
	.w5(32'hbb83141d),
	.w6(32'h3c0dc6b1),
	.w7(32'hbb977423),
	.w8(32'hbbecaaeb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85c9e6),
	.w1(32'hbbbc7256),
	.w2(32'hba83f3b9),
	.w3(32'h3befb027),
	.w4(32'h3bfc3889),
	.w5(32'hbc785ccc),
	.w6(32'h3c397fd8),
	.w7(32'hbcd6c706),
	.w8(32'h3c9133ef),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc508e2),
	.w1(32'hbcbb19ab),
	.w2(32'hbdaca0d7),
	.w3(32'hbc1eb523),
	.w4(32'hbd3bf5e3),
	.w5(32'h3989545c),
	.w6(32'hbc873819),
	.w7(32'h3caec75d),
	.w8(32'hbd194463),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd304a5e),
	.w1(32'hbcbf97fd),
	.w2(32'hbb71c0b6),
	.w3(32'h3caacb2c),
	.w4(32'h3c4f0998),
	.w5(32'h3d53edaf),
	.w6(32'h3d1f15cb),
	.w7(32'h3c706703),
	.w8(32'hbcc7a4e5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d70be41),
	.w1(32'hbaab4c31),
	.w2(32'h3c3a690c),
	.w3(32'hbd100377),
	.w4(32'h3bc05046),
	.w5(32'h3b6799ee),
	.w6(32'h3bcf225f),
	.w7(32'h3ce80864),
	.w8(32'hbc298fff),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce89266),
	.w1(32'hbcc3d77f),
	.w2(32'h3d557dab),
	.w3(32'hbc8a29b6),
	.w4(32'hbc4f62dd),
	.w5(32'hbce90f5f),
	.w6(32'hbca37e71),
	.w7(32'hbd1830fa),
	.w8(32'hbd073157),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68a2be),
	.w1(32'h3c35d178),
	.w2(32'hbd1675c8),
	.w3(32'hbd75c907),
	.w4(32'hbd29c8db),
	.w5(32'hba89e67f),
	.w6(32'hbc0f8fc2),
	.w7(32'hbc859c2d),
	.w8(32'hbbd443a3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c7ea8),
	.w1(32'h3aae8213),
	.w2(32'h3d9492a8),
	.w3(32'h3be79b58),
	.w4(32'hbc56f105),
	.w5(32'hbcf8aae7),
	.w6(32'hbc83118c),
	.w7(32'hbc807a76),
	.w8(32'hbd1a97f7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b46d0),
	.w1(32'h3ceffa30),
	.w2(32'hbd06dedd),
	.w3(32'hbc351ac2),
	.w4(32'hbd52c023),
	.w5(32'h3d0116eb),
	.w6(32'hbcd1abc5),
	.w7(32'h3d131daf),
	.w8(32'hbc6d29f8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd092076),
	.w1(32'hb81405a8),
	.w2(32'hb8cedf91),
	.w3(32'h3d166c0b),
	.w4(32'h38a1888a),
	.w5(32'h38216b33),
	.w6(32'h38ac3488),
	.w7(32'hb66be402),
	.w8(32'hb5ff6609),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d668),
	.w1(32'h3a74f655),
	.w2(32'h3b2b23d5),
	.w3(32'h3b30c0a5),
	.w4(32'h3b0ecb45),
	.w5(32'h3b86ff2a),
	.w6(32'h3bacda38),
	.w7(32'h3b7505f3),
	.w8(32'h3acc2070),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5d652),
	.w1(32'hba901701),
	.w2(32'hba649d91),
	.w3(32'hbaabb980),
	.w4(32'hba8bf6dc),
	.w5(32'hba6e2891),
	.w6(32'hba997b9d),
	.w7(32'hba7da5de),
	.w8(32'hba437461),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0f450),
	.w1(32'hb9548332),
	.w2(32'hb94dc7b2),
	.w3(32'hb99d6886),
	.w4(32'hb939f2b0),
	.w5(32'hb982ca3b),
	.w6(32'hb984a07c),
	.w7(32'hb94f3aa1),
	.w8(32'hb95dae64),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cac989),
	.w1(32'hb9aeceaf),
	.w2(32'hb9da2959),
	.w3(32'hba2bc5ee),
	.w4(32'hb9acb51a),
	.w5(32'hba6b4d1e),
	.w6(32'hb9509942),
	.w7(32'hb995fe5a),
	.w8(32'hba0e88d2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81b1c6),
	.w1(32'h3b8da4db),
	.w2(32'h3a7d4674),
	.w3(32'hbb157156),
	.w4(32'hb9c6d4a0),
	.w5(32'h3b50d13c),
	.w6(32'h3b5446e1),
	.w7(32'h3b7314a6),
	.w8(32'hbb85b66f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa145f),
	.w1(32'hbaa4c0eb),
	.w2(32'hbaf0d804),
	.w3(32'hba4a758a),
	.w4(32'hba94bc52),
	.w5(32'hbac12550),
	.w6(32'hba3651ee),
	.w7(32'hba98fdf1),
	.w8(32'hba93419c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eb70c),
	.w1(32'h3bbcf189),
	.w2(32'h3b20f595),
	.w3(32'hbaf93cb4),
	.w4(32'h38142e17),
	.w5(32'hbab4f75e),
	.w6(32'h3aed69ca),
	.w7(32'h3a816b82),
	.w8(32'hbac39abf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384864bf),
	.w1(32'hb8d0d283),
	.w2(32'h39c102f4),
	.w3(32'h39e7d8bc),
	.w4(32'h3a6a4961),
	.w5(32'h39ddbf3c),
	.w6(32'hb973030a),
	.w7(32'h38a50163),
	.w8(32'h398691c1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1fec7),
	.w1(32'hbbbb7a27),
	.w2(32'h3cb24d50),
	.w3(32'h3bac082f),
	.w4(32'hbb7d71cb),
	.w5(32'hbc94e7f6),
	.w6(32'h3c2fac54),
	.w7(32'hbc36861f),
	.w8(32'hbb1d98b0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0de09),
	.w1(32'h3c12a558),
	.w2(32'h3bf8bea3),
	.w3(32'h3bd0077a),
	.w4(32'h3c010b20),
	.w5(32'h3ba5ff38),
	.w6(32'h3c318ed6),
	.w7(32'h3c2ce803),
	.w8(32'h3ba51a86),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5c11),
	.w1(32'h3bdd2254),
	.w2(32'h3b603cda),
	.w3(32'h3a9c906a),
	.w4(32'h3b3a31b7),
	.w5(32'h3b7641fa),
	.w6(32'h3b58193c),
	.w7(32'h3ba69278),
	.w8(32'h3a243fae),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5803590),
	.w1(32'hb8016566),
	.w2(32'hb68e8082),
	.w3(32'h3797b544),
	.w4(32'hb7a82340),
	.w5(32'hb780147d),
	.w6(32'hb6ded829),
	.w7(32'hb84a1359),
	.w8(32'hb8328d75),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba54ea),
	.w1(32'h3c821f26),
	.w2(32'hbcc12cce),
	.w3(32'hbc2e3157),
	.w4(32'hbc6e0d7b),
	.w5(32'h3be01480),
	.w6(32'hbc25a130),
	.w7(32'h3c20aba9),
	.w8(32'hbca27917),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c13e3),
	.w1(32'hbc576a6a),
	.w2(32'h39f6026f),
	.w3(32'h39f35866),
	.w4(32'hbb2f0ac1),
	.w5(32'hbc332093),
	.w6(32'h3be85439),
	.w7(32'hbb887e5b),
	.w8(32'hbc084a76),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0ffb0),
	.w1(32'h38b54626),
	.w2(32'h38da662f),
	.w3(32'h38696fad),
	.w4(32'h3833f539),
	.w5(32'h381e923e),
	.w6(32'h3891f704),
	.w7(32'h37fffda0),
	.w8(32'hb6bf5917),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8737631),
	.w1(32'hb884f8b0),
	.w2(32'hb85e558c),
	.w3(32'hb8929f7a),
	.w4(32'hb8b76544),
	.w5(32'hb82717c0),
	.w6(32'hb81e8667),
	.w7(32'hb85fe214),
	.w8(32'hb88abf70),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb423f35),
	.w1(32'hbba378ee),
	.w2(32'hbc2dc5a8),
	.w3(32'hbbac6fef),
	.w4(32'hbbb8bc6e),
	.w5(32'hbbbf5bdb),
	.w6(32'hbb233b26),
	.w7(32'hbb9340c0),
	.w8(32'hbc2b260f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20e364),
	.w1(32'h3b6d3c81),
	.w2(32'h3bbbabb2),
	.w3(32'h3aab4fca),
	.w4(32'h3991e2de),
	.w5(32'h3b3cf0fe),
	.w6(32'h3b8a57a4),
	.w7(32'h3b97b9a2),
	.w8(32'h3c02cd45),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b291106),
	.w1(32'hbacd3e4b),
	.w2(32'hbba756dd),
	.w3(32'h3b426e25),
	.w4(32'hbb90d987),
	.w5(32'hbc1aac4f),
	.w6(32'hba9ac2ba),
	.w7(32'hbbbe72aa),
	.w8(32'hbc13af93),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db3db),
	.w1(32'h3b5ca775),
	.w2(32'h3b26d35d),
	.w3(32'h3b224970),
	.w4(32'h3b5dc0bf),
	.w5(32'h3acc428b),
	.w6(32'h3bd14538),
	.w7(32'h3b948fc7),
	.w8(32'hbb22eeb5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbc2d0),
	.w1(32'h3c253621),
	.w2(32'h3bcd508d),
	.w3(32'h3ba9e54d),
	.w4(32'h3baf84ed),
	.w5(32'h3b383fe1),
	.w6(32'h3bcce2c1),
	.w7(32'h3bdd3948),
	.w8(32'h3b5836d4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57f72f),
	.w1(32'hbc824a34),
	.w2(32'hbbdb33fc),
	.w3(32'hbb8d34a8),
	.w4(32'hbc1ae752),
	.w5(32'hbcb11d64),
	.w6(32'h3a9e9b08),
	.w7(32'hbc638823),
	.w8(32'hbcb305dc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f4218),
	.w1(32'hbad76912),
	.w2(32'hbb7fec18),
	.w3(32'h396b8495),
	.w4(32'hbb6ca1fc),
	.w5(32'hbb250cfb),
	.w6(32'h3b27fd80),
	.w7(32'h3a0535a4),
	.w8(32'h3bad5157),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39890eef),
	.w1(32'hbaa0d359),
	.w2(32'hba9f1fb3),
	.w3(32'h3ac0ecd2),
	.w4(32'hba8561c1),
	.w5(32'h3916f19a),
	.w6(32'h3a756d80),
	.w7(32'hb93e54de),
	.w8(32'h3aa7e84e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48204a),
	.w1(32'h3c760271),
	.w2(32'h3bf73460),
	.w3(32'h3bd09c8f),
	.w4(32'h3c7603cf),
	.w5(32'h3c908698),
	.w6(32'h3c21fd43),
	.w7(32'h3c4d35ba),
	.w8(32'h3b67326e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc2296),
	.w1(32'hba96aa54),
	.w2(32'h3a42a929),
	.w3(32'hbb9916af),
	.w4(32'hbbced680),
	.w5(32'hbba2a751),
	.w6(32'hb820e9b3),
	.w7(32'hb9ad850c),
	.w8(32'h3a85a110),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20a5e0),
	.w1(32'hbc0d8c5c),
	.w2(32'hbc1eaf91),
	.w3(32'hbc36cad8),
	.w4(32'hbc0d36e6),
	.w5(32'hbbfe94d5),
	.w6(32'hbc308c76),
	.w7(32'hbc20aaca),
	.w8(32'hbc1cc1e8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b675f7b),
	.w1(32'h3b17d323),
	.w2(32'h3b6a38ce),
	.w3(32'hb84b18a4),
	.w4(32'h3a8bc007),
	.w5(32'h3a948b72),
	.w6(32'h3b0520ea),
	.w7(32'h3b6adc13),
	.w8(32'h3b0cccb9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c46e4),
	.w1(32'h3c446f0e),
	.w2(32'h3c992c96),
	.w3(32'h3c10e24c),
	.w4(32'h3c69e9cf),
	.w5(32'h3bbf2cc7),
	.w6(32'h3cc7f4d7),
	.w7(32'h3c618a64),
	.w8(32'h3a568c3d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfff581),
	.w1(32'h3b967d47),
	.w2(32'h3b18c7e1),
	.w3(32'h3c05fdb7),
	.w4(32'h3c2a69b4),
	.w5(32'h3b46fad9),
	.w6(32'h3afc6660),
	.w7(32'h3b70afb6),
	.w8(32'hbc03cd23),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be315ad),
	.w1(32'h3b94605a),
	.w2(32'h3c01bc11),
	.w3(32'hba08b28c),
	.w4(32'h3ac448a8),
	.w5(32'h3b27a9a2),
	.w6(32'h3c46cb62),
	.w7(32'h3c1dfd6c),
	.w8(32'hbb5acb8a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f51ed),
	.w1(32'h3cb15df1),
	.w2(32'hbd78ab13),
	.w3(32'hbc2fd255),
	.w4(32'h3c0a038c),
	.w5(32'h3c9c6e0f),
	.w6(32'h3b725c40),
	.w7(32'h3ce270cd),
	.w8(32'hbb1b381c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb252647),
	.w1(32'h3aa194fe),
	.w2(32'hbd64881e),
	.w3(32'h3a85b544),
	.w4(32'h3c6c0b5e),
	.w5(32'hbd358990),
	.w6(32'h3d2c711f),
	.w7(32'h3c2d7847),
	.w8(32'hbbb45008),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule