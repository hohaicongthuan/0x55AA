module layer_8_featuremap_21(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f805fca),
	.w1(32'h3e299fd5),
	.w2(32'h3e52f32f),
	.w3(32'h3e1e5360),
	.w4(32'h3f649101),
	.w5(32'h3922a30c),
	.w6(32'h3e62e825),
	.w7(32'h3f05be4d),
	.w8(32'h3e73827b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb711538b),
	.w1(32'h3e16d97a),
	.w2(32'h3f930ce4),
	.w3(32'h3fa90a7e),
	.w4(32'h3e43b331),
	.w5(32'h3f8432d7),
	.w6(32'h3e310d5b),
	.w7(32'h3f9d3a02),
	.w8(32'h3f82d412),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e9e730f),
	.w1(32'h3d990f40),
	.w2(32'h3d926202),
	.w3(32'h3d353c73),
	.w4(32'h3f0873d7),
	.w5(32'hb83fece6),
	.w6(32'h3e84b4f7),
	.w7(32'h3f0ba153),
	.w8(32'h3e204732),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fb3bfc8),
	.w1(32'h3e49695e),
	.w2(32'h38374fba),
	.w3(32'h3f927bb3),
	.w4(32'h3d7d3830),
	.w5(32'h3d04f189),
	.w6(32'hb7c90c70),
	.w7(32'h3daf22bf),
	.w8(32'h3e24975a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e8b0a62),
	.w1(32'h3e43f499),
	.w2(32'h3e9206fa),
	.w3(32'h3f63a4ae),
	.w4(32'h3e965351),
	.w5(32'h3f5aedcf),
	.w6(32'hb843001c),
	.w7(32'hb896904b),
	.w8(32'h3ed52411),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6417f),
	.w1(32'h3f8cd45d),
	.w2(32'h3e0f22a8),
	.w3(32'h3f6ecdcd),
	.w4(32'h3e9e56bf),
	.w5(32'h3e378958),
	.w6(32'h3faf28b6),
	.w7(32'h3ee73aa0),
	.w8(32'hb8a32528),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5cabdcc),
	.w1(32'h3d865c92),
	.w2(32'h3f9ba484),
	.w3(32'h3d3cecba),
	.w4(32'hb4b50c68),
	.w5(32'h3d6f1d23),
	.w6(32'h3fbca632),
	.w7(32'h3f9074d7),
	.w8(32'h3f71a5b6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f616586),
	.w1(32'h3e8eb296),
	.w2(32'h3e4c6aa2),
	.w3(32'h3fae5d0e),
	.w4(32'h3deb4b8f),
	.w5(32'h3ecda35d),
	.w6(32'hb7b665b3),
	.w7(32'h3e45a1c0),
	.w8(32'h3e0bcf5d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2d1028),
	.w1(32'h3ec991dd),
	.w2(32'h3e9ad5a8),
	.w3(32'h3fab2535),
	.w4(32'hb7b0c743),
	.w5(32'h3f11811a),
	.w6(32'h3f5fd633),
	.w7(32'h3e36bf80),
	.w8(32'h3f5af50c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f1c9fde),
	.w1(32'h3e0ebeb2),
	.w2(32'h3f804646),
	.w3(32'h3dc1e022),
	.w4(32'h3f68c94a),
	.w5(32'h3e06430c),
	.w6(32'hb80b13b1),
	.w7(32'h3e27d12f),
	.w8(32'h3e1086e7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e6aa04d),
	.w1(32'h3fa43526),
	.w2(32'h3d1c4afb),
	.w3(32'h3d3d74bd),
	.w4(32'h3f492a6f),
	.w5(32'h3e8111f2),
	.w6(32'h3f9610c2),
	.w7(32'h3ed8c0b7),
	.w8(32'h38ebde70),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e823ada),
	.w1(32'h38596363),
	.w2(32'h3f653aac),
	.w3(32'h3f7c2a4a),
	.w4(32'h383d92fc),
	.w5(32'h3dcf291f),
	.w6(32'hbec23fe4),
	.w7(32'h3d28823a),
	.w8(32'h3ed95532),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ebcca90),
	.w1(32'h3dfd56c9),
	.w2(32'h3c515499),
	.w3(32'h375633d6),
	.w4(32'hb8615eac),
	.w5(32'h3de9ce21),
	.w6(32'h3e5becf2),
	.w7(32'h3d840013),
	.w8(32'h3e374f0a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7a6fc),
	.w1(32'h3d9380e4),
	.w2(32'h3f075f5e),
	.w3(32'hbe0fb312),
	.w4(32'h3ddc91ef),
	.w5(32'hbee1a358),
	.w6(32'h3e0b13b8),
	.w7(32'hbf44a150),
	.w8(32'h3e427bde),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d89bb8f),
	.w1(32'h3b8a5d08),
	.w2(32'h3ef5deb2),
	.w3(32'hb6257721),
	.w4(32'h3d0b8dd3),
	.w5(32'h3c800670),
	.w6(32'h3d012874),
	.w7(32'h3db3d91f),
	.w8(32'h3c00c1bd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3540e004),
	.w1(32'h3e011118),
	.w2(32'h3d84f835),
	.w3(32'h3e2e60a2),
	.w4(32'hbc20b025),
	.w5(32'h3e850799),
	.w6(32'h36938208),
	.w7(32'h3d1df869),
	.w8(32'hbffbfeb7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e838bfd),
	.w1(32'h3d78c75d),
	.w2(32'h3cce54d8),
	.w3(32'h3c9dc4ae),
	.w4(32'h3e201806),
	.w5(32'h3e8c3ae1),
	.w6(32'h3e426371),
	.w7(32'h3d69e0c8),
	.w8(32'h3da3b531),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38040afd),
	.w1(32'h3e3bb3ce),
	.w2(32'hbc1cb837),
	.w3(32'h3c9f08c5),
	.w4(32'h3781f610),
	.w5(32'h3e1d6845),
	.w6(32'h3ec877b1),
	.w7(32'hbd19017d),
	.w8(32'h386741db),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d165fd5),
	.w1(32'hbdd783e5),
	.w2(32'hbd62ed48),
	.w3(32'h3d685f31),
	.w4(32'h39b34c72),
	.w5(32'h39f540a5),
	.w6(32'h3df8cf70),
	.w7(32'h3cbbee85),
	.w8(32'h3e06a858),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e8b3e2e),
	.w1(32'h3eee2654),
	.w2(32'h3e18252c),
	.w3(32'h3e3bb39a),
	.w4(32'hbcf16e4f),
	.w5(32'h3eaed037),
	.w6(32'h3cfc8918),
	.w7(32'hbf141269),
	.w8(32'h3df7f883),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c15f4),
	.w1(32'h3d5de6a0),
	.w2(32'h387dcacc),
	.w3(32'hb6546d87),
	.w4(32'h3d063103),
	.w5(32'h3d9efdb6),
	.w6(32'hb8cb4862),
	.w7(32'h3da49317),
	.w8(32'h3ed1667d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d75a1cf),
	.w1(32'h3edd433f),
	.w2(32'h3ba6373f),
	.w3(32'h3e50cce0),
	.w4(32'hb8bc3520),
	.w5(32'h3d8dc576),
	.w6(32'h3dc3df3e),
	.w7(32'h3dbf04b7),
	.w8(32'h3e0eb062),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd969d6a),
	.w1(32'h3eaa169b),
	.w2(32'h3906a5cc),
	.w3(32'h3ab635db),
	.w4(32'h3e84d173),
	.w5(32'h3dbe42aa),
	.w6(32'h3ad1af04),
	.w7(32'h3e71ea97),
	.w8(32'h3d14afa4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dfa8870),
	.w1(32'h3da04d1f),
	.w2(32'h3f2304a3),
	.w3(32'h3e651cc6),
	.w4(32'hb8539f19),
	.w5(32'hbd295555),
	.w6(32'h3e053e21),
	.w7(32'h3e22bb88),
	.w8(32'h3f60a0cd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab213d9),
	.w1(32'h3d044418),
	.w2(32'h3d0f69f6),
	.w3(32'h3b82f960),
	.w4(32'h3dab4609),
	.w5(32'h3e3b9a83),
	.w6(32'h3d82468a),
	.w7(32'h3e887345),
	.w8(32'hbcbc4cb5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd64f087),
	.w1(32'h3dd765b0),
	.w2(32'h3942b8c8),
	.w3(32'h3a7381d2),
	.w4(32'hbd9afa40),
	.w5(32'h3d46520a),
	.w6(32'h3dc332b1),
	.w7(32'hb78f455e),
	.w8(32'hbdda55e8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c6dda),
	.w1(32'h385ffbe4),
	.w2(32'hb689b487),
	.w3(32'h3edf1ab7),
	.w4(32'h3d53ce19),
	.w5(32'h3df41b88),
	.w6(32'h3e0823ab),
	.w7(32'h3d823497),
	.w8(32'h3a4061c9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6b40e),
	.w1(32'h3c953f91),
	.w2(32'h3a9af48f),
	.w3(32'h3b3cf500),
	.w4(32'h3aa14fe8),
	.w5(32'h3ef2690c),
	.w6(32'h3a8227eb),
	.w7(32'h3c2c9f97),
	.w8(32'h3c9e43a0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4ed537),
	.w1(32'h3897a9ba),
	.w2(32'h3b239fd0),
	.w3(32'h3b2520af),
	.w4(32'h3d68a90c),
	.w5(32'h3ad6d222),
	.w6(32'h3ca17fbf),
	.w7(32'h3a04a415),
	.w8(32'h3ce6264b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d96c3df),
	.w1(32'h3ab0df73),
	.w2(32'h3a236629),
	.w3(32'h3ac02f67),
	.w4(32'hb6e4c555),
	.w5(32'h3a4d09b3),
	.w6(32'hb6fc9785),
	.w7(32'h3d8cf18e),
	.w8(32'h3a963b2e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dafcd9e),
	.w1(32'h3d7e257d),
	.w2(32'h3bcc9eff),
	.w3(32'h3d108443),
	.w4(32'h3b3e9ce0),
	.w5(32'h3a76b53f),
	.w6(32'h3d232748),
	.w7(32'h3a2ff7fc),
	.w8(32'h3d4603b2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e88e586),
	.w1(32'h3b8ce353),
	.w2(32'h372a53c4),
	.w3(32'h3aa847c3),
	.w4(32'h3dbed940),
	.w5(32'h3a5d2e37),
	.w6(32'hb816f300),
	.w7(32'h3d4f1893),
	.w8(32'h3ae5683f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1426c),
	.w1(32'h3a805d6a),
	.w2(32'hb62942fc),
	.w3(32'hb5ff6e07),
	.w4(32'h3b8ca220),
	.w5(32'h3a3f20c2),
	.w6(32'h3a0125e2),
	.w7(32'h3d464f25),
	.w8(32'h3bee6846),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e75438),
	.w1(32'h3c02a4ac),
	.w2(32'h3dc8e09c),
	.w3(32'h3b5820b7),
	.w4(32'h3a109fc4),
	.w5(32'h3e5014de),
	.w6(32'h3de2ce81),
	.w7(32'h3cc7669b),
	.w8(32'h3c818896),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dfbc3a5),
	.w1(32'hb92456d7),
	.w2(32'h3df46aae),
	.w3(32'h3b203650),
	.w4(32'hb90de737),
	.w5(32'h3a822176),
	.w6(32'h3a29fb18),
	.w7(32'h3988a8e6),
	.w8(32'hb8ebc386),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a6109),
	.w1(32'h3d1d2a75),
	.w2(32'h37e52a28),
	.w3(32'h3e0037f7),
	.w4(32'h3d93feb3),
	.w5(32'h3abc5996),
	.w6(32'h39e00880),
	.w7(32'h3d999f6e),
	.w8(32'h3b21ad94),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ee2b),
	.w1(32'h39e1bc7d),
	.w2(32'h3dae0e77),
	.w3(32'h3a684eef),
	.w4(32'h3d4d854b),
	.w5(32'h3c1b51e9),
	.w6(32'h3be53e72),
	.w7(32'h3dbef915),
	.w8(32'h358f314c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8152fd),
	.w1(32'h3cd3e8aa),
	.w2(32'hb76b4d56),
	.w3(32'h3b83d736),
	.w4(32'h3d801e86),
	.w5(32'h3b32748b),
	.w6(32'h3c1babd6),
	.w7(32'h3a64e302),
	.w8(32'h3c90cfb3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17b8ef),
	.w1(32'h3a580969),
	.w2(32'h3d5def5d),
	.w3(32'h3cd9c388),
	.w4(32'h3a71fd3f),
	.w5(32'h3dadff75),
	.w6(32'h3b098e76),
	.w7(32'h3b4291f4),
	.w8(32'h3cfe0575),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd84ac4),
	.w1(32'h3635db89),
	.w2(32'h3c8fb200),
	.w3(32'h3a05f94a),
	.w4(32'h3acbe2f8),
	.w5(32'h34bd66af),
	.w6(32'h3c7beb1c),
	.w7(32'h3db5553f),
	.w8(32'h35eaeecd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a157e2f),
	.w1(32'h3c847350),
	.w2(32'h3abb11dd),
	.w3(32'h3cffcc43),
	.w4(32'h3d66791c),
	.w5(32'h3b1b5228),
	.w6(32'h3b124f17),
	.w7(32'h39249825),
	.w8(32'h39b13d55),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3865c0eb),
	.w1(32'h370f114d),
	.w2(32'hb7a99013),
	.w3(32'h384bd7d5),
	.w4(32'h37229232),
	.w5(32'hb7ca1980),
	.w6(32'h37eef3d2),
	.w7(32'hb7f3987b),
	.w8(32'hb809bf31),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a03866),
	.w1(32'hb7e55d11),
	.w2(32'hb7dbe7be),
	.w3(32'hb75f037c),
	.w4(32'hb78011b5),
	.w5(32'hb7acaf0d),
	.w6(32'hb80dd940),
	.w7(32'hb811525e),
	.w8(32'hb8295a44),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38db1d97),
	.w1(32'h38ce006c),
	.w2(32'h38ed8185),
	.w3(32'h38b9febf),
	.w4(32'h3880b999),
	.w5(32'h38b026d5),
	.w6(32'h38857a08),
	.w7(32'h378474bf),
	.w8(32'h3841a7d8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395bf9e6),
	.w1(32'h397e639b),
	.w2(32'h397db71d),
	.w3(32'h38dd0a4f),
	.w4(32'h38faacca),
	.w5(32'h394328b6),
	.w6(32'hb6652b09),
	.w7(32'hb7c4eba2),
	.w8(32'h38b87c2f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36833aff),
	.w1(32'hb6e9d200),
	.w2(32'hb82f6fa0),
	.w3(32'h37a50759),
	.w4(32'hb795caad),
	.w5(32'hb8013823),
	.w6(32'hb829438b),
	.w7(32'hb8be31b7),
	.w8(32'hb8c623a1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb544fda7),
	.w1(32'hb3802ec3),
	.w2(32'hb51fb3e1),
	.w3(32'hb52608ef),
	.w4(32'hb1aa9aa7),
	.w5(32'hb4f90e6a),
	.w6(32'h32d6d422),
	.w7(32'h3534d577),
	.w8(32'h3448ddb0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ccda03),
	.w1(32'h38d04852),
	.w2(32'h38d3250a),
	.w3(32'h38be23b0),
	.w4(32'h38bb9063),
	.w5(32'h38bd3053),
	.w6(32'hb7d4b894),
	.w7(32'hb7cfba67),
	.w8(32'h3728ce9e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382430f7),
	.w1(32'h378fc3fe),
	.w2(32'h383284b8),
	.w3(32'h37cc3396),
	.w4(32'h370240e6),
	.w5(32'h382524f4),
	.w6(32'hb76b77e3),
	.w7(32'hb802c208),
	.w8(32'hb53a4b8e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e1c2c),
	.w1(32'h389f0506),
	.w2(32'h38d20820),
	.w3(32'h38b46778),
	.w4(32'h3857545c),
	.w5(32'h390dcb44),
	.w6(32'h3801643e),
	.w7(32'h3821af5c),
	.w8(32'h38c19428),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37966693),
	.w1(32'hb8777ccf),
	.w2(32'hb8d33e7e),
	.w3(32'hb3e35390),
	.w4(32'hb8a2963e),
	.w5(32'hb8cfe18f),
	.w6(32'hb8ad35db),
	.w7(32'hb92cacfb),
	.w8(32'hb91ed399),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3f5e6),
	.w1(32'h39d47b81),
	.w2(32'h39dae6ee),
	.w3(32'h39be8308),
	.w4(32'h39aab69d),
	.w5(32'h39e85d87),
	.w6(32'h396c374c),
	.w7(32'h3904245e),
	.w8(32'h399ab4a5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a4c71),
	.w1(32'h385564c3),
	.w2(32'h38c93c2e),
	.w3(32'h38413833),
	.w4(32'h385d5c43),
	.w5(32'h38ba9593),
	.w6(32'h374db098),
	.w7(32'h3769446f),
	.w8(32'h38408747),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807caa2),
	.w1(32'h38732feb),
	.w2(32'h389e43d5),
	.w3(32'h389d57f3),
	.w4(32'h388f81f5),
	.w5(32'h392f596b),
	.w6(32'hb644a193),
	.w7(32'hb830dfad),
	.w8(32'h38710d17),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5553c11),
	.w1(32'h35261027),
	.w2(32'hb59aba2b),
	.w3(32'hb4ca9981),
	.w4(32'h3596203c),
	.w5(32'h330bcda2),
	.w6(32'h358b5421),
	.w7(32'h3620db08),
	.w8(32'h35d8fc26),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d5b7bd),
	.w1(32'h39317e5e),
	.w2(32'h39349d30),
	.w3(32'hb5a7e909),
	.w4(32'h382f7086),
	.w5(32'h38a0f984),
	.w6(32'hb8f1ea4e),
	.w7(32'hb91fb2df),
	.w8(32'hb89b222b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382aa117),
	.w1(32'h3772410a),
	.w2(32'h360b79dc),
	.w3(32'h36f13691),
	.w4(32'hb6d27ceb),
	.w5(32'h376b54e6),
	.w6(32'h366094c1),
	.w7(32'hb7d433f6),
	.w8(32'hb5deb970),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39353d8c),
	.w1(32'h389018ad),
	.w2(32'h383b9e5e),
	.w3(32'h38eef4d2),
	.w4(32'h38600e89),
	.w5(32'h38864bb7),
	.w6(32'h3814b4e1),
	.w7(32'hb809b9da),
	.w8(32'h367e2232),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b0f74a),
	.w1(32'h38c54f99),
	.w2(32'h38cac3ce),
	.w3(32'h38464b1e),
	.w4(32'h386ed893),
	.w5(32'h3838063a),
	.w6(32'h36657edb),
	.w7(32'h37185981),
	.w8(32'h37c1d09a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d85539),
	.w1(32'h38579b7f),
	.w2(32'h38b0ec03),
	.w3(32'h376191a3),
	.w4(32'h37f380b1),
	.w5(32'h38c00b31),
	.w6(32'hb6c49fc3),
	.w7(32'hb6684aae),
	.w8(32'h388bb91a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3594dd48),
	.w1(32'h36c5fbac),
	.w2(32'h369d15ed),
	.w3(32'hb5877c58),
	.w4(32'h36af9707),
	.w5(32'h367b802d),
	.w6(32'h3255e3da),
	.w7(32'h3664c193),
	.w8(32'h36826cbe),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62c3ac7),
	.w1(32'h3602a3aa),
	.w2(32'h365fc690),
	.w3(32'hb6b93da3),
	.w4(32'hb60b9744),
	.w5(32'hb539e512),
	.w6(32'hb68a153b),
	.w7(32'h352459d7),
	.w8(32'hb5773766),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e8e54),
	.w1(32'h391b0801),
	.w2(32'h395e9a19),
	.w3(32'h3966091a),
	.w4(32'h3917e462),
	.w5(32'h3995e4bb),
	.w6(32'h382872d8),
	.w7(32'hb89ea725),
	.w8(32'h38f7f467),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d17439),
	.w1(32'hb739f4cf),
	.w2(32'hb76f6f31),
	.w3(32'h37d6db41),
	.w4(32'hb732629d),
	.w5(32'hb72af7c4),
	.w6(32'h38273d7f),
	.w7(32'hb68230cc),
	.w8(32'h34efc0b5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37254ee9),
	.w1(32'h36b1cb4c),
	.w2(32'h370b03fa),
	.w3(32'hb50a72ac),
	.w4(32'h34f9907d),
	.w5(32'h3609cab8),
	.w6(32'h371f85d6),
	.w7(32'h35e85704),
	.w8(32'h36ceb078),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3813fff9),
	.w1(32'h36dac20b),
	.w2(32'hb7e07af3),
	.w3(32'h380962fb),
	.w4(32'h371b1393),
	.w5(32'hb6b90c5c),
	.w6(32'h37478af0),
	.w7(32'hb79cc9d8),
	.w8(32'hb791d33c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3857773a),
	.w1(32'h378ef191),
	.w2(32'h3858f3ad),
	.w3(32'h3867326c),
	.w4(32'h375a201a),
	.w5(32'h382cfa1d),
	.w6(32'hb6ef3618),
	.w7(32'hb822a737),
	.w8(32'hb77a5703),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3857d532),
	.w1(32'h38044b91),
	.w2(32'h37ebb630),
	.w3(32'h37ca4e2c),
	.w4(32'h370f215a),
	.w5(32'h37acc210),
	.w6(32'hb88947b7),
	.w7(32'hb8fbc596),
	.w8(32'hb89a95d9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb42566cd),
	.w1(32'hb67a463c),
	.w2(32'hb690aa24),
	.w3(32'h3556f4df),
	.w4(32'hb6474070),
	.w5(32'hb673f4c5),
	.w6(32'h356e9696),
	.w7(32'hb61f30ed),
	.w8(32'hb63d4ebd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397651a8),
	.w1(32'h39b1310b),
	.w2(32'h39e43ec3),
	.w3(32'h392cf8e7),
	.w4(32'h39641301),
	.w5(32'h399a2f60),
	.w6(32'h365a3feb),
	.w7(32'h383968e0),
	.w8(32'h3930fa0c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h343870b5),
	.w1(32'hb66600c4),
	.w2(32'hb682a953),
	.w3(32'h3511239a),
	.w4(32'hb625571c),
	.w5(32'hb642343c),
	.w6(32'hb52a6d55),
	.w7(32'hb62b5588),
	.w8(32'hb647e730),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38112a70),
	.w1(32'h36fb5701),
	.w2(32'h380f4be4),
	.w3(32'h385ca8d9),
	.w4(32'h380b85b3),
	.w5(32'h3898df1b),
	.w6(32'h3739c051),
	.w7(32'hb7d803d2),
	.w8(32'h380f73ca),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36600c80),
	.w1(32'h3501c0ef),
	.w2(32'hb6a5bf54),
	.w3(32'h36cc97ee),
	.w4(32'h368f2b84),
	.w5(32'hb6622e69),
	.w6(32'h36a82419),
	.w7(32'h36802001),
	.w8(32'hb50208ba),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361ebf71),
	.w1(32'hb7bcb10d),
	.w2(32'h375e8643),
	.w3(32'h3712484f),
	.w4(32'hb7916422),
	.w5(32'h36fb735f),
	.w6(32'hb7a80623),
	.w7(32'hb89dc9c2),
	.w8(32'hb809f65d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4dc2a61),
	.w1(32'hb476ab04),
	.w2(32'hb50ad175),
	.w3(32'hb49b14f4),
	.w4(32'h33576ae9),
	.w5(32'hb45a70c9),
	.w6(32'h34a72bb2),
	.w7(32'h34dbcb5d),
	.w8(32'h351bc7f4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a931e2),
	.w1(32'h3892839a),
	.w2(32'h38d542c2),
	.w3(32'h3854409d),
	.w4(32'h384d2fbe),
	.w5(32'h389b9290),
	.w6(32'h35c67692),
	.w7(32'h371d7281),
	.w8(32'h38189157),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3391b96a),
	.w1(32'hb4dc7d3e),
	.w2(32'hb58cb9f2),
	.w3(32'h350c2be8),
	.w4(32'h33762441),
	.w5(32'hb51f0846),
	.w6(32'h354da42b),
	.w7(32'h3518db00),
	.w8(32'h34898a41),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956964f),
	.w1(32'h39409d6a),
	.w2(32'h39636ea7),
	.w3(32'h3959ad89),
	.w4(32'h3929d2ee),
	.w5(32'h3977e87c),
	.w6(32'h38a24f7a),
	.w7(32'h37cb7e1e),
	.w8(32'h39027e51),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ea0abe),
	.w1(32'hb7442b1d),
	.w2(32'hb8835dc4),
	.w3(32'hb68d5ec8),
	.w4(32'hb83214df),
	.w5(32'hb8c0e0d6),
	.w6(32'hb81d4851),
	.w7(32'hb8dd3c74),
	.w8(32'hb8d5b8f7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d677af),
	.w1(32'hb55e7bb9),
	.w2(32'h362c00b3),
	.w3(32'h372018ab),
	.w4(32'h34f8072d),
	.w5(32'h3658dd39),
	.w6(32'h37069d6b),
	.w7(32'h35d6346c),
	.w8(32'h3595f8cd),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb547d709),
	.w1(32'hb573fb99),
	.w2(32'hb59b03ee),
	.w3(32'hb5853395),
	.w4(32'hb5596fe1),
	.w5(32'hb54dbba7),
	.w6(32'h33890b91),
	.w7(32'hb2a0dccb),
	.w8(32'h34a3f161),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880a275),
	.w1(32'h37bf8d75),
	.w2(32'h38ba2004),
	.w3(32'h3829da29),
	.w4(32'h380a7331),
	.w5(32'h38a1b337),
	.w6(32'hb82a6db7),
	.w7(32'hb811a587),
	.w8(32'h378cc217),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944d26f),
	.w1(32'h39259794),
	.w2(32'h393778b7),
	.w3(32'h39503f3f),
	.w4(32'h391a5888),
	.w5(32'h395a406d),
	.w6(32'h388d628f),
	.w7(32'h37561b2b),
	.w8(32'h38cba479),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c4bf0),
	.w1(32'h39877a90),
	.w2(32'h399a5d32),
	.w3(32'h39a2d1ac),
	.w4(32'h39113bab),
	.w5(32'h39f8aa0f),
	.w6(32'h39246712),
	.w7(32'hb4bae84b),
	.w8(32'h3997b05f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a11752),
	.w1(32'h39a86aff),
	.w2(32'h39b1643c),
	.w3(32'h3990a9a4),
	.w4(32'h395e6108),
	.w5(32'h399b39fa),
	.w6(32'h38d6766a),
	.w7(32'h35e92157),
	.w8(32'h390e9b10),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b18752),
	.w1(32'h39032f9b),
	.w2(32'h3952da56),
	.w3(32'h37f60a42),
	.w4(32'h38a65237),
	.w5(32'h395733df),
	.w6(32'hb7819acd),
	.w7(32'h3861e973),
	.w8(32'h392f50d9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ad60b5),
	.w1(32'hb61eb39a),
	.w2(32'hb6f2d4e7),
	.w3(32'hb6af5352),
	.w4(32'hb4130c89),
	.w5(32'hb6a693a3),
	.w6(32'h3480c8df),
	.w7(32'h36bc1db8),
	.w8(32'hb40196cf),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a1cd88),
	.w1(32'h34667b6a),
	.w2(32'hb5879fbb),
	.w3(32'hb56afae9),
	.w4(32'h34b9e1b0),
	.w5(32'hb5129b23),
	.w6(32'h34c0021d),
	.w7(32'h35b10eea),
	.w8(32'h35163168),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6334424),
	.w1(32'hb5db7dcf),
	.w2(32'hb5d0e28c),
	.w3(32'hb543ad10),
	.w4(32'h35202992),
	.w5(32'h35b03d59),
	.w6(32'h349fb652),
	.w7(32'h35aa3b1d),
	.w8(32'h35f287e4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3741647e),
	.w1(32'h37d724ae),
	.w2(32'h38111087),
	.w3(32'h37039d7f),
	.w4(32'h37cde6e0),
	.w5(32'h37d7df84),
	.w6(32'hb5a8fdcb),
	.w7(32'h3750a003),
	.w8(32'h37b44e7b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38966b15),
	.w1(32'h3885f5f1),
	.w2(32'h390078a1),
	.w3(32'h38768ae9),
	.w4(32'h3874653f),
	.w5(32'h38bcea68),
	.w6(32'hb81d7bfe),
	.w7(32'hb7b48c70),
	.w8(32'h37ba2f71),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34e9277f),
	.w1(32'hb68d0ba6),
	.w2(32'h371a5f55),
	.w3(32'h36c990dc),
	.w4(32'h366a8173),
	.w5(32'h36a05a2d),
	.w6(32'hb667289e),
	.w7(32'hb64eebef),
	.w8(32'h36864fb3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380c9a2d),
	.w1(32'hb8021206),
	.w2(32'h37b4020b),
	.w3(32'h389fbdd1),
	.w4(32'hb702a859),
	.w5(32'h37a73399),
	.w6(32'h376ec4dc),
	.w7(32'hb86c31d9),
	.w8(32'hb80c6744),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389e03a5),
	.w1(32'h380e8031),
	.w2(32'h38830602),
	.w3(32'h38a20e02),
	.w4(32'h37ca7fcd),
	.w5(32'h389c71d5),
	.w6(32'h38038e60),
	.w7(32'hb7d94f15),
	.w8(32'h37bf5dac),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80589f8),
	.w1(32'hb824c12c),
	.w2(32'hb847824b),
	.w3(32'hb7e6f90a),
	.w4(32'hb84d9402),
	.w5(32'hb84c0edd),
	.w6(32'hb7c8a9af),
	.w7(32'hb8916389),
	.w8(32'hb87fd92f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382d14c8),
	.w1(32'h37dfe8ca),
	.w2(32'h383518ca),
	.w3(32'h380bf69e),
	.w4(32'h365ca939),
	.w5(32'h37df458f),
	.w6(32'hb629443b),
	.w7(32'hb81cc3b9),
	.w8(32'h36d59ffc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39475c01),
	.w1(32'h38d7cb4a),
	.w2(32'h3917a676),
	.w3(32'h3938b3bb),
	.w4(32'h38dbaa78),
	.w5(32'h3918d912),
	.w6(32'h38672acb),
	.w7(32'hb7a0ac7a),
	.w8(32'h38464eee),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb600e775),
	.w1(32'hb5352eaf),
	.w2(32'hb625d9f6),
	.w3(32'hb5df6efe),
	.w4(32'hb4276921),
	.w5(32'hb5eec618),
	.w6(32'hb4bd6f97),
	.w7(32'h35481e13),
	.w8(32'hb54b22d0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fe47c6),
	.w1(32'hb63b0a40),
	.w2(32'hb6df4b2c),
	.w3(32'hb6c94290),
	.w4(32'hb55a082a),
	.w5(32'hb6a7881c),
	.w6(32'hb5f14005),
	.w7(32'h3636945e),
	.w8(32'hb557959f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb631a777),
	.w1(32'hb5689070),
	.w2(32'hb6489b50),
	.w3(32'hb60f94d0),
	.w4(32'h34d043dd),
	.w5(32'hb5d95c4c),
	.w6(32'h34e97245),
	.w7(32'h36149be9),
	.w8(32'h348137f2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dccc5c),
	.w1(32'h368bc34e),
	.w2(32'h36d8f2b6),
	.w3(32'h3663587c),
	.w4(32'h361f4c34),
	.w5(32'h3696ddd4),
	.w6(32'h37197b0a),
	.w7(32'h36d06d29),
	.w8(32'h371d5653),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377f0b6e),
	.w1(32'hb6944035),
	.w2(32'h36310dc9),
	.w3(32'h371bbb21),
	.w4(32'hb7a8fad8),
	.w5(32'hb7ade6c7),
	.w6(32'h3719b597),
	.w7(32'hb7621a1e),
	.w8(32'hb70b08e9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7886a82),
	.w1(32'hb716812d),
	.w2(32'hb6f7489e),
	.w3(32'hb6c9fef3),
	.w4(32'hb6df7329),
	.w5(32'hb6aa6db4),
	.w6(32'hb6ee6e44),
	.w7(32'hb72b4126),
	.w8(32'h33a9b025),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379ff5e4),
	.w1(32'hb7db28de),
	.w2(32'h37a1f950),
	.w3(32'h38063671),
	.w4(32'hb7f714bb),
	.w5(32'h35c1a080),
	.w6(32'hb78e87c1),
	.w7(32'hb8a36999),
	.w8(32'hb8836d04),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80a8c39),
	.w1(32'hb85b0fff),
	.w2(32'hb703296b),
	.w3(32'hb7cf1cd0),
	.w4(32'hb8406df8),
	.w5(32'hb7087717),
	.w6(32'hb8291869),
	.w7(32'hb881bf3b),
	.w8(32'hbb0fad77),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb800764),
	.w1(32'hbaece278),
	.w2(32'hbb480db8),
	.w3(32'h3a83614a),
	.w4(32'h3b1d8e3e),
	.w5(32'h3b448795),
	.w6(32'hb9a298d1),
	.w7(32'h3b32c16c),
	.w8(32'hbb9eb500),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc527d7),
	.w1(32'hbbbc25d7),
	.w2(32'hbc5f45e0),
	.w3(32'h3b5f1ad8),
	.w4(32'hbc73d971),
	.w5(32'hbc77ac05),
	.w6(32'hbc9f264a),
	.w7(32'hbc9d6931),
	.w8(32'h3ab31b8e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e30dc),
	.w1(32'hbacc4f2b),
	.w2(32'hbc0ffe01),
	.w3(32'h39f6b28b),
	.w4(32'hbb6af752),
	.w5(32'hbb68f425),
	.w6(32'hba3ea616),
	.w7(32'hbb102ca9),
	.w8(32'hbc5ce116),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4aa5cb),
	.w1(32'hbb9885f8),
	.w2(32'hbaa063cd),
	.w3(32'hbc01aabb),
	.w4(32'hbb025829),
	.w5(32'h3b2bdcaf),
	.w6(32'hbbb2c4b7),
	.w7(32'h3b20be64),
	.w8(32'hbc89376b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9454b4),
	.w1(32'hbc5d83f1),
	.w2(32'h3c420613),
	.w3(32'hbb5cc534),
	.w4(32'h3b9b6b81),
	.w5(32'h3ca46796),
	.w6(32'hbc88127b),
	.w7(32'h3bf1826d),
	.w8(32'h3c4905ae),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd043083),
	.w1(32'hbd030a01),
	.w2(32'hbc10344a),
	.w3(32'hbc658234),
	.w4(32'hbbe9bc12),
	.w5(32'hbb91cd71),
	.w6(32'hbc27e50e),
	.w7(32'hbc34a967),
	.w8(32'hbc0501f8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a5e25),
	.w1(32'hbbadda8e),
	.w2(32'h3c19bac4),
	.w3(32'hbb06bab0),
	.w4(32'hbb43cb06),
	.w5(32'h3c405f94),
	.w6(32'hbb7f6b73),
	.w7(32'h3c944bd4),
	.w8(32'hbc69705d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fcc9d),
	.w1(32'h3b210f94),
	.w2(32'h3d1981ac),
	.w3(32'h3a5ed519),
	.w4(32'h3c094c4c),
	.w5(32'h3cd8ac4f),
	.w6(32'hbc1ad28b),
	.w7(32'h3c515ff9),
	.w8(32'hbc626ef2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e3f62),
	.w1(32'hbb858733),
	.w2(32'h3a878fc9),
	.w3(32'hbc04c9f1),
	.w4(32'h39d86998),
	.w5(32'h3bb51410),
	.w6(32'hbbbc3d75),
	.w7(32'h3b8d66fa),
	.w8(32'h3a9bac74),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18ed32),
	.w1(32'hb8a6ec01),
	.w2(32'hbbd300e4),
	.w3(32'h392d6175),
	.w4(32'hbb0123b5),
	.w5(32'hbb6029a5),
	.w6(32'h3a20d60f),
	.w7(32'hbb0d9abe),
	.w8(32'h3b36e591),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987eab),
	.w1(32'hbaf39430),
	.w2(32'hbc641bb5),
	.w3(32'h3b03b966),
	.w4(32'hbb9c3eda),
	.w5(32'hbba7b9d7),
	.w6(32'h3681cc81),
	.w7(32'hbb89d9ed),
	.w8(32'hbbf34430),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0ed8c),
	.w1(32'h3c09b025),
	.w2(32'h3b1ceefa),
	.w3(32'h3c77ded6),
	.w4(32'hbc88ffb3),
	.w5(32'hbabd2187),
	.w6(32'hbc84d96f),
	.w7(32'h3b93e2c7),
	.w8(32'hbd190de1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced5a90),
	.w1(32'h3c35c42f),
	.w2(32'h3d433047),
	.w3(32'hbc0ae5b8),
	.w4(32'h3cd5af00),
	.w5(32'h3d2df773),
	.w6(32'hbb5f98a3),
	.w7(32'h3cbc8fe5),
	.w8(32'hbc27546c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c914e),
	.w1(32'hbd15435c),
	.w2(32'h3b2df515),
	.w3(32'hbcc59642),
	.w4(32'hbd00ff2c),
	.w5(32'hbc0a4d8d),
	.w6(32'hbd17ec8c),
	.w7(32'hbbfcbca6),
	.w8(32'h3b3a3f45),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d7224),
	.w1(32'hbb8ac4bc),
	.w2(32'hba081225),
	.w3(32'hb8054131),
	.w4(32'h3b63095c),
	.w5(32'h3b279856),
	.w6(32'h3b12ce9a),
	.w7(32'hbb461d1c),
	.w8(32'hba48300a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6def1),
	.w1(32'h3ae7ab07),
	.w2(32'hbb9337ee),
	.w3(32'hbb87446a),
	.w4(32'hbb3a224b),
	.w5(32'h3bfdc5a4),
	.w6(32'hbad249d8),
	.w7(32'hbbeaba98),
	.w8(32'hbc9e9d92),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf109a),
	.w1(32'hbc9c05ce),
	.w2(32'hbc23eeca),
	.w3(32'h3ba14ea7),
	.w4(32'hbc00edf5),
	.w5(32'hbbe14774),
	.w6(32'hbce13456),
	.w7(32'hbb99e6fa),
	.w8(32'h3c746a4e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f3f02),
	.w1(32'hbacdffcf),
	.w2(32'hbbd89bd9),
	.w3(32'h3c13b9b9),
	.w4(32'hbc4bf70c),
	.w5(32'hbc3925e4),
	.w6(32'hbb9b8053),
	.w7(32'hbba8e8a5),
	.w8(32'hbbaa85a0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2daffb),
	.w1(32'h3b5b8fd7),
	.w2(32'h3c6eac1e),
	.w3(32'h3bac2c96),
	.w4(32'h3bd2f442),
	.w5(32'h3c40f659),
	.w6(32'hbbb99a71),
	.w7(32'h3ab994b8),
	.w8(32'h3b3857e6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe54668),
	.w1(32'hbbec812e),
	.w2(32'hbc5bab5d),
	.w3(32'hba7c58de),
	.w4(32'hbc9ae37a),
	.w5(32'h3c0820ce),
	.w6(32'hbc33f183),
	.w7(32'hbc568711),
	.w8(32'hbc6f222e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65638c),
	.w1(32'hba49f1d1),
	.w2(32'h3b88d396),
	.w3(32'h3bb24c1e),
	.w4(32'h3c579e1e),
	.w5(32'h3cdc4adb),
	.w6(32'hbbb0cc82),
	.w7(32'h3c1a4beb),
	.w8(32'hbc392f94),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfc8f9),
	.w1(32'h39b00dd8),
	.w2(32'hbbc720cb),
	.w3(32'hbb9907df),
	.w4(32'h3acd5c62),
	.w5(32'hbb054d05),
	.w6(32'hbb685b14),
	.w7(32'hbbc09289),
	.w8(32'hbc1673ee),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac962f),
	.w1(32'h3c16463e),
	.w2(32'hbb80e047),
	.w3(32'h3bca315c),
	.w4(32'hbbd77e25),
	.w5(32'hbc1477ec),
	.w6(32'hbc09559a),
	.w7(32'h3a251859),
	.w8(32'hbb8f64b5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule