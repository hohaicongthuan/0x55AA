module layer_10_featuremap_165(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5537bfe),
	.w1(32'hb6b7f16f),
	.w2(32'h366ef1e8),
	.w3(32'hb572428a),
	.w4(32'h36c03243),
	.w5(32'h37532b38),
	.w6(32'hb582199b),
	.w7(32'hb5363a50),
	.w8(32'h33abd04d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e7742c),
	.w1(32'h39aefa5e),
	.w2(32'h394073e3),
	.w3(32'h399e0ddb),
	.w4(32'h39c837e1),
	.w5(32'h394ff109),
	.w6(32'h37e94be3),
	.w7(32'h39201631),
	.w8(32'h386ce811),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fed250),
	.w1(32'h351daef8),
	.w2(32'h369d28ea),
	.w3(32'h36d17658),
	.w4(32'hb6517e58),
	.w5(32'h3642e7f7),
	.w6(32'hb57d4bde),
	.w7(32'h35326423),
	.w8(32'h3693a5a5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68af2c0),
	.w1(32'hb801b2b8),
	.w2(32'hb83121bb),
	.w3(32'hb808e393),
	.w4(32'hb84a6c1b),
	.w5(32'hb86890ea),
	.w6(32'hb8027502),
	.w7(32'hb841b7ff),
	.w8(32'hb8953c5f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f7889a),
	.w1(32'hb881c632),
	.w2(32'hb919c379),
	.w3(32'h38275fda),
	.w4(32'hb7c9c51c),
	.w5(32'hb8f07b0e),
	.w6(32'h3881da0e),
	.w7(32'hb5ff4bf7),
	.w8(32'hb8a07f4e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c00494),
	.w1(32'hb74cb752),
	.w2(32'hb790678b),
	.w3(32'h35ff8f91),
	.w4(32'hb74acb64),
	.w5(32'hb72c082f),
	.w6(32'h38030580),
	.w7(32'h374669e9),
	.w8(32'h36c10aaa),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd90ed),
	.w1(32'h382da635),
	.w2(32'hb704c129),
	.w3(32'hb80a8592),
	.w4(32'h392644f0),
	.w5(32'h38d43831),
	.w6(32'h374e4986),
	.w7(32'h3947bca1),
	.w8(32'h3975e72e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aec610),
	.w1(32'hba014120),
	.w2(32'hba2a35a8),
	.w3(32'hba4769c9),
	.w4(32'hba5d1daf),
	.w5(32'hba66e465),
	.w6(32'hba342b1e),
	.w7(32'hba84b213),
	.w8(32'hba2885ad),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90fc379),
	.w1(32'hb94d543a),
	.w2(32'hb922f110),
	.w3(32'hb869899b),
	.w4(32'hb95d4a26),
	.w5(32'hb96525f5),
	.w6(32'h3715dfca),
	.w7(32'hb96e2fde),
	.w8(32'hb961a29a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba797870),
	.w1(32'hba2d369e),
	.w2(32'hbb0a3075),
	.w3(32'hb906334a),
	.w4(32'hb9cbd7da),
	.w5(32'hbb079c5b),
	.w6(32'h3a0d9a5a),
	.w7(32'h388090d9),
	.w8(32'hbb127213),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa5fc2),
	.w1(32'hb9488c53),
	.w2(32'hb9b8bda1),
	.w3(32'hb848e036),
	.w4(32'hb761b49b),
	.w5(32'hb98808d9),
	.w6(32'hb8b8d6ec),
	.w7(32'hb8615cba),
	.w8(32'hb9798b02),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba082c1f),
	.w1(32'h3a5ce166),
	.w2(32'hb95e9557),
	.w3(32'hba85dc6e),
	.w4(32'h3a2abe15),
	.w5(32'h372fb3b5),
	.w6(32'hba7098f8),
	.w7(32'h3a59dd06),
	.w8(32'h391db489),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14c2c6),
	.w1(32'hba8a5f5c),
	.w2(32'hbb2e3fa8),
	.w3(32'h395fe9ef),
	.w4(32'hba34dc9e),
	.w5(32'hbb3230a5),
	.w6(32'h3a068f20),
	.w7(32'hba1c96c3),
	.w8(32'hbb29cb37),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23b036),
	.w1(32'h3a0e8f8f),
	.w2(32'h38a2a501),
	.w3(32'h3a5028db),
	.w4(32'h3a37d84f),
	.w5(32'h399d320d),
	.w6(32'h3a39c066),
	.w7(32'h3a3e800f),
	.w8(32'h3a00a870),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998ee12),
	.w1(32'hb7c763f7),
	.w2(32'hba623212),
	.w3(32'h3a1208fc),
	.w4(32'h3a46a57c),
	.w5(32'hb9d0c34e),
	.w6(32'h3a0f922b),
	.w7(32'h3a30e256),
	.w8(32'hb9226a58),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cfd61),
	.w1(32'hb9540ea1),
	.w2(32'hba491faf),
	.w3(32'h3960297f),
	.w4(32'hb9221ac7),
	.w5(32'hba83dc9b),
	.w6(32'h399a2ecd),
	.w7(32'hb9a6ace2),
	.w8(32'hbad49a1e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe5c93),
	.w1(32'h37ee38a6),
	.w2(32'hb818a34f),
	.w3(32'hb8f2ea46),
	.w4(32'hb9173584),
	.w5(32'hb9223d41),
	.w6(32'hb9532224),
	.w7(32'hb94b6722),
	.w8(32'hb906b977),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944c805),
	.w1(32'hba2695e8),
	.w2(32'hba92acbc),
	.w3(32'h38fbb696),
	.w4(32'hba104594),
	.w5(32'hbacef9d5),
	.w6(32'hb9b186e1),
	.w7(32'hba46c37b),
	.w8(32'hba8928ea),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c93bbe),
	.w1(32'h3937c8e0),
	.w2(32'hba1553aa),
	.w3(32'h3a6fc12e),
	.w4(32'hb8ffb5bb),
	.w5(32'hbaa2502d),
	.w6(32'h39cb6412),
	.w7(32'hb9e58902),
	.w8(32'hba8073e5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3746bb03),
	.w1(32'h375f3d46),
	.w2(32'h379e5413),
	.w3(32'h36e77b9d),
	.w4(32'h370d3d9e),
	.w5(32'h3776859e),
	.w6(32'h36b1c875),
	.w7(32'h363a8b2f),
	.w8(32'h376ad337),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372a0989),
	.w1(32'h37530167),
	.w2(32'h37cc9670),
	.w3(32'h36f5e908),
	.w4(32'h3704eb03),
	.w5(32'h37ae050e),
	.w6(32'h376618bd),
	.w7(32'h365a84bf),
	.w8(32'h37b8e814),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3941b01f),
	.w1(32'h3a078cb8),
	.w2(32'h393816b5),
	.w3(32'hb8c0a904),
	.w4(32'h39b2e508),
	.w5(32'h39569844),
	.w6(32'hb9823895),
	.w7(32'h39456893),
	.w8(32'h37ef384d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa5a6b),
	.w1(32'hb9677a98),
	.w2(32'hbb3ca0fb),
	.w3(32'hb9e4b89f),
	.w4(32'h3a5a4c2b),
	.w5(32'hbb412e72),
	.w6(32'h39b49cfb),
	.w7(32'h3a78e715),
	.w8(32'hbb61c82e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38d134),
	.w1(32'hb9d6c6af),
	.w2(32'hbac80281),
	.w3(32'h389bf8ad),
	.w4(32'h38884cfa),
	.w5(32'hbae0e187),
	.w6(32'h3912d365),
	.w7(32'hb79ed8eb),
	.w8(32'hbaf6c004),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4be032),
	.w1(32'hb9ba9b1f),
	.w2(32'hbac1b6e1),
	.w3(32'hb9ca7310),
	.w4(32'hb82d511b),
	.w5(32'hbaa33c81),
	.w6(32'hba65569b),
	.w7(32'hb9f76060),
	.w8(32'hbacd3886),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ed78e),
	.w1(32'hb787f2bb),
	.w2(32'hb97b6d55),
	.w3(32'h3803de28),
	.w4(32'h3814cb5f),
	.w5(32'hb9a3fdf2),
	.w6(32'h38388a9e),
	.w7(32'h38a76524),
	.w8(32'hb9a310cf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372dc771),
	.w1(32'h37cb91e2),
	.w2(32'h383eb78d),
	.w3(32'h3473c22e),
	.w4(32'h374e87bd),
	.w5(32'h384ac9b6),
	.w6(32'hb65b3706),
	.w7(32'h37b6a1f9),
	.w8(32'h3854c325),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ed0a2),
	.w1(32'h3995f5ed),
	.w2(32'h38ab47c5),
	.w3(32'h39395f97),
	.w4(32'h39b64f46),
	.w5(32'h388b18a3),
	.w6(32'h372d2bf1),
	.w7(32'h39b96eeb),
	.w8(32'h38d3a9ef),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0691ec),
	.w1(32'h3a11153c),
	.w2(32'h399de99b),
	.w3(32'hba4415ca),
	.w4(32'h39c94e34),
	.w5(32'h393c20b4),
	.w6(32'hba5b975b),
	.w7(32'h39c94d62),
	.w8(32'h39360e03),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc7dee),
	.w1(32'hb9b56208),
	.w2(32'hba8d27e6),
	.w3(32'h3947fe48),
	.w4(32'hb89bacac),
	.w5(32'hbaa988a7),
	.w6(32'h3a127acc),
	.w7(32'h38ccf9a2),
	.w8(32'hbacc02ef),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7187655),
	.w1(32'h36c8ea7a),
	.w2(32'h362e6fd9),
	.w3(32'hb776fceb),
	.w4(32'h35c51de2),
	.w5(32'hb596b92c),
	.w6(32'h3564cbae),
	.w7(32'hb62d5604),
	.w8(32'hb650ca1a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb600def6),
	.w1(32'h37335c69),
	.w2(32'h38192550),
	.w3(32'hb5bb9c85),
	.w4(32'h36891cb7),
	.w5(32'h37ad164b),
	.w6(32'h37a4258c),
	.w7(32'h3799236d),
	.w8(32'h37f291e6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9c3ff),
	.w1(32'hb9a3e164),
	.w2(32'hba397edd),
	.w3(32'h3883dbab),
	.w4(32'hb84aa0ec),
	.w5(32'hba5542f3),
	.w6(32'h38f4f8a1),
	.w7(32'h37720834),
	.w8(32'hba5c6871),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9104706),
	.w1(32'h37bea6ec),
	.w2(32'hb9cb945d),
	.w3(32'hb820512c),
	.w4(32'h391607cb),
	.w5(32'hb955e20e),
	.w6(32'hb8f1e10a),
	.w7(32'h38e0cbbf),
	.w8(32'hb97e8cef),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883a24b),
	.w1(32'hb8468c3b),
	.w2(32'hb7b0087e),
	.w3(32'hb8c64f63),
	.w4(32'hb8ee39e8),
	.w5(32'hb91eb9c4),
	.w6(32'h374edadd),
	.w7(32'hb8488663),
	.w8(32'hb88d59be),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9942d97),
	.w1(32'hb93f8fbb),
	.w2(32'hb958fca3),
	.w3(32'hb91c0883),
	.w4(32'hb8881d82),
	.w5(32'hb8baabe3),
	.w6(32'hb8a52c1e),
	.w7(32'hb8ae8084),
	.w8(32'hb8cd9ea4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8c2e2),
	.w1(32'h398f175d),
	.w2(32'hba29691e),
	.w3(32'hb9a7e43a),
	.w4(32'h398dafa1),
	.w5(32'hba501634),
	.w6(32'hb7dc51b7),
	.w7(32'h39fc5f54),
	.w8(32'hbaa6518a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18ad02),
	.w1(32'h3a8bb40c),
	.w2(32'hb9f48c7b),
	.w3(32'hbab7f36e),
	.w4(32'h3a3f7dc5),
	.w5(32'hb98cd81e),
	.w6(32'hbb284507),
	.w7(32'h3a2b908c),
	.w8(32'hb95bba46),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba775ac9),
	.w1(32'h3a00c7f3),
	.w2(32'hba42e22b),
	.w3(32'hbb0c6728),
	.w4(32'hba4f7fe9),
	.w5(32'hba616a1c),
	.w6(32'hbb322c77),
	.w7(32'hba601136),
	.w8(32'hbaa420a1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c14ca),
	.w1(32'hb9910ea5),
	.w2(32'h37dfdb35),
	.w3(32'hb9b411a5),
	.w4(32'h37b93107),
	.w5(32'h39b8bc7b),
	.w6(32'hb8c6fa08),
	.w7(32'h3949a5c2),
	.w8(32'h3a174d47),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383e9cd8),
	.w1(32'h381f8be8),
	.w2(32'h37734780),
	.w3(32'h3817a465),
	.w4(32'h37ba3e69),
	.w5(32'h37476100),
	.w6(32'h388a46ce),
	.w7(32'hb65b6a3a),
	.w8(32'h3840006a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a6446b),
	.w1(32'h362b4610),
	.w2(32'h38101e18),
	.w3(32'hb8378d75),
	.w4(32'hb7cd711f),
	.w5(32'h380435d6),
	.w6(32'hb7bf2c72),
	.w7(32'hb765147a),
	.w8(32'h37f0fac9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78bd812),
	.w1(32'h3a91f30b),
	.w2(32'h39dddf8a),
	.w3(32'hb90534df),
	.w4(32'h3a634011),
	.w5(32'h38c4d249),
	.w6(32'h38dcbcfb),
	.w7(32'h3aa81ac9),
	.w8(32'hb9dab85c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f1372),
	.w1(32'hb9f84782),
	.w2(32'hba9e7e22),
	.w3(32'h399c8e92),
	.w4(32'hb9668ec0),
	.w5(32'hbaa59466),
	.w6(32'h3a6d97a8),
	.w7(32'hba02bff3),
	.w8(32'hbb0532c8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed422c),
	.w1(32'hb95c58e2),
	.w2(32'hbaab61f2),
	.w3(32'h39c8956c),
	.w4(32'h39b30dd4),
	.w5(32'hbab47190),
	.w6(32'h39e3d826),
	.w7(32'h39c3f04f),
	.w8(32'hbac7dbaf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b0b75),
	.w1(32'hb9e29a3d),
	.w2(32'hbaf96ade),
	.w3(32'h38a32196),
	.w4(32'h39860b6a),
	.w5(32'hbafeeb43),
	.w6(32'h3947cde6),
	.w7(32'h391bfe8c),
	.w8(32'hbb11fe25),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7676c),
	.w1(32'hb9067b5e),
	.w2(32'hba6bfd6a),
	.w3(32'hb8c830dd),
	.w4(32'h38afc51a),
	.w5(32'hba48a455),
	.w6(32'hb8cc7811),
	.w7(32'h39169a97),
	.w8(32'hba697f4f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fc0d2a),
	.w1(32'hbaadfd9e),
	.w2(32'hbb0f59d2),
	.w3(32'h37593d03),
	.w4(32'hbae1c188),
	.w5(32'hbb31d5fd),
	.w6(32'hb9c62029),
	.w7(32'hbb0884d7),
	.w8(32'hbb490a30),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81a4304),
	.w1(32'h3566ea9d),
	.w2(32'h38244453),
	.w3(32'hb88be3d3),
	.w4(32'h372cc011),
	.w5(32'h385c4fa8),
	.w6(32'hb78d47c7),
	.w7(32'hb4c556cf),
	.w8(32'h381446a6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38930ff7),
	.w1(32'hb7865e14),
	.w2(32'hb9649d92),
	.w3(32'h37c9a1eb),
	.w4(32'h38e8ca82),
	.w5(32'hb91ae30a),
	.w6(32'h39582e40),
	.w7(32'h388fbfc4),
	.w8(32'hb72165db),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb865e07c),
	.w1(32'hb88f6983),
	.w2(32'h383904a0),
	.w3(32'hb8042a18),
	.w4(32'hb8d5540c),
	.w5(32'hb74356fb),
	.w6(32'h37dae9af),
	.w7(32'hb83e6b72),
	.w8(32'h36493d79),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00a60d),
	.w1(32'h396da7ee),
	.w2(32'hba23d237),
	.w3(32'hb8fd4ea5),
	.w4(32'h39d8047b),
	.w5(32'hba5307d0),
	.w6(32'hb9717f3b),
	.w7(32'h396591f1),
	.w8(32'hba7156eb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb871c813),
	.w1(32'hb801c5f9),
	.w2(32'hb933cec9),
	.w3(32'h389a51ff),
	.w4(32'h38e115d6),
	.w5(32'hb909f286),
	.w6(32'h394324cc),
	.w7(32'h38f30cf3),
	.w8(32'hb89a4053),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b8b6b),
	.w1(32'hba600d9f),
	.w2(32'hbaec93f2),
	.w3(32'h3a79eb71),
	.w4(32'hb9b06e37),
	.w5(32'hbae6b61d),
	.w6(32'h39cbb640),
	.w7(32'hb976339c),
	.w8(32'hba87495a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba864c),
	.w1(32'h3903a7f0),
	.w2(32'hb79fa762),
	.w3(32'hb7b19eea),
	.w4(32'h388f7de6),
	.w5(32'hb721c368),
	.w6(32'hb8ab5887),
	.w7(32'h3895cf6e),
	.w8(32'h37b3999f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c4bfe6),
	.w1(32'h341d1728),
	.w2(32'hb858cd9b),
	.w3(32'h37dda7a2),
	.w4(32'hb7b24845),
	.w5(32'hb8bed9e4),
	.w6(32'h3852ac5a),
	.w7(32'hb8172dc8),
	.w8(32'hb8d5c4a7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c9a206),
	.w1(32'h375078c5),
	.w2(32'h373c8a6a),
	.w3(32'hb789c550),
	.w4(32'h36acbb1e),
	.w5(32'h36c523c6),
	.w6(32'h375dda99),
	.w7(32'h37055258),
	.w8(32'h3795de32),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3684df6e),
	.w1(32'hb771b519),
	.w2(32'hb7352f1e),
	.w3(32'hb6abd817),
	.w4(32'hb79487c6),
	.w5(32'hb6fa150f),
	.w6(32'hb638ecb3),
	.w7(32'hb58acda3),
	.w8(32'hb592b480),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb9a44),
	.w1(32'h398f58bc),
	.w2(32'hb82146f7),
	.w3(32'hb9a55138),
	.w4(32'h391dce15),
	.w5(32'hb88ce46c),
	.w6(32'hb9ab5504),
	.w7(32'h392b295d),
	.w8(32'hb91cfcb4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ed3a01),
	.w1(32'h38748a6b),
	.w2(32'h38cc93e7),
	.w3(32'hb862c509),
	.w4(32'h3833eb0d),
	.w5(32'h35f5cb4f),
	.w6(32'hb8c0e084),
	.w7(32'h37dfc493),
	.w8(32'hb800b13c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ecb8f),
	.w1(32'hb99b9169),
	.w2(32'hb92b8a22),
	.w3(32'hb9624c14),
	.w4(32'hb9075024),
	.w5(32'h3760c5eb),
	.w6(32'hb92df495),
	.w7(32'hba28972c),
	.w8(32'hba289f6f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb22dc),
	.w1(32'hb7ecbb7d),
	.w2(32'h38b0481a),
	.w3(32'hb9139585),
	.w4(32'hb6c1d195),
	.w5(32'hb8bcabc7),
	.w6(32'hb97f1a99),
	.w7(32'h38e8be5e),
	.w8(32'hb982b40e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37847e5b),
	.w1(32'hb6d9c188),
	.w2(32'h3747e494),
	.w3(32'h3784cb13),
	.w4(32'h369c7aa2),
	.w5(32'h379ff4f2),
	.w6(32'h3617759c),
	.w7(32'hb6a4eb63),
	.w8(32'h33ed1568),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb676b4aa),
	.w1(32'hb6c453b5),
	.w2(32'h376e0210),
	.w3(32'h3733fa7c),
	.w4(32'hb75ff870),
	.w5(32'h3506ad6b),
	.w6(32'hb69efa1a),
	.w7(32'hb6c6d86c),
	.w8(32'h372b70fe),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803dd76),
	.w1(32'hb6200e99),
	.w2(32'h38a784f4),
	.w3(32'h38a56cfd),
	.w4(32'h383c5a3f),
	.w5(32'h3896d530),
	.w6(32'h3894f124),
	.w7(32'h3889fe89),
	.w8(32'h38c6b164),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379bbc6e),
	.w1(32'h3786078c),
	.w2(32'h37b6a165),
	.w3(32'h371ab7e0),
	.w4(32'h368c78f9),
	.w5(32'h37b676e0),
	.w6(32'h377585ff),
	.w7(32'h378f24e5),
	.w8(32'h37ec0776),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8917829),
	.w1(32'hb9d05509),
	.w2(32'hb9110aba),
	.w3(32'h39bc845f),
	.w4(32'h397be299),
	.w5(32'hb893b45c),
	.w6(32'hba0960a9),
	.w7(32'hb9f25901),
	.w8(32'hba251106),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93df5cd),
	.w1(32'h391bc33f),
	.w2(32'hbaba5184),
	.w3(32'hb5072a73),
	.w4(32'h39c01668),
	.w5(32'hbab0817b),
	.w6(32'hb9b4506b),
	.w7(32'h387f7ce7),
	.w8(32'hbacd6522),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba833f7d),
	.w1(32'hb9820088),
	.w2(32'hbaa7f515),
	.w3(32'hba72de84),
	.w4(32'h388d70da),
	.w5(32'hba6334b8),
	.w6(32'hba909926),
	.w7(32'hb6c8dae3),
	.w8(32'hba5757c2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993435c),
	.w1(32'h39915677),
	.w2(32'hbaf8ebd1),
	.w3(32'h39ddbfc7),
	.w4(32'h3a51e4e8),
	.w5(32'hbacbc19a),
	.w6(32'hb90afaa6),
	.w7(32'h39e756e2),
	.w8(32'hbae9cdbe),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7819eb4),
	.w1(32'h37057b97),
	.w2(32'h37e9bbe8),
	.w3(32'hb7cb7faa),
	.w4(32'h35004f08),
	.w5(32'h3794e5ed),
	.w6(32'h36c3ae51),
	.w7(32'h37020da8),
	.w8(32'h379fcedc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3784e0db),
	.w1(32'h368ec55e),
	.w2(32'h384dd82a),
	.w3(32'h37543229),
	.w4(32'hb4b64394),
	.w5(32'h38402e1a),
	.w6(32'h37834f3b),
	.w7(32'h3745bcc4),
	.w8(32'h384d1c66),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37335031),
	.w1(32'hb68a55a9),
	.w2(32'h37f03286),
	.w3(32'h37cf6c2f),
	.w4(32'hb69fdcf5),
	.w5(32'h37cf883e),
	.w6(32'h37962733),
	.w7(32'hb6965666),
	.w8(32'h3749c8ce),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f06b8),
	.w1(32'h37c086cc),
	.w2(32'h388f07f2),
	.w3(32'hb95016f5),
	.w4(32'hb7dd3cbe),
	.w5(32'h3949cdcc),
	.w6(32'hb95ef892),
	.w7(32'hb8ac714e),
	.w8(32'h3933968d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370d5d7f),
	.w1(32'h36151f59),
	.w2(32'h37ab3940),
	.w3(32'hb6d2b671),
	.w4(32'hb69ef514),
	.w5(32'h37a2002c),
	.w6(32'hb66c9ecc),
	.w7(32'hb587dbaf),
	.w8(32'h37fecc25),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85845ec),
	.w1(32'hb971e411),
	.w2(32'h37de51bc),
	.w3(32'hb8554f36),
	.w4(32'hb94d507d),
	.w5(32'hb80c555d),
	.w6(32'hb99e81ed),
	.w7(32'hb9c3f55c),
	.w8(32'h397b5616),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e4c03),
	.w1(32'hb98b184b),
	.w2(32'hb9afb220),
	.w3(32'h39cfae9a),
	.w4(32'hb9702835),
	.w5(32'hba03cdb3),
	.w6(32'h393d6952),
	.w7(32'hba41d75d),
	.w8(32'hba7415e9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1cbb3),
	.w1(32'hb9f5626d),
	.w2(32'hbac9ad6e),
	.w3(32'hb96d3e5e),
	.w4(32'hb9da024e),
	.w5(32'hbaf74f9f),
	.w6(32'hb9423f78),
	.w7(32'hba7f6af0),
	.w8(32'hbb145fe4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9709af8),
	.w1(32'hb89a3d4a),
	.w2(32'hba75f09c),
	.w3(32'h3955e2da),
	.w4(32'h38f3b231),
	.w5(32'hba716f66),
	.w6(32'h37ef4d41),
	.w7(32'hb7a65e01),
	.w8(32'hba617612),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c36cc),
	.w1(32'h37580996),
	.w2(32'hb9962763),
	.w3(32'h396ac897),
	.w4(32'h38d1870f),
	.w5(32'hba0666f9),
	.w6(32'h39754295),
	.w7(32'h38a1b675),
	.w8(32'hba0b44d0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e5e1a),
	.w1(32'h38dfa124),
	.w2(32'hb9dabdd4),
	.w3(32'hb7c5541f),
	.w4(32'h39551b34),
	.w5(32'hb9f38197),
	.w6(32'h39b49157),
	.w7(32'h39bd1541),
	.w8(32'hba052993),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f4d8a7),
	.w1(32'hb9dce006),
	.w2(32'hba4530fc),
	.w3(32'hb963ad42),
	.w4(32'hb9ff86db),
	.w5(32'hba85b267),
	.w6(32'hb967c921),
	.w7(32'hba1c6724),
	.w8(32'hba92b258),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb730bd2d),
	.w1(32'h365c43e3),
	.w2(32'h37886f46),
	.w3(32'hb616343d),
	.w4(32'h36b15e18),
	.w5(32'h37882b9b),
	.w6(32'h375d0749),
	.w7(32'h37142b95),
	.w8(32'h37b73b02),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36da3ebb),
	.w1(32'h3707fdf3),
	.w2(32'h3781f6c7),
	.w3(32'hb670e016),
	.w4(32'h35d51eb6),
	.w5(32'h3795aa42),
	.w6(32'h362f052f),
	.w7(32'h3739ea83),
	.w8(32'h37cc220f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6066d97),
	.w1(32'h381edb5b),
	.w2(32'h36ec01ab),
	.w3(32'h373df8a7),
	.w4(32'h37ce1e2f),
	.w5(32'hb744ac74),
	.w6(32'h38284749),
	.w7(32'h370d4f94),
	.w8(32'hb53cd1ce),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3695dc3e),
	.w1(32'h36a21f79),
	.w2(32'h36b08389),
	.w3(32'hb788ed83),
	.w4(32'h35e786b4),
	.w5(32'h3600e27e),
	.w6(32'h3697a54f),
	.w7(32'h35b70be4),
	.w8(32'h36ff8c61),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cd559),
	.w1(32'hb8fdd773),
	.w2(32'hb9c46094),
	.w3(32'hba673c77),
	.w4(32'h39204c81),
	.w5(32'h39185cb9),
	.w6(32'h38d3b1f3),
	.w7(32'h3a86e4bf),
	.w8(32'h3a45a509),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b5480),
	.w1(32'h39d4b1ab),
	.w2(32'h38a30dec),
	.w3(32'hb762329d),
	.w4(32'h38cd61c9),
	.w5(32'hb8b82fdc),
	.w6(32'hb89c2531),
	.w7(32'h393f6686),
	.w8(32'hb87eee5b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0150d),
	.w1(32'h3901d120),
	.w2(32'hb98d8451),
	.w3(32'h39ee2bb0),
	.w4(32'h3a13a7fc),
	.w5(32'hb9aa9f55),
	.w6(32'h3a5b0c4e),
	.w7(32'h3a11daaa),
	.w8(32'hba027d41),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a5f8c),
	.w1(32'hba19ab12),
	.w2(32'hba82960e),
	.w3(32'hba0f8afe),
	.w4(32'hba2e83df),
	.w5(32'hba7c50b8),
	.w6(32'hba8a60aa),
	.w7(32'hba8876f5),
	.w8(32'hba87bebb),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a66a6),
	.w1(32'h3a00506e),
	.w2(32'hba158863),
	.w3(32'hba42ea0e),
	.w4(32'hb8671a66),
	.w5(32'hba017bc3),
	.w6(32'hba4bdcc9),
	.w7(32'h39aefd90),
	.w8(32'hb9a271e2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82f73b),
	.w1(32'hbaa17c62),
	.w2(32'hbb0c1539),
	.w3(32'hb9cbc88b),
	.w4(32'hba6a28f8),
	.w5(32'hbafa6016),
	.w6(32'h39b845da),
	.w7(32'hb9810f3d),
	.w8(32'hbad1420c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907fe40),
	.w1(32'h381c4ec8),
	.w2(32'hb9b35b4d),
	.w3(32'h39bfb54f),
	.w4(32'h39e78893),
	.w5(32'hb7898bba),
	.w6(32'h3998086d),
	.w7(32'h3a005255),
	.w8(32'h39ec29c8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba108610),
	.w1(32'hb8c2aa84),
	.w2(32'hbaaf0b9c),
	.w3(32'h3a5d2176),
	.w4(32'h3aa89a4f),
	.w5(32'hb969ce57),
	.w6(32'h3aab81cb),
	.w7(32'h3acf15c8),
	.w8(32'h39cd35ce),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c8655),
	.w1(32'h38d7f919),
	.w2(32'h33f1ebae),
	.w3(32'h362bcd95),
	.w4(32'h396ea32b),
	.w5(32'h39b8be0f),
	.w6(32'h3a389d48),
	.w7(32'h3a3a0bde),
	.w8(32'h3a14ad9e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22e5a6),
	.w1(32'hba0afb00),
	.w2(32'hba7c2ccc),
	.w3(32'hb978776b),
	.w4(32'hb6022414),
	.w5(32'hba3715c7),
	.w6(32'hb8942631),
	.w7(32'h387ab520),
	.w8(32'hb9849f59),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e43475),
	.w1(32'hb8e4b73f),
	.w2(32'hb901f2d4),
	.w3(32'h39065bbb),
	.w4(32'hb99968aa),
	.w5(32'hb80e0616),
	.w6(32'h3894ad94),
	.w7(32'hb99b4d94),
	.w8(32'hb88aa952),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cbc5f),
	.w1(32'hba280d3c),
	.w2(32'hbae3f402),
	.w3(32'h39a7c876),
	.w4(32'h391b6a1a),
	.w5(32'hbb08fa67),
	.w6(32'h3992419b),
	.w7(32'hb8f32f00),
	.w8(32'hbaf3e048),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67b08e),
	.w1(32'hb8d5c038),
	.w2(32'hb9d911ea),
	.w3(32'hba923ee5),
	.w4(32'h39ab263c),
	.w5(32'h3936acb6),
	.w6(32'hb91c327f),
	.w7(32'h3a443bdd),
	.w8(32'h37119ab2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3812f0),
	.w1(32'h3aae9d10),
	.w2(32'h3946fc76),
	.w3(32'h39f51b1f),
	.w4(32'h3a00da2f),
	.w5(32'hb8f4dae8),
	.w6(32'hba4de23d),
	.w7(32'hba3b72df),
	.w8(32'hb98030da),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac05e16),
	.w1(32'h39ed0687),
	.w2(32'hba435c51),
	.w3(32'hbb7b703c),
	.w4(32'h3acc5245),
	.w5(32'h39a79894),
	.w6(32'h3a25a380),
	.w7(32'h3b8fb4b9),
	.w8(32'h3a6dd385),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b21d6),
	.w1(32'hba0a8cf0),
	.w2(32'hbab8a995),
	.w3(32'h397ad585),
	.w4(32'h36c22509),
	.w5(32'hbae53efc),
	.w6(32'h3a2b96ef),
	.w7(32'hb8c12b6a),
	.w8(32'hbb0ef83c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba344722),
	.w1(32'hb9f4a15e),
	.w2(32'hba924e78),
	.w3(32'hb9388476),
	.w4(32'hb8b3dd59),
	.w5(32'hba04e693),
	.w6(32'h3aa8538e),
	.w7(32'h3a595c79),
	.w8(32'hba1eee84),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb966337c),
	.w1(32'hb949ab07),
	.w2(32'h3940bb63),
	.w3(32'hb94cb8f5),
	.w4(32'hb8dea64f),
	.w5(32'h38b15715),
	.w6(32'hb7e2ab7c),
	.w7(32'h38819fad),
	.w8(32'h389e65c2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba378983),
	.w1(32'hb9f27075),
	.w2(32'hbaa64601),
	.w3(32'hb9d8b813),
	.w4(32'hba106ee2),
	.w5(32'hba5360bb),
	.w6(32'hba0c01b3),
	.w7(32'hba43d91b),
	.w8(32'hba207201),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8fd9d),
	.w1(32'h39db4c9a),
	.w2(32'hb909d8ed),
	.w3(32'hb94ddab4),
	.w4(32'h3a43e245),
	.w5(32'hb8d36024),
	.w6(32'h38af5816),
	.w7(32'h39ff4c0d),
	.w8(32'h36eedab5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351111bb),
	.w1(32'h36622122),
	.w2(32'hb82cc252),
	.w3(32'hb80c7085),
	.w4(32'hb81edd22),
	.w5(32'hb89e0834),
	.w6(32'hb68a19ce),
	.w7(32'h37fe1482),
	.w8(32'hb70daf5b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8754714),
	.w1(32'hb7cb8670),
	.w2(32'hb800bac1),
	.w3(32'hb883536d),
	.w4(32'hb888b73a),
	.w5(32'hb8799f94),
	.w6(32'hb8c165b7),
	.w7(32'hb7f5d368),
	.w8(32'hb837416f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba362d78),
	.w1(32'hba4327b2),
	.w2(32'hbaac080d),
	.w3(32'hb93eea40),
	.w4(32'hba43c358),
	.w5(32'hbad433d3),
	.w6(32'h3987a805),
	.w7(32'hba747836),
	.w8(32'hbb0b9ecd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbba7b),
	.w1(32'hb7477ab1),
	.w2(32'hba306855),
	.w3(32'h39b74c69),
	.w4(32'h39af46f4),
	.w5(32'hba613216),
	.w6(32'h39e133ef),
	.w7(32'h395f3af9),
	.w8(32'hbaa1020b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d140ff),
	.w1(32'h38b9094b),
	.w2(32'hb9706829),
	.w3(32'h39a273d8),
	.w4(32'h3a869f69),
	.w5(32'hb879dacd),
	.w6(32'h3a0a3718),
	.w7(32'h3a3b4f34),
	.w8(32'hb99c4646),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9935395),
	.w1(32'h39a8962f),
	.w2(32'hb9c35867),
	.w3(32'hb92891c6),
	.w4(32'h39461ada),
	.w5(32'hba088c79),
	.w6(32'hb79d16c8),
	.w7(32'h378f7c72),
	.w8(32'hba247888),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f4ed5),
	.w1(32'h3968124e),
	.w2(32'hb9b96148),
	.w3(32'hb9a777e9),
	.w4(32'h391dff1c),
	.w5(32'hb933edc4),
	.w6(32'hb9c0123c),
	.w7(32'h38b7ff62),
	.w8(32'hb9c03e06),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7b0c6),
	.w1(32'hb9c2b203),
	.w2(32'hba64fd0b),
	.w3(32'hb92908b5),
	.w4(32'hb98abf30),
	.w5(32'hba8b1406),
	.w6(32'hb7dd06b3),
	.w7(32'hb986e093),
	.w8(32'hbaa0d38d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b9b81),
	.w1(32'hb88ff7f6),
	.w2(32'hba748be3),
	.w3(32'h392fa3bf),
	.w4(32'h38986fd5),
	.w5(32'hba75906c),
	.w6(32'h39585490),
	.w7(32'hb8195fe7),
	.w8(32'hba8cb38f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8caf8fe),
	.w1(32'hb7a2b786),
	.w2(32'hb79ae991),
	.w3(32'hb88b2b85),
	.w4(32'hb7ae1b59),
	.w5(32'hb7cbd6b9),
	.w6(32'hb82e3fe1),
	.w7(32'hb7ca2f60),
	.w8(32'hb78699fc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c58b75),
	.w1(32'h3274403b),
	.w2(32'h370ba102),
	.w3(32'hb507f96b),
	.w4(32'hb6e92ee0),
	.w5(32'h350ec095),
	.w6(32'hb6d713b1),
	.w7(32'hb6d09862),
	.w8(32'h36894f0d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb851c6b5),
	.w1(32'h37fcb047),
	.w2(32'h370d1a2d),
	.w3(32'hb84acb5f),
	.w4(32'h3837c533),
	.w5(32'h37583e56),
	.w6(32'hb8068336),
	.w7(32'h382440a7),
	.w8(32'h383b0039),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b3f0a),
	.w1(32'h39166677),
	.w2(32'hb78b9a93),
	.w3(32'h392ead8e),
	.w4(32'h390360cd),
	.w5(32'h388b6ee9),
	.w6(32'h38839aa0),
	.w7(32'h37d3eecb),
	.w8(32'h377da981),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2a035),
	.w1(32'hb890a641),
	.w2(32'hba057946),
	.w3(32'h389d286a),
	.w4(32'h39d60cb5),
	.w5(32'hba530d3e),
	.w6(32'h3a0dccf2),
	.w7(32'h39d3cdf7),
	.w8(32'hba685440),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e45c97),
	.w1(32'hb9152a0a),
	.w2(32'hb9f3b31f),
	.w3(32'h38c3da80),
	.w4(32'hb7a51dda),
	.w5(32'hb9974427),
	.w6(32'h3936e635),
	.w7(32'hb83b5416),
	.w8(32'hb92da9bd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c7d8a),
	.w1(32'hb9b85679),
	.w2(32'hba264139),
	.w3(32'hb96838d3),
	.w4(32'hb9bfc978),
	.w5(32'hba31dd48),
	.w6(32'h399d611a),
	.w7(32'hb94da42f),
	.w8(32'hba088470),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6514133),
	.w1(32'h3a1c50a0),
	.w2(32'hb8da143e),
	.w3(32'hb82115fa),
	.w4(32'h3a059ae1),
	.w5(32'hb97474ae),
	.w6(32'hb8db7158),
	.w7(32'hb979ce2a),
	.w8(32'hba06a8fe),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f58d65),
	.w1(32'h373aeaa7),
	.w2(32'hb6f7dda2),
	.w3(32'h37cba395),
	.w4(32'h3723d4f8),
	.w5(32'h37b4acf9),
	.w6(32'h38188b86),
	.w7(32'h3648014d),
	.w8(32'h378fc1ce),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dac193),
	.w1(32'h393e67a7),
	.w2(32'h390288b7),
	.w3(32'h38608826),
	.w4(32'h37e6b5e3),
	.w5(32'h38a768d5),
	.w6(32'hb896bd22),
	.w7(32'hb8467c99),
	.w8(32'h38312eee),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cc8b06),
	.w1(32'h3716fb3e),
	.w2(32'h37878aca),
	.w3(32'h36172e78),
	.w4(32'h35e58ca2),
	.w5(32'h372693c1),
	.w6(32'h36d89b58),
	.w7(32'h3670fb3d),
	.w8(32'h3743c367),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c403a),
	.w1(32'h399a0538),
	.w2(32'h37b6ee0d),
	.w3(32'h395157ae),
	.w4(32'h39aed240),
	.w5(32'h36bea01e),
	.w6(32'h393737a8),
	.w7(32'h39c4cd98),
	.w8(32'hb7149d3e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39746522),
	.w1(32'h3a2d208d),
	.w2(32'h3927765b),
	.w3(32'h387da83a),
	.w4(32'h3a1a2b46),
	.w5(32'hb891f98c),
	.w6(32'h3839b0c0),
	.w7(32'h39c98892),
	.w8(32'hb85e7a94),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379e52a2),
	.w1(32'hba90853c),
	.w2(32'hba83abc4),
	.w3(32'h3a37abe1),
	.w4(32'hb9e0b247),
	.w5(32'hbad5e1d2),
	.w6(32'h38117448),
	.w7(32'hba97df23),
	.w8(32'hba8ca964),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8639ede),
	.w1(32'h3690b6a2),
	.w2(32'hb91777c7),
	.w3(32'hba32838d),
	.w4(32'hb5de8588),
	.w5(32'hb91d1f17),
	.w6(32'h38afb43b),
	.w7(32'hb90faa15),
	.w8(32'h37f19ea2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38850d54),
	.w1(32'hba02862b),
	.w2(32'hba20dfb6),
	.w3(32'hb6ce941f),
	.w4(32'hb9cc227a),
	.w5(32'hb9e79f02),
	.w6(32'hba207be2),
	.w7(32'hba07437e),
	.w8(32'hba00e3fd),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10809f),
	.w1(32'h3a38e7ef),
	.w2(32'h3a16502f),
	.w3(32'hb98c407b),
	.w4(32'h399786fc),
	.w5(32'hb8867351),
	.w6(32'hba457e98),
	.w7(32'hba5cba19),
	.w8(32'hb9c22182),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1c5bb),
	.w1(32'hb89e26eb),
	.w2(32'hba40065b),
	.w3(32'h38eb1a21),
	.w4(32'hb8d57584),
	.w5(32'hba479f0c),
	.w6(32'hb98df2ef),
	.w7(32'h387d453e),
	.w8(32'hba2df52d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38973a26),
	.w1(32'h3a3697da),
	.w2(32'h39ca98bd),
	.w3(32'h393f8955),
	.w4(32'h3a165247),
	.w5(32'h39f25c01),
	.w6(32'h398a0d80),
	.w7(32'h397ce2f8),
	.w8(32'h394bc3e8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8598502),
	.w1(32'hba1adeb0),
	.w2(32'hba9b5b3d),
	.w3(32'h3998a06f),
	.w4(32'h3807c1ba),
	.w5(32'hba8ee46c),
	.w6(32'hb8f72c68),
	.w7(32'hb908bf56),
	.w8(32'hbaab7bb3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d5efa1),
	.w1(32'h398deb45),
	.w2(32'hb99348e5),
	.w3(32'h39689e98),
	.w4(32'h3958bc34),
	.w5(32'hba44b62a),
	.w6(32'h3a3c17d1),
	.w7(32'h39d97e36),
	.w8(32'hb9f8226b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c7ce1),
	.w1(32'hb9a988d2),
	.w2(32'hb9e31499),
	.w3(32'hba4497b1),
	.w4(32'hba0e580e),
	.w5(32'hb9840aea),
	.w6(32'h3a5e6161),
	.w7(32'h3a803e98),
	.w8(32'h370fafe9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d0520),
	.w1(32'hba18b641),
	.w2(32'hba944887),
	.w3(32'h39ec35d3),
	.w4(32'h3898bce2),
	.w5(32'hba89dc2c),
	.w6(32'h37cc3d32),
	.w7(32'h39cb1174),
	.w8(32'hb97343d6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974ab73),
	.w1(32'hb9119aa2),
	.w2(32'hba1186f9),
	.w3(32'h391d4d4f),
	.w4(32'h39cec50c),
	.w5(32'hb96b7afa),
	.w6(32'hba22571e),
	.w7(32'hb9e896e7),
	.w8(32'hba5bf93c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c95c93),
	.w1(32'hba05b686),
	.w2(32'hb8814f33),
	.w3(32'h39824025),
	.w4(32'hb933ac9f),
	.w5(32'hba6f96b4),
	.w6(32'h3a2ff1a6),
	.w7(32'h3a139352),
	.w8(32'hb9dfbd41),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aba80c),
	.w1(32'h38bcd7cf),
	.w2(32'hb96ebb3d),
	.w3(32'hb9b0ebef),
	.w4(32'h37c8d436),
	.w5(32'hb98f8b6f),
	.w6(32'h39699b47),
	.w7(32'h383ecba3),
	.w8(32'hb9c4f41b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba102da9),
	.w1(32'h389c803f),
	.w2(32'hba8b758e),
	.w3(32'hb91f72c6),
	.w4(32'h3927166a),
	.w5(32'hbab08f2b),
	.w6(32'h3a4feb3a),
	.w7(32'h39fe3526),
	.w8(32'hba832749),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ade7f),
	.w1(32'hb9009e5d),
	.w2(32'h3a154463),
	.w3(32'hb9345322),
	.w4(32'h395705a5),
	.w5(32'h3811aae6),
	.w6(32'hba0a5e7a),
	.w7(32'hb7e6b17e),
	.w8(32'h39f8eaf3),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905e582),
	.w1(32'h3983032f),
	.w2(32'h39bb7342),
	.w3(32'hb985e8dd),
	.w4(32'h38a584e4),
	.w5(32'h39656839),
	.w6(32'h3972030a),
	.w7(32'h39aad5e1),
	.w8(32'h39e18cc2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39baca20),
	.w1(32'hb9d49195),
	.w2(32'h38a6efad),
	.w3(32'h3939db65),
	.w4(32'h39ba0fcf),
	.w5(32'h3a97c859),
	.w6(32'hb9367e15),
	.w7(32'hb91126ee),
	.w8(32'h37647731),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fce7b),
	.w1(32'hb98fc686),
	.w2(32'hba4b29a9),
	.w3(32'h3a51bb47),
	.w4(32'hb9985aba),
	.w5(32'hba17d6be),
	.w6(32'hb9c80d5e),
	.w7(32'hb9d79a18),
	.w8(32'hb9e206e6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a31b2),
	.w1(32'hb9ac99e6),
	.w2(32'hba1e02b7),
	.w3(32'hba09c381),
	.w4(32'h395fcfc5),
	.w5(32'hb909626b),
	.w6(32'h394eb6a5),
	.w7(32'h39fafc45),
	.w8(32'h39515455),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3848acd4),
	.w1(32'hb9af9538),
	.w2(32'hbaab2ef5),
	.w3(32'h38c4234d),
	.w4(32'hba496627),
	.w5(32'hbadba174),
	.w6(32'hb90cb960),
	.w7(32'hbabb37ab),
	.w8(32'hbb0c875d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386e6abf),
	.w1(32'h3a352ebb),
	.w2(32'h3a1a5d3a),
	.w3(32'h3808496c),
	.w4(32'h3a16e91f),
	.w5(32'h3a272542),
	.w6(32'h3a04afbe),
	.w7(32'h3a0fa01c),
	.w8(32'h39ebf369),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8883bbd),
	.w1(32'hba86dbf6),
	.w2(32'hba566983),
	.w3(32'h3a278300),
	.w4(32'hbaadc298),
	.w5(32'hbb2229fd),
	.w6(32'hb9cb2e63),
	.w7(32'hba8e1e64),
	.w8(32'hbb04421c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba083ee5),
	.w1(32'hb8c1b1fb),
	.w2(32'hb9d2aa14),
	.w3(32'hba5be213),
	.w4(32'hba4198ac),
	.w5(32'hba5ff5f6),
	.w6(32'hb8a47d45),
	.w7(32'hba6e66ad),
	.w8(32'hbaf20d7d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb4638),
	.w1(32'h3961e788),
	.w2(32'hba14cffd),
	.w3(32'hb8f84691),
	.w4(32'h39a05a7a),
	.w5(32'hba13710e),
	.w6(32'h3a970914),
	.w7(32'h396dfe14),
	.w8(32'hba26167e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d94611),
	.w1(32'h3a3fe407),
	.w2(32'hb919b03d),
	.w3(32'h3a0199c4),
	.w4(32'h3a459283),
	.w5(32'hb9bf701a),
	.w6(32'hb7a4b95d),
	.w7(32'h3903d556),
	.w8(32'hba0ef31b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02b0ed),
	.w1(32'h3a365ad2),
	.w2(32'h3a66d86e),
	.w3(32'h399c00ec),
	.w4(32'h3a67546e),
	.w5(32'h3a80e62c),
	.w6(32'h39ce4c32),
	.w7(32'h3a626c53),
	.w8(32'h3a5ef6a0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938aaa9),
	.w1(32'hb852ebf6),
	.w2(32'h3941e06a),
	.w3(32'hb882e981),
	.w4(32'hb897bc23),
	.w5(32'h3984c172),
	.w6(32'hb972b9ba),
	.w7(32'hb80d30c5),
	.w8(32'hb9197837),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987c4bb),
	.w1(32'h3971a06c),
	.w2(32'hb998b129),
	.w3(32'h38b6da2f),
	.w4(32'h3982baec),
	.w5(32'hba589e30),
	.w6(32'hb87b9786),
	.w7(32'h3993000c),
	.w8(32'hb97d1c46),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b20670),
	.w1(32'h3837c814),
	.w2(32'h3a57ee6d),
	.w3(32'h379c458b),
	.w4(32'h3a1c09b0),
	.w5(32'h3b07a441),
	.w6(32'hb901dcb8),
	.w7(32'h3aa4deaf),
	.w8(32'h3acc7c40),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9903b35),
	.w1(32'h3942ace4),
	.w2(32'hb9bc44a9),
	.w3(32'hb9e7ab80),
	.w4(32'h3a1dfdb4),
	.w5(32'h3a166713),
	.w6(32'hba93c9c4),
	.w7(32'hb722c7fb),
	.w8(32'h3967fcec),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c3bb85),
	.w1(32'h39880ac9),
	.w2(32'h3980c8cb),
	.w3(32'h3a660fd2),
	.w4(32'h397c926a),
	.w5(32'h39b6d5f8),
	.w6(32'h384f224e),
	.w7(32'h389cf228),
	.w8(32'h38b0d5d7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39904228),
	.w1(32'h39967173),
	.w2(32'h3994c7dd),
	.w3(32'h3993e513),
	.w4(32'h393c3480),
	.w5(32'h398b2b39),
	.w6(32'h37b9fea2),
	.w7(32'h38a68d9a),
	.w8(32'hb8070097),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ad8c4),
	.w1(32'hba36fc17),
	.w2(32'hbab2e46a),
	.w3(32'h38c6f42e),
	.w4(32'hb91a6e95),
	.w5(32'hba5ad181),
	.w6(32'hba64e1b2),
	.w7(32'hba360f5e),
	.w8(32'hbab00acd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968efa9),
	.w1(32'hba8d39bc),
	.w2(32'hb990c14e),
	.w3(32'hb9e0d2ff),
	.w4(32'hba8e805f),
	.w5(32'h391e5fa9),
	.w6(32'hba720cb4),
	.w7(32'h385ec7b8),
	.w8(32'hba78398b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3f1aa),
	.w1(32'h39e25bd1),
	.w2(32'h37a63611),
	.w3(32'hba3f837e),
	.w4(32'h3a0dda59),
	.w5(32'hb8c3137f),
	.w6(32'h3a213d58),
	.w7(32'h3a6b19d1),
	.w8(32'hb8bac0cc),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6807c),
	.w1(32'h39582c67),
	.w2(32'h38f52d85),
	.w3(32'h38ea9755),
	.w4(32'h3836ada7),
	.w5(32'h3943bb5d),
	.w6(32'hb8c8dc9f),
	.w7(32'hb73e7bb4),
	.w8(32'hb93495ca),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba369960),
	.w1(32'h3a81a664),
	.w2(32'hb7066143),
	.w3(32'hbac31cf0),
	.w4(32'h38090377),
	.w5(32'hb976cfe3),
	.w6(32'hba9a3b2e),
	.w7(32'hb9c5cf42),
	.w8(32'hba332ede),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be889a),
	.w1(32'hb8db3148),
	.w2(32'hb9822c90),
	.w3(32'h39082ebe),
	.w4(32'hb9017bd1),
	.w5(32'hb965c08e),
	.w6(32'hb65b95fa),
	.w7(32'hb93fe177),
	.w8(32'hb8ae6637),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db0ac1),
	.w1(32'h398cbaf7),
	.w2(32'h39bad0da),
	.w3(32'hb9bb2086),
	.w4(32'h391e178e),
	.w5(32'h39674a75),
	.w6(32'h389a111c),
	.w7(32'h38da2d13),
	.w8(32'h394edd05),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b5424),
	.w1(32'hb9c8dade),
	.w2(32'hba1c7bc1),
	.w3(32'h3a639674),
	.w4(32'h3a1ebbdb),
	.w5(32'hb99c1a3f),
	.w6(32'h3a3f5487),
	.w7(32'h3a786e3d),
	.w8(32'h37c017e3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ef98e),
	.w1(32'hba38e236),
	.w2(32'hbac527c2),
	.w3(32'h3802a052),
	.w4(32'h388f2d0c),
	.w5(32'hba463f73),
	.w6(32'h3a1f9b76),
	.w7(32'hb74eaed9),
	.w8(32'hba8e9bc3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ef3c0),
	.w1(32'h39226572),
	.w2(32'hb92390d8),
	.w3(32'hb9d551c4),
	.w4(32'hb868e05b),
	.w5(32'hb9bc552b),
	.w6(32'hbabf4c48),
	.w7(32'hb99bed81),
	.w8(32'hba1f4053),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba794610),
	.w1(32'hb904f2f0),
	.w2(32'hba8a8c79),
	.w3(32'hba207697),
	.w4(32'hb52b4eac),
	.w5(32'hba9a8cf3),
	.w6(32'h3946f647),
	.w7(32'h38f1f9f3),
	.w8(32'hbabc49b5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39860854),
	.w1(32'hba1d6450),
	.w2(32'hba641b79),
	.w3(32'h393ff888),
	.w4(32'hba283b79),
	.w5(32'hba51bd47),
	.w6(32'hb9a16c14),
	.w7(32'hba0674e2),
	.w8(32'hb893b5fe),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933ace0),
	.w1(32'h395e4ae8),
	.w2(32'hbaa32237),
	.w3(32'h3ac6c0da),
	.w4(32'h3a163b71),
	.w5(32'hba9b87b4),
	.w6(32'h3a96e9da),
	.w7(32'h39f55f97),
	.w8(32'hba289775),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1e908),
	.w1(32'hba09ee31),
	.w2(32'hbaafc8e5),
	.w3(32'hba091416),
	.w4(32'hba34229e),
	.w5(32'hbab90dfd),
	.w6(32'hba54c29a),
	.w7(32'hb9f19d93),
	.w8(32'hba9835cb),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17123d),
	.w1(32'hba838c68),
	.w2(32'hb9dbfdc3),
	.w3(32'hb94c36cc),
	.w4(32'hba5779a9),
	.w5(32'hbaf6b602),
	.w6(32'h39a4efc9),
	.w7(32'hb9dd6ccc),
	.w8(32'hbaa219ee),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8906607),
	.w1(32'hba5db2ec),
	.w2(32'h3976e902),
	.w3(32'hb9d19dd4),
	.w4(32'hba386283),
	.w5(32'h3a3487a7),
	.w6(32'hba9d4dad),
	.w7(32'hb97da646),
	.w8(32'hb93dfc05),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3911951b),
	.w1(32'hb82aa3a0),
	.w2(32'h3871c343),
	.w3(32'h3a8b86b7),
	.w4(32'h39b1b61c),
	.w5(32'h39d6cedf),
	.w6(32'h3a58c481),
	.w7(32'h39f3fdf2),
	.w8(32'h3a0c5811),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b7ae37),
	.w1(32'h39a80da5),
	.w2(32'h39b2bdd5),
	.w3(32'h36d518a3),
	.w4(32'h39389e66),
	.w5(32'h3944e3b9),
	.w6(32'h39654149),
	.w7(32'h3919ca58),
	.w8(32'h39a39e38),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d55d04),
	.w1(32'hb9d61021),
	.w2(32'hba75d14d),
	.w3(32'h399d9609),
	.w4(32'hba11e548),
	.w5(32'hba8d17be),
	.w6(32'hba667b75),
	.w7(32'hba768eb2),
	.w8(32'hbab821bc),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba196f09),
	.w1(32'hba09d837),
	.w2(32'hba056558),
	.w3(32'hba282c86),
	.w4(32'hba244262),
	.w5(32'hbaa29af8),
	.w6(32'hba05f2dd),
	.w7(32'hb9dbd3f0),
	.w8(32'hb99908df),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bdcd9),
	.w1(32'h3a836296),
	.w2(32'hb7c0720b),
	.w3(32'hbaa69fd5),
	.w4(32'h3a5397c4),
	.w5(32'h3554a803),
	.w6(32'h3a1f5a63),
	.w7(32'hb799617b),
	.w8(32'hb9b91b28),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12e928),
	.w1(32'h3a475e9a),
	.w2(32'h38da194a),
	.w3(32'h3a0fef2e),
	.w4(32'h3a05ea1a),
	.w5(32'h39ae9a61),
	.w6(32'h3a07e164),
	.w7(32'h3a2da432),
	.w8(32'h393da679),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a372f21),
	.w1(32'h394c46d1),
	.w2(32'h39639ec7),
	.w3(32'h3a2c0176),
	.w4(32'h39a781ae),
	.w5(32'h39d57939),
	.w6(32'h39a0ecd1),
	.w7(32'h397ddd2f),
	.w8(32'h397a5d7c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7654f3f),
	.w1(32'hb9ee3b5b),
	.w2(32'hba74ee98),
	.w3(32'hb823e9f6),
	.w4(32'hb93967c2),
	.w5(32'hb9c84ad1),
	.w6(32'hba64546a),
	.w7(32'hb9f7f055),
	.w8(32'hb9d97de0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f8a56),
	.w1(32'hb9eaac3d),
	.w2(32'hbacb129c),
	.w3(32'hba009a32),
	.w4(32'hb9081b37),
	.w5(32'hbab08676),
	.w6(32'hb9f42419),
	.w7(32'h39ae6910),
	.w8(32'hba57bb69),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e448a3),
	.w1(32'hb9f8731c),
	.w2(32'hbaacca33),
	.w3(32'hb9f8c19a),
	.w4(32'hba2f50ad),
	.w5(32'hb9fb0d3b),
	.w6(32'hba131ad7),
	.w7(32'hb9f9adbe),
	.w8(32'hba1d3bb4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9553b8a),
	.w1(32'hb86f9e24),
	.w2(32'hb9da09f1),
	.w3(32'hb9f6f2a8),
	.w4(32'hb98025c7),
	.w5(32'hba11f45f),
	.w6(32'hb89fe42a),
	.w7(32'hb9d581f0),
	.w8(32'hb8fc793d),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c764c),
	.w1(32'hba2084bd),
	.w2(32'hba73a049),
	.w3(32'hb995a0bf),
	.w4(32'h39ba6432),
	.w5(32'hbab47bcd),
	.w6(32'h3a1d408b),
	.w7(32'hba2ebb26),
	.w8(32'hbb129d19),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93b7df),
	.w1(32'hba3bde1e),
	.w2(32'h39138d90),
	.w3(32'h39677788),
	.w4(32'h3997c27f),
	.w5(32'h3a9e9d16),
	.w6(32'h39601b1e),
	.w7(32'h3a73bf9d),
	.w8(32'h3ab0cff9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9249577),
	.w1(32'h397b507e),
	.w2(32'h3a077bb1),
	.w3(32'hb99fe962),
	.w4(32'h396f0f02),
	.w5(32'h398518fb),
	.w6(32'h381f697f),
	.w7(32'hb84abe71),
	.w8(32'hb7ce4c9a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396cec99),
	.w1(32'hb99f00bd),
	.w2(32'hba90fbeb),
	.w3(32'h39331bfb),
	.w4(32'h389b0edb),
	.w5(32'hba03625a),
	.w6(32'hb98ab298),
	.w7(32'hba1e148f),
	.w8(32'hba75e7b1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba641f20),
	.w1(32'hb9cab25b),
	.w2(32'hb9c9cb1c),
	.w3(32'hba6f72fb),
	.w4(32'hb9d6e54a),
	.w5(32'hb9afea11),
	.w6(32'hb946de98),
	.w7(32'hb98ab0a0),
	.w8(32'h38ecb28f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f31d30),
	.w1(32'hb934f4b6),
	.w2(32'hb97c5a6d),
	.w3(32'h36f9a78c),
	.w4(32'hb9a20e15),
	.w5(32'hb9455280),
	.w6(32'hb9aa66a7),
	.w7(32'hb9a622f7),
	.w8(32'hb9a9d9e5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9078392),
	.w1(32'hb9ce7626),
	.w2(32'hbaac4f82),
	.w3(32'h3898d47f),
	.w4(32'hb9cea7d5),
	.w5(32'hba22cd82),
	.w6(32'hb8e30f87),
	.w7(32'hb829bdf1),
	.w8(32'hb9d5dea3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c354a),
	.w1(32'hb968f9c8),
	.w2(32'hbaaca805),
	.w3(32'hb90c41c7),
	.w4(32'h3a89293e),
	.w5(32'h3a18e885),
	.w6(32'h3a1f5214),
	.w7(32'h39483535),
	.w8(32'h38eb2a65),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba967b81),
	.w1(32'hb9ae2d21),
	.w2(32'hba9a6e3d),
	.w3(32'h38a45218),
	.w4(32'hb9dcdd2e),
	.w5(32'hba9d4bc3),
	.w6(32'hba57d6d5),
	.w7(32'hba6f6511),
	.w8(32'hbaea8eb5),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a43a7c),
	.w1(32'h39e295c3),
	.w2(32'h38274d7a),
	.w3(32'hb91e4ad8),
	.w4(32'h3980d0ce),
	.w5(32'hb9df3957),
	.w6(32'h399323e7),
	.w7(32'h399c28fe),
	.w8(32'hb93b6043),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391441bf),
	.w1(32'hba91dfa4),
	.w2(32'hbb34f48d),
	.w3(32'h39d4dda5),
	.w4(32'hba94cdf9),
	.w5(32'hbb38c7a2),
	.w6(32'hba4c37b6),
	.w7(32'hbab6063f),
	.w8(32'hbb48bbf0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd6982),
	.w1(32'h394eb5b6),
	.w2(32'hb9fb5b54),
	.w3(32'hba161e6c),
	.w4(32'hb8c52bab),
	.w5(32'hba1486a7),
	.w6(32'hb905f895),
	.w7(32'hb9d755b3),
	.w8(32'hba08d978),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fdb884),
	.w1(32'h395bcd1c),
	.w2(32'h39609ad2),
	.w3(32'hb7477957),
	.w4(32'h394cfa51),
	.w5(32'h3956dc26),
	.w6(32'h396809f0),
	.w7(32'h392526f3),
	.w8(32'h391ee263),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a988cf),
	.w1(32'h39895fbd),
	.w2(32'h39db1a66),
	.w3(32'h3991a57f),
	.w4(32'h3941d0fd),
	.w5(32'h39aa7d1b),
	.w6(32'h39359879),
	.w7(32'h393c78c6),
	.w8(32'h399d9e1d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb7936),
	.w1(32'h3983efe9),
	.w2(32'h39b1d985),
	.w3(32'h39906be6),
	.w4(32'h39281169),
	.w5(32'h39bb3e87),
	.w6(32'hb784c98a),
	.w7(32'hb7aab229),
	.w8(32'hb817b345),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01bba2),
	.w1(32'hba1724b9),
	.w2(32'hbab10874),
	.w3(32'hb9a0c764),
	.w4(32'hba10025a),
	.w5(32'hbadbe292),
	.w6(32'hba461fd3),
	.w7(32'hba87d7ae),
	.w8(32'hbac0ba47),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a09c3),
	.w1(32'hba0f0cb8),
	.w2(32'h3a39f597),
	.w3(32'hba168a16),
	.w4(32'h38837f9e),
	.w5(32'h3a686586),
	.w6(32'hb983df8c),
	.w7(32'h3838d2d4),
	.w8(32'h3a66419c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f95b1),
	.w1(32'h389c12c2),
	.w2(32'hba38dbfa),
	.w3(32'hb98bc590),
	.w4(32'h3986c210),
	.w5(32'hba4a72e1),
	.w6(32'h3931244b),
	.w7(32'h391dd76a),
	.w8(32'hba7f0294),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39756cf6),
	.w1(32'h38cdc725),
	.w2(32'hba1985eb),
	.w3(32'hb787fdf6),
	.w4(32'hb93a58d0),
	.w5(32'hba26a9aa),
	.w6(32'hb9afa447),
	.w7(32'hb9b5e415),
	.w8(32'hb99baa4f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380d5798),
	.w1(32'h38c4379d),
	.w2(32'hba784003),
	.w3(32'h38c9838f),
	.w4(32'h3a108dd1),
	.w5(32'hba34693f),
	.w6(32'h3a3c8085),
	.w7(32'h3a346b8f),
	.w8(32'hba3ef237),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf3d1a),
	.w1(32'h39deff13),
	.w2(32'h365a01b5),
	.w3(32'h3a1115a1),
	.w4(32'h3a31f952),
	.w5(32'h39a3cf01),
	.w6(32'h3a5c2e20),
	.w7(32'h3a411e3d),
	.w8(32'hb95e1bd8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39168667),
	.w1(32'hb8dfce06),
	.w2(32'hbac9a7ec),
	.w3(32'h3a0f30f0),
	.w4(32'hba21b4d8),
	.w5(32'hbac2b770),
	.w6(32'hba0e8617),
	.w7(32'hba95059b),
	.w8(32'hbb1a049c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c79e04),
	.w1(32'hb9c4d0ea),
	.w2(32'hb98cfc19),
	.w3(32'hb93c1007),
	.w4(32'hb9d90728),
	.w5(32'hba160950),
	.w6(32'hb95225eb),
	.w7(32'hb9e6f1da),
	.w8(32'hb983f189),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fac1c),
	.w1(32'h38087b39),
	.w2(32'h397d1bd9),
	.w3(32'hb9d4ee57),
	.w4(32'h39331374),
	.w5(32'h39db0325),
	.w6(32'hb945e9c3),
	.w7(32'hb91f303f),
	.w8(32'h38e16562),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b320e),
	.w1(32'h3761fe88),
	.w2(32'hba8a00ea),
	.w3(32'h39804bf7),
	.w4(32'h38b02f66),
	.w5(32'hba7a6421),
	.w6(32'hba3808aa),
	.w7(32'hb95bddd3),
	.w8(32'hba492dd2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b8a54),
	.w1(32'hba00c074),
	.w2(32'hba431d23),
	.w3(32'hb8759ebf),
	.w4(32'h388a45a7),
	.w5(32'hba19a368),
	.w6(32'hb8c585d3),
	.w7(32'h3a20ded3),
	.w8(32'hbad130d7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956d558),
	.w1(32'hba7bcb1f),
	.w2(32'hbaeb6694),
	.w3(32'h38041eb9),
	.w4(32'hb9b1ffce),
	.w5(32'hbad66853),
	.w6(32'hb9912acb),
	.w7(32'hba163c24),
	.w8(32'hbabb93ad),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16c069),
	.w1(32'hb9fcdbe9),
	.w2(32'hba3666e4),
	.w3(32'hb984534a),
	.w4(32'hba0d812b),
	.w5(32'hba1f4622),
	.w6(32'hb98f286d),
	.w7(32'hb9e2f86a),
	.w8(32'hb9732ee4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9965be3),
	.w1(32'h39d82a43),
	.w2(32'h39d57fd6),
	.w3(32'hb9cc5f89),
	.w4(32'h39d0bd10),
	.w5(32'h39e3b0c1),
	.w6(32'h399887a0),
	.w7(32'h39a10731),
	.w8(32'h39969935),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be3f8a),
	.w1(32'h3a13b64f),
	.w2(32'h3a14b2a9),
	.w3(32'h39ad8f75),
	.w4(32'h3a0fa93a),
	.w5(32'h3a1983d7),
	.w6(32'h39e66ca7),
	.w7(32'h39b083b0),
	.w8(32'h39d13149),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c46b96),
	.w1(32'h3a541ba8),
	.w2(32'h39aa89b9),
	.w3(32'h39999607),
	.w4(32'h3a33679f),
	.w5(32'h397f91b4),
	.w6(32'h39668f63),
	.w7(32'h39f9137b),
	.w8(32'hb9132d81),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8834cc),
	.w1(32'hb9bad21d),
	.w2(32'hb9d831d4),
	.w3(32'hba0c9a81),
	.w4(32'hb994826a),
	.w5(32'hba1d3dda),
	.w6(32'hba836d94),
	.w7(32'hba556a56),
	.w8(32'hba8066cd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c61afb),
	.w1(32'hb9373f43),
	.w2(32'hba3ca763),
	.w3(32'hb9963ec9),
	.w4(32'hb9d0cdd2),
	.w5(32'hba713f7a),
	.w6(32'h383adeca),
	.w7(32'h39891b1b),
	.w8(32'hb9df18fb),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47f8d7),
	.w1(32'h3a87307c),
	.w2(32'h3999e5b4),
	.w3(32'hba58e198),
	.w4(32'h3a3ff4e4),
	.w5(32'h39f5e315),
	.w6(32'hb9985d13),
	.w7(32'h3a29fdad),
	.w8(32'h3a50e49a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d50022),
	.w1(32'hba04aeda),
	.w2(32'hbaacc99e),
	.w3(32'h39a350d6),
	.w4(32'h37f7aa0c),
	.w5(32'hba31ea9b),
	.w6(32'hba56272f),
	.w7(32'h3989ecbf),
	.w8(32'hba875f38),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94099a5),
	.w1(32'hb9a32bbc),
	.w2(32'hb99822c1),
	.w3(32'hb8887315),
	.w4(32'hb9a0e7cc),
	.w5(32'hb9955d6e),
	.w6(32'hb9b7c427),
	.w7(32'hb9d1c923),
	.w8(32'hb977b650),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c08718),
	.w1(32'h38ed57f7),
	.w2(32'hb68c7a33),
	.w3(32'hb9ce0a8e),
	.w4(32'h3936fc9c),
	.w5(32'h3929850b),
	.w6(32'h392ca97c),
	.w7(32'h38a12b99),
	.w8(32'hb85fed10),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397cd017),
	.w1(32'hb9609457),
	.w2(32'h38195867),
	.w3(32'h39937cfc),
	.w4(32'hba0c7de2),
	.w5(32'hb78ca6b3),
	.w6(32'hb9ef1fb8),
	.w7(32'hb98efb2f),
	.w8(32'hba86ba84),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ab706),
	.w1(32'h3821f22b),
	.w2(32'hba56d35b),
	.w3(32'hba51f43e),
	.w4(32'h39f3ee55),
	.w5(32'hb9c901fe),
	.w6(32'hb891d20b),
	.w7(32'hb9e2707b),
	.w8(32'hb9ba83ae),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972bdaf),
	.w1(32'h37ef1b9d),
	.w2(32'h3780a759),
	.w3(32'hb9ef275e),
	.w4(32'h389a11a0),
	.w5(32'hb851dd40),
	.w6(32'hb8b7b4cb),
	.w7(32'hb781c870),
	.w8(32'hb8a58b96),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48ece2),
	.w1(32'h3a41b405),
	.w2(32'h39590cc9),
	.w3(32'hb8b1d10f),
	.w4(32'h3a60654a),
	.w5(32'h39366df4),
	.w6(32'h3a717049),
	.w7(32'h3a9cffdb),
	.w8(32'h39089609),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b46604),
	.w1(32'hba3459ee),
	.w2(32'hbb4c3d1a),
	.w3(32'h3a159526),
	.w4(32'hba43dda6),
	.w5(32'hbb0c5414),
	.w6(32'hba2347ec),
	.w7(32'hbac1edc5),
	.w8(32'hbb1f7c33),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba733728),
	.w1(32'h391324a7),
	.w2(32'hba492d27),
	.w3(32'hba8b8666),
	.w4(32'hba0764a9),
	.w5(32'hba5163c2),
	.w6(32'hb4b1a256),
	.w7(32'hb9830751),
	.w8(32'hb9ce3bfd),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e28220),
	.w1(32'h39ba074d),
	.w2(32'hba056168),
	.w3(32'hb9fca532),
	.w4(32'h39d91f1c),
	.w5(32'hba36cacb),
	.w6(32'hb9fa2462),
	.w7(32'hb96e828f),
	.w8(32'hba49862e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b5b01),
	.w1(32'h39825225),
	.w2(32'hb829f0f2),
	.w3(32'h3a619e74),
	.w4(32'h394998e3),
	.w5(32'hb9985d92),
	.w6(32'h3a0080b8),
	.w7(32'hb8f32bd4),
	.w8(32'hb9c3d34f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caa26e),
	.w1(32'h394db21f),
	.w2(32'h3899909a),
	.w3(32'h3984cfdc),
	.w4(32'h39733f08),
	.w5(32'h391bbd2f),
	.w6(32'h37a63bb4),
	.w7(32'h38afbda7),
	.w8(32'h38874a81),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39784650),
	.w1(32'h38ebc485),
	.w2(32'hb89185cf),
	.w3(32'h39341b9a),
	.w4(32'hb8a6b67b),
	.w5(32'hb8ab3d92),
	.w6(32'h381a7724),
	.w7(32'h38c783cd),
	.w8(32'hb9ece289),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39118bed),
	.w1(32'hb9d0a091),
	.w2(32'hb9e24cb1),
	.w3(32'h38f228f8),
	.w4(32'hb9f285ef),
	.w5(32'hb9dcb23d),
	.w6(32'hba060fd6),
	.w7(32'hba139553),
	.w8(32'hb98df473),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac7f2f),
	.w1(32'h39ea52d0),
	.w2(32'h3a0643f9),
	.w3(32'hb9ed0b49),
	.w4(32'h39b226da),
	.w5(32'h3a0278cc),
	.w6(32'h39a22aa8),
	.w7(32'h39748feb),
	.w8(32'h396f5005),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ace09),
	.w1(32'h394a6be7),
	.w2(32'h394b7073),
	.w3(32'h399d40e3),
	.w4(32'h3910bf5d),
	.w5(32'h3947d4b7),
	.w6(32'hb7685946),
	.w7(32'h3897fa21),
	.w8(32'h3912efea),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398161a8),
	.w1(32'hb9d4d4d7),
	.w2(32'hb9d4c2e4),
	.w3(32'h397756aa),
	.w4(32'hba286551),
	.w5(32'hba6421c9),
	.w6(32'hb97219e6),
	.w7(32'hb9925a48),
	.w8(32'hb8f817d2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8e816),
	.w1(32'h398766e8),
	.w2(32'h3866afe8),
	.w3(32'hba05bd10),
	.w4(32'h38b8e887),
	.w5(32'hb980154e),
	.w6(32'hb9458124),
	.w7(32'h39c2308e),
	.w8(32'h38ebb28f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9504a37),
	.w1(32'hb9ac5ce8),
	.w2(32'hbaffd568),
	.w3(32'h38a59fa4),
	.w4(32'hb94ff2f6),
	.w5(32'hbb1ae823),
	.w6(32'h3a9b90e1),
	.w7(32'h39221db8),
	.w8(32'hbad8cf78),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a78a8),
	.w1(32'hb900683a),
	.w2(32'hba10eab4),
	.w3(32'hb99620c9),
	.w4(32'hb8ed2716),
	.w5(32'hba96ffe5),
	.w6(32'h39fa3dbe),
	.w7(32'h37fd1452),
	.w8(32'hba395279),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb31f4),
	.w1(32'hba61d103),
	.w2(32'hbac351d2),
	.w3(32'h39f7b6da),
	.w4(32'hb960a4d2),
	.w5(32'hba70eb87),
	.w6(32'hb90c8f73),
	.w7(32'hba23813a),
	.w8(32'hba93d9d2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f4163),
	.w1(32'h3a9201cf),
	.w2(32'h3a546bb1),
	.w3(32'hba24727f),
	.w4(32'h3a92d2cb),
	.w5(32'h3a6848db),
	.w6(32'h3a73f239),
	.w7(32'h3a64b17d),
	.w8(32'h3a867304),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90e8f4),
	.w1(32'h399231f9),
	.w2(32'h3997f875),
	.w3(32'h3a6dceeb),
	.w4(32'h3963aef3),
	.w5(32'h399b62f8),
	.w6(32'hb78b5341),
	.w7(32'h38fb208c),
	.w8(32'h39601dac),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d22631),
	.w1(32'h3995afc9),
	.w2(32'h398a1e83),
	.w3(32'h39c54388),
	.w4(32'h3991115e),
	.w5(32'h399dca21),
	.w6(32'h3916d101),
	.w7(32'h3904c0ea),
	.w8(32'h3899e001),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397937cc),
	.w1(32'h39b93d87),
	.w2(32'h3987136a),
	.w3(32'h3994b4ba),
	.w4(32'h39abfbf0),
	.w5(32'h39af73f8),
	.w6(32'h394bb8ed),
	.w7(32'h39556b8f),
	.w8(32'h392c4d53),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c0618),
	.w1(32'h35e5c5a0),
	.w2(32'h3a29f27e),
	.w3(32'h3a5d66bd),
	.w4(32'h3995a240),
	.w5(32'hba08efc4),
	.w6(32'h38867d03),
	.w7(32'hb9055133),
	.w8(32'hb78be02c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca64d8),
	.w1(32'hb9152a78),
	.w2(32'hba4cd5f1),
	.w3(32'hb86d33d6),
	.w4(32'hb9d678f2),
	.w5(32'hb9dadd1b),
	.w6(32'hb9ad3791),
	.w7(32'hb9da30db),
	.w8(32'hb9c7391e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3c423),
	.w1(32'h3a0d8364),
	.w2(32'h39308ce1),
	.w3(32'hba540a3d),
	.w4(32'h3988e931),
	.w5(32'hb8cab4e2),
	.w6(32'hb9cff150),
	.w7(32'h393eb035),
	.w8(32'hb9936faf),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89802d3),
	.w1(32'h397199cd),
	.w2(32'h38ee7e0a),
	.w3(32'hb97a96f6),
	.w4(32'h38d3fe3c),
	.w5(32'h39508d5a),
	.w6(32'hb981d350),
	.w7(32'h39041e2d),
	.w8(32'hb9089d91),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39968305),
	.w1(32'h39f10b3c),
	.w2(32'h3a0109a9),
	.w3(32'h39a09bde),
	.w4(32'h39c9db40),
	.w5(32'h39d2187a),
	.w6(32'h398f082e),
	.w7(32'h3986748f),
	.w8(32'h39a9085f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc89bf),
	.w1(32'hb9fe179b),
	.w2(32'h3a3fac71),
	.w3(32'h3a1a85f9),
	.w4(32'hba56693e),
	.w5(32'hba5a8889),
	.w6(32'hb8ef734e),
	.w7(32'hba9100a1),
	.w8(32'hba8ba43d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e73493),
	.w1(32'h3a8a6808),
	.w2(32'h3a6376b2),
	.w3(32'hb9e285d9),
	.w4(32'h3a9df502),
	.w5(32'h3a8a5531),
	.w6(32'h3a5498c7),
	.w7(32'h3a4eb491),
	.w8(32'h3a712a80),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6df424),
	.w1(32'h37f72ac5),
	.w2(32'hba1f2b38),
	.w3(32'h3a8c6554),
	.w4(32'hb94cc550),
	.w5(32'hb9170f45),
	.w6(32'h39d99dae),
	.w7(32'h38333c5d),
	.w8(32'hba16c0fb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc888d),
	.w1(32'h3989e960),
	.w2(32'hb90c80de),
	.w3(32'h39edfdc6),
	.w4(32'h3974ef1a),
	.w5(32'hb86a5f96),
	.w6(32'h3966e601),
	.w7(32'hb889ed4b),
	.w8(32'h399a08da),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a571436),
	.w1(32'hb9cf2faa),
	.w2(32'hba3658c0),
	.w3(32'h3a81fcfc),
	.w4(32'hb909289d),
	.w5(32'hba64f466),
	.w6(32'h3a71eb6f),
	.w7(32'h3911091e),
	.w8(32'h38b14720),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule