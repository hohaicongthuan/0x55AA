module layer_10_featuremap_166(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a31a23),
	.w1(32'h391f092a),
	.w2(32'hbaab1bd8),
	.w3(32'hb9cdaa9d),
	.w4(32'h3a94c05c),
	.w5(32'h38fcf080),
	.w6(32'h398697c6),
	.w7(32'h39fcc47f),
	.w8(32'h3955e583),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecd60c),
	.w1(32'h388fb325),
	.w2(32'hb9acb81f),
	.w3(32'hbae97a96),
	.w4(32'hb96c3898),
	.w5(32'hb9013f7a),
	.w6(32'hb9b45058),
	.w7(32'h387666dc),
	.w8(32'hb9ef713f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba210e),
	.w1(32'hb71db2f9),
	.w2(32'hb826352b),
	.w3(32'hb8871807),
	.w4(32'hba032229),
	.w5(32'hba2b705d),
	.w6(32'hb8aa74d2),
	.w7(32'hb8754a27),
	.w8(32'hb842ef4e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b92d57),
	.w1(32'hb9af0ada),
	.w2(32'hba2185e4),
	.w3(32'hbace0cd9),
	.w4(32'hba4d4617),
	.w5(32'hba6f1dd2),
	.w6(32'hb95f4dc2),
	.w7(32'h39320ca0),
	.w8(32'h3911de21),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e57e7c),
	.w1(32'h38dfbd7c),
	.w2(32'hb9e464a2),
	.w3(32'hb9417400),
	.w4(32'h39aeeab3),
	.w5(32'hb81a4102),
	.w6(32'hb7a55431),
	.w7(32'hb9796310),
	.w8(32'h39bfbebd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ff93a),
	.w1(32'hba1948d6),
	.w2(32'hba2d0c1a),
	.w3(32'h39347be0),
	.w4(32'hba08ebae),
	.w5(32'hba32ae2a),
	.w6(32'hb9bdd269),
	.w7(32'hba292b33),
	.w8(32'hba043fe8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b2991),
	.w1(32'h3ab76e3f),
	.w2(32'hb9ef859e),
	.w3(32'h3af956f6),
	.w4(32'hb98fb328),
	.w5(32'hbb8bcf11),
	.w6(32'h3a3114aa),
	.w7(32'hba95ca4e),
	.w8(32'hbb0987b7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31d2d7),
	.w1(32'hbba26693),
	.w2(32'hbbb464b1),
	.w3(32'hbb9795af),
	.w4(32'hbbb95095),
	.w5(32'hba62ba37),
	.w6(32'hbb0bc2f4),
	.w7(32'h3ad7e532),
	.w8(32'h3a593cbb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f58d0),
	.w1(32'h397089a3),
	.w2(32'h39735b0e),
	.w3(32'h39e98c50),
	.w4(32'h390d7ddd),
	.w5(32'h38d0bf3b),
	.w6(32'h3a6c77a5),
	.w7(32'h3a0e6539),
	.w8(32'h39dc261d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c882d),
	.w1(32'h3b715d13),
	.w2(32'h3a11c617),
	.w3(32'hba921656),
	.w4(32'hba0eb947),
	.w5(32'hbb2516bd),
	.w6(32'hbb025828),
	.w7(32'hbafefa77),
	.w8(32'hbaa046fb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f12ceb),
	.w1(32'hb8fa65f3),
	.w2(32'h391d0c29),
	.w3(32'h39b3b3c1),
	.w4(32'h37a3d1be),
	.w5(32'h3a2be792),
	.w6(32'h399b0df4),
	.w7(32'h39af065c),
	.w8(32'h38d93166),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e4523),
	.w1(32'h3b5f327d),
	.w2(32'hba83f586),
	.w3(32'h3b64dda2),
	.w4(32'h3b190b5c),
	.w5(32'hbba075d2),
	.w6(32'hb96e4310),
	.w7(32'hbac42433),
	.w8(32'hbb833a37),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fb04c),
	.w1(32'h39fae611),
	.w2(32'hbb00eccf),
	.w3(32'hbb5c61fd),
	.w4(32'hbb756418),
	.w5(32'hbb859e9b),
	.w6(32'hbb5e603a),
	.w7(32'hbb48f86c),
	.w8(32'hbb338a2d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f30a8),
	.w1(32'hbaca47cf),
	.w2(32'hbb2da8b8),
	.w3(32'h3a1f67cb),
	.w4(32'hb9450198),
	.w5(32'hbacf5d4b),
	.w6(32'h39df0186),
	.w7(32'hba21d2a9),
	.w8(32'hb917d368),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995e59d),
	.w1(32'h3a5c6c99),
	.w2(32'h39ea6bf0),
	.w3(32'h3920260e),
	.w4(32'h3afc4b9d),
	.w5(32'h3ad6ae77),
	.w6(32'h3a68e1b6),
	.w7(32'h3ada1633),
	.w8(32'h3a7b0990),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13e0dc),
	.w1(32'h39c1522c),
	.w2(32'hbb3853bc),
	.w3(32'hbb1a5cd2),
	.w4(32'hbb93e977),
	.w5(32'hbb81e77f),
	.w6(32'hbb00086f),
	.w7(32'hbb27bbd7),
	.w8(32'hb8e43a5a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a51a1c),
	.w1(32'h3829fa15),
	.w2(32'h3a277613),
	.w3(32'h38b5121f),
	.w4(32'hb9a15fc5),
	.w5(32'hb9ea6361),
	.w6(32'h391a1b8c),
	.w7(32'h399d07e2),
	.w8(32'hba69a031),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf7aaf),
	.w1(32'h3a1d7cc9),
	.w2(32'hbb61dcfd),
	.w3(32'hbba60f7d),
	.w4(32'hbbc5c375),
	.w5(32'hbbfd9bda),
	.w6(32'hbb4785a5),
	.w7(32'h3a88cdcf),
	.w8(32'h3a978643),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeed13f),
	.w1(32'hb987748a),
	.w2(32'hbad89924),
	.w3(32'hbad79dd0),
	.w4(32'hbb49ee0b),
	.w5(32'hbb6cbfa7),
	.w6(32'hbade96b7),
	.w7(32'hb9292fe6),
	.w8(32'hb9d3cf06),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fa8b7),
	.w1(32'hb98d69a8),
	.w2(32'hb80e05c6),
	.w3(32'hb9c7843e),
	.w4(32'hb9b8caeb),
	.w5(32'hb93bb4ba),
	.w6(32'hb9884919),
	.w7(32'hb905c254),
	.w8(32'hb8e9877b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81bc022),
	.w1(32'h3979e308),
	.w2(32'hb83259b6),
	.w3(32'hb912aa42),
	.w4(32'h397323e4),
	.w5(32'h39012d44),
	.w6(32'h39ea746b),
	.w7(32'h3987a073),
	.w8(32'h3a0b6aeb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe7022),
	.w1(32'h3a0c1402),
	.w2(32'h3638030d),
	.w3(32'h395c7588),
	.w4(32'h3a8d768d),
	.w5(32'h3a13be23),
	.w6(32'h39ce3f93),
	.w7(32'h3ae33600),
	.w8(32'hb861c2a4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00d289),
	.w1(32'h3b0fb991),
	.w2(32'h3b06e91b),
	.w3(32'hbb1c3dbb),
	.w4(32'hbbaafa83),
	.w5(32'hbbc32fd6),
	.w6(32'hba656ff8),
	.w7(32'h3acdd8b8),
	.w8(32'h3bac0fe3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f4181),
	.w1(32'h3b006789),
	.w2(32'h3aa24877),
	.w3(32'hbabd7b3f),
	.w4(32'hba10e5ce),
	.w5(32'hba56bb28),
	.w6(32'hba87ea56),
	.w7(32'hba3ea1be),
	.w8(32'hb8eab8c0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c9b0b),
	.w1(32'h3abd03fd),
	.w2(32'h3aa62d97),
	.w3(32'hbb922686),
	.w4(32'hba24ffcd),
	.w5(32'h3a82f8da),
	.w6(32'hbadbf992),
	.w7(32'h3a1d0c03),
	.w8(32'h3a5a8bdd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39135c1e),
	.w1(32'h378d0314),
	.w2(32'h3a3fc4b8),
	.w3(32'h389a533f),
	.w4(32'hb9c4cfd8),
	.w5(32'hb9ef3ca9),
	.w6(32'hb9695a99),
	.w7(32'hb9281563),
	.w8(32'h38ccf6f9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb855fc68),
	.w1(32'hba016fa1),
	.w2(32'hb9d61eeb),
	.w3(32'hb95c0f4e),
	.w4(32'hba0b9ae0),
	.w5(32'hb9b5ad29),
	.w6(32'hb9af7b27),
	.w7(32'hb9c29cea),
	.w8(32'hb996c0ab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4b7f1),
	.w1(32'h3ac5c421),
	.w2(32'h3ad8b7a2),
	.w3(32'hbb9a7511),
	.w4(32'hb9e1626f),
	.w5(32'hb9e50605),
	.w6(32'hbba1b753),
	.w7(32'hbb9eaedf),
	.w8(32'h39a0f31e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87eb37),
	.w1(32'hba4f4d4d),
	.w2(32'hba492c95),
	.w3(32'hba597847),
	.w4(32'hba30843c),
	.w5(32'hba3e3888),
	.w6(32'hba1ec940),
	.w7(32'hbabc2156),
	.w8(32'hba74b8c9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba874c15),
	.w1(32'h3b394b8f),
	.w2(32'h3b9fb05f),
	.w3(32'hbb32cfc7),
	.w4(32'hba036511),
	.w5(32'h3a8a8060),
	.w6(32'hba98b8aa),
	.w7(32'hbaa316ab),
	.w8(32'h39c0038d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8657b01),
	.w1(32'h37e9d9c3),
	.w2(32'hb8f19db2),
	.w3(32'h3885ed1b),
	.w4(32'h380b9925),
	.w5(32'hb81b977f),
	.w6(32'h396657a2),
	.w7(32'h38194bfd),
	.w8(32'h391214c5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a31b72),
	.w1(32'hb957d303),
	.w2(32'hb998770b),
	.w3(32'h399f91a7),
	.w4(32'hb8c6d386),
	.w5(32'hb9a75720),
	.w6(32'hb8722b57),
	.w7(32'hb99687f8),
	.w8(32'hb99846ed),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00bff2),
	.w1(32'h3ade3a50),
	.w2(32'h39e22c39),
	.w3(32'hb98b42a4),
	.w4(32'hba07ea91),
	.w5(32'hba965294),
	.w6(32'h38a20860),
	.w7(32'h38431bd8),
	.w8(32'h38f79cbd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a187b14),
	.w1(32'h3a538d7e),
	.w2(32'h391e1e92),
	.w3(32'h39f6d385),
	.w4(32'h3a2509f0),
	.w5(32'hb7fee63d),
	.w6(32'h3aac244b),
	.w7(32'h3abdce39),
	.w8(32'hb7eaee8d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a202c1e),
	.w1(32'h3a515527),
	.w2(32'h3a27a05a),
	.w3(32'hb9ca4ece),
	.w4(32'h38b3e8ca),
	.w5(32'hb9fab017),
	.w6(32'h3992984c),
	.w7(32'h39907d1e),
	.w8(32'h39f58d70),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b026aca),
	.w1(32'h3a43ecbb),
	.w2(32'hbaa9f385),
	.w3(32'hba9856bf),
	.w4(32'hbae815a6),
	.w5(32'hbb371812),
	.w6(32'hb923c451),
	.w7(32'hb9e2a4a7),
	.w8(32'hba01c7fd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cb0e8),
	.w1(32'h3ba1bf9b),
	.w2(32'h3a26f09c),
	.w3(32'hbb819a47),
	.w4(32'h3b9ec52a),
	.w5(32'hbb689871),
	.w6(32'hbb5b5c8b),
	.w7(32'hb9ae42ce),
	.w8(32'h3a0c4da2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5bd54),
	.w1(32'h3bf5047c),
	.w2(32'h3bc1b6bd),
	.w3(32'hbb2f2cfa),
	.w4(32'h3bc211ed),
	.w5(32'h3ba2dcd8),
	.w6(32'hbb6e8fa2),
	.w7(32'h3b05cb1b),
	.w8(32'hbb0d6bed),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98d34f),
	.w1(32'h3b6d2911),
	.w2(32'h3bf8a1a9),
	.w3(32'hbb027e03),
	.w4(32'h3b45422c),
	.w5(32'h3b8dd486),
	.w6(32'hbb0ed6a7),
	.w7(32'h39574f7a),
	.w8(32'h3b006f5c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6e123),
	.w1(32'h3a04eacc),
	.w2(32'h394f8ad9),
	.w3(32'hbaf5d856),
	.w4(32'hb917b3f2),
	.w5(32'hb9c31178),
	.w6(32'hbad03ceb),
	.w7(32'hb98c792a),
	.w8(32'hba1a9aeb),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f084a6),
	.w1(32'h398bab28),
	.w2(32'hb93b2fcd),
	.w3(32'hb9394d1d),
	.w4(32'h399120f0),
	.w5(32'hb7dd0650),
	.w6(32'h39c0e14e),
	.w7(32'h398743ae),
	.w8(32'h39c0500d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7e356),
	.w1(32'h3929e3a8),
	.w2(32'h3a14e681),
	.w3(32'hb99a1300),
	.w4(32'h39751129),
	.w5(32'h39bcfe77),
	.w6(32'h37fe121e),
	.w7(32'h3949f27f),
	.w8(32'h380ccfd4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa0067),
	.w1(32'h3a1f6df9),
	.w2(32'h3a8498c4),
	.w3(32'h3aa99add),
	.w4(32'h3a1ce196),
	.w5(32'h3a1aa5db),
	.w6(32'h3a857071),
	.w7(32'h397fd7a9),
	.w8(32'h3929201b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b423b58),
	.w1(32'h3b85fce4),
	.w2(32'h3a087638),
	.w3(32'hbb18eae4),
	.w4(32'hbaf1fec9),
	.w5(32'hbb41dada),
	.w6(32'hbb37eaca),
	.w7(32'hbaa64b93),
	.w8(32'h3a2e95be),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95db47),
	.w1(32'h3b46a9d1),
	.w2(32'h3b25c57c),
	.w3(32'hb9babc6e),
	.w4(32'h3ab17bf1),
	.w5(32'h3ac0bfd1),
	.w6(32'h3a56163f),
	.w7(32'h3b210cda),
	.w8(32'h3ae54b07),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab71c01),
	.w1(32'h3b11c580),
	.w2(32'h3abd242e),
	.w3(32'hbb2751dd),
	.w4(32'hbad9840e),
	.w5(32'hb9ed7996),
	.w6(32'h39215ead),
	.w7(32'h3ae88233),
	.w8(32'h3a806ccc),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3094b4),
	.w1(32'h3b30b7c2),
	.w2(32'h3b19868c),
	.w3(32'h3a518f1a),
	.w4(32'h3ac55605),
	.w5(32'h3ab1190b),
	.w6(32'h3b5233cf),
	.w7(32'h3b587271),
	.w8(32'h3b836891),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be996f8),
	.w1(32'h3b46a95a),
	.w2(32'hbb59f0e4),
	.w3(32'hba2cf6b9),
	.w4(32'hbba5d34b),
	.w5(32'hbc0beba2),
	.w6(32'hbafaf2a0),
	.w7(32'hb8f1a88f),
	.w8(32'h39ac6673),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1218a4),
	.w1(32'hba1b18c8),
	.w2(32'hb8800ffb),
	.w3(32'hb9da8e99),
	.w4(32'hba3ccd14),
	.w5(32'hb9989994),
	.w6(32'hba1a2aac),
	.w7(32'hba1a3e28),
	.w8(32'hb9a0fab4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba099a70),
	.w1(32'h393bc6e3),
	.w2(32'h3a378e28),
	.w3(32'hb9bc7a62),
	.w4(32'h3a163d8a),
	.w5(32'h3a63b9d1),
	.w6(32'h3a260ba7),
	.w7(32'h3a93ad4a),
	.w8(32'h3ac1a769),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba363320),
	.w1(32'h3929a7fa),
	.w2(32'h3a440e25),
	.w3(32'hba3f6eb0),
	.w4(32'h390d0a72),
	.w5(32'h39f09bcc),
	.w6(32'h381bb349),
	.w7(32'h399cc70f),
	.w8(32'h3a40e0c0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9da2e),
	.w1(32'hb82d7ba1),
	.w2(32'h3a06011d),
	.w3(32'hbaa17cd4),
	.w4(32'hbb1f1134),
	.w5(32'hba86bffc),
	.w6(32'hbac5cd80),
	.w7(32'hba8eb41a),
	.w8(32'hb7733766),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940c723),
	.w1(32'h3980e3a2),
	.w2(32'h39264f9f),
	.w3(32'hb91c106c),
	.w4(32'hb9f87f83),
	.w5(32'hb98c5e03),
	.w6(32'h3a0c25ff),
	.w7(32'h3a69067f),
	.w8(32'h3ac81f74),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d15a),
	.w1(32'h3ac9d9b0),
	.w2(32'hbb345111),
	.w3(32'hbaf88c8d),
	.w4(32'hbb4fc330),
	.w5(32'hbbf351e8),
	.w6(32'hbb8cbcb8),
	.w7(32'hbb138bdf),
	.w8(32'hbab06823),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30ecae),
	.w1(32'h383b804a),
	.w2(32'hb9a25c0c),
	.w3(32'hba1c54a1),
	.w4(32'hba7b3ad3),
	.w5(32'hba1362d8),
	.w6(32'h3a6b0988),
	.w7(32'h3a71c70d),
	.w8(32'h3aa56829),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e160a),
	.w1(32'h3a22e286),
	.w2(32'hb97f90fb),
	.w3(32'hb8eae836),
	.w4(32'h39908707),
	.w5(32'hb940f250),
	.w6(32'h3a5b17f4),
	.w7(32'h39e16965),
	.w8(32'h39e99622),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d02aba),
	.w1(32'h3a59d059),
	.w2(32'h3a5bff08),
	.w3(32'h37b69a53),
	.w4(32'h3a08f32a),
	.w5(32'h39dc87e8),
	.w6(32'h3a470ae9),
	.w7(32'h3a49df88),
	.w8(32'h3a49dcda),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cf111),
	.w1(32'h399df2e0),
	.w2(32'hb9ad40e5),
	.w3(32'h39943ea6),
	.w4(32'h385aeef2),
	.w5(32'hb9527471),
	.w6(32'hb8f3bdd7),
	.w7(32'hba2a0a5b),
	.w8(32'hb9844024),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9264984),
	.w1(32'h39d78a95),
	.w2(32'h39e6f1df),
	.w3(32'h392193fc),
	.w4(32'h39ea5c11),
	.w5(32'h393be95d),
	.w6(32'h3a6d93ce),
	.w7(32'h3a45f6d7),
	.w8(32'h3a1c5a22),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a13bd8),
	.w1(32'hb9f222a9),
	.w2(32'hb92be5db),
	.w3(32'h3888e3aa),
	.w4(32'hba06f4b8),
	.w5(32'hba17f2ee),
	.w6(32'hb99058ea),
	.w7(32'hba564cd1),
	.w8(32'hb9bdf9b6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6af8c8),
	.w1(32'h381e23a6),
	.w2(32'hba9c77ea),
	.w3(32'hbaa02593),
	.w4(32'hbb02d3dd),
	.w5(32'hbb5365d5),
	.w6(32'hba8e99ca),
	.w7(32'hb9b1c2d5),
	.w8(32'hb9a94f23),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae40f13),
	.w1(32'h3b14c967),
	.w2(32'hb905e25e),
	.w3(32'hbb1d6f25),
	.w4(32'hba36fb86),
	.w5(32'hb90f8343),
	.w6(32'hba28cd19),
	.w7(32'h3a8192a9),
	.w8(32'h3b2597de),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa5be2),
	.w1(32'h3a89194d),
	.w2(32'h39ddb787),
	.w3(32'h3990cddc),
	.w4(32'h3a107d0a),
	.w5(32'h39ec9714),
	.w6(32'h3a17388d),
	.w7(32'h3a4b8cf3),
	.w8(32'h3aac53ba),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a1706),
	.w1(32'h3a3eca3c),
	.w2(32'h3a0983c5),
	.w3(32'h3a881e22),
	.w4(32'h3a460a50),
	.w5(32'h3a0123c6),
	.w6(32'h3a3484d9),
	.w7(32'h3a058f57),
	.w8(32'h3a012c1c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997b0cd),
	.w1(32'hb9b7ddca),
	.w2(32'hb90309d6),
	.w3(32'h39345067),
	.w4(32'hb9ee154e),
	.w5(32'hb989aa58),
	.w6(32'hb9c03c2b),
	.w7(32'hb9b9516b),
	.w8(32'hb94f337b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88933c1),
	.w1(32'h39dc5e9f),
	.w2(32'h3990ab57),
	.w3(32'hb9828002),
	.w4(32'h39f6b4b5),
	.w5(32'h38a07df3),
	.w6(32'hb7a55b15),
	.w7(32'h3865b435),
	.w8(32'hb99d1a0e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc5940),
	.w1(32'h3b842437),
	.w2(32'hba85d66d),
	.w3(32'h3b2bc446),
	.w4(32'hbaadebd6),
	.w5(32'hbbc4dd55),
	.w6(32'hbb8f29e2),
	.w7(32'hbba3de5b),
	.w8(32'hb9b5cda7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addf45b),
	.w1(32'h3afc9680),
	.w2(32'hbb1468f5),
	.w3(32'hbbb7e75a),
	.w4(32'hbba06b4d),
	.w5(32'hbbb49353),
	.w6(32'h3b297fc8),
	.w7(32'h3b246fae),
	.w8(32'h3ac818ec),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39aa76),
	.w1(32'hb936f954),
	.w2(32'hbb0d4e82),
	.w3(32'hbb8558e1),
	.w4(32'hbba7324e),
	.w5(32'hbb8deed4),
	.w6(32'h3a87385a),
	.w7(32'h3ac7e22c),
	.w8(32'h3b1564d7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba24bc9),
	.w1(32'h3b8aa30b),
	.w2(32'h3b4e8599),
	.w3(32'hbbdc48b5),
	.w4(32'h39be2a3b),
	.w5(32'h3a4e1121),
	.w6(32'hbb74746a),
	.w7(32'h392ebdb2),
	.w8(32'hbb11a862),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37be4222),
	.w1(32'h39cd442a),
	.w2(32'h3a16da13),
	.w3(32'h39602aa0),
	.w4(32'h39f1f6b9),
	.w5(32'h39ae6c02),
	.w6(32'h39977878),
	.w7(32'h39db34c5),
	.w8(32'h39e3e11a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39765f43),
	.w1(32'hb94e3ac8),
	.w2(32'hb98c73fa),
	.w3(32'h388eec6f),
	.w4(32'hb8c4ab8e),
	.w5(32'hb929a9f6),
	.w6(32'hb894fcf1),
	.w7(32'hb9001ea2),
	.w8(32'h38b95737),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905c651),
	.w1(32'hb9935075),
	.w2(32'hb9abb138),
	.w3(32'hb8aa1813),
	.w4(32'hb94b8405),
	.w5(32'hb978d233),
	.w6(32'hb9380704),
	.w7(32'hb9947c83),
	.w8(32'hb8910bd4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3eb44f),
	.w1(32'h38de696c),
	.w2(32'hba535b60),
	.w3(32'hb9c95720),
	.w4(32'hba57e9f9),
	.w5(32'hbabf1865),
	.w6(32'hba07ace8),
	.w7(32'hb95c69a1),
	.w8(32'hba58a421),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97031f3),
	.w1(32'h38077a05),
	.w2(32'h39306894),
	.w3(32'hb969f6f9),
	.w4(32'hb823a93e),
	.w5(32'hb8e408f2),
	.w6(32'hb960853c),
	.w7(32'h38ecd9be),
	.w8(32'h380d3716),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b329995),
	.w1(32'h3b13e359),
	.w2(32'h3aace7dd),
	.w3(32'hb8d38fd2),
	.w4(32'h39b15c08),
	.w5(32'hbaa1ae9b),
	.w6(32'h39cd96da),
	.w7(32'hb9807f84),
	.w8(32'h3883cc43),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91e95d),
	.w1(32'h3b3f1f65),
	.w2(32'hbb5eb83f),
	.w3(32'hba92b43a),
	.w4(32'hb95ffecd),
	.w5(32'hbbbbddcf),
	.w6(32'hbaea9d01),
	.w7(32'hb9dbda87),
	.w8(32'hb94199d3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f779cd),
	.w1(32'h3a1cc473),
	.w2(32'h3882a119),
	.w3(32'hbaf989e8),
	.w4(32'hba803540),
	.w5(32'hba6c5d1e),
	.w6(32'hbac50340),
	.w7(32'hb88a3d32),
	.w8(32'hbaa511c9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa398ac),
	.w1(32'h3a3ebe1b),
	.w2(32'hb99e13b1),
	.w3(32'hba7fbc43),
	.w4(32'hbac23d3f),
	.w5(32'hbae6f112),
	.w6(32'hba9c56fb),
	.w7(32'hb9300d2c),
	.w8(32'hb9e09cac),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69c966),
	.w1(32'h3b151683),
	.w2(32'hba0463dc),
	.w3(32'hb8381f07),
	.w4(32'hb9e9ed42),
	.w5(32'hbb3be633),
	.w6(32'hba925318),
	.w7(32'hbaf216f1),
	.w8(32'h39213768),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33d0ea),
	.w1(32'h3ac8b21b),
	.w2(32'h3904ad0b),
	.w3(32'h3aab0338),
	.w4(32'h3a753f07),
	.w5(32'h39d43fd5),
	.w6(32'h3a9c7f4d),
	.w7(32'h3a5e07b4),
	.w8(32'h3a881adc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bae06),
	.w1(32'h3abe60c3),
	.w2(32'hb9bae12c),
	.w3(32'hb9beb74b),
	.w4(32'hbad07e37),
	.w5(32'hbb2dce7d),
	.w6(32'hb8d40db8),
	.w7(32'hb9bbe2c8),
	.w8(32'hb97b91b2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39242d4f),
	.w1(32'h3a2ad553),
	.w2(32'h3a19e04f),
	.w3(32'hb913aa3c),
	.w4(32'h39ef3ae5),
	.w5(32'h39701cca),
	.w6(32'h3a076c63),
	.w7(32'h3a28e6d8),
	.w8(32'h3a24e1da),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b846ff),
	.w1(32'hb893e506),
	.w2(32'h372a97bc),
	.w3(32'h3993434d),
	.w4(32'h377dfaf0),
	.w5(32'h37889fae),
	.w6(32'hb75dbfb1),
	.w7(32'h398c2e3d),
	.w8(32'h3903c5df),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b13f9e),
	.w1(32'hb78780a8),
	.w2(32'h38aec80b),
	.w3(32'hb9965b93),
	.w4(32'hb916522a),
	.w5(32'hb9016f10),
	.w6(32'hb90a52e4),
	.w7(32'h39afaa69),
	.w8(32'hb98710d5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5125f),
	.w1(32'h39e7896b),
	.w2(32'h3a44e8c5),
	.w3(32'hb9f1ae2e),
	.w4(32'h39f365b0),
	.w5(32'h3a110870),
	.w6(32'h39c1d8b8),
	.w7(32'h3a2ed314),
	.w8(32'h3a1a5ece),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4b863),
	.w1(32'h3b52609d),
	.w2(32'h3ab32213),
	.w3(32'hba3e5c32),
	.w4(32'h3b22da3f),
	.w5(32'h3ab2108c),
	.w6(32'h370744a8),
	.w7(32'h3b1f7de7),
	.w8(32'h39d7f0aa),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24a6ff),
	.w1(32'h38ffef43),
	.w2(32'h382e4135),
	.w3(32'h3a2b3094),
	.w4(32'h3964fc3b),
	.w5(32'h393b59d5),
	.w6(32'h3a0ba97c),
	.w7(32'h39b71bb1),
	.w8(32'h39ff536f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2102e),
	.w1(32'hba86c168),
	.w2(32'hb8d9a040),
	.w3(32'hbb63636d),
	.w4(32'hbafe8cd1),
	.w5(32'hb7db16e4),
	.w6(32'hbace9052),
	.w7(32'h39d39a59),
	.w8(32'h3a57977b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ff88),
	.w1(32'h3b41148f),
	.w2(32'hba8253dd),
	.w3(32'h3a5a6dbc),
	.w4(32'hbace8fbf),
	.w5(32'hbbaec718),
	.w6(32'h37c51e8e),
	.w7(32'h3a96347b),
	.w8(32'h3b0377ac),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f2627),
	.w1(32'h3aca9844),
	.w2(32'h3b78a3e3),
	.w3(32'hb8a6b00f),
	.w4(32'h3a9d13dd),
	.w5(32'h3af11afc),
	.w6(32'hb99cb2e1),
	.w7(32'h3a3c56af),
	.w8(32'h3a99650a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e94e5),
	.w1(32'h3b97392c),
	.w2(32'h3aa7c0fd),
	.w3(32'h3ab0e5c5),
	.w4(32'h3b15bd49),
	.w5(32'hbb317d1c),
	.w6(32'hbab0d5c2),
	.w7(32'hbb367ace),
	.w8(32'hbae94bd5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd78e2),
	.w1(32'h3b131002),
	.w2(32'h3b35ed70),
	.w3(32'hbafce01a),
	.w4(32'h3a4871de),
	.w5(32'h3a8fc626),
	.w6(32'hbb02f242),
	.w7(32'hb9b006d6),
	.w8(32'hb9cc3287),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4f367),
	.w1(32'hba734123),
	.w2(32'hbb77378a),
	.w3(32'hbb59e3f7),
	.w4(32'hbb8e6796),
	.w5(32'hbbad916d),
	.w6(32'hbb1a41b9),
	.w7(32'hbac485e8),
	.w8(32'hb8c53eb2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a800ddb),
	.w1(32'hb928890a),
	.w2(32'h389e0713),
	.w3(32'hbab462c3),
	.w4(32'hbab259d3),
	.w5(32'hbab1e41c),
	.w6(32'hba2d9e64),
	.w7(32'hba5bf6cc),
	.w8(32'h3a5032c9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb631666),
	.w1(32'hba6ec91b),
	.w2(32'h3a706212),
	.w3(32'hbb9c297f),
	.w4(32'hbb00a9a0),
	.w5(32'h3948735c),
	.w6(32'hbb846683),
	.w7(32'hba9fdfb8),
	.w8(32'hbaa0f45c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba567c35),
	.w1(32'hb9fb68d6),
	.w2(32'hb80b16ac),
	.w3(32'hba1fec3f),
	.w4(32'hba30af08),
	.w5(32'hba6ee70c),
	.w6(32'hb9914de1),
	.w7(32'hb9e70acb),
	.w8(32'hb98e5d6f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c5946),
	.w1(32'h3a8126b8),
	.w2(32'hba53d01c),
	.w3(32'hbb69b5ab),
	.w4(32'hbb257249),
	.w5(32'hbb7e09cb),
	.w6(32'hba918e3f),
	.w7(32'h3a4f151c),
	.w8(32'h3a93e8dd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9abb81),
	.w1(32'h3b5e1b4e),
	.w2(32'h3b0745f6),
	.w3(32'h39f08cdd),
	.w4(32'h3ac7097e),
	.w5(32'hbb1e69df),
	.w6(32'hbaebdb84),
	.w7(32'hbb16e1bb),
	.w8(32'hb8d2a9da),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39776ac6),
	.w1(32'h3b23970a),
	.w2(32'hbb1b9e97),
	.w3(32'hbbaa825d),
	.w4(32'h39f6238f),
	.w5(32'hbb95df8f),
	.w6(32'h3ab847d9),
	.w7(32'h3bbfd955),
	.w8(32'h3ba7df46),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fe8c8),
	.w1(32'h3c0b84de),
	.w2(32'h3b767cbb),
	.w3(32'hbb1cebfb),
	.w4(32'h3ba7fade),
	.w5(32'h3b0738b5),
	.w6(32'hba71157b),
	.w7(32'h3b5c0954),
	.w8(32'h3b1552c5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2cee8),
	.w1(32'h3aa178ff),
	.w2(32'h3b04cdc9),
	.w3(32'hbb824395),
	.w4(32'hb72e7ce6),
	.w5(32'h3aa7a09b),
	.w6(32'hbb240545),
	.w7(32'h3a2b7cdd),
	.w8(32'hb99562f9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b658a10),
	.w1(32'h3b01157d),
	.w2(32'hba20d85b),
	.w3(32'hbaca88a7),
	.w4(32'hb7e77cda),
	.w5(32'hbba31153),
	.w6(32'hbb1e5115),
	.w7(32'hbb099d74),
	.w8(32'hba11c254),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83334e),
	.w1(32'hbaff690f),
	.w2(32'hba144c62),
	.w3(32'hb95f0688),
	.w4(32'hbb0cc4c0),
	.w5(32'hbaceeebb),
	.w6(32'hb87a0731),
	.w7(32'hb925b5eb),
	.w8(32'h3a370d1f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f6cd0),
	.w1(32'hba90502a),
	.w2(32'h3a864e06),
	.w3(32'hbbb4be76),
	.w4(32'hb9c991cb),
	.w5(32'hbb81e2de),
	.w6(32'h3a0a8dce),
	.w7(32'h3b32e1b5),
	.w8(32'h3b224e2d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f078a),
	.w1(32'h3ad3a3a8),
	.w2(32'h3a8f48d6),
	.w3(32'h3aa1cc7e),
	.w4(32'h3aecaf82),
	.w5(32'hbb0cab1f),
	.w6(32'hb89f5f43),
	.w7(32'hb951fb55),
	.w8(32'hbb166c4c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949a3ea),
	.w1(32'hb9368578),
	.w2(32'h377ef54a),
	.w3(32'hb92f4aaf),
	.w4(32'hb9b94149),
	.w5(32'hba07fca1),
	.w6(32'h38250e1a),
	.w7(32'h39b4e911),
	.w8(32'h392a5260),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8299baf),
	.w1(32'h36df8ab8),
	.w2(32'hba8986df),
	.w3(32'hba57bb85),
	.w4(32'hb9dfdc8f),
	.w5(32'hba4020d5),
	.w6(32'h3a303db9),
	.w7(32'h3a1798ec),
	.w8(32'hb845ed5d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa58f69),
	.w1(32'h39e5f0dc),
	.w2(32'hba05f0a6),
	.w3(32'hbb17dfa6),
	.w4(32'hbb030912),
	.w5(32'hbb45a94f),
	.w6(32'hbb272cb7),
	.w7(32'hba3dbb25),
	.w8(32'hba47598a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10b0ed),
	.w1(32'h3abe26f9),
	.w2(32'h3b26380c),
	.w3(32'hbb6e25a9),
	.w4(32'h37f305b1),
	.w5(32'h3a9690bf),
	.w6(32'hbb27f438),
	.w7(32'h3a5a7884),
	.w8(32'h3aaf87c9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6655f3),
	.w1(32'hb8965743),
	.w2(32'h3ad2c18d),
	.w3(32'hbb1517d7),
	.w4(32'hba5cc104),
	.w5(32'hb7750a90),
	.w6(32'hbb297410),
	.w7(32'hba9ad640),
	.w8(32'h3a1a9043),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fab2d),
	.w1(32'hb9fdf809),
	.w2(32'h3900ae66),
	.w3(32'hbb0552d2),
	.w4(32'hba0f851a),
	.w5(32'h39b148b1),
	.w6(32'h39dd1491),
	.w7(32'h3a8a3b07),
	.w8(32'h3ab506f3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b242b8a),
	.w1(32'h3b1276cd),
	.w2(32'hba813959),
	.w3(32'hbb476cd2),
	.w4(32'hbb0f8fa7),
	.w5(32'hbaf561a1),
	.w6(32'hb9a6c82c),
	.w7(32'h3a881089),
	.w8(32'h3a2d082f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c2a29),
	.w1(32'hbaa0f214),
	.w2(32'hbb19e053),
	.w3(32'hb88313f6),
	.w4(32'hbb02f15e),
	.w5(32'hbb57c70d),
	.w6(32'hba35aba5),
	.w7(32'hbad56980),
	.w8(32'hba1b8e03),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39996b04),
	.w1(32'h3ae3ee17),
	.w2(32'h3aed707a),
	.w3(32'hbaa03353),
	.w4(32'h3a0ca23d),
	.w5(32'h3a31bacb),
	.w6(32'h39e01751),
	.w7(32'h3aab8e69),
	.w8(32'h3a9ea9eb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73a436),
	.w1(32'hb8982141),
	.w2(32'hb9a6a29e),
	.w3(32'h3a3a6318),
	.w4(32'h3939532e),
	.w5(32'hb9331155),
	.w6(32'h382f5531),
	.w7(32'hb92dcaa5),
	.w8(32'h38db4bcd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886f33e),
	.w1(32'hba2d1761),
	.w2(32'hba809c15),
	.w3(32'h38ca5721),
	.w4(32'hb9f89f2d),
	.w5(32'hba494e9f),
	.w6(32'hb78a9a72),
	.w7(32'hb9b280fd),
	.w8(32'hba025e17),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b59d91),
	.w1(32'hb9ec2441),
	.w2(32'hba10f8d5),
	.w3(32'hb9938c8a),
	.w4(32'hb9ac8733),
	.w5(32'hb9ecbd97),
	.w6(32'hb9a9f0c7),
	.w7(32'hb9db4182),
	.w8(32'hb99eb926),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba6e2d),
	.w1(32'hb9b5f98f),
	.w2(32'hba3f9d7b),
	.w3(32'hb984dfca),
	.w4(32'h3988442a),
	.w5(32'h395ce4c9),
	.w6(32'hb9d553e0),
	.w7(32'hb88c35d8),
	.w8(32'hb9e2ca72),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb855c6ee),
	.w1(32'h3ad49050),
	.w2(32'h3a7b1d6a),
	.w3(32'hba7a2a92),
	.w4(32'hb98ccfe8),
	.w5(32'hba24ec4e),
	.w6(32'hba22cb93),
	.w7(32'hb94fbbe4),
	.w8(32'hba7c170c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba173037),
	.w1(32'hba1adc59),
	.w2(32'hba5833f4),
	.w3(32'hb9e61898),
	.w4(32'hba543df5),
	.w5(32'hba5b4e05),
	.w6(32'hb90ca27c),
	.w7(32'hb9d9a57d),
	.w8(32'hb95f0fbb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedc294),
	.w1(32'h3a8be745),
	.w2(32'hb9910702),
	.w3(32'hba96faa7),
	.w4(32'hbaeaa376),
	.w5(32'hbb042969),
	.w6(32'hbab6ceb1),
	.w7(32'hbab531a0),
	.w8(32'hb98f0b00),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb161860),
	.w1(32'h3a7d5b2d),
	.w2(32'h3af3c6c8),
	.w3(32'hbb3c3640),
	.w4(32'hba0bdb31),
	.w5(32'h3aa9996d),
	.w6(32'hbb0fa688),
	.w7(32'h38e845da),
	.w8(32'h386ed9e8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e68e6),
	.w1(32'hba66de09),
	.w2(32'hba8f6577),
	.w3(32'hb9109b08),
	.w4(32'h39c7273e),
	.w5(32'h394bfa24),
	.w6(32'hb9250406),
	.w7(32'h38d84607),
	.w8(32'hba80c9cd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6eb111),
	.w1(32'h37d9e078),
	.w2(32'h399e747f),
	.w3(32'h3806ae51),
	.w4(32'h3993413e),
	.w5(32'h39aada28),
	.w6(32'h3a2a525e),
	.w7(32'h39239728),
	.w8(32'h3a0fc1c4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49d205),
	.w1(32'hb98d0b55),
	.w2(32'hb9a61915),
	.w3(32'h3a164de4),
	.w4(32'hb9477eb5),
	.w5(32'hb93c4912),
	.w6(32'h38ef9266),
	.w7(32'hb8e249f4),
	.w8(32'h39455132),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf3140),
	.w1(32'hb9eec5b8),
	.w2(32'hb8c8d7d7),
	.w3(32'hb910b1f2),
	.w4(32'hba08a124),
	.w5(32'h38374a63),
	.w6(32'hb9958512),
	.w7(32'hb9db734b),
	.w8(32'h388b218d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e22d7),
	.w1(32'h3af7d345),
	.w2(32'hbb905684),
	.w3(32'hbb6ee18f),
	.w4(32'hbba14ac9),
	.w5(32'hbc024aa7),
	.w6(32'hb98bd70e),
	.w7(32'hb905b005),
	.w8(32'hba5e92b0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0568e8),
	.w1(32'h3ad0386f),
	.w2(32'hb9c41117),
	.w3(32'hba9bea94),
	.w4(32'hbae8fcd7),
	.w5(32'hbb4ee0ec),
	.w6(32'hbb362e51),
	.w7(32'hba8888ce),
	.w8(32'hba3aab40),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e4250),
	.w1(32'h3a0d5e08),
	.w2(32'h38cf866f),
	.w3(32'h39ae6a23),
	.w4(32'h374cdf53),
	.w5(32'hba09d218),
	.w6(32'hb8f1646a),
	.w7(32'hb96a18d8),
	.w8(32'hb8bb5503),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965507a),
	.w1(32'hba4d666f),
	.w2(32'hbac5b031),
	.w3(32'hba7ad097),
	.w4(32'hba4194e3),
	.w5(32'hba46120e),
	.w6(32'h3a2a53a2),
	.w7(32'h3a495e98),
	.w8(32'hb94ef0e0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b91518),
	.w1(32'h3a3b7921),
	.w2(32'h3a322f37),
	.w3(32'hb92b1c3f),
	.w4(32'h3a099b90),
	.w5(32'h394411db),
	.w6(32'h373ef5d4),
	.w7(32'h3a1f66cf),
	.w8(32'h392a6e7f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961aaa2),
	.w1(32'h3852520a),
	.w2(32'hba833c8e),
	.w3(32'hbaae09ad),
	.w4(32'hbad5e0c9),
	.w5(32'hbab0590d),
	.w6(32'hba873d24),
	.w7(32'hba082917),
	.w8(32'hb8a70d67),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1220a),
	.w1(32'hbabadfe6),
	.w2(32'hba75c5a4),
	.w3(32'h3982930e),
	.w4(32'hba84b6d1),
	.w5(32'h3940c602),
	.w6(32'h3a895102),
	.w7(32'h38f44bc1),
	.w8(32'h39f6f10d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8679f5),
	.w1(32'h3b21e7d8),
	.w2(32'hba81a421),
	.w3(32'hba096e39),
	.w4(32'hbb4d31e3),
	.w5(32'hbbbde0c7),
	.w6(32'hbb41e80c),
	.w7(32'hbaf706c6),
	.w8(32'h38a0e1bc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c9039),
	.w1(32'h3a9aa4db),
	.w2(32'h3abaa860),
	.w3(32'hbb0bc805),
	.w4(32'h3a14231b),
	.w5(32'h3a361d4b),
	.w6(32'hba96cfda),
	.w7(32'h3a1127f9),
	.w8(32'h397a199b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a826a29),
	.w1(32'h388d33b8),
	.w2(32'hb9b5970a),
	.w3(32'hb937f43a),
	.w4(32'hba9066d6),
	.w5(32'hbae58ef1),
	.w6(32'hbb1e7557),
	.w7(32'hba923cff),
	.w8(32'h398ed8f4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72418b),
	.w1(32'h3b048fc5),
	.w2(32'hb99decbe),
	.w3(32'hba04c416),
	.w4(32'hbaae2135),
	.w5(32'hbb736e84),
	.w6(32'hba5e338d),
	.w7(32'hb9ecdc07),
	.w8(32'h3a63a225),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad44ea),
	.w1(32'h3a5b2cc6),
	.w2(32'hba41621a),
	.w3(32'hbb1efa52),
	.w4(32'h39a00bf3),
	.w5(32'hb9f3d7f8),
	.w6(32'h39d09ac1),
	.w7(32'h3aed6127),
	.w8(32'h391e3028),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b157a30),
	.w1(32'h3aacf65b),
	.w2(32'hb960c8ad),
	.w3(32'hb8a7d0bf),
	.w4(32'hb8d5e787),
	.w5(32'hbae97cda),
	.w6(32'hba93a447),
	.w7(32'hba77cbb5),
	.w8(32'hba151cb5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370296d8),
	.w1(32'hb6c7984a),
	.w2(32'hb9356969),
	.w3(32'hba08a167),
	.w4(32'hb9ce3a1a),
	.w5(32'hb9c9fc50),
	.w6(32'hb9d5d800),
	.w7(32'hb94890e7),
	.w8(32'hb960d2d2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f9f07),
	.w1(32'h3a53f1e8),
	.w2(32'h3b62bf6a),
	.w3(32'hbbc73088),
	.w4(32'hbb3283bf),
	.w5(32'hb6b50df2),
	.w6(32'hbba58292),
	.w7(32'hbaed5b2f),
	.w8(32'hba43268c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3566e),
	.w1(32'h3989c972),
	.w2(32'hb9e02ac4),
	.w3(32'hbac3c495),
	.w4(32'hba66cd5a),
	.w5(32'hba3e45de),
	.w6(32'hba4ede02),
	.w7(32'h36bba9d1),
	.w8(32'h39da753b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387ddf24),
	.w1(32'h37b15aed),
	.w2(32'hb84d7b09),
	.w3(32'hb797fa98),
	.w4(32'hb852d595),
	.w5(32'hb84e0f1b),
	.w6(32'h380aa80e),
	.w7(32'hb7d2156d),
	.w8(32'hb8713fe2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e9a98),
	.w1(32'hb7fff3df),
	.w2(32'h37c6088e),
	.w3(32'hb7d32083),
	.w4(32'hb6d455a5),
	.w5(32'h36adf593),
	.w6(32'hb7f32a88),
	.w7(32'hb737b34a),
	.w8(32'hb76b78b0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab58d66),
	.w1(32'h3a61b1b7),
	.w2(32'h3a79cc29),
	.w3(32'h39acfe21),
	.w4(32'h3a84cf6f),
	.w5(32'hb8795689),
	.w6(32'hb80fad3b),
	.w7(32'hb82f848a),
	.w8(32'h3847d666),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75afb8),
	.w1(32'h39970cea),
	.w2(32'hb9123fb0),
	.w3(32'hbb1b8e41),
	.w4(32'hba0887c7),
	.w5(32'hbab376ef),
	.w6(32'hbb244cb8),
	.w7(32'h388ce4ef),
	.w8(32'hbabe9841),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3369a),
	.w1(32'h3a78b33e),
	.w2(32'hba85cbe0),
	.w3(32'hbb14518c),
	.w4(32'hbb09c3a4),
	.w5(32'hbb394e9f),
	.w6(32'hbb30efc9),
	.w7(32'hbad5c61a),
	.w8(32'hbb30749b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74dc2ba),
	.w1(32'hb7324872),
	.w2(32'hb70f8235),
	.w3(32'h3792397f),
	.w4(32'hb63024fd),
	.w5(32'h3658f7d5),
	.w6(32'h36f430a0),
	.w7(32'h35abfa89),
	.w8(32'h37664253),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b477027),
	.w1(32'h3b1b8631),
	.w2(32'h396a86f9),
	.w3(32'hba8c3141),
	.w4(32'hba18f472),
	.w5(32'hbb069505),
	.w6(32'hbb0918cb),
	.w7(32'hba8809a0),
	.w8(32'hbaa9e4f3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9850936),
	.w1(32'h399173f4),
	.w2(32'h3a90cb4b),
	.w3(32'hbae2ee51),
	.w4(32'hb9da254f),
	.w5(32'h3a293641),
	.w6(32'hbac854a6),
	.w7(32'h3902778a),
	.w8(32'h3a711ec5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cde22),
	.w1(32'h3af27b5c),
	.w2(32'hba44732e),
	.w3(32'hba2580db),
	.w4(32'hbabc6ac1),
	.w5(32'hbb68a862),
	.w6(32'hbae208c7),
	.w7(32'hbb15ab7d),
	.w8(32'hba912ca4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5557d7),
	.w1(32'h3a77eb77),
	.w2(32'h3b548ea0),
	.w3(32'hbb928c2b),
	.w4(32'h389061a1),
	.w5(32'h3ac90432),
	.w6(32'hbb42b6e3),
	.w7(32'hbb370265),
	.w8(32'hba2623ca),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9acd3),
	.w1(32'hb8118e96),
	.w2(32'hbac58c5b),
	.w3(32'hba103527),
	.w4(32'hb92543a5),
	.w5(32'hba5abfda),
	.w6(32'hb90c94df),
	.w7(32'h39d312e2),
	.w8(32'hb61edf7a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7f003),
	.w1(32'hbaa232f7),
	.w2(32'hba767cc8),
	.w3(32'hbb134451),
	.w4(32'hbb10c76d),
	.w5(32'hbacef47a),
	.w6(32'hbad235fd),
	.w7(32'hba704fda),
	.w8(32'hba85c482),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a733f7f),
	.w1(32'h3b2f0dc9),
	.w2(32'h3b32e6fd),
	.w3(32'h3a6ec5ea),
	.w4(32'h3af61485),
	.w5(32'h3b1ed369),
	.w6(32'h3aeec1eb),
	.w7(32'h3b2fb7c6),
	.w8(32'h3b321245),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffdb34),
	.w1(32'h3ac35254),
	.w2(32'h3a3b5398),
	.w3(32'hbaf1266c),
	.w4(32'h39daa008),
	.w5(32'h399e9e94),
	.w6(32'hba86e826),
	.w7(32'h3a51fcc7),
	.w8(32'h39bd0d46),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96e769),
	.w1(32'h3a77002f),
	.w2(32'h3a6f59b6),
	.w3(32'hba03a995),
	.w4(32'h3a69cf8c),
	.w5(32'h3a5dae55),
	.w6(32'hb85c218c),
	.w7(32'h3a46874d),
	.w8(32'h395b49ed),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e6829),
	.w1(32'h3a5f9e2f),
	.w2(32'h37a4874f),
	.w3(32'h39408dcf),
	.w4(32'hb9432a37),
	.w5(32'hba6a1af5),
	.w6(32'hb94a56a5),
	.w7(32'hb9d1eac4),
	.w8(32'hba07671c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3888a1a2),
	.w1(32'h38d37119),
	.w2(32'h382b3cf6),
	.w3(32'h386ac166),
	.w4(32'hb755c061),
	.w5(32'hb8ac05f9),
	.w6(32'h3917a99c),
	.w7(32'h38f22daa),
	.w8(32'hb8aacd3c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b2748),
	.w1(32'h39a6beeb),
	.w2(32'hba274b10),
	.w3(32'hba819101),
	.w4(32'hbac34d4d),
	.w5(32'hbb2ea020),
	.w6(32'hba8796e1),
	.w7(32'hba18bda9),
	.w8(32'h3a0df4e9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a976e88),
	.w1(32'h3a7b5211),
	.w2(32'hb971f978),
	.w3(32'h3a41fccb),
	.w4(32'h39e07578),
	.w5(32'hba811cd8),
	.w6(32'hb98b4306),
	.w7(32'hb9a59ab4),
	.w8(32'hba328571),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a253e),
	.w1(32'h395504b3),
	.w2(32'h3a9a085d),
	.w3(32'hbab87a63),
	.w4(32'hba86783b),
	.w5(32'h3a7d7190),
	.w6(32'h38e589ef),
	.w7(32'h39243f7d),
	.w8(32'h3aa1616f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38108fa7),
	.w1(32'hb8ca12f2),
	.w2(32'h391132ed),
	.w3(32'h394055aa),
	.w4(32'h3852d1af),
	.w5(32'h35a7afd1),
	.w6(32'hb8a208e3),
	.w7(32'hb9995d65),
	.w8(32'hb9dad112),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad43c8),
	.w1(32'hb997c821),
	.w2(32'hba826afc),
	.w3(32'hb9c2ff9a),
	.w4(32'hbb42d01f),
	.w5(32'hbb4923ae),
	.w6(32'hba425e52),
	.w7(32'hbb1bf67e),
	.w8(32'hba910ee3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82c4109),
	.w1(32'hb974dc3a),
	.w2(32'hb948dc07),
	.w3(32'hb8f61718),
	.w4(32'hb994e232),
	.w5(32'hb990d548),
	.w6(32'hb9090ae5),
	.w7(32'hb95db41d),
	.w8(32'hb937f65a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6f7f6),
	.w1(32'hb957dd36),
	.w2(32'hb8e16bb2),
	.w3(32'hb9b271af),
	.w4(32'hb9a33535),
	.w5(32'hb9263ba8),
	.w6(32'hb94fe627),
	.w7(32'hb9481525),
	.w8(32'hb8cb69a6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe2099),
	.w1(32'hb925ab38),
	.w2(32'h39fc004e),
	.w3(32'hbad3ea26),
	.w4(32'hb9ad854e),
	.w5(32'h392ad92b),
	.w6(32'hba6d98bc),
	.w7(32'h39939168),
	.w8(32'h3a01f9fc),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e09a4),
	.w1(32'h3b92eccb),
	.w2(32'h3aaae306),
	.w3(32'hbaf4a4cc),
	.w4(32'hb9670936),
	.w5(32'hbb1158f2),
	.w6(32'h3a69717e),
	.w7(32'h3b2a36f6),
	.w8(32'h3b3afb10),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e42295),
	.w1(32'hb8d38209),
	.w2(32'h39dabed3),
	.w3(32'h39325cea),
	.w4(32'h38e87bb8),
	.w5(32'h39aa0609),
	.w6(32'h38da83de),
	.w7(32'hb9b7ca83),
	.w8(32'hb9cf1811),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6546f),
	.w1(32'h391ce8d1),
	.w2(32'h3996a459),
	.w3(32'hbb143680),
	.w4(32'hbaad2b62),
	.w5(32'hb9e7c75c),
	.w6(32'hbad44487),
	.w7(32'hb9ba4502),
	.w8(32'hb9bbb866),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dca1d),
	.w1(32'h3a8aa2c1),
	.w2(32'h3a48117c),
	.w3(32'h373917fa),
	.w4(32'hb8ecb644),
	.w5(32'hba1c54a1),
	.w6(32'h398aadb5),
	.w7(32'hb98f9ff0),
	.w8(32'h3a19d25a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2af589),
	.w1(32'h3ac381bc),
	.w2(32'hbaf91a4b),
	.w3(32'hbb5958fe),
	.w4(32'hbb129d4c),
	.w5(32'hbb82ce49),
	.w6(32'hbb5298b7),
	.w7(32'hbae99206),
	.w8(32'hbacc3322),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b6796),
	.w1(32'h3aa3d05a),
	.w2(32'h38df0a24),
	.w3(32'h3a51c0b2),
	.w4(32'hba5675b1),
	.w5(32'hbad29794),
	.w6(32'h3a030d46),
	.w7(32'h373347b5),
	.w8(32'h3877ec46),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b447785),
	.w1(32'h3a9ec9ca),
	.w2(32'hb954c3f3),
	.w3(32'hba8bb035),
	.w4(32'hbaf1a041),
	.w5(32'hbb173a3f),
	.w6(32'hbac1b112),
	.w7(32'hb9457b91),
	.w8(32'h3a6cbd45),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984b70e),
	.w1(32'hba13b406),
	.w2(32'hb9eb0db9),
	.w3(32'hb9f67c5b),
	.w4(32'hba2a4727),
	.w5(32'hba18190e),
	.w6(32'hba1472bd),
	.w7(32'hba59ac4f),
	.w8(32'hba549fd8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f31c4),
	.w1(32'hb9a48ca0),
	.w2(32'hba223fa2),
	.w3(32'hba9a89b8),
	.w4(32'hba999db1),
	.w5(32'hbac144c9),
	.w6(32'hbaa065a5),
	.w7(32'hb9dcd50f),
	.w8(32'h3a2fc32a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79630e2),
	.w1(32'hb857d122),
	.w2(32'hb827a4ec),
	.w3(32'hb7710f3e),
	.w4(32'hb80e56c6),
	.w5(32'hb531e8ae),
	.w6(32'hb794e083),
	.w7(32'hb7924d98),
	.w8(32'hb72f0abe),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddbf3f),
	.w1(32'h3a335692),
	.w2(32'h3a47382a),
	.w3(32'hb976a025),
	.w4(32'h3866fbbc),
	.w5(32'hb8396af1),
	.w6(32'hb95f07e4),
	.w7(32'hb93e94f0),
	.w8(32'h394917d7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11cc29),
	.w1(32'hba18901f),
	.w2(32'hb96a0403),
	.w3(32'hb98aaef5),
	.w4(32'hb9657de4),
	.w5(32'h39291853),
	.w6(32'hb765838e),
	.w7(32'h383e7b67),
	.w8(32'hb98254d4),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf60ca),
	.w1(32'h36ff1d9d),
	.w2(32'hbb063f47),
	.w3(32'hba384855),
	.w4(32'hbace2e6e),
	.w5(32'hbb179b07),
	.w6(32'hbad37447),
	.w7(32'hba8bc7f3),
	.w8(32'h394a93b5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb770f882),
	.w1(32'hb72d5d86),
	.w2(32'hb73899a5),
	.w3(32'hb6edf28d),
	.w4(32'h363720f4),
	.w5(32'h366db30a),
	.w6(32'hb70ac415),
	.w7(32'hb705f05b),
	.w8(32'hb6838000),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4d7a2),
	.w1(32'hb898bf21),
	.w2(32'h3691030d),
	.w3(32'hb8833467),
	.w4(32'hb8869094),
	.w5(32'h37792a6c),
	.w6(32'hb7c34a47),
	.w7(32'h382313c0),
	.w8(32'h39232e9f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8eba03),
	.w1(32'hba2546c6),
	.w2(32'hb9b37868),
	.w3(32'hbaa6ae0c),
	.w4(32'hba856efa),
	.w5(32'h39693b86),
	.w6(32'h3a4d6604),
	.w7(32'h39f07d30),
	.w8(32'h3aa2902e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac43d6f),
	.w1(32'hba5fcf3b),
	.w2(32'hbaa86c17),
	.w3(32'hb9c0db5d),
	.w4(32'hbb0dbabb),
	.w5(32'hbb4e08b6),
	.w6(32'h3a48aabb),
	.w7(32'hb905b177),
	.w8(32'h3a98691b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ee6d3),
	.w1(32'h3aea51e8),
	.w2(32'h391fb93c),
	.w3(32'hbb470e28),
	.w4(32'h3a88cbdc),
	.w5(32'hbaa8dd3e),
	.w6(32'hbb4d72c9),
	.w7(32'h3a3a2247),
	.w8(32'hb9daf206),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ac94f6),
	.w1(32'hb940c52e),
	.w2(32'hb8cbcd7c),
	.w3(32'hb9bc1679),
	.w4(32'hb9b4d3f5),
	.w5(32'hba1d7e9d),
	.w6(32'hb76040e8),
	.w7(32'hb994e05d),
	.w8(32'hb9be77ec),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc165a4),
	.w1(32'h3ad40dd4),
	.w2(32'hbb982239),
	.w3(32'hbb56f542),
	.w4(32'hbb9605d4),
	.w5(32'hbbd81405),
	.w6(32'hba92b112),
	.w7(32'hbaad1e6c),
	.w8(32'hba9091d4),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0824eb),
	.w1(32'h3ba760fd),
	.w2(32'h3b4e1dfc),
	.w3(32'hba573cd0),
	.w4(32'h3b3907b5),
	.w5(32'h3a50bf0c),
	.w6(32'hbadd3808),
	.w7(32'h3830fd62),
	.w8(32'h3abb4323),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7ad4d),
	.w1(32'h3a89e795),
	.w2(32'h379cc384),
	.w3(32'h3a246f40),
	.w4(32'h3a0259c9),
	.w5(32'hba9a86b5),
	.w6(32'hba18bed6),
	.w7(32'hba7b5828),
	.w8(32'hba9f1d36),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b517c2),
	.w1(32'hb81e724c),
	.w2(32'hb84ba406),
	.w3(32'h3759fc10),
	.w4(32'hb828d14e),
	.w5(32'hb7e211fa),
	.w6(32'hb69d3b01),
	.w7(32'h35cb9f5d),
	.w8(32'h353d09b5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910f636),
	.w1(32'hb81b65bf),
	.w2(32'h39751721),
	.w3(32'hb9431052),
	.w4(32'hb8633bef),
	.w5(32'h399365fe),
	.w6(32'h3845a561),
	.w7(32'h398401de),
	.w8(32'h3a199255),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80b414c),
	.w1(32'hb7dc1b2e),
	.w2(32'hb819bc9b),
	.w3(32'hb7d91fb8),
	.w4(32'hb7be0340),
	.w5(32'hb7ac0946),
	.w6(32'h379ce6b4),
	.w7(32'h36f34a8b),
	.w8(32'hb8029a28),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d5b31),
	.w1(32'h3a864e71),
	.w2(32'hba5445e3),
	.w3(32'hb8ed6b75),
	.w4(32'hb992bfca),
	.w5(32'hbb1e9ed2),
	.w6(32'hba82d52e),
	.w7(32'hb9c42b8e),
	.w8(32'hba216674),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f6f30),
	.w1(32'h3a0739f1),
	.w2(32'hb8a731b4),
	.w3(32'hbae9a6e6),
	.w4(32'hbac6e894),
	.w5(32'hbab041bc),
	.w6(32'hb9bd6753),
	.w7(32'h39010aba),
	.w8(32'h39b42b0d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab781cf),
	.w1(32'h38b5eb38),
	.w2(32'hbaba2ec6),
	.w3(32'hbb4b50ed),
	.w4(32'hbaa03fcd),
	.w5(32'hba927477),
	.w6(32'hbb38321a),
	.w7(32'hba911f4d),
	.w8(32'hbaf6709e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b0f43),
	.w1(32'h39968597),
	.w2(32'hb903bf2f),
	.w3(32'hb9d24303),
	.w4(32'h366503a4),
	.w5(32'h38dc8345),
	.w6(32'h39ff62b4),
	.w7(32'h3a0b9a82),
	.w8(32'h39c64341),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b000b92),
	.w1(32'h3a48be40),
	.w2(32'hba0e5cc7),
	.w3(32'hbaa282b5),
	.w4(32'hbb24090b),
	.w5(32'hbb4de3c5),
	.w6(32'hbb08f322),
	.w7(32'hbac08e56),
	.w8(32'hba2641a1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d46bf),
	.w1(32'h3a63c7bb),
	.w2(32'h38db5b76),
	.w3(32'hb960fb54),
	.w4(32'h3a37c0ee),
	.w5(32'hba3ae86f),
	.w6(32'h39773c13),
	.w7(32'h3a5a78ed),
	.w8(32'hba99c006),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb747abe2),
	.w1(32'hb791782a),
	.w2(32'hb7220ec8),
	.w3(32'h37875e1a),
	.w4(32'h36adc8a7),
	.w5(32'h36dab7c1),
	.w6(32'hb7286778),
	.w7(32'hb6c5295d),
	.w8(32'hb7168816),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a28d2),
	.w1(32'hbb147575),
	.w2(32'hba9cb997),
	.w3(32'hb9fa5254),
	.w4(32'hbaa237fe),
	.w5(32'hba82077a),
	.w6(32'h394ab5b5),
	.w7(32'hb9282c04),
	.w8(32'h39c5b225),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb837ab47),
	.w1(32'hb7fdcd11),
	.w2(32'hb76599da),
	.w3(32'h377ffe3b),
	.w4(32'h37c62dfa),
	.w5(32'h38035bc6),
	.w6(32'hb791f334),
	.w7(32'hb617e21d),
	.w8(32'hb72d47bd),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a999321),
	.w1(32'h3a434fe7),
	.w2(32'hb96cd587),
	.w3(32'hbab11397),
	.w4(32'hbacae030),
	.w5(32'hbb191be2),
	.w6(32'hbaac9790),
	.w7(32'hba25b2b3),
	.w8(32'hba451fb8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae70d82),
	.w1(32'h3ac02a87),
	.w2(32'h3a3fc247),
	.w3(32'hba6a50ad),
	.w4(32'h3a37b8f1),
	.w5(32'h3a7bafd9),
	.w6(32'hb909cb7c),
	.w7(32'h3ab179d5),
	.w8(32'hba0eb675),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97d89d7),
	.w1(32'h3a703753),
	.w2(32'h3a68801f),
	.w3(32'hbabb5278),
	.w4(32'hb925a267),
	.w5(32'hb86b3823),
	.w6(32'hb9fed0c1),
	.w7(32'h3a0ca284),
	.w8(32'h389d9397),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904a2e8),
	.w1(32'h3956b997),
	.w2(32'h3864ac08),
	.w3(32'h39fc5b06),
	.w4(32'h39d49c22),
	.w5(32'h3982dd0b),
	.w6(32'h3a082656),
	.w7(32'h39be6cc3),
	.w8(32'h39820a13),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac97565),
	.w1(32'hb9690291),
	.w2(32'h3a0bb207),
	.w3(32'hbb385e23),
	.w4(32'hbaa65a22),
	.w5(32'h3936252e),
	.w6(32'hba22f9ac),
	.w7(32'h39cb176c),
	.w8(32'h39e19a59),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a5c9c),
	.w1(32'h3a2bb433),
	.w2(32'hb9856b0d),
	.w3(32'hba85a200),
	.w4(32'hba3d84a5),
	.w5(32'hbab5f76c),
	.w6(32'hbabfe270),
	.w7(32'hba49dd22),
	.w8(32'hb94603ca),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3833f6),
	.w1(32'h3ade0052),
	.w2(32'hbaa7fdf9),
	.w3(32'hbae42931),
	.w4(32'hbaced39b),
	.w5(32'hbb544dfa),
	.w6(32'hbb2eb3d4),
	.w7(32'hbafff141),
	.w8(32'hbb1fc042),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb725788f),
	.w1(32'hb7983c9a),
	.w2(32'h37889b9e),
	.w3(32'hb7d79ded),
	.w4(32'hb77b86c0),
	.w5(32'h373514f6),
	.w6(32'hb8038ec9),
	.w7(32'h3594dafc),
	.w8(32'h3829527a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3831cc61),
	.w1(32'h37660599),
	.w2(32'h3826dc69),
	.w3(32'h37acb0c3),
	.w4(32'hb8ac2065),
	.w5(32'hb9180960),
	.w6(32'hb7cd3da6),
	.w7(32'h36758ea2),
	.w8(32'hb87742c9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09ab32),
	.w1(32'h3b271cf1),
	.w2(32'h390b1888),
	.w3(32'hbb0e670f),
	.w4(32'hbafb27bb),
	.w5(32'hbb2aa3bc),
	.w6(32'h3aab8f85),
	.w7(32'h3ad48b68),
	.w8(32'h3a925ed8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fcfd8),
	.w1(32'h3ab7ec1b),
	.w2(32'h39bdea69),
	.w3(32'hbb25d792),
	.w4(32'hbaaff140),
	.w5(32'hbadf5776),
	.w6(32'h3b00a7a6),
	.w7(32'h3b331413),
	.w8(32'h3b407d69),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98936d8),
	.w1(32'h3acb7457),
	.w2(32'h3aaba00c),
	.w3(32'hbaf6dbe5),
	.w4(32'h3884657c),
	.w5(32'h3a384644),
	.w6(32'h39343097),
	.w7(32'h3a94dd16),
	.w8(32'h3ab85507),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb60202),
	.w1(32'h3b632fa5),
	.w2(32'h39957aa3),
	.w3(32'h3a885cdf),
	.w4(32'hb9a44495),
	.w5(32'hbb96f576),
	.w6(32'hbac2c70c),
	.w7(32'hbb384452),
	.w8(32'hbae1afcb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398df4d6),
	.w1(32'hb92218d0),
	.w2(32'hb9f6c57a),
	.w3(32'h3689ef5c),
	.w4(32'hb9e7cb78),
	.w5(32'hb9ca3bd7),
	.w6(32'hb93c7b35),
	.w7(32'hb8bc226d),
	.w8(32'hb6e28a18),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63985c),
	.w1(32'hb81dc2c5),
	.w2(32'hba839b3b),
	.w3(32'h389edac7),
	.w4(32'hb9d5da29),
	.w5(32'hba33139e),
	.w6(32'h3a0a3596),
	.w7(32'h399834ca),
	.w8(32'h38906e42),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bb4ee),
	.w1(32'h3bf3e36c),
	.w2(32'hbadd4fba),
	.w3(32'hb9f311f8),
	.w4(32'h3b745ece),
	.w5(32'hbbbd6661),
	.w6(32'h39fb32b4),
	.w7(32'h3b323485),
	.w8(32'hbac6893c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b663fa6),
	.w1(32'h3964522d),
	.w2(32'hbba5d6eb),
	.w3(32'hbb5476e8),
	.w4(32'hbb7cca79),
	.w5(32'hbbcbf722),
	.w6(32'hba9488e3),
	.w7(32'hba76b8a3),
	.w8(32'hba97c4cc),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b611b29),
	.w1(32'h3b502a7b),
	.w2(32'hb98ebc62),
	.w3(32'hbaff4b4d),
	.w4(32'hba8a149a),
	.w5(32'hbb5066ca),
	.w6(32'hbb240a20),
	.w7(32'hb9e2ab2a),
	.w8(32'h39e7fc4e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0441e1),
	.w1(32'h3ab401b0),
	.w2(32'h3afc9b25),
	.w3(32'hbaf2426b),
	.w4(32'h3aa75f4f),
	.w5(32'h3ac0e873),
	.w6(32'hba96b361),
	.w7(32'h3a7290e9),
	.w8(32'hb9740875),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79383a),
	.w1(32'h3abf768d),
	.w2(32'h3b090fc1),
	.w3(32'hba0183a5),
	.w4(32'h3a863da6),
	.w5(32'h3b1309b3),
	.w6(32'hb82f8307),
	.w7(32'h3ac93055),
	.w8(32'h3ac72a01),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb773b638),
	.w1(32'hb69585bd),
	.w2(32'hb702461b),
	.w3(32'hb7220544),
	.w4(32'hb66f8f09),
	.w5(32'h340ad6f2),
	.w6(32'hb704da28),
	.w7(32'hb7516806),
	.w8(32'hb7969038),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bb9cd4),
	.w1(32'hb716e760),
	.w2(32'hb74ba51d),
	.w3(32'h36f56576),
	.w4(32'h36fd6811),
	.w5(32'h36e6ffc5),
	.w6(32'hb6cb6ed9),
	.w7(32'hb6ac577f),
	.w8(32'hb51017d8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c4a5b),
	.w1(32'h3a6f2e71),
	.w2(32'h394dd40e),
	.w3(32'hba079da2),
	.w4(32'hba6dd12f),
	.w5(32'hba9a1d88),
	.w6(32'h3820abc9),
	.w7(32'h39af41e9),
	.w8(32'h39d57c36),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7729a6b),
	.w1(32'hb7b97076),
	.w2(32'hb78ad808),
	.w3(32'h37473efc),
	.w4(32'hb7a784d2),
	.w5(32'hb719d990),
	.w6(32'h372c0c78),
	.w7(32'hb6f12040),
	.w8(32'hb7a175ed),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada0106),
	.w1(32'h3a23276a),
	.w2(32'hbab74da3),
	.w3(32'h3aa249d9),
	.w4(32'hba10c691),
	.w5(32'hbb2319b8),
	.w6(32'h3a66fd30),
	.w7(32'hb9aa39af),
	.w8(32'hba7cc642),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997cea4),
	.w1(32'h3a419898),
	.w2(32'hba6c766d),
	.w3(32'hbb1b7acd),
	.w4(32'hba15daf0),
	.w5(32'hbac323b8),
	.w6(32'h3a38fa56),
	.w7(32'h3af9d037),
	.w8(32'h3ad4f534),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f629fa),
	.w1(32'h3a8e3594),
	.w2(32'h3a2d6a96),
	.w3(32'hba4688db),
	.w4(32'hb9e04a41),
	.w5(32'hb9aad731),
	.w6(32'hb9a2df95),
	.w7(32'h3998f1b1),
	.w8(32'h3a40a275),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ab1473),
	.w1(32'hb81f0d69),
	.w2(32'hb765a6c8),
	.w3(32'h34da9ca8),
	.w4(32'hb7aab16e),
	.w5(32'h345d4f68),
	.w6(32'hb6ad1e64),
	.w7(32'hb530043f),
	.w8(32'h3604708a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babd38e),
	.w1(32'h3b7eb684),
	.w2(32'hba6c5d34),
	.w3(32'hbb2a871d),
	.w4(32'hbb17b55e),
	.w5(32'hbb926513),
	.w6(32'hbaf1c8c6),
	.w7(32'hb7f6cfff),
	.w8(32'h3b0a8144),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3cba7),
	.w1(32'h3a8a7f31),
	.w2(32'hb9419068),
	.w3(32'hba3ba7e6),
	.w4(32'hba1c9fd7),
	.w5(32'hbaf28bef),
	.w6(32'hba57e9dd),
	.w7(32'hb9911cf9),
	.w8(32'hb95fe6b2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f75a0),
	.w1(32'hb87fb403),
	.w2(32'hb811c617),
	.w3(32'hb838961c),
	.w4(32'hb83a130c),
	.w5(32'h36c64fef),
	.w6(32'hb85473db),
	.w7(32'hb7d21e55),
	.w8(32'hb76afd62),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b339dee),
	.w1(32'h3acd9180),
	.w2(32'hba15a26a),
	.w3(32'hb8801592),
	.w4(32'hba94679c),
	.w5(32'hbb1881ec),
	.w6(32'hba9b325a),
	.w7(32'hba75e3b5),
	.w8(32'hb913888d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97977ed),
	.w1(32'hb93e020b),
	.w2(32'hb8d3a262),
	.w3(32'hb96f7e18),
	.w4(32'hb92a15cb),
	.w5(32'hb867111b),
	.w6(32'hb90878d6),
	.w7(32'hb88fff0c),
	.w8(32'h367cda4f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e167a),
	.w1(32'h3952dfa9),
	.w2(32'h38e35351),
	.w3(32'h37481f43),
	.w4(32'h376c91ed),
	.w5(32'hb706f048),
	.w6(32'h38a0b921),
	.w7(32'h36956093),
	.w8(32'h382099a4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73b79b5),
	.w1(32'hb7bcf7bf),
	.w2(32'hb7b2bf01),
	.w3(32'hb4f881a9),
	.w4(32'hb6884b72),
	.w5(32'h367fda58),
	.w6(32'h372490c8),
	.w7(32'h3733962f),
	.w8(32'hb77c9888),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f2f7d4),
	.w1(32'hb6d56b1d),
	.w2(32'h3703fffa),
	.w3(32'hb7bb50bc),
	.w4(32'hb826824c),
	.w5(32'hb5e2295f),
	.w6(32'hb888dffc),
	.w7(32'hb860f5cb),
	.w8(32'hb84f687c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4390ac),
	.w1(32'h3a983533),
	.w2(32'h3a0c14e1),
	.w3(32'hba1159f3),
	.w4(32'h39db7416),
	.w5(32'h396756ab),
	.w6(32'hb93b131a),
	.w7(32'h3a0d2870),
	.w8(32'h386f65ba),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf5292),
	.w1(32'h3b50daa3),
	.w2(32'hb9e085bf),
	.w3(32'h3b39e1c0),
	.w4(32'h39eee4e0),
	.w5(32'hbb56778a),
	.w6(32'hbaa49bad),
	.w7(32'hbb406119),
	.w8(32'hba2eae11),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26c225),
	.w1(32'h3ac60057),
	.w2(32'hba0a1b0a),
	.w3(32'hba2a0315),
	.w4(32'hba75c53d),
	.w5(32'hbb1529e9),
	.w6(32'hbaaf71b3),
	.w7(32'hb9cf962b),
	.w8(32'hb673e800),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44c542),
	.w1(32'h3abb8c00),
	.w2(32'hba03b987),
	.w3(32'hb9357f5e),
	.w4(32'hbada1331),
	.w5(32'hbb75bf78),
	.w6(32'hbb47ae10),
	.w7(32'hbb251a44),
	.w8(32'hba794d8f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8934a6c),
	.w1(32'hb7bd1960),
	.w2(32'hb83185eb),
	.w3(32'hb7fc91cb),
	.w4(32'h372fd07b),
	.w5(32'hb7b51d8d),
	.w6(32'h369ac43e),
	.w7(32'hb6b96939),
	.w8(32'hb818f751),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39048bb2),
	.w1(32'hb9985153),
	.w2(32'hba1309ff),
	.w3(32'hb7857a46),
	.w4(32'hb9858916),
	.w5(32'hb9916071),
	.w6(32'h38c4658a),
	.w7(32'h3790bf2a),
	.w8(32'h388ec52a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370a317c),
	.w1(32'hb5f25283),
	.w2(32'hb7d338fa),
	.w3(32'h37a61e69),
	.w4(32'hb74d504d),
	.w5(32'hb7df3a76),
	.w6(32'h376255f2),
	.w7(32'hb5cecf4e),
	.w8(32'hb807adc3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb726252d),
	.w1(32'hb785ed2b),
	.w2(32'hb6be3c2d),
	.w3(32'h36794080),
	.w4(32'hb686bac2),
	.w5(32'h364d6026),
	.w6(32'h357ae772),
	.w7(32'hb607f94a),
	.w8(32'hb68acb35),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390adf80),
	.w1(32'hbab147e5),
	.w2(32'hbb15a3db),
	.w3(32'hbb21be12),
	.w4(32'hbb3137d6),
	.w5(32'hbb286d69),
	.w6(32'hbaa35aaa),
	.w7(32'hb91e570c),
	.w8(32'h38a67802),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d25576),
	.w1(32'h39ea0b41),
	.w2(32'h39cd5525),
	.w3(32'h3986f676),
	.w4(32'h39c448a8),
	.w5(32'h39fa7711),
	.w6(32'h39fca826),
	.w7(32'h3a236ac4),
	.w8(32'h3a491750),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8789430),
	.w1(32'hb58d60b3),
	.w2(32'h38823d1c),
	.w3(32'h387b5441),
	.w4(32'h37b7a372),
	.w5(32'hb827c9e4),
	.w6(32'h39054854),
	.w7(32'hb8ccc7cf),
	.w8(32'hb90117a7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7970471),
	.w1(32'hb9e3789d),
	.w2(32'hba302a55),
	.w3(32'hb9c9eeaa),
	.w4(32'hba92fe53),
	.w5(32'hba37a41e),
	.w6(32'hb9c0c7b8),
	.w7(32'hb8e5eb55),
	.w8(32'hb932eb38),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c91f0),
	.w1(32'h36e607be),
	.w2(32'h380f786c),
	.w3(32'hb8513b36),
	.w4(32'h37efdc66),
	.w5(32'h3892d49d),
	.w6(32'hb790e0f2),
	.w7(32'h38d83fdc),
	.w8(32'h38e2b77a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a263aa7),
	.w1(32'h38285e24),
	.w2(32'hba01fd45),
	.w3(32'hba7461d7),
	.w4(32'hba7478dd),
	.w5(32'hba98a738),
	.w6(32'hba22954f),
	.w7(32'hba1595c0),
	.w8(32'hb988d1a6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd2a0a),
	.w1(32'hb95dbf65),
	.w2(32'hb9bdb997),
	.w3(32'hb9101bb9),
	.w4(32'hb97d1cad),
	.w5(32'hb994076f),
	.w6(32'hb8bbbc4b),
	.w7(32'hb92b269a),
	.w8(32'hb9209c3f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3490f4),
	.w1(32'hb9615335),
	.w2(32'hbb72b6d1),
	.w3(32'hbaa03a5b),
	.w4(32'hbb7e8c65),
	.w5(32'hbba6d3c3),
	.w6(32'hbb512109),
	.w7(32'hbb49164a),
	.w8(32'hb919b8bc),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7afd1e4),
	.w1(32'hb90aebef),
	.w2(32'hb7750d2a),
	.w3(32'hb60c647a),
	.w4(32'hb8b804b5),
	.w5(32'hb88e4bed),
	.w6(32'h3841b92f),
	.w7(32'h38664c30),
	.w8(32'h38f71fd3),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2a1f6),
	.w1(32'h3a1f4146),
	.w2(32'hba6b386c),
	.w3(32'hbb65007b),
	.w4(32'hba6ccdc5),
	.w5(32'hba0ef8b6),
	.w6(32'h3b02b0a9),
	.w7(32'h3b4f534d),
	.w8(32'h3adf8d3a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule