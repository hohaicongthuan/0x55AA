module layer_10_featuremap_436(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96dd888),
	.w1(32'hbb728676),
	.w2(32'h3b76a3de),
	.w3(32'h3acb1dbf),
	.w4(32'hbb5d286e),
	.w5(32'h3b49934f),
	.w6(32'h3b2804bc),
	.w7(32'hbae70f5d),
	.w8(32'h3b12d852),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7346c1),
	.w1(32'hbb9479a8),
	.w2(32'hbb324987),
	.w3(32'hb92df3b4),
	.w4(32'hba86a698),
	.w5(32'h3b407d16),
	.w6(32'hba1d92b3),
	.w7(32'hba41deed),
	.w8(32'h3a956d49),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4255),
	.w1(32'h3bcf23f5),
	.w2(32'h3b4adb61),
	.w3(32'hbb9d1549),
	.w4(32'h3baf0f5d),
	.w5(32'h3b831b08),
	.w6(32'hbbba3b30),
	.w7(32'h3b57a421),
	.w8(32'h39deb8d6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85d62c),
	.w1(32'hbc0cee51),
	.w2(32'hbb3f7c6a),
	.w3(32'hba384fde),
	.w4(32'hbbf68533),
	.w5(32'hbb63f887),
	.w6(32'h39446ca4),
	.w7(32'hbbbeb1b3),
	.w8(32'hbbaa5c7e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb470662),
	.w1(32'hb98cf5d8),
	.w2(32'h3a89ec2c),
	.w3(32'hbb9a4f3d),
	.w4(32'hbaca117d),
	.w5(32'hba9123de),
	.w6(32'hbb909f3f),
	.w7(32'hba64298d),
	.w8(32'hba1e74ca),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4daafd),
	.w1(32'hbac2f76c),
	.w2(32'hbb8d6201),
	.w3(32'hb924592f),
	.w4(32'h3a217347),
	.w5(32'hbb121f59),
	.w6(32'h38c7f50d),
	.w7(32'h3ad84537),
	.w8(32'hba7d27e1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cbec2),
	.w1(32'hbb7b08c2),
	.w2(32'h3aeffea9),
	.w3(32'hbb72e231),
	.w4(32'hbb22501c),
	.w5(32'h3b6e219f),
	.w6(32'hbb765217),
	.w7(32'hba45b9e9),
	.w8(32'h3bf3ec8e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3da2e4),
	.w1(32'h3c1dfd10),
	.w2(32'h3c413f5b),
	.w3(32'h3c01b166),
	.w4(32'h3c31e7ba),
	.w5(32'h3bb66c49),
	.w6(32'h3ba0a23a),
	.w7(32'h3be40966),
	.w8(32'h3bfafcf8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dc599),
	.w1(32'h3a12fe30),
	.w2(32'h3b03f96e),
	.w3(32'hba217ecc),
	.w4(32'hba720623),
	.w5(32'hb9284f2d),
	.w6(32'hb9a2e847),
	.w7(32'hb99c53c9),
	.w8(32'hba8fbc3b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf18273),
	.w1(32'h3c390203),
	.w2(32'h3ba50de4),
	.w3(32'h3bb4a926),
	.w4(32'h3c42929f),
	.w5(32'h3b93b0e2),
	.w6(32'h3b797228),
	.w7(32'h3c547e3d),
	.w8(32'h3b9408d1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a385ff6),
	.w1(32'h38bb2f35),
	.w2(32'hba5bd964),
	.w3(32'h39868d78),
	.w4(32'hba810251),
	.w5(32'hbb1d2b88),
	.w6(32'h38bf762e),
	.w7(32'h3a9f39f3),
	.w8(32'hba9d7757),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb622),
	.w1(32'hbb0eeec0),
	.w2(32'h3aefb136),
	.w3(32'hbc20a301),
	.w4(32'hbbaafc12),
	.w5(32'hbb301a60),
	.w6(32'hbc3356e5),
	.w7(32'hbbb50787),
	.w8(32'h3b991087),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c308dc7),
	.w1(32'h3b95e6bc),
	.w2(32'h3bb2b0dc),
	.w3(32'h3be38741),
	.w4(32'h3b26e45a),
	.w5(32'h3b20c827),
	.w6(32'h3bcaf0a8),
	.w7(32'hbb53a960),
	.w8(32'hba92959f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f80bc),
	.w1(32'h3bab8857),
	.w2(32'h3bc3840d),
	.w3(32'hba18125a),
	.w4(32'h3c030a2b),
	.w5(32'h3bb90b76),
	.w6(32'hbab9a5a3),
	.w7(32'h3b96744d),
	.w8(32'h3b2624bd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b125cee),
	.w1(32'hbaae3bb4),
	.w2(32'h3a3712a0),
	.w3(32'h3b32f71e),
	.w4(32'hbb021c55),
	.w5(32'h3b0caf69),
	.w6(32'h3599c604),
	.w7(32'hba0fdf61),
	.w8(32'h3b0c1997),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbfa1e),
	.w1(32'h3ac21d33),
	.w2(32'h3b80d17b),
	.w3(32'h3a9bb0ca),
	.w4(32'h3ae8657b),
	.w5(32'h3bc41308),
	.w6(32'h3b2f3f5b),
	.w7(32'h3ab7311e),
	.w8(32'h3b83d362),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b89c5),
	.w1(32'h3a8f65d9),
	.w2(32'h3b3cec97),
	.w3(32'hbac7a0e3),
	.w4(32'hb9f8c040),
	.w5(32'h3aa3ca11),
	.w6(32'hbaa9dbbf),
	.w7(32'h3a4a0fdf),
	.w8(32'h3a4d55d9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf09e19),
	.w1(32'h3c3edbc6),
	.w2(32'h3c8633db),
	.w3(32'h3bc9da52),
	.w4(32'h3c23467b),
	.w5(32'h3c2d7fba),
	.w6(32'hb79a02e2),
	.w7(32'h3c26a64f),
	.w8(32'h3c177fa9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1576a),
	.w1(32'h3bab8e4d),
	.w2(32'h3b40c29c),
	.w3(32'h3bd319b5),
	.w4(32'h3b9c6093),
	.w5(32'hbac85b1e),
	.w6(32'h3b5710f6),
	.w7(32'h3b54d783),
	.w8(32'h399a050d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918b3c0),
	.w1(32'h39c0fd8d),
	.w2(32'h3926a009),
	.w3(32'hba93469e),
	.w4(32'h3aef9c16),
	.w5(32'h36411123),
	.w6(32'hb902983b),
	.w7(32'h3aca63c8),
	.w8(32'hb90d805d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0aa4c),
	.w1(32'h3adcbfc7),
	.w2(32'hbb0b2252),
	.w3(32'hbabaae87),
	.w4(32'h3b388701),
	.w5(32'hbb10ace1),
	.w6(32'hba8738d6),
	.w7(32'h3a5f9f31),
	.w8(32'hbafe5d4a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30294b),
	.w1(32'hbb9727c2),
	.w2(32'hbb10a1d8),
	.w3(32'hbacaffaa),
	.w4(32'hbbb79326),
	.w5(32'hbaa0a3f2),
	.w6(32'hba0e94de),
	.w7(32'hbb7b3808),
	.w8(32'hbb200a34),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7cb03),
	.w1(32'h39de098a),
	.w2(32'h3c81b683),
	.w3(32'hbbea5167),
	.w4(32'hbc192d9b),
	.w5(32'h3c162075),
	.w6(32'hbc2d8cb0),
	.w7(32'hba3eb8c7),
	.w8(32'h3c823143),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb122e38),
	.w1(32'hbb4abd1e),
	.w2(32'hba0d117f),
	.w3(32'hbb46b4ae),
	.w4(32'hba895fb2),
	.w5(32'h3a9f87a2),
	.w6(32'hba99a628),
	.w7(32'h3b67ad67),
	.w8(32'h3b85ae47),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba30390),
	.w1(32'hbc0214ea),
	.w2(32'hbc182c44),
	.w3(32'h3ba559ec),
	.w4(32'hbb50b807),
	.w5(32'hb9ebf659),
	.w6(32'h3c7c15ab),
	.w7(32'h3a1e6332),
	.w8(32'hb9105cb6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dcf9b),
	.w1(32'h3b9368da),
	.w2(32'h3b91202c),
	.w3(32'hba157700),
	.w4(32'h3b84adaf),
	.w5(32'h3b64a982),
	.w6(32'h3a1385a0),
	.w7(32'h3b773224),
	.w8(32'h3bab6df3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebe796),
	.w1(32'hb9d2deba),
	.w2(32'h3b7b1440),
	.w3(32'h3b981c77),
	.w4(32'h3b883182),
	.w5(32'h3b350c82),
	.w6(32'h3b8bda9f),
	.w7(32'hbac25d8f),
	.w8(32'h39ba739f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ead27),
	.w1(32'h3c2115fd),
	.w2(32'hb9f2b128),
	.w3(32'hbc34672f),
	.w4(32'h3c474db8),
	.w5(32'h3b6a3d0b),
	.w6(32'hbbb542df),
	.w7(32'h3c62e974),
	.w8(32'h3a8c91a7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e63ec),
	.w1(32'hbabc8227),
	.w2(32'hba3b322b),
	.w3(32'h3aff3c40),
	.w4(32'hbb41f81e),
	.w5(32'hbb4827ca),
	.w6(32'h3a96432d),
	.w7(32'hbb02be3c),
	.w8(32'hbb036290),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcab7c),
	.w1(32'h3af5a7e3),
	.w2(32'hbb2259c8),
	.w3(32'h398b3b3b),
	.w4(32'h3c43e91c),
	.w5(32'h3bb5aa30),
	.w6(32'h3ace3097),
	.w7(32'h3c64f9f1),
	.w8(32'h3bf2e8d9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e9597),
	.w1(32'h3b2adc40),
	.w2(32'h3b635ac0),
	.w3(32'h3b328185),
	.w4(32'hba23bb41),
	.w5(32'h3a4dd428),
	.w6(32'h3b8ac6e1),
	.w7(32'hba0392d6),
	.w8(32'h3ad98cd4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ab332),
	.w1(32'hb86624db),
	.w2(32'h3a5fbe44),
	.w3(32'h3956f411),
	.w4(32'hba03475c),
	.w5(32'h3b392a29),
	.w6(32'h37f36247),
	.w7(32'hba1adb15),
	.w8(32'h3acf15e5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcecfee),
	.w1(32'h3b54f13c),
	.w2(32'h3b8e9119),
	.w3(32'hbbd97693),
	.w4(32'h3b1261b8),
	.w5(32'h3ae820d9),
	.w6(32'hbbec4a65),
	.w7(32'h39572e3c),
	.w8(32'h3aaba51c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac405b9),
	.w1(32'hba126b8c),
	.w2(32'hbac94ff7),
	.w3(32'hbb7ac4a9),
	.w4(32'hba86a4b9),
	.w5(32'hba829533),
	.w6(32'hbb1f75b2),
	.w7(32'h390fc62d),
	.w8(32'h3a9a9dd0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9621e),
	.w1(32'h3a366add),
	.w2(32'h39967ae5),
	.w3(32'hbacfb4a3),
	.w4(32'h3b85e1a8),
	.w5(32'h3a2b713a),
	.w6(32'hbb08355d),
	.w7(32'h3bd91fd1),
	.w8(32'h3b428dc8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66d08f),
	.w1(32'hbb734f21),
	.w2(32'hbaa28cf5),
	.w3(32'hbb899465),
	.w4(32'hbb4d0ca9),
	.w5(32'hba1f319e),
	.w6(32'hbbc5454d),
	.w7(32'hbb40a403),
	.w8(32'hbae1d08b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9de8b),
	.w1(32'hbc36ad69),
	.w2(32'h3c4ea4b5),
	.w3(32'hbbd02744),
	.w4(32'hbc4ec2aa),
	.w5(32'h3b853b2a),
	.w6(32'hbbbb567a),
	.w7(32'hbc2334a2),
	.w8(32'h3b1401c4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dc876),
	.w1(32'hbc11c915),
	.w2(32'hbc38175e),
	.w3(32'hb9bfdc9c),
	.w4(32'hbbd8dcc5),
	.w5(32'hbb3bdc90),
	.w6(32'h3b7a3092),
	.w7(32'hbb10fd0f),
	.w8(32'hba93bca0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c10fb),
	.w1(32'hbbd8bfa6),
	.w2(32'hbbe4971a),
	.w3(32'hbbbbbbda),
	.w4(32'hbba6862c),
	.w5(32'hbb24f8d0),
	.w6(32'hbb4fc9b3),
	.w7(32'h3b087842),
	.w8(32'h3af67ace),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ef1f3),
	.w1(32'hb94b26a7),
	.w2(32'h3a0350bf),
	.w3(32'h39a76f5b),
	.w4(32'h3ac99ed0),
	.w5(32'h3942779d),
	.w6(32'h3a8062b1),
	.w7(32'h3b1da673),
	.w8(32'hb9430752),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81a68a),
	.w1(32'h3b12aa11),
	.w2(32'h3bb5e8c0),
	.w3(32'h3b8bf650),
	.w4(32'h3a95f79a),
	.w5(32'h399e6009),
	.w6(32'h3b2be324),
	.w7(32'h3b95828b),
	.w8(32'hba03c39f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0802f0),
	.w1(32'hbb40b00e),
	.w2(32'hba0028cf),
	.w3(32'hbb899196),
	.w4(32'hbb8d155b),
	.w5(32'hbae5df87),
	.w6(32'hbbb0a566),
	.w7(32'hbbba991c),
	.w8(32'hbb298c4c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab6b5b),
	.w1(32'hbbbdf4be),
	.w2(32'hbaa2a347),
	.w3(32'hbb9ab6a0),
	.w4(32'hbbbbbd5d),
	.w5(32'h3b24eee9),
	.w6(32'hbb3787fe),
	.w7(32'hbb635ea4),
	.w8(32'h3a80cce9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba97a14),
	.w1(32'h3bb80985),
	.w2(32'h3c24cbec),
	.w3(32'h3b4baaa6),
	.w4(32'h3be7c9c4),
	.w5(32'h3c026ac8),
	.w6(32'h3a82004a),
	.w7(32'h3c090055),
	.w8(32'h3bbefb1c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60a8fa),
	.w1(32'h3b5aee47),
	.w2(32'hbbb5d12f),
	.w3(32'h3b57cdd8),
	.w4(32'h3be06166),
	.w5(32'hba607f0a),
	.w6(32'h3b1d3819),
	.w7(32'h3bcb2e74),
	.w8(32'hbb9663e4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9fb93),
	.w1(32'hba6df105),
	.w2(32'hbb21c94d),
	.w3(32'h3bc40e77),
	.w4(32'h39ab99b5),
	.w5(32'h3ba6e5af),
	.w6(32'h3bbc0b1d),
	.w7(32'hbacd55cc),
	.w8(32'h3b31beaa),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85070a),
	.w1(32'hbb575724),
	.w2(32'h3929797b),
	.w3(32'hbba2f1ad),
	.w4(32'hbb962222),
	.w5(32'hbb1ab7f6),
	.w6(32'hbadbe0de),
	.w7(32'hbb8b8a21),
	.w8(32'hbbb13e4d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2349c8),
	.w1(32'h3c2f820e),
	.w2(32'h3c6b7aa7),
	.w3(32'h3c0aaf41),
	.w4(32'h3bfed35c),
	.w5(32'h3bf1264d),
	.w6(32'hba88ffc3),
	.w7(32'h3a9fe668),
	.w8(32'h3b709f47),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d799a),
	.w1(32'h3b6baf30),
	.w2(32'h3810d41f),
	.w3(32'hba7d0410),
	.w4(32'h3b3aca9e),
	.w5(32'hba79e94c),
	.w6(32'hba08ff9c),
	.w7(32'h3b14eda8),
	.w8(32'hba30b3b2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba883310),
	.w1(32'h3b212be7),
	.w2(32'hba473424),
	.w3(32'hbaf087e3),
	.w4(32'h3ab7c85a),
	.w5(32'h3a633708),
	.w6(32'hbb2970ae),
	.w7(32'h3afcc3a2),
	.w8(32'h3a9a5b75),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf35f54),
	.w1(32'hbaa39ffd),
	.w2(32'hbba19911),
	.w3(32'hbba5329f),
	.w4(32'hbb09437e),
	.w5(32'hbbf6da15),
	.w6(32'hbb906ebb),
	.w7(32'hbb4f245d),
	.w8(32'hbbbf541c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c1f70),
	.w1(32'hbaf2ee05),
	.w2(32'h3b0dce79),
	.w3(32'hbb30fd7d),
	.w4(32'hba357f74),
	.w5(32'h3b9ea879),
	.w6(32'hbb0e4c2a),
	.w7(32'hbb2e4172),
	.w8(32'h3b64d961),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb154b38),
	.w1(32'h3b982113),
	.w2(32'h3bcac2df),
	.w3(32'hbb9858dd),
	.w4(32'h3bcbf163),
	.w5(32'h3be857ce),
	.w6(32'hbbb627ff),
	.w7(32'h3bd538c1),
	.w8(32'h3c1490e9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dc95e),
	.w1(32'h3c171b89),
	.w2(32'h3c064119),
	.w3(32'h3c2821ad),
	.w4(32'h3c292d70),
	.w5(32'h3b2faef9),
	.w6(32'h3b772858),
	.w7(32'hb8983328),
	.w8(32'h39968906),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb457521),
	.w1(32'h3ba6f58e),
	.w2(32'hbb3c35f3),
	.w3(32'hbb341745),
	.w4(32'h3bcaf6ef),
	.w5(32'hbae5c09b),
	.w6(32'hbb59cb5b),
	.w7(32'h3beb4540),
	.w8(32'hba918735),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d1c67),
	.w1(32'h39a34a3a),
	.w2(32'h3af063ee),
	.w3(32'h3afabddc),
	.w4(32'hba4072fb),
	.w5(32'h3b0dd399),
	.w6(32'h3af4f359),
	.w7(32'hbad6859a),
	.w8(32'h3a1cc454),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ad271),
	.w1(32'hba08c859),
	.w2(32'hbacd4ad1),
	.w3(32'hbabbdbbd),
	.w4(32'hbb365e30),
	.w5(32'hbb7e0e3c),
	.w6(32'hbb2b32fd),
	.w7(32'hbb379c27),
	.w8(32'hbaa74deb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7f9f7),
	.w1(32'hbabc22c7),
	.w2(32'hba20a42a),
	.w3(32'hbafaf961),
	.w4(32'h37fc44e2),
	.w5(32'h3a1e14a7),
	.w6(32'hbaca6bcd),
	.w7(32'hba4fc6c6),
	.w8(32'hbb4b4f99),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b907b0e),
	.w1(32'h3900ee64),
	.w2(32'h3ab6eae9),
	.w3(32'h3b1e6f5e),
	.w4(32'h3a57522c),
	.w5(32'h3a370201),
	.w6(32'h3aecc596),
	.w7(32'h3a6c2c54),
	.w8(32'h3a961a65),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae467f6),
	.w1(32'h3b2c11f8),
	.w2(32'h380fae0f),
	.w3(32'h3aa3fc20),
	.w4(32'h38cf5484),
	.w5(32'hb974c792),
	.w6(32'h3a7614e9),
	.w7(32'hbaec4fdd),
	.w8(32'hbb32aad3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a855a8a),
	.w1(32'h3bee2cd1),
	.w2(32'h3b421db9),
	.w3(32'hba8a05dd),
	.w4(32'h3afe4bc4),
	.w5(32'hbb9915a1),
	.w6(32'hbb91328f),
	.w7(32'hba9512f3),
	.w8(32'hbbb320ce),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37213c),
	.w1(32'h3c39ba2f),
	.w2(32'h3ba38239),
	.w3(32'hba7ff0c9),
	.w4(32'h3c1902b9),
	.w5(32'h3b03619c),
	.w6(32'h3b128d88),
	.w7(32'h3c57ec7e),
	.w8(32'h3bc80c31),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa38749),
	.w1(32'h3aa734a6),
	.w2(32'h39e1cbfc),
	.w3(32'h3a6395b0),
	.w4(32'hb9162632),
	.w5(32'h3a89ed7f),
	.w6(32'h3b2883b3),
	.w7(32'h3ad7ff90),
	.w8(32'hba1fee1e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0dd0),
	.w1(32'h3b32c558),
	.w2(32'hbad2b340),
	.w3(32'h3b4b0c86),
	.w4(32'h398a639a),
	.w5(32'hbb67b447),
	.w6(32'h3b4f6624),
	.w7(32'hba96cf17),
	.w8(32'hb8ea9f8a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48b069),
	.w1(32'h3b71bab7),
	.w2(32'h3b586642),
	.w3(32'h3ab53f35),
	.w4(32'h3b8a1032),
	.w5(32'h3b57d832),
	.w6(32'h3b0c2d7e),
	.w7(32'h3b872734),
	.w8(32'h3b32f525),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9a127),
	.w1(32'hb916ed55),
	.w2(32'hb9010472),
	.w3(32'h3ab24c32),
	.w4(32'hbaa01ea5),
	.w5(32'h3983591e),
	.w6(32'h3b1e6489),
	.w7(32'hbaa3d114),
	.w8(32'h3b13fadc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39688388),
	.w1(32'h3b3fd041),
	.w2(32'h3bb1b8a9),
	.w3(32'hb9f35be3),
	.w4(32'h3adb772a),
	.w5(32'hbb0d897a),
	.w6(32'hbb468972),
	.w7(32'hbac0515b),
	.w8(32'hbb117ce4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb974773),
	.w1(32'hbb195399),
	.w2(32'h3b207e03),
	.w3(32'hbb9ff288),
	.w4(32'hbb00eb9d),
	.w5(32'h3b79dad0),
	.w6(32'hbb7752a1),
	.w7(32'hbadb7e29),
	.w8(32'h3b3f2d93),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb135e9c),
	.w1(32'h3b94fab6),
	.w2(32'h3b680382),
	.w3(32'hbbb9b554),
	.w4(32'hb9a6c16f),
	.w5(32'hb96289bb),
	.w6(32'hbb60bce3),
	.w7(32'h3abe9690),
	.w8(32'hbaf4e1bc),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51db5a),
	.w1(32'hbc2268da),
	.w2(32'hbbe47955),
	.w3(32'hbb8f5757),
	.w4(32'hbc64a613),
	.w5(32'h3b5467a6),
	.w6(32'h3aae52d4),
	.w7(32'hba2b50c5),
	.w8(32'h3aaea174),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44df77),
	.w1(32'hbb3128b2),
	.w2(32'hbaee1d49),
	.w3(32'hbac8f75a),
	.w4(32'h3c12d836),
	.w5(32'hba3413a8),
	.w6(32'hbb82636c),
	.w7(32'hba9e25b2),
	.w8(32'hbbb73af9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90297b),
	.w1(32'h3b297760),
	.w2(32'h3ab5af2b),
	.w3(32'h3b83fb40),
	.w4(32'hbc10810a),
	.w5(32'hbc883780),
	.w6(32'h3b7301a2),
	.w7(32'hbbf0ecf9),
	.w8(32'h3bd0984d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f871c),
	.w1(32'h3a0c849b),
	.w2(32'hb93ae2fd),
	.w3(32'h3ade5d0d),
	.w4(32'hbbc582d8),
	.w5(32'hbbe34d8b),
	.w6(32'h3b950a8d),
	.w7(32'h3ae45494),
	.w8(32'hbb7f3cb5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e990f),
	.w1(32'h3c8d8de1),
	.w2(32'h3ca07440),
	.w3(32'hbba630dc),
	.w4(32'h3cdef235),
	.w5(32'h3d0430f4),
	.w6(32'hbb06344a),
	.w7(32'h3c827226),
	.w8(32'hbcd31061),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78aa51),
	.w1(32'h3c5b86cf),
	.w2(32'h3c661736),
	.w3(32'hbce0f728),
	.w4(32'hb9a53d4f),
	.w5(32'h3c0d6605),
	.w6(32'hbc2aa521),
	.w7(32'h3c414faf),
	.w8(32'h3c1a14b4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c9758),
	.w1(32'hbcbbb2a3),
	.w2(32'h3c1ca10b),
	.w3(32'hbba5dea9),
	.w4(32'hbc60d314),
	.w5(32'h3cdf079d),
	.w6(32'h3a2221f4),
	.w7(32'h39836533),
	.w8(32'hbaeb0adf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06e61d),
	.w1(32'h3c1eb0d2),
	.w2(32'h3c65fc98),
	.w3(32'hbd04efaf),
	.w4(32'h3c0df89e),
	.w5(32'h3b5064df),
	.w6(32'h37832965),
	.w7(32'hbad28480),
	.w8(32'hb860d9b4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c7ea9),
	.w1(32'hbaa73009),
	.w2(32'hbb963d77),
	.w3(32'h3c1f835c),
	.w4(32'hbad719d8),
	.w5(32'h3b8b7be7),
	.w6(32'h3baaa457),
	.w7(32'hbc474cdc),
	.w8(32'h3c63b40a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f9cc0),
	.w1(32'h3b711918),
	.w2(32'hbc101c3b),
	.w3(32'hba8db368),
	.w4(32'h3ccf6417),
	.w5(32'hbc052334),
	.w6(32'h3a08adb2),
	.w7(32'h3c03f280),
	.w8(32'hbb715c8a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bd86b),
	.w1(32'h3b2c31d7),
	.w2(32'hbbf4c2c2),
	.w3(32'hbd089ef1),
	.w4(32'h3b7bd24e),
	.w5(32'hbc187334),
	.w6(32'hbc6f46b3),
	.w7(32'h3b82183c),
	.w8(32'h3c00414f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b2a58),
	.w1(32'h3c36f3e5),
	.w2(32'h3c9540ca),
	.w3(32'hbc316918),
	.w4(32'hbb13894b),
	.w5(32'h3c8d821c),
	.w6(32'hbba7f49b),
	.w7(32'h3be8f1ed),
	.w8(32'h3c765ddd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb29ad6),
	.w1(32'h395b68a5),
	.w2(32'h3c3ca747),
	.w3(32'h3c8a8839),
	.w4(32'hbc10780e),
	.w5(32'h3b50de48),
	.w6(32'h3c7fa2da),
	.w7(32'hbbfb03b3),
	.w8(32'h3b7ecf93),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05b2c3),
	.w1(32'hbb8389ed),
	.w2(32'hbc53528b),
	.w3(32'hbb8519a0),
	.w4(32'hbc10c292),
	.w5(32'hbbc5cfee),
	.w6(32'hbb8c8533),
	.w7(32'h3bc55fc7),
	.w8(32'h3d3c8410),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b17c5),
	.w1(32'h3bb1eafd),
	.w2(32'hbbf4ba4f),
	.w3(32'h3c94cfbe),
	.w4(32'h3896025e),
	.w5(32'hbc8b9bd7),
	.w6(32'h3c359a19),
	.w7(32'hbbc1b737),
	.w8(32'hbb489d11),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8219b3),
	.w1(32'h3b53cfab),
	.w2(32'hbb1fca3d),
	.w3(32'hbbfbd4f5),
	.w4(32'h3ac7bc03),
	.w5(32'hbc6a3a6a),
	.w6(32'h3aec40a3),
	.w7(32'hbb382343),
	.w8(32'hbb17a4fd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cadd6c7),
	.w1(32'h3b0c1ea2),
	.w2(32'hbb301442),
	.w3(32'hbbc1498d),
	.w4(32'hbb567c90),
	.w5(32'hba92e0bd),
	.w6(32'h3acf64de),
	.w7(32'h3b25a2d5),
	.w8(32'h3a0f620e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bbf95),
	.w1(32'hbc946701),
	.w2(32'hbbbe8a48),
	.w3(32'hbb02a278),
	.w4(32'hbb644856),
	.w5(32'hbc739a59),
	.w6(32'h3c0deec4),
	.w7(32'hbbf2c36a),
	.w8(32'hb8813b88),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30af93),
	.w1(32'hbc305e36),
	.w2(32'hbc05b220),
	.w3(32'hbc1f9396),
	.w4(32'hbc0e7723),
	.w5(32'hbca42b97),
	.w6(32'hbc42b30e),
	.w7(32'hbb9306c9),
	.w8(32'h3c23a214),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba9c93),
	.w1(32'hb9f199d8),
	.w2(32'hba719695),
	.w3(32'hbc2a14b5),
	.w4(32'hbb64a40a),
	.w5(32'hbb800bb9),
	.w6(32'hbb49e053),
	.w7(32'hbc24deb0),
	.w8(32'hbae028ce),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96ebd5),
	.w1(32'h3c1f5654),
	.w2(32'h3b2b318c),
	.w3(32'h3c006c9a),
	.w4(32'h3c2e28b6),
	.w5(32'hbcbdbf21),
	.w6(32'hb89e50fe),
	.w7(32'h3ad8ec84),
	.w8(32'hbc28a0c8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d894),
	.w1(32'hbc33bcde),
	.w2(32'hbb025668),
	.w3(32'hbc1b78da),
	.w4(32'hbc0640c7),
	.w5(32'hbb298ed4),
	.w6(32'hbc2707e6),
	.w7(32'hbc390ca0),
	.w8(32'hbbf4cef9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91b2f0),
	.w1(32'hb9b3d8d2),
	.w2(32'hb934733f),
	.w3(32'h3b935616),
	.w4(32'h39a8976a),
	.w5(32'hbaa653a2),
	.w6(32'hbbf14d6e),
	.w7(32'hbaae4085),
	.w8(32'h3b84cd20),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca325d),
	.w1(32'h3b0afb28),
	.w2(32'h3b9650e1),
	.w3(32'h39506803),
	.w4(32'h3c1c40ab),
	.w5(32'h3c71d791),
	.w6(32'h3bdaface),
	.w7(32'h3b23806f),
	.w8(32'h3b3fea14),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38121481),
	.w1(32'hbb1d0b91),
	.w2(32'h3d0232ce),
	.w3(32'h3a60e628),
	.w4(32'hbc6d1489),
	.w5(32'h3c153180),
	.w6(32'h3aed28cc),
	.w7(32'hbca3d1b3),
	.w8(32'hbd5c401e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb214ae1),
	.w1(32'h3b4c2394),
	.w2(32'h3a9d17e5),
	.w3(32'h3c1a41e6),
	.w4(32'hbbbd1326),
	.w5(32'hbc630b5a),
	.w6(32'h3b5a9722),
	.w7(32'hbae3b49d),
	.w8(32'hbba15ca4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd14393),
	.w1(32'hbba10ce0),
	.w2(32'hbb8c0c60),
	.w3(32'hbb1c60de),
	.w4(32'h3c381bf2),
	.w5(32'h3c2b5a76),
	.w6(32'h39966539),
	.w7(32'h3b7c3f96),
	.w8(32'hbc630a23),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10f191),
	.w1(32'hbc544d56),
	.w2(32'hbc4f7db1),
	.w3(32'hbbef81ca),
	.w4(32'hbc2ad2d9),
	.w5(32'h3a20de96),
	.w6(32'hbc92c5f5),
	.w7(32'h3b78a96d),
	.w8(32'h3b02777c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fc4d0),
	.w1(32'h3aca30b0),
	.w2(32'h3b940741),
	.w3(32'hbb017c6e),
	.w4(32'h3c131ad1),
	.w5(32'hbc469759),
	.w6(32'h3bae7d73),
	.w7(32'h3bada501),
	.w8(32'hbc0cedbf),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0a1b1),
	.w1(32'hbc0eec3c),
	.w2(32'h3bf678b5),
	.w3(32'hbbee890d),
	.w4(32'hbc886f85),
	.w5(32'hbc58637b),
	.w6(32'hbc3a7496),
	.w7(32'hbbb59c02),
	.w8(32'h3bf26bf9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2a4a0),
	.w1(32'hbaea122a),
	.w2(32'h3c4c7694),
	.w3(32'h3ac745bb),
	.w4(32'hbae48667),
	.w5(32'h3ab92b56),
	.w6(32'hb904e509),
	.w7(32'hbbdd48b7),
	.w8(32'hbc0c23c5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdafc60),
	.w1(32'hbc3d5b2b),
	.w2(32'hba722636),
	.w3(32'hbbe5e328),
	.w4(32'hbc8f1cc5),
	.w5(32'h3c4da280),
	.w6(32'h39efa6d6),
	.w7(32'hbac83f5d),
	.w8(32'hbc668e11),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8c040),
	.w1(32'hbb9750c5),
	.w2(32'hbae602eb),
	.w3(32'hbbf30e37),
	.w4(32'hbbe6fda1),
	.w5(32'h3bc65cd7),
	.w6(32'h3c9398a6),
	.w7(32'hbc1c3c17),
	.w8(32'hbb360c27),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf55cc),
	.w1(32'h3c2404c7),
	.w2(32'h3c5e2964),
	.w3(32'h3bc2a235),
	.w4(32'hba9aeb9f),
	.w5(32'hbc865ea1),
	.w6(32'hbb0a2979),
	.w7(32'hbc7726ec),
	.w8(32'h3d062547),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf096e),
	.w1(32'hbbd3b5d1),
	.w2(32'hbbe6df0d),
	.w3(32'h3c2433d0),
	.w4(32'h3cf23e1d),
	.w5(32'hbc429476),
	.w6(32'hbca957ca),
	.w7(32'hbabbb9d5),
	.w8(32'h3c7f2d05),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d13edc5),
	.w1(32'h3bb7d9ca),
	.w2(32'h3c4d202e),
	.w3(32'h3bc3e740),
	.w4(32'hbb7289ad),
	.w5(32'h3c85a3b1),
	.w6(32'h39c1eb0d),
	.w7(32'hbc1194d2),
	.w8(32'hbb99c0cf),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b041d77),
	.w1(32'hbbe77aa4),
	.w2(32'hbaad565b),
	.w3(32'hb8680d44),
	.w4(32'hbc8a8063),
	.w5(32'hbb312442),
	.w6(32'hbbf322e5),
	.w7(32'h3b083faf),
	.w8(32'h3c62f338),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b913eda),
	.w1(32'h3c4fcf7f),
	.w2(32'h3c10bea6),
	.w3(32'h3c348a4a),
	.w4(32'h3c691de4),
	.w5(32'h3cbeea6f),
	.w6(32'h3b9aaf8e),
	.w7(32'h3b36857d),
	.w8(32'hbc2e75d0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb64f49),
	.w1(32'hbb966c4b),
	.w2(32'h3a8329cd),
	.w3(32'hbd0f1dcf),
	.w4(32'hbc011baf),
	.w5(32'hbbe8d248),
	.w6(32'hbc9f2e01),
	.w7(32'h3b2af1e4),
	.w8(32'hbbe5c92c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec91a8),
	.w1(32'h3b96d0b3),
	.w2(32'h3b601550),
	.w3(32'h3c23f32f),
	.w4(32'h3a6de570),
	.w5(32'hbb7bc8ec),
	.w6(32'h3b8c9089),
	.w7(32'h3c01e1ab),
	.w8(32'h3c7e01a6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b733274),
	.w1(32'hbb4f8a60),
	.w2(32'hbbb40639),
	.w3(32'hbb38e792),
	.w4(32'hbb26ed8c),
	.w5(32'h3c9015b3),
	.w6(32'h3b71caee),
	.w7(32'h3c1baa0d),
	.w8(32'h3b1db609),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2e0b7),
	.w1(32'h3be4e786),
	.w2(32'h3c5ca48e),
	.w3(32'hbb81e3b9),
	.w4(32'h3b508635),
	.w5(32'hbc0a752f),
	.w6(32'hbae1e991),
	.w7(32'h3bf1e676),
	.w8(32'h3b2a53b6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb729ccc),
	.w1(32'h3b8a8640),
	.w2(32'h3bb53858),
	.w3(32'hbbef42a8),
	.w4(32'hbc316527),
	.w5(32'hbba8699f),
	.w6(32'h3a6f8e6f),
	.w7(32'h3b70f614),
	.w8(32'h3a87f9da),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e90b9b),
	.w1(32'hbc790956),
	.w2(32'hbc95547c),
	.w3(32'h3c3a3b34),
	.w4(32'hbcc69f79),
	.w5(32'hbbf34e05),
	.w6(32'hbb0a25c7),
	.w7(32'hbb8b094a),
	.w8(32'h3c93b10a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8befa),
	.w1(32'hbc8439b3),
	.w2(32'hbc02dab4),
	.w3(32'h3ccfbc8e),
	.w4(32'h3a325478),
	.w5(32'h3df1478a),
	.w6(32'h3bf2974a),
	.w7(32'hbcc67ea3),
	.w8(32'hbcbc7684),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce1b28d),
	.w1(32'h3b803b47),
	.w2(32'hba4b4c0c),
	.w3(32'hbd7bca2f),
	.w4(32'hba5e4573),
	.w5(32'hb90b8b1f),
	.w6(32'hbca9da2b),
	.w7(32'hbac57181),
	.w8(32'h3a21c1c8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06ce99),
	.w1(32'h3adbac06),
	.w2(32'h3c25560d),
	.w3(32'h3c017408),
	.w4(32'hbbfd803e),
	.w5(32'h3bd307e0),
	.w6(32'h3c10f8b2),
	.w7(32'h3a95962a),
	.w8(32'h3bb9f1af),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30900b),
	.w1(32'hbb6c85a5),
	.w2(32'h3bfc7ca4),
	.w3(32'h3c2a5ae2),
	.w4(32'hbbc08935),
	.w5(32'h3d048471),
	.w6(32'h3bce63df),
	.w7(32'hbb11fe11),
	.w8(32'hbae5ff48),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a4d8d),
	.w1(32'hbb0b5587),
	.w2(32'h3cb132b0),
	.w3(32'hb9f6d1ad),
	.w4(32'h3bcf16c2),
	.w5(32'h3ba87716),
	.w6(32'hbc2e18ed),
	.w7(32'hbbf23a03),
	.w8(32'hbd11759b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94bd53),
	.w1(32'hbc51ebd0),
	.w2(32'hbc72af68),
	.w3(32'hbb5a4ded),
	.w4(32'hbbc8b10c),
	.w5(32'h3c118d1f),
	.w6(32'h3af6edbf),
	.w7(32'h3bbef314),
	.w8(32'h3c75928f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc314928),
	.w1(32'hba620dc6),
	.w2(32'h3bcca0d1),
	.w3(32'hbb968414),
	.w4(32'hbc7c028b),
	.w5(32'h3cca06ea),
	.w6(32'h3b2d9a4b),
	.w7(32'hb998946d),
	.w8(32'h3ca4e369),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc128c8),
	.w1(32'h3b22c055),
	.w2(32'h3a8f0101),
	.w3(32'h3d93122b),
	.w4(32'h3c12133b),
	.w5(32'h3c799649),
	.w6(32'hbb823ebc),
	.w7(32'hba7fa315),
	.w8(32'hbb7b8177),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba506d55),
	.w1(32'h3bd3d652),
	.w2(32'h3acc3458),
	.w3(32'h3a2fbe77),
	.w4(32'hbbb12bd2),
	.w5(32'hbc04bc88),
	.w6(32'hbbb08f6b),
	.w7(32'hbc04d60c),
	.w8(32'hba99ca13),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38febb8b),
	.w1(32'hbc673b04),
	.w2(32'hbc8caeca),
	.w3(32'hb9460d51),
	.w4(32'hbba74ecf),
	.w5(32'hbc19b4ec),
	.w6(32'h3c252718),
	.w7(32'hbbbb88f7),
	.w8(32'h3c2f8cb0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30fff8),
	.w1(32'h3be88fbb),
	.w2(32'h3b828bd3),
	.w3(32'h3c391b6e),
	.w4(32'hbc1042dd),
	.w5(32'h3c4c507b),
	.w6(32'hbb40d0ca),
	.w7(32'hbb0428e4),
	.w8(32'h3bd8a4e2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adb133),
	.w1(32'hbc059894),
	.w2(32'h3c51d8b5),
	.w3(32'h3c62375a),
	.w4(32'hbc0189de),
	.w5(32'h3c046def),
	.w6(32'h3bb18f32),
	.w7(32'hbc3c5374),
	.w8(32'hbc93e81c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42fd5),
	.w1(32'hbc24c02b),
	.w2(32'h3ae7fd1d),
	.w3(32'hbc5b976c),
	.w4(32'h3b1b1ff2),
	.w5(32'h3ceff643),
	.w6(32'hbc60a081),
	.w7(32'h3b751cf6),
	.w8(32'h3a1ba0f0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c6c0e),
	.w1(32'h3a954c27),
	.w2(32'h3bb2f7f2),
	.w3(32'hbc080d8d),
	.w4(32'h3acad86b),
	.w5(32'hbc87e1eb),
	.w6(32'h3c51aed7),
	.w7(32'h3b55ea6f),
	.w8(32'hbae44cf7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0ce2c),
	.w1(32'h3b149b19),
	.w2(32'h3bc8ef14),
	.w3(32'hbc312d22),
	.w4(32'hbc129e44),
	.w5(32'hbbdeed22),
	.w6(32'hbc131e71),
	.w7(32'hbc5ec1b6),
	.w8(32'h3b78d33f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6c814),
	.w1(32'h3ab13e8f),
	.w2(32'h3b3c2c25),
	.w3(32'hbc96ab15),
	.w4(32'h38c909e5),
	.w5(32'hbb2e4227),
	.w6(32'hbc17289c),
	.w7(32'h3bb8cc68),
	.w8(32'h3be68ca5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22e822),
	.w1(32'hbab3cad3),
	.w2(32'hbb776f0c),
	.w3(32'hbaabe14a),
	.w4(32'h3ad6456f),
	.w5(32'hbb09123b),
	.w6(32'h3a965009),
	.w7(32'hbb2c4ad2),
	.w8(32'hbbdaf307),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12fc2c),
	.w1(32'hbbcf0011),
	.w2(32'h3c8988fa),
	.w3(32'h3aecca3c),
	.w4(32'hbaa739bc),
	.w5(32'h3d96d701),
	.w6(32'hbb608050),
	.w7(32'h3ca78426),
	.w8(32'hbce45b9d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdcd288),
	.w1(32'hbb35739a),
	.w2(32'hbbb55976),
	.w3(32'hbc20c0cc),
	.w4(32'h3b027323),
	.w5(32'hbbf35304),
	.w6(32'hbc22d26d),
	.w7(32'hbab3d663),
	.w8(32'hbc8408a8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53e68c),
	.w1(32'h3c07a523),
	.w2(32'hbb224f96),
	.w3(32'hbbe60313),
	.w4(32'h3c100f25),
	.w5(32'hbb44dcd3),
	.w6(32'h3bd1cc56),
	.w7(32'h3c041724),
	.w8(32'h3b365f5a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf2e06),
	.w1(32'h39fcd2c9),
	.w2(32'h3b08b16d),
	.w3(32'h3bb42a4a),
	.w4(32'hbb2e0b5e),
	.w5(32'h3b8fce05),
	.w6(32'h3c167236),
	.w7(32'hbbe5d1f7),
	.w8(32'hba9f68f8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bb8d5),
	.w1(32'h3af56800),
	.w2(32'h3c6462cc),
	.w3(32'hbb67db09),
	.w4(32'h3c3c31ed),
	.w5(32'h3ce42d2c),
	.w6(32'hbb8b831b),
	.w7(32'h3b51547f),
	.w8(32'hbbde5197),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04668e),
	.w1(32'h3c120b0a),
	.w2(32'h3d1f6210),
	.w3(32'h3b03d387),
	.w4(32'hbb7e1c7b),
	.w5(32'h3ce8ae07),
	.w6(32'hba65b28f),
	.w7(32'hbc7cda37),
	.w8(32'hbd596d12),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0dccf),
	.w1(32'h3a046149),
	.w2(32'hbc456213),
	.w3(32'h3c28d1b5),
	.w4(32'h3cf48a29),
	.w5(32'hbbb3ef67),
	.w6(32'hbbc7522f),
	.w7(32'h3b9d3a17),
	.w8(32'hbc633158),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc03a54),
	.w1(32'h3c52d0c8),
	.w2(32'h3c08ae22),
	.w3(32'hbc871182),
	.w4(32'h3a827601),
	.w5(32'hbbbb4d3f),
	.w6(32'h3b9165ed),
	.w7(32'h3ba3a2b4),
	.w8(32'h3b9e5c3f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0b9ba),
	.w1(32'h3c4760d4),
	.w2(32'h3bb739ff),
	.w3(32'h39d64aaa),
	.w4(32'hbb5a8e73),
	.w5(32'hba1c64ee),
	.w6(32'h3bca298b),
	.w7(32'hbc212db1),
	.w8(32'hbc0e8bd2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf0d51),
	.w1(32'hbac5c618),
	.w2(32'h3c0e6beb),
	.w3(32'hbc0df6ef),
	.w4(32'hbc0f4b09),
	.w5(32'h3cd89ccf),
	.w6(32'hbc2cd5a6),
	.w7(32'hbb7f7973),
	.w8(32'h3c38492c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8582d),
	.w1(32'hbc723989),
	.w2(32'hbb10b439),
	.w3(32'h3bad9c1b),
	.w4(32'hbc81a872),
	.w5(32'h3c23af05),
	.w6(32'hbb347b32),
	.w7(32'hbc3169e6),
	.w8(32'h3b1cc240),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe47771),
	.w1(32'hbbed5ef6),
	.w2(32'hbc63e641),
	.w3(32'hbad20cfa),
	.w4(32'h3c97a8f9),
	.w5(32'hbc952cb8),
	.w6(32'hba58a1b0),
	.w7(32'h3c42e178),
	.w8(32'h3d27add2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1458c),
	.w1(32'hbbce6b42),
	.w2(32'hbb35f5b3),
	.w3(32'h3ae24fc3),
	.w4(32'hbc0451a1),
	.w5(32'h3b6f8ed8),
	.w6(32'hbb7b613f),
	.w7(32'hbad81ea0),
	.w8(32'hbc1b881c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf87a63),
	.w1(32'hbb27d2ec),
	.w2(32'h38e5070c),
	.w3(32'h3be9750b),
	.w4(32'hb9da942e),
	.w5(32'h3ca65502),
	.w6(32'hbc0326f9),
	.w7(32'hb93733ce),
	.w8(32'h3b04c8fe),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc305e59),
	.w1(32'hbbac7b55),
	.w2(32'hbab6257d),
	.w3(32'hbc3e246a),
	.w4(32'h3b4cd91c),
	.w5(32'h3952110b),
	.w6(32'hbc1ec61f),
	.w7(32'h3b61ccfb),
	.w8(32'hbc17421f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7eb81e),
	.w1(32'hbaa2a4dd),
	.w2(32'h39e11b46),
	.w3(32'h3a1403da),
	.w4(32'h3c02ce6b),
	.w5(32'hbbda9d43),
	.w6(32'hbbdb301e),
	.w7(32'hbb8a1953),
	.w8(32'hbb58c1c3),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe07caa),
	.w1(32'h3afddf2f),
	.w2(32'hba9ade96),
	.w3(32'hbc47069c),
	.w4(32'h3c01743d),
	.w5(32'h3c5d2813),
	.w6(32'hbc307de1),
	.w7(32'h3aad1546),
	.w8(32'hbbbefba2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8f501),
	.w1(32'h3c3a0e65),
	.w2(32'h3b0237de),
	.w3(32'hbc62be68),
	.w4(32'h3bc34483),
	.w5(32'hbc2b25c9),
	.w6(32'hbaef709b),
	.w7(32'h3c162d0e),
	.w8(32'hbc4b02cd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08a94b),
	.w1(32'h3b991430),
	.w2(32'h3b0ba5f2),
	.w3(32'h3b59c351),
	.w4(32'h3c85d25d),
	.w5(32'h3cb7af29),
	.w6(32'hbbd7e6cd),
	.w7(32'h3b8be344),
	.w8(32'hbbc5f13e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f1deb),
	.w1(32'h3b59ea3a),
	.w2(32'h3c0a021b),
	.w3(32'hbca1e794),
	.w4(32'h3be3b4eb),
	.w5(32'h3c44e0e4),
	.w6(32'hbc960b5a),
	.w7(32'h3c08e6d9),
	.w8(32'h3b2db0a9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33dd8f),
	.w1(32'h3c0e1ca6),
	.w2(32'h3baae880),
	.w3(32'h3c026c4f),
	.w4(32'h3b582089),
	.w5(32'h3b362d36),
	.w6(32'h3bc7e8c3),
	.w7(32'h3b258a88),
	.w8(32'hbb470866),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb75c1),
	.w1(32'h3c4d4adf),
	.w2(32'h3b8d3032),
	.w3(32'h39e3d6b2),
	.w4(32'h3ae03500),
	.w5(32'hbc69226c),
	.w6(32'hbb3902cb),
	.w7(32'h3c15dac7),
	.w8(32'hbb8b8d4a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43b29f),
	.w1(32'h3becc2c0),
	.w2(32'hbada67f2),
	.w3(32'hb807f9f2),
	.w4(32'h3c394282),
	.w5(32'hbc827eab),
	.w6(32'h3c39ac1d),
	.w7(32'h3c291a9d),
	.w8(32'hbb584531),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4c8f7),
	.w1(32'h3b8940b4),
	.w2(32'h3bff2bb0),
	.w3(32'hbb63ef58),
	.w4(32'h3ab9d6b3),
	.w5(32'hbc5f4507),
	.w6(32'h37bcdd22),
	.w7(32'h3be82bf7),
	.w8(32'h3b8d0e1e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06296d),
	.w1(32'hba76310d),
	.w2(32'hbb8337d1),
	.w3(32'h3b99dff6),
	.w4(32'h3b97333d),
	.w5(32'hbbb900dc),
	.w6(32'h3b6880c9),
	.w7(32'h3c0538cb),
	.w8(32'hb9e12ceb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5785c),
	.w1(32'hbbb25690),
	.w2(32'hbb84a819),
	.w3(32'h3a9d8ef3),
	.w4(32'hbc36baeb),
	.w5(32'hbc067a2e),
	.w6(32'h3c3aebbe),
	.w7(32'hbc211943),
	.w8(32'hbb18b6f8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5333c),
	.w1(32'h3afd2ce1),
	.w2(32'h3b95fb97),
	.w3(32'hbbd35345),
	.w4(32'hb9563a82),
	.w5(32'hbc7d74d9),
	.w6(32'hbc4fe652),
	.w7(32'hbba0b73c),
	.w8(32'hbb8c97a1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabaefa),
	.w1(32'hbb528da8),
	.w2(32'hbc328d91),
	.w3(32'hbc04c025),
	.w4(32'h3bdd4134),
	.w5(32'hbbb4b8e1),
	.w6(32'h3bc0a41f),
	.w7(32'h3b71d9dd),
	.w8(32'h3c120265),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f8397),
	.w1(32'h3ba857f0),
	.w2(32'h388ac990),
	.w3(32'hbcc29eb3),
	.w4(32'hbbbcde89),
	.w5(32'hbb82baa5),
	.w6(32'hbbb21287),
	.w7(32'h3b00eb2e),
	.w8(32'h3b901b0c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb270fc3),
	.w1(32'h3b157726),
	.w2(32'h3c989522),
	.w3(32'h3b82e27a),
	.w4(32'hbd08bd11),
	.w5(32'h3ceb165b),
	.w6(32'hbae649d9),
	.w7(32'hbc44c5de),
	.w8(32'hbc33fc02),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d3194),
	.w1(32'h3b7664dc),
	.w2(32'h3c4410c0),
	.w3(32'h3d6d6909),
	.w4(32'hbc0c9e94),
	.w5(32'hbbc6efee),
	.w6(32'h3bb14103),
	.w7(32'hbb709623),
	.w8(32'h3c45375e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf929),
	.w1(32'h3b33bec8),
	.w2(32'hbb7149b3),
	.w3(32'hbc34ca54),
	.w4(32'hbc5a9b02),
	.w5(32'hbc95a270),
	.w6(32'hbc09a975),
	.w7(32'h3b530482),
	.w8(32'h3c9444bd),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2777ec),
	.w1(32'hbc427d8a),
	.w2(32'hbd51091c),
	.w3(32'h3bfaf3ab),
	.w4(32'h3c465647),
	.w5(32'hbcc9b286),
	.w6(32'h3a812ec0),
	.w7(32'h3ca121da),
	.w8(32'h3da3c6a5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2704f),
	.w1(32'hbb6a42bb),
	.w2(32'h3b286fb5),
	.w3(32'hbc4b82d1),
	.w4(32'h3bdd4d7c),
	.w5(32'h3ad2f1a4),
	.w6(32'hba6adab6),
	.w7(32'hbb723fd6),
	.w8(32'hbc0b59ed),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d08e),
	.w1(32'hbc6b267d),
	.w2(32'hbc0072a7),
	.w3(32'hbcd73dab),
	.w4(32'hbc9f1ff9),
	.w5(32'hbcb51ba2),
	.w6(32'hbbc42c1d),
	.w7(32'hbcbb4403),
	.w8(32'hbc562637),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8be6e6),
	.w1(32'h3adbaf5d),
	.w2(32'hb8b8289d),
	.w3(32'hbab78df2),
	.w4(32'hbbc1fda8),
	.w5(32'h3a2dab4f),
	.w6(32'hb9ec64e8),
	.w7(32'hbbf2c655),
	.w8(32'hba88d0ce),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d7a76),
	.w1(32'hbb74f1ce),
	.w2(32'h3c0f4761),
	.w3(32'h398dde51),
	.w4(32'hbce859b4),
	.w5(32'h3c0bb98e),
	.w6(32'hbb04c4f5),
	.w7(32'hbcb2bd56),
	.w8(32'hbaab97ed),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88ff6b),
	.w1(32'hb98e18cb),
	.w2(32'h3ae85880),
	.w3(32'h3cac9a51),
	.w4(32'hb9f22054),
	.w5(32'hbc4cbab0),
	.w6(32'hbb0aa1f1),
	.w7(32'h3b64212d),
	.w8(32'h3b04fcdb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab25ad8),
	.w1(32'h3c89fa8b),
	.w2(32'h3c7b22d9),
	.w3(32'hbb515f0a),
	.w4(32'h3c96b0d4),
	.w5(32'hbd4b5a0a),
	.w6(32'hbb8290ab),
	.w7(32'h3c475125),
	.w8(32'h3cb048a5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4864f),
	.w1(32'h3b5f1262),
	.w2(32'hbaccfe34),
	.w3(32'h3d4244c3),
	.w4(32'h3bf01058),
	.w5(32'hbaf0895b),
	.w6(32'hb97a8f32),
	.w7(32'hbafbf631),
	.w8(32'hbc65b1a1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d8b0b),
	.w1(32'h3b095f82),
	.w2(32'hbb35e771),
	.w3(32'h3c88142e),
	.w4(32'h3c004892),
	.w5(32'hbac3ba71),
	.w6(32'hbbc478fb),
	.w7(32'h3b061ca5),
	.w8(32'hbb9126f3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b9402),
	.w1(32'hbb013262),
	.w2(32'h3ac86c07),
	.w3(32'hbbe6d375),
	.w4(32'hbb79dfe8),
	.w5(32'hbb3a0fa3),
	.w6(32'hb940c65d),
	.w7(32'h3b9f5440),
	.w8(32'hba9a67ba),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fba0a),
	.w1(32'h3c84e54a),
	.w2(32'h3bbddaed),
	.w3(32'h3c2211d0),
	.w4(32'h3cb59a90),
	.w5(32'hbb99622a),
	.w6(32'hbaa07abc),
	.w7(32'h3bb3cb95),
	.w8(32'hbb41d0e2),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e8284),
	.w1(32'h3ba3b10a),
	.w2(32'h3b6ac4e8),
	.w3(32'hba2fbf07),
	.w4(32'hbb510fc8),
	.w5(32'hbc1e6ec4),
	.w6(32'h3c7e8246),
	.w7(32'hbb7cf19f),
	.w8(32'hbb2bb7de),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56a7d4),
	.w1(32'h3c25ed78),
	.w2(32'h3c9e7dfc),
	.w3(32'hbb0cc788),
	.w4(32'hbb31c4a4),
	.w5(32'h3c2fe9e3),
	.w6(32'hbafd4ffc),
	.w7(32'hbc4c0890),
	.w8(32'hbc3ad194),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b329e6e),
	.w1(32'h3b50ac01),
	.w2(32'hbad2e883),
	.w3(32'hbb88709c),
	.w4(32'hbc328bf5),
	.w5(32'hbcc0a256),
	.w6(32'hbbc53581),
	.w7(32'h3b2ce302),
	.w8(32'h3b0a844a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98eaf93),
	.w1(32'h3b249aeb),
	.w2(32'hbc1bbaec),
	.w3(32'h3c8960dd),
	.w4(32'h3d18a923),
	.w5(32'hbcb172ba),
	.w6(32'hba419030),
	.w7(32'h3bc717c3),
	.w8(32'hbbf10ed4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ffe6a),
	.w1(32'hbc0cd740),
	.w2(32'h3c8c54be),
	.w3(32'hbd5b4520),
	.w4(32'hbd792694),
	.w5(32'h3c87c5c7),
	.w6(32'hbcd9d6a9),
	.w7(32'hbcc562b6),
	.w8(32'h3c0c1d81),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba85013),
	.w1(32'h3c04ef8f),
	.w2(32'hbc0529ed),
	.w3(32'h3d5169cb),
	.w4(32'hba670e10),
	.w5(32'hbbccf433),
	.w6(32'h3bec0787),
	.w7(32'h3b99672b),
	.w8(32'hbb418026),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1c089),
	.w1(32'hbb5ccf1c),
	.w2(32'hbb993063),
	.w3(32'h3b7aadd3),
	.w4(32'h3b4c871f),
	.w5(32'hbb00e284),
	.w6(32'hbb90742a),
	.w7(32'h3b681299),
	.w8(32'h3b5cbd36),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c241809),
	.w1(32'h3b893906),
	.w2(32'hba90a5c3),
	.w3(32'h3b82eccc),
	.w4(32'hbc03e739),
	.w5(32'h397bb813),
	.w6(32'h3c6f5746),
	.w7(32'h3b884e9f),
	.w8(32'h3c905567),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2888d5),
	.w1(32'hbaf68bc6),
	.w2(32'hbcf48b1b),
	.w3(32'h3c71ff78),
	.w4(32'h3c5d4e25),
	.w5(32'hbc973655),
	.w6(32'h3bce1864),
	.w7(32'h3c3c173e),
	.w8(32'h3cba13a0),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74b49d),
	.w1(32'h3befa2a5),
	.w2(32'hb7d6861d),
	.w3(32'hbcdca514),
	.w4(32'h3bf5fe9c),
	.w5(32'h3b82e000),
	.w6(32'hbc11ad30),
	.w7(32'h3c3d9e21),
	.w8(32'h3c09cf59),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f9e35),
	.w1(32'hbb620452),
	.w2(32'hbc6dad3b),
	.w3(32'hbb9c117e),
	.w4(32'h3cf4e728),
	.w5(32'h3c5b2684),
	.w6(32'h3aedcbc9),
	.w7(32'hbbaec7b8),
	.w8(32'h3b8726e7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0434cf),
	.w1(32'h3b7fa5c0),
	.w2(32'h3bc1a628),
	.w3(32'hbb7d1125),
	.w4(32'hba6719ef),
	.w5(32'h3b250591),
	.w6(32'hbc17bff6),
	.w7(32'h3be1887a),
	.w8(32'h3bd8679f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c613f),
	.w1(32'h398cffc6),
	.w2(32'h3b63cc9c),
	.w3(32'hbc16b787),
	.w4(32'hba9f633e),
	.w5(32'h3b205b2e),
	.w6(32'hba34c601),
	.w7(32'hbc5fe299),
	.w8(32'hbab8d690),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ce9c4),
	.w1(32'h3c2db807),
	.w2(32'hbc061c54),
	.w3(32'h3bf40aa2),
	.w4(32'h3c0dcae0),
	.w5(32'h3b1e09d4),
	.w6(32'hbac74ef0),
	.w7(32'h3c24f8ef),
	.w8(32'hbadc3c71),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1378ca),
	.w1(32'h3b9ff342),
	.w2(32'h3bdf3bd8),
	.w3(32'hbc148f5a),
	.w4(32'hbaee698e),
	.w5(32'hbbffa353),
	.w6(32'hbbd9850d),
	.w7(32'hbbbf21bf),
	.w8(32'hbbdb69de),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40b445),
	.w1(32'hb9a0a0e3),
	.w2(32'h3b141a19),
	.w3(32'hbc32d4c5),
	.w4(32'hbbbad3fd),
	.w5(32'hbc11f7c5),
	.w6(32'h3992af5f),
	.w7(32'h3bf6b688),
	.w8(32'hbb2262d7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99e479),
	.w1(32'hbb72e178),
	.w2(32'hbbc9849e),
	.w3(32'hb9d6d0b1),
	.w4(32'hbc1008f1),
	.w5(32'h3aef329d),
	.w6(32'h3985ed78),
	.w7(32'hbbad8076),
	.w8(32'hbc6b4d8a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc504159),
	.w1(32'h3c26a4f4),
	.w2(32'h3c0cb794),
	.w3(32'h3c926652),
	.w4(32'h3c7326f3),
	.w5(32'hbbf7c1b3),
	.w6(32'hbbd51bed),
	.w7(32'h3b802f92),
	.w8(32'hbb7e45b0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1706cc),
	.w1(32'h3bbf6a6a),
	.w2(32'h3bb72965),
	.w3(32'hbcd7f451),
	.w4(32'h3a40a9c1),
	.w5(32'h3c373d84),
	.w6(32'hbc87c807),
	.w7(32'h3b9ace85),
	.w8(32'h3b2c85bc),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae27b7e),
	.w1(32'h39d52d68),
	.w2(32'h3c19cfd8),
	.w3(32'h3bb7e2a4),
	.w4(32'hba3b5715),
	.w5(32'hbacef1f7),
	.w6(32'h3ab4cda1),
	.w7(32'hbb6fbdb9),
	.w8(32'h3b0c0074),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16f6b0),
	.w1(32'hbae11ad9),
	.w2(32'h3ba4f055),
	.w3(32'hbba22e48),
	.w4(32'hbbeeae4a),
	.w5(32'h3bdcef15),
	.w6(32'h3bba859e),
	.w7(32'hbc482809),
	.w8(32'h3a2db11c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9fd94),
	.w1(32'hbb461bec),
	.w2(32'hbbd484f1),
	.w3(32'hbafabe1b),
	.w4(32'hbcaaa1bb),
	.w5(32'hbd231893),
	.w6(32'h3b0d999a),
	.w7(32'h3b20b5b5),
	.w8(32'hb9e15ed3),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb4ec),
	.w1(32'h3bd3f61b),
	.w2(32'h3c5330a3),
	.w3(32'h3b868177),
	.w4(32'h3befe1b1),
	.w5(32'hbcd9bc8c),
	.w6(32'h3c18e981),
	.w7(32'h3b99eae7),
	.w8(32'hbb97fb61),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31b7e8),
	.w1(32'h3ad29a21),
	.w2(32'hbc29d601),
	.w3(32'hbb46559e),
	.w4(32'h3b8b294a),
	.w5(32'hbccfda34),
	.w6(32'h38e257a0),
	.w7(32'h3b90362b),
	.w8(32'hbc557216),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eb5996),
	.w1(32'hba33841d),
	.w2(32'h3b9bc7fc),
	.w3(32'h3b619d3b),
	.w4(32'hba031150),
	.w5(32'h3c3c9f3c),
	.w6(32'hbc292fd6),
	.w7(32'hbb22f846),
	.w8(32'h3a94f938),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9f24b),
	.w1(32'hbb4fa656),
	.w2(32'hba0abd8c),
	.w3(32'hbbbf52f1),
	.w4(32'hbbf2514b),
	.w5(32'hbb95ea14),
	.w6(32'hbb220c0d),
	.w7(32'hbbd8fc0d),
	.w8(32'hbbb470f0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85ae47),
	.w1(32'h3a96af9e),
	.w2(32'hbbb76bee),
	.w3(32'hbbf85a24),
	.w4(32'hbc287a37),
	.w5(32'h3aa3d5be),
	.w6(32'hbc1c5654),
	.w7(32'h3b19ebf6),
	.w8(32'hbbe91cd2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97808a),
	.w1(32'hbb328d51),
	.w2(32'h3bb20b3a),
	.w3(32'h393d87ab),
	.w4(32'hbb13d696),
	.w5(32'hb990d90b),
	.w6(32'h3b46518e),
	.w7(32'hbb749edf),
	.w8(32'hba8a8b83),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e7d88),
	.w1(32'h3a5aded1),
	.w2(32'h3b3d4bf0),
	.w3(32'hbbf42aa8),
	.w4(32'h3aa351b2),
	.w5(32'hbad31160),
	.w6(32'h3b16eac1),
	.w7(32'hbb92b594),
	.w8(32'hbb4a1a8a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb421475),
	.w1(32'hbaff9b5d),
	.w2(32'hbb8bae24),
	.w3(32'h3a4ebab6),
	.w4(32'hbb8ef6e2),
	.w5(32'h3c0875e6),
	.w6(32'hb73b4e8c),
	.w7(32'hbb84b35a),
	.w8(32'hbb6a41b2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdac481),
	.w1(32'hbb615222),
	.w2(32'hbb8ffaa9),
	.w3(32'hbbe40bc5),
	.w4(32'hbb35b538),
	.w5(32'h3b928a21),
	.w6(32'hbc1051da),
	.w7(32'hb9811921),
	.w8(32'hbaa1c82b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf14e07),
	.w1(32'hbbb27dc8),
	.w2(32'hbb9125b4),
	.w3(32'h3b702059),
	.w4(32'h3a963324),
	.w5(32'h3adc2ac7),
	.w6(32'h3bcc76e1),
	.w7(32'hbba7ec6d),
	.w8(32'hba1e97c9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06c9b9),
	.w1(32'h3b4505e8),
	.w2(32'hbab09eae),
	.w3(32'hbb2b31d5),
	.w4(32'hbbf1ba0f),
	.w5(32'hbc39133e),
	.w6(32'h3a5050ab),
	.w7(32'hbba790b6),
	.w8(32'hbad9a439),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8079f0),
	.w1(32'hbb0c313d),
	.w2(32'hba6e9d11),
	.w3(32'h3baa1589),
	.w4(32'hbb17ae91),
	.w5(32'h3a2899fc),
	.w6(32'h3c09c2bc),
	.w7(32'h3b3f5819),
	.w8(32'h3b57060b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59929),
	.w1(32'h3b27c039),
	.w2(32'hbadc76d8),
	.w3(32'h3b713094),
	.w4(32'hbae3ed8d),
	.w5(32'hbb92e98a),
	.w6(32'h3b5075a2),
	.w7(32'hbb4b4044),
	.w8(32'h3a49645b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60e0e5),
	.w1(32'h3bc6749a),
	.w2(32'hba825393),
	.w3(32'h3c17a18a),
	.w4(32'hba6fdbfb),
	.w5(32'hbc0c6801),
	.w6(32'h3b89c2fc),
	.w7(32'hba5352ea),
	.w8(32'h3ad17766),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1367),
	.w1(32'hbb1c75f7),
	.w2(32'hbb7988fe),
	.w3(32'hbc14fb8e),
	.w4(32'hbba065a6),
	.w5(32'hbb68d346),
	.w6(32'hba10bd42),
	.w7(32'hbb8bed7f),
	.w8(32'h3a217432),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc03a89),
	.w1(32'hb99c54c3),
	.w2(32'hba6b6960),
	.w3(32'h39ce6a0c),
	.w4(32'hbb09af1f),
	.w5(32'hbb0c52ea),
	.w6(32'h3b99c330),
	.w7(32'hbaa1cfb0),
	.w8(32'hbafb77c1),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ae2ed3),
	.w1(32'hbc02bc3c),
	.w2(32'h3beef5ec),
	.w3(32'hba6d6da1),
	.w4(32'hbb32af7c),
	.w5(32'h3bc62c0d),
	.w6(32'h3ae20dcc),
	.w7(32'hbb81fb6a),
	.w8(32'h3b73b428),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49f0e6),
	.w1(32'hb9c9ef44),
	.w2(32'h3b946beb),
	.w3(32'hbb81785c),
	.w4(32'hbb5ea538),
	.w5(32'h3b11db5d),
	.w6(32'hba7b03f8),
	.w7(32'hbae899fc),
	.w8(32'h3a89b3a1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb511e99),
	.w1(32'hbba211bd),
	.w2(32'h3a41cd8d),
	.w3(32'h3a4a7aa5),
	.w4(32'h3bfea2ac),
	.w5(32'hbb2f933d),
	.w6(32'h3b080c1b),
	.w7(32'hbb4e351d),
	.w8(32'h3b495c55),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba48901),
	.w1(32'h3b7d7f25),
	.w2(32'h3bd9cfaa),
	.w3(32'h3c41afc7),
	.w4(32'hbb3d1b78),
	.w5(32'hbc8ae1d3),
	.w6(32'hb9d79ac6),
	.w7(32'hbbe69f89),
	.w8(32'hbaeb4cc9),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c557f5e),
	.w1(32'h3b4f46fb),
	.w2(32'h3c0e35dd),
	.w3(32'h3b3002f5),
	.w4(32'h3beffe0d),
	.w5(32'hbc88afde),
	.w6(32'hbc24f1cd),
	.w7(32'h3c0fc903),
	.w8(32'h3c11ef49),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe49d3),
	.w1(32'hbc074a1f),
	.w2(32'hbb303b3a),
	.w3(32'h3b0ac4a6),
	.w4(32'h3b89dc05),
	.w5(32'h3bf743da),
	.w6(32'h3a802355),
	.w7(32'hb9be5f2f),
	.w8(32'hba15599f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e153f),
	.w1(32'hbb6bc530),
	.w2(32'h3ba4d573),
	.w3(32'h3977ce1f),
	.w4(32'h3b6b510f),
	.w5(32'h3c25d15e),
	.w6(32'hbba26df1),
	.w7(32'hbc0936ef),
	.w8(32'h3b5b5692),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c480da9),
	.w1(32'h3be48cda),
	.w2(32'h3bd52655),
	.w3(32'h3b44439a),
	.w4(32'h37491d0e),
	.w5(32'h3b835104),
	.w6(32'h3b835452),
	.w7(32'hbb5290ba),
	.w8(32'h3c09dc29),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d1f2f),
	.w1(32'h3ad0f8e8),
	.w2(32'h3c64424f),
	.w3(32'h3b39122e),
	.w4(32'hbac344f0),
	.w5(32'hbbde9fda),
	.w6(32'h39a4ebdc),
	.w7(32'hba18c942),
	.w8(32'h3c8c564d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e4464),
	.w1(32'hbb5860bf),
	.w2(32'hbb138ea7),
	.w3(32'h3b3a32be),
	.w4(32'h39e105e5),
	.w5(32'hbb5b8ec5),
	.w6(32'h3bb6c1fc),
	.w7(32'h3bcdc23e),
	.w8(32'h3b86d36d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba519aa1),
	.w1(32'hb9530540),
	.w2(32'h376adad8),
	.w3(32'h3b978738),
	.w4(32'h3b99e3f8),
	.w5(32'hbbbc3483),
	.w6(32'h3b9ed874),
	.w7(32'h3c028d59),
	.w8(32'hba58d5e1),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac01299),
	.w1(32'hbbfde10a),
	.w2(32'hbc169b53),
	.w3(32'hbb67318b),
	.w4(32'hbbb9ccd5),
	.w5(32'hbb0cde30),
	.w6(32'h3b49cfdd),
	.w7(32'hbadba05a),
	.w8(32'hba3d8916),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382856d1),
	.w1(32'hbaf28749),
	.w2(32'h3a72cc95),
	.w3(32'h3c3af514),
	.w4(32'hbb1f5364),
	.w5(32'h3c491b33),
	.w6(32'hbbb24ebc),
	.w7(32'h3b8e32e4),
	.w8(32'hbb50c6bc),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e8a45),
	.w1(32'h3af9719d),
	.w2(32'h3b02c8db),
	.w3(32'hbba65780),
	.w4(32'h3a9b599d),
	.w5(32'hbc15965e),
	.w6(32'hbc0060ce),
	.w7(32'hba6c8d9f),
	.w8(32'hba42cf41),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c88a1),
	.w1(32'h3a9be512),
	.w2(32'hbb72dd23),
	.w3(32'h39b89ccd),
	.w4(32'hb9b0e000),
	.w5(32'hbbafebd0),
	.w6(32'hbaa0a6de),
	.w7(32'h3adcf2e4),
	.w8(32'hbbc46372),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b966e71),
	.w1(32'hbb6e1ca4),
	.w2(32'hba4cfb6e),
	.w3(32'h3ab1fd90),
	.w4(32'h3a604058),
	.w5(32'h3c38b352),
	.w6(32'h3ada0bae),
	.w7(32'hbbe34b2c),
	.w8(32'h3aed4907),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b200),
	.w1(32'h3bb391e7),
	.w2(32'h3b4ac11e),
	.w3(32'hba33e212),
	.w4(32'h3b2505e4),
	.w5(32'h3ca63a7f),
	.w6(32'hbc3f5661),
	.w7(32'hbb5f4e86),
	.w8(32'hbc101d41),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5ffbc),
	.w1(32'h3935aad5),
	.w2(32'hb892324d),
	.w3(32'h3ba492ff),
	.w4(32'h3aa4b6a6),
	.w5(32'hbb2bed8a),
	.w6(32'hbb369a47),
	.w7(32'hbb6f12f8),
	.w8(32'hbb9a65aa),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f88d4),
	.w1(32'h3b07b68f),
	.w2(32'hbbac1e4a),
	.w3(32'h3acd7f43),
	.w4(32'h3ba3a9d8),
	.w5(32'h3bbcd2d8),
	.w6(32'hbb9b222e),
	.w7(32'h37d7b8f4),
	.w8(32'hbbaa59ca),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00abfb),
	.w1(32'hbb9d7f9c),
	.w2(32'h3c113a68),
	.w3(32'h3b13dc86),
	.w4(32'hbbe37312),
	.w5(32'h3c0d80e3),
	.w6(32'hbad2345f),
	.w7(32'hbbf594ce),
	.w8(32'hbb00fedb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdd00a),
	.w1(32'h3b1676cd),
	.w2(32'hba570c54),
	.w3(32'h3b6cb950),
	.w4(32'hbb0f75d2),
	.w5(32'h3a3d1839),
	.w6(32'h3983c34a),
	.w7(32'hba860489),
	.w8(32'h3b844e79),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50225a),
	.w1(32'h3b0bf0b7),
	.w2(32'hba9d42cb),
	.w3(32'h39ee413b),
	.w4(32'hb9c71135),
	.w5(32'hbb65a859),
	.w6(32'h3b6bb7b9),
	.w7(32'h3b0e2a32),
	.w8(32'h3bc5f4c0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3348dd),
	.w1(32'h3b94f09f),
	.w2(32'h3b239ffd),
	.w3(32'h3bc070fb),
	.w4(32'h3b21b91e),
	.w5(32'hbad63dc0),
	.w6(32'h3ad22f4a),
	.w7(32'h3b7cbeb8),
	.w8(32'hb8181388),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafea9a2),
	.w1(32'h3a595b51),
	.w2(32'hb91edba1),
	.w3(32'h3b0c63b7),
	.w4(32'hb9ac4893),
	.w5(32'hba306b8c),
	.w6(32'h3b07f55e),
	.w7(32'hbb2a39ec),
	.w8(32'hb91eb2dd),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75c5f6),
	.w1(32'h3a992d95),
	.w2(32'hba84777d),
	.w3(32'h3b4b0c0f),
	.w4(32'h391ea476),
	.w5(32'hba17d86d),
	.w6(32'h3b5d1669),
	.w7(32'h3a959739),
	.w8(32'h3bc183ca),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c448199),
	.w1(32'hbb4c50d5),
	.w2(32'hbbba9de4),
	.w3(32'hba9c057d),
	.w4(32'hbbcf7781),
	.w5(32'h3985d8fd),
	.w6(32'h3b555b06),
	.w7(32'h3b5d35b5),
	.w8(32'hbaac8897),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3e5ee),
	.w1(32'h3ba74cb5),
	.w2(32'h3ad904d0),
	.w3(32'h3b9148b7),
	.w4(32'h3b519da0),
	.w5(32'hbc6c1c2d),
	.w6(32'hb98f5eb5),
	.w7(32'h37c5d87d),
	.w8(32'hbb9d1c4e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c106143),
	.w1(32'hbb2eb950),
	.w2(32'hbc12b701),
	.w3(32'h3a188bcf),
	.w4(32'hbb4548f6),
	.w5(32'hbb5ddf41),
	.w6(32'hbb690cff),
	.w7(32'hbb80ce88),
	.w8(32'hbb6794cb),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b028954),
	.w1(32'h3bc638f5),
	.w2(32'h3bef1be8),
	.w3(32'hbb139206),
	.w4(32'h3a13348a),
	.w5(32'h3b8d5c20),
	.w6(32'h3a2f6bdd),
	.w7(32'hbb0221b7),
	.w8(32'hbb7499b3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6dae3),
	.w1(32'h3b68af78),
	.w2(32'h3c3d6938),
	.w3(32'h3aa743e5),
	.w4(32'h3aefc8f3),
	.w5(32'hbb42faf0),
	.w6(32'hba8dd21d),
	.w7(32'hbbd2889b),
	.w8(32'hbb7e0931),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a20cd),
	.w1(32'h3c5966c8),
	.w2(32'h3c0954f5),
	.w3(32'h3a84b6ce),
	.w4(32'h3c050beb),
	.w5(32'h3ae06c5b),
	.w6(32'h3ac170ea),
	.w7(32'hbb49baa2),
	.w8(32'hbb91ddd2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa6d02),
	.w1(32'hbb5a68d8),
	.w2(32'h3c301ef3),
	.w3(32'hbafd9d93),
	.w4(32'h3c3b8806),
	.w5(32'h3b760ee0),
	.w6(32'h39de333a),
	.w7(32'h3c16a295),
	.w8(32'hbb7fd6f8),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd86c6),
	.w1(32'hbb6656be),
	.w2(32'hbb2c93ee),
	.w3(32'h3b9ab574),
	.w4(32'hbbdddfb0),
	.w5(32'hbb14f1ac),
	.w6(32'h3ba5cb50),
	.w7(32'hbbe65ce0),
	.w8(32'hbbd02799),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90abfba),
	.w1(32'hbb649fec),
	.w2(32'h3c001b81),
	.w3(32'hbb9a930f),
	.w4(32'h3a8d6137),
	.w5(32'hb99a356a),
	.w6(32'hbb8f7002),
	.w7(32'h3a66b79b),
	.w8(32'h3a149648),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3c810),
	.w1(32'hba0a935a),
	.w2(32'hbaf8a345),
	.w3(32'h3b93ba29),
	.w4(32'hbacea403),
	.w5(32'hbb9842c8),
	.w6(32'h3ae61822),
	.w7(32'hbb0cb396),
	.w8(32'hbb5577a7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aea0a),
	.w1(32'h3bce11fb),
	.w2(32'h3c0e33a9),
	.w3(32'h3b464120),
	.w4(32'h3b90bdb8),
	.w5(32'h3b8ecf86),
	.w6(32'h3b94ebdd),
	.w7(32'hb96100eb),
	.w8(32'h3b8a30e2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5754d8),
	.w1(32'h3b805ec6),
	.w2(32'h3b415727),
	.w3(32'h3ba6707d),
	.w4(32'hbbc2d6b6),
	.w5(32'h3b04fa6e),
	.w6(32'h3b5d1b08),
	.w7(32'hbb4674f8),
	.w8(32'hbb9cd393),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c299476),
	.w1(32'hbba70a6d),
	.w2(32'hbab5ad39),
	.w3(32'hb792c4d4),
	.w4(32'hbaf39b55),
	.w5(32'hba877c42),
	.w6(32'hbacb13cf),
	.w7(32'hbbaad259),
	.w8(32'hbaa42eea),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58d83f),
	.w1(32'hb82ff0c3),
	.w2(32'hbafb38b1),
	.w3(32'hbb24267c),
	.w4(32'hbc24502d),
	.w5(32'h3c8701a2),
	.w6(32'hbb798c66),
	.w7(32'h3babf5fc),
	.w8(32'h3c2eca2b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12e72b),
	.w1(32'hbb8b6052),
	.w2(32'h3b29fbca),
	.w3(32'h3be0a417),
	.w4(32'hba8d4946),
	.w5(32'hbb909fc6),
	.w6(32'hbb885c48),
	.w7(32'hbb74c143),
	.w8(32'h3aa3c7a7),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908da1f),
	.w1(32'h3a7b1b3c),
	.w2(32'h3a33c2f3),
	.w3(32'hbae89dcf),
	.w4(32'h3b930088),
	.w5(32'h3c001358),
	.w6(32'hbbe21db1),
	.w7(32'hbb6e53ad),
	.w8(32'h3b849ea7),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb633c08),
	.w1(32'hb91f1e5f),
	.w2(32'hbbf8bcc1),
	.w3(32'h3b8466f4),
	.w4(32'hbbe4253d),
	.w5(32'h3b4413b0),
	.w6(32'h3b8b7174),
	.w7(32'h3b7addea),
	.w8(32'hbb07f833),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63bd4e),
	.w1(32'h3bc29762),
	.w2(32'h3c4badb8),
	.w3(32'h3bcb81a5),
	.w4(32'h3b2f7c68),
	.w5(32'h3ba7a9cb),
	.w6(32'h3bf4451b),
	.w7(32'h3b387816),
	.w8(32'hbbe1138f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8da49db),
	.w1(32'h3b84b718),
	.w2(32'h3bebd342),
	.w3(32'hbb254a40),
	.w4(32'h3be7eb2a),
	.w5(32'h3c09f9fe),
	.w6(32'hbbb419ef),
	.w7(32'h3a4dff26),
	.w8(32'hba7da133),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd18825),
	.w1(32'hbbb457bc),
	.w2(32'hba7133c1),
	.w3(32'h3b93e9f1),
	.w4(32'hbbf06965),
	.w5(32'h3aebe0ff),
	.w6(32'h3b11d12f),
	.w7(32'hbb918c84),
	.w8(32'hbb8aec29),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule