module layer_10_featuremap_451(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b083196),
	.w1(32'h3b7c5124),
	.w2(32'hbb082d3a),
	.w3(32'hbaa863e8),
	.w4(32'h3b83085d),
	.w5(32'hbb338e89),
	.w6(32'hbc1eb226),
	.w7(32'hb9b26733),
	.w8(32'hbbc6e1ca),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea18b5),
	.w1(32'h3bca8922),
	.w2(32'h3c2cb663),
	.w3(32'h3b542396),
	.w4(32'h3b26bd31),
	.w5(32'h3c2d9d1f),
	.w6(32'hba9c3446),
	.w7(32'h399eef1e),
	.w8(32'h3beeddeb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15b3ae),
	.w1(32'hbb8952a8),
	.w2(32'h392d9d4f),
	.w3(32'h3c1b94ec),
	.w4(32'hbb6d9c2a),
	.w5(32'hb7636f23),
	.w6(32'h3be8f2f1),
	.w7(32'h3b754162),
	.w8(32'hba175c32),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adedcfe),
	.w1(32'hbb9254e8),
	.w2(32'hbae03f0c),
	.w3(32'h39b25481),
	.w4(32'hba8d1cf1),
	.w5(32'hbaf37e65),
	.w6(32'hbab79d70),
	.w7(32'hbae5f797),
	.w8(32'hba5f59e5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1353b0),
	.w1(32'h3acc3895),
	.w2(32'h3b9962e4),
	.w3(32'h3af75b0c),
	.w4(32'h3aa2e5b9),
	.w5(32'h3c882dc1),
	.w6(32'h3a9cc95c),
	.w7(32'h39e4d77a),
	.w8(32'h3ba38178),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f8137),
	.w1(32'h3b951dc1),
	.w2(32'h3b3c4b05),
	.w3(32'h3c133f82),
	.w4(32'h38fbfe81),
	.w5(32'h3bca8e11),
	.w6(32'h3bece231),
	.w7(32'h3aac252b),
	.w8(32'h3b9050cf),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0abf29),
	.w1(32'hb9e983b5),
	.w2(32'hbae46485),
	.w3(32'h3bbd89b9),
	.w4(32'hbb09e782),
	.w5(32'hbbfc5b7b),
	.w6(32'hb9e1919a),
	.w7(32'hbb919ab5),
	.w8(32'hbb70eba9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb713ba),
	.w1(32'hbbb90be2),
	.w2(32'hbb737093),
	.w3(32'hbc5cfcad),
	.w4(32'hbba620f7),
	.w5(32'h3b93b7ad),
	.w6(32'hbc0b342f),
	.w7(32'hbb92f491),
	.w8(32'hbb6c69c7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c6943),
	.w1(32'hbb96f23b),
	.w2(32'hbaa636e2),
	.w3(32'hb7fa45ab),
	.w4(32'hba60ba27),
	.w5(32'h3b047c3b),
	.w6(32'hbb857312),
	.w7(32'hbb955f73),
	.w8(32'hbae931e7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d70c3),
	.w1(32'hb93328f7),
	.w2(32'hba3d67c9),
	.w3(32'h3affe0e4),
	.w4(32'h3b9e690d),
	.w5(32'h3b307c38),
	.w6(32'hbb2ca1ed),
	.w7(32'hba76903c),
	.w8(32'hbb634159),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a1796),
	.w1(32'h3b0c6a69),
	.w2(32'h3b402cb6),
	.w3(32'h3b7d2995),
	.w4(32'h3accbdf3),
	.w5(32'h3b587314),
	.w6(32'hba24d195),
	.w7(32'hb9f32da8),
	.w8(32'h3b2e6c64),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae35827),
	.w1(32'h3bb1d16f),
	.w2(32'h3b226fd1),
	.w3(32'h3bfa75be),
	.w4(32'h3b86cd9e),
	.w5(32'h3ac168ad),
	.w6(32'h3c08395d),
	.w7(32'h39f34fff),
	.w8(32'hb9a7aa62),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb128e22),
	.w1(32'h3a520340),
	.w2(32'hbbf4c65d),
	.w3(32'hbb919cca),
	.w4(32'h38b56644),
	.w5(32'hbc16c67c),
	.w6(32'hbb52ed15),
	.w7(32'hbb05d81d),
	.w8(32'hbc22dbd3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c3e1f),
	.w1(32'h3b620182),
	.w2(32'hbae52aa9),
	.w3(32'hbba88c07),
	.w4(32'hb94b703f),
	.w5(32'hbace158e),
	.w6(32'hbbda3b1f),
	.w7(32'hbb831f32),
	.w8(32'hb895a1ad),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ac84d),
	.w1(32'hbb0faad6),
	.w2(32'hbb00c9f8),
	.w3(32'hbac19f09),
	.w4(32'hbb6ca373),
	.w5(32'hbace881c),
	.w6(32'hbb1ee6bb),
	.w7(32'h3a96feb4),
	.w8(32'hba6d09aa),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb517f77),
	.w1(32'h39f1006d),
	.w2(32'hbb25f71d),
	.w3(32'hbb90dc4b),
	.w4(32'hbbb8fc62),
	.w5(32'hbbc9f1b7),
	.w6(32'hbc0b0383),
	.w7(32'hbb7bbf13),
	.w8(32'hbc010803),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fab0d),
	.w1(32'h3a0c3005),
	.w2(32'h395232ab),
	.w3(32'hba8cd5aa),
	.w4(32'h3bc1aedb),
	.w5(32'h3a42ef34),
	.w6(32'hbb72db81),
	.w7(32'hb9a8bca1),
	.w8(32'h39b9673c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05cc14),
	.w1(32'hbc02a431),
	.w2(32'hbc4605a0),
	.w3(32'hbc97632c),
	.w4(32'hbbc1cd5d),
	.w5(32'hba67bdd0),
	.w6(32'hbc3a6e8d),
	.w7(32'hbbbf1175),
	.w8(32'h39182ac2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39688dd1),
	.w1(32'hbb061389),
	.w2(32'hbaa5efd8),
	.w3(32'hbb00c4d1),
	.w4(32'hb9d60308),
	.w5(32'h3b7cde98),
	.w6(32'hbb6a036c),
	.w7(32'hbb8c7e7e),
	.w8(32'hbb306e41),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ce5e6),
	.w1(32'hbbaf5f38),
	.w2(32'hbc1ed603),
	.w3(32'h39428b19),
	.w4(32'h3ba310f9),
	.w5(32'hbb8c4434),
	.w6(32'h394954e5),
	.w7(32'hb8bec57b),
	.w8(32'hbb320e35),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22b3a3),
	.w1(32'hbb9bad4b),
	.w2(32'hbb14fb8b),
	.w3(32'hbc015379),
	.w4(32'hbbc16f44),
	.w5(32'h3b1b5746),
	.w6(32'hbae556ad),
	.w7(32'hbb2aff9e),
	.w8(32'h39c084f7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb7073),
	.w1(32'hbacb2f84),
	.w2(32'hbb3f401e),
	.w3(32'h3b26fbc6),
	.w4(32'h3a32ec4e),
	.w5(32'hbb8289e9),
	.w6(32'hba172c05),
	.w7(32'h3b69ec92),
	.w8(32'hb98a7a73),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e64d7),
	.w1(32'hbc7c3ca2),
	.w2(32'hbbf5c35b),
	.w3(32'hbccb7885),
	.w4(32'hbb64e574),
	.w5(32'hbbe90af9),
	.w6(32'hbc83c412),
	.w7(32'hbc317401),
	.w8(32'hbc276063),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a029d),
	.w1(32'h3aa2a7b4),
	.w2(32'h3b814e2c),
	.w3(32'hbb9eb789),
	.w4(32'h3992e6ff),
	.w5(32'h3b62e5a5),
	.w6(32'hbc23a34f),
	.w7(32'hb9949066),
	.w8(32'h3bec176c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39837ca5),
	.w1(32'h3ba1fc9d),
	.w2(32'h3b449290),
	.w3(32'h3bfef1ee),
	.w4(32'h3b307547),
	.w5(32'hbae62869),
	.w6(32'h3c279dfa),
	.w7(32'hbb266a6f),
	.w8(32'h3aad1871),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f29dc),
	.w1(32'hbc13215e),
	.w2(32'hbbc21bbb),
	.w3(32'hbaf42a50),
	.w4(32'hbc3adec8),
	.w5(32'hba4e6cdb),
	.w6(32'hbb27c78c),
	.w7(32'hbc274c6c),
	.w8(32'hbae5184a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2524c),
	.w1(32'hbbc0e82a),
	.w2(32'hb9e6c824),
	.w3(32'hbbd9fe03),
	.w4(32'h3ba99a2a),
	.w5(32'h3c4c5519),
	.w6(32'hbb4f6c7c),
	.w7(32'h3b8bfed7),
	.w8(32'h3ae90b01),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c198115),
	.w1(32'h3b8a3839),
	.w2(32'h3b878c86),
	.w3(32'h3c126ceb),
	.w4(32'h3bc1ce92),
	.w5(32'h3b061e19),
	.w6(32'hbb685816),
	.w7(32'h3bb41b73),
	.w8(32'h3b8dca75),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42adfc),
	.w1(32'hbbb69c9f),
	.w2(32'hbbf224f6),
	.w3(32'h3b69a8b9),
	.w4(32'hba82750b),
	.w5(32'hb9c5f1c8),
	.w6(32'h3b871bcc),
	.w7(32'hbb01fede),
	.w8(32'hb7cfff1f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989245),
	.w1(32'h3afac85e),
	.w2(32'h3b36c833),
	.w3(32'h3b859428),
	.w4(32'hbaa0520b),
	.w5(32'hba2e0c78),
	.w6(32'h3b5ae6ca),
	.w7(32'hba8f1097),
	.w8(32'hbb2fac03),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd8952),
	.w1(32'hbb554b16),
	.w2(32'hbb215a5a),
	.w3(32'h3b8b5b69),
	.w4(32'h3ab5004c),
	.w5(32'h3af0912d),
	.w6(32'h3b0abb04),
	.w7(32'hbaadf10b),
	.w8(32'hb971db36),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dedb8),
	.w1(32'h3a18a321),
	.w2(32'hbaa58aa9),
	.w3(32'hbae10d64),
	.w4(32'hba169fdc),
	.w5(32'hbb70b8da),
	.w6(32'hbb3195c4),
	.w7(32'h3b6b5fa8),
	.w8(32'hbad484da),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a325dfc),
	.w1(32'hba9d5db5),
	.w2(32'hbbb8300a),
	.w3(32'hbad07c0d),
	.w4(32'h3be3cc5c),
	.w5(32'h3b21d940),
	.w6(32'hbb0d5826),
	.w7(32'h37a0b11c),
	.w8(32'hb8c26596),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb929e57),
	.w1(32'h3c164af3),
	.w2(32'h3c347407),
	.w3(32'h3b3e14c3),
	.w4(32'h3be7ef8c),
	.w5(32'h3bf1aa94),
	.w6(32'h39ca43c6),
	.w7(32'hbb136a77),
	.w8(32'hbadb8555),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c91a4),
	.w1(32'h3a5c1bbe),
	.w2(32'hbb70052c),
	.w3(32'h3b55e516),
	.w4(32'hbaeacbaf),
	.w5(32'h3a8171a8),
	.w6(32'hb9ccbfae),
	.w7(32'hbb518da7),
	.w8(32'h3aa87774),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb966dd5),
	.w1(32'h3b98a8f8),
	.w2(32'h3accf524),
	.w3(32'hbb9008e6),
	.w4(32'h3b11c222),
	.w5(32'hbb586e3b),
	.w6(32'hbb4dec2e),
	.w7(32'hb98b62e1),
	.w8(32'hba7d0e4a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fe757),
	.w1(32'hbb9a80be),
	.w2(32'h3bf6cefa),
	.w3(32'hbb996e72),
	.w4(32'hbbf023db),
	.w5(32'h3bfa6671),
	.w6(32'hbba22478),
	.w7(32'hbbb10852),
	.w8(32'hbb2cec2f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87fbae),
	.w1(32'h3bb49b4e),
	.w2(32'h3b87439c),
	.w3(32'h3c324eee),
	.w4(32'h3c2f4401),
	.w5(32'h3aca4af8),
	.w6(32'hbb0e26ff),
	.w7(32'h3bdcffd6),
	.w8(32'h3bd0e6db),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e0c89),
	.w1(32'h3a81c888),
	.w2(32'hbb72c472),
	.w3(32'h3c7ee7d9),
	.w4(32'h3a81ce2b),
	.w5(32'hbbd3173b),
	.w6(32'h3c81b925),
	.w7(32'h3b7cedf2),
	.w8(32'hbb53422b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab8966),
	.w1(32'h3aa445af),
	.w2(32'hbab055d2),
	.w3(32'hba21f986),
	.w4(32'h3b481f87),
	.w5(32'h3a72baa6),
	.w6(32'h3a0b4cc8),
	.w7(32'hbadfb74f),
	.w8(32'hb98e32c4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53f723),
	.w1(32'h3a585108),
	.w2(32'hbb66bbae),
	.w3(32'h3ae18a8f),
	.w4(32'h3b67b2a2),
	.w5(32'hbbb2099b),
	.w6(32'h3b60b3d1),
	.w7(32'h39f14698),
	.w8(32'h3aaa43fb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f0e6c),
	.w1(32'hb9a4a50e),
	.w2(32'h3b47c2eb),
	.w3(32'h3babc9f0),
	.w4(32'hba5fefe7),
	.w5(32'h3ba486f5),
	.w6(32'h3904c175),
	.w7(32'h3b024f28),
	.w8(32'h3b7b8853),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eceff),
	.w1(32'h3a4d5eac),
	.w2(32'h39996222),
	.w3(32'hbae11dfb),
	.w4(32'h3b94185a),
	.w5(32'hbaae09d0),
	.w6(32'hbb2ec43b),
	.w7(32'hbb1ef67a),
	.w8(32'hbb60152b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf24bba),
	.w1(32'hba0810de),
	.w2(32'hbc1f711b),
	.w3(32'hbbfb96f1),
	.w4(32'hb9977ac5),
	.w5(32'hbc0a3291),
	.w6(32'hbc41cce2),
	.w7(32'h3aa440c4),
	.w8(32'hbb896985),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba93ebf),
	.w1(32'h3b8dd04a),
	.w2(32'h3ab3a20d),
	.w3(32'hbb6c8279),
	.w4(32'h3ac6cce6),
	.w5(32'h3b1f88ff),
	.w6(32'hbb93449b),
	.w7(32'h3ab7febe),
	.w8(32'h3b16d2ff),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084e58),
	.w1(32'hbafaa301),
	.w2(32'hbaf0da13),
	.w3(32'h3b583f1e),
	.w4(32'hbb9640fb),
	.w5(32'hbbe62a76),
	.w6(32'hbaf59a8b),
	.w7(32'hb9ff39ac),
	.w8(32'hbbb9f5e7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6b6f4),
	.w1(32'hbbbd2115),
	.w2(32'hbb644b1a),
	.w3(32'hbbbf25ee),
	.w4(32'hbbbcdd8a),
	.w5(32'h3a157275),
	.w6(32'hbbf5c558),
	.w7(32'h3ace992f),
	.w8(32'h3a5976f8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bd2ce),
	.w1(32'hbc71bb94),
	.w2(32'hbca6be1f),
	.w3(32'hbc06005e),
	.w4(32'hbc46f1f4),
	.w5(32'hbc401e3a),
	.w6(32'hbafc53db),
	.w7(32'hbc2237b6),
	.w8(32'hbc12a06e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae92b2b),
	.w1(32'hb91350ad),
	.w2(32'h39ce393f),
	.w3(32'hba77c83f),
	.w4(32'h3a2a3a51),
	.w5(32'h3af48b02),
	.w6(32'h3b0e17f8),
	.w7(32'hbb679102),
	.w8(32'hb99d64de),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96370d),
	.w1(32'hb8f5c64d),
	.w2(32'hbb9ff4ca),
	.w3(32'hbbaf1416),
	.w4(32'hba0eed98),
	.w5(32'hbb95d968),
	.w6(32'hbb606df8),
	.w7(32'h3b7695a8),
	.w8(32'hba9407a1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36edd2),
	.w1(32'h3aa8a20c),
	.w2(32'h3a75cd6a),
	.w3(32'hb9120219),
	.w4(32'hbb19131b),
	.w5(32'h3c346844),
	.w6(32'hb9be791b),
	.w7(32'hbb55a140),
	.w8(32'h3b82ca3d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e5389),
	.w1(32'hbb231705),
	.w2(32'h3b591065),
	.w3(32'hbb35ca5f),
	.w4(32'hbbb770dd),
	.w5(32'hbaa9fc52),
	.w6(32'h3ad8e5dc),
	.w7(32'hbb5bdd33),
	.w8(32'hba1e259a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2e3f5),
	.w1(32'h3aecac55),
	.w2(32'h3b0e9aa4),
	.w3(32'h3be72c31),
	.w4(32'h3931bb59),
	.w5(32'h3adcb3d6),
	.w6(32'h3ba33011),
	.w7(32'h3aad2bbc),
	.w8(32'h3affaf86),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfcc90),
	.w1(32'hbc100651),
	.w2(32'hbbc5c5af),
	.w3(32'hbc1d5c4b),
	.w4(32'hbc07ae6f),
	.w5(32'hbabde6db),
	.w6(32'hbbeccb75),
	.w7(32'hbc0afa3a),
	.w8(32'hba5bc07d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb207f7e),
	.w1(32'h3bbed727),
	.w2(32'h3b34598c),
	.w3(32'hbab07bc1),
	.w4(32'h3c3dfc12),
	.w5(32'h3c093050),
	.w6(32'hbb8aa9d3),
	.w7(32'h3b05af1f),
	.w8(32'h3b740be6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1856e5),
	.w1(32'h3aa92126),
	.w2(32'hba8bdcd3),
	.w3(32'h3a58822c),
	.w4(32'h3b83b4ad),
	.w5(32'h3afeaf51),
	.w6(32'h3b8504d0),
	.w7(32'hb9cebd4d),
	.w8(32'h3b43ae58),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc6f02),
	.w1(32'h3ba00caf),
	.w2(32'h388f0af6),
	.w3(32'hbb617202),
	.w4(32'h3bfc1b01),
	.w5(32'h3bd7637d),
	.w6(32'hbb3d5f03),
	.w7(32'h3b5962ff),
	.w8(32'h3b63be03),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a254c91),
	.w1(32'h3a375697),
	.w2(32'h3b2f477f),
	.w3(32'h3aed68d8),
	.w4(32'hbb76113e),
	.w5(32'h3c4b4104),
	.w6(32'hba1dda11),
	.w7(32'h3a8c1bd9),
	.w8(32'h3bce1726),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14141e),
	.w1(32'hba20e25f),
	.w2(32'hbab667f9),
	.w3(32'h3b483418),
	.w4(32'h3aad7f85),
	.w5(32'h3b34a382),
	.w6(32'h3bb0371d),
	.w7(32'h3b3a99e0),
	.w8(32'h3b6040c9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb885ed7),
	.w1(32'h3b47d769),
	.w2(32'hbb992e86),
	.w3(32'hbbcfeac3),
	.w4(32'hb9f9711c),
	.w5(32'h3accedce),
	.w6(32'hbbb02bd3),
	.w7(32'hbbb71be4),
	.w8(32'h3a92a307),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94a386),
	.w1(32'h3ac235ac),
	.w2(32'hbbbee6ac),
	.w3(32'hbc316fa2),
	.w4(32'h3c383506),
	.w5(32'h3d036c57),
	.w6(32'hbad0d4ff),
	.w7(32'h3a71ed29),
	.w8(32'h3c053466),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed113b),
	.w1(32'hbb37fcfa),
	.w2(32'hbb0354a4),
	.w3(32'h3a3ca9ac),
	.w4(32'hbb8500be),
	.w5(32'hba463a12),
	.w6(32'hba18bdb1),
	.w7(32'hbabada9b),
	.w8(32'hba898d94),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec428d),
	.w1(32'hbae6d4fc),
	.w2(32'hbaea3a74),
	.w3(32'hbafc2b63),
	.w4(32'hba3b3fe2),
	.w5(32'hb674bb4f),
	.w6(32'h38b29d5e),
	.w7(32'hbb582985),
	.w8(32'h3b6e9c22),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae22d23),
	.w1(32'h3b9f7ae0),
	.w2(32'h3bb26c91),
	.w3(32'hba8c6dfb),
	.w4(32'h3c01ab8f),
	.w5(32'h3c0793e0),
	.w6(32'hbaa867e5),
	.w7(32'h3a5b0d5f),
	.w8(32'hb9d3ea0b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966e55d),
	.w1(32'h3baf83b0),
	.w2(32'hbad1a971),
	.w3(32'hbb0e29dc),
	.w4(32'h3b7162e4),
	.w5(32'hbb88fd39),
	.w6(32'hba9e3c7a),
	.w7(32'h3ae8b048),
	.w8(32'hbb4c5140),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaca3a),
	.w1(32'h3a70d5ca),
	.w2(32'h3a61b860),
	.w3(32'hbbcc4076),
	.w4(32'hbbc34305),
	.w5(32'hbb708831),
	.w6(32'hbbd868b3),
	.w7(32'hbb7e5704),
	.w8(32'hbb688eaa),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf49cc),
	.w1(32'hbb24b411),
	.w2(32'hbb9381e5),
	.w3(32'hbad6b301),
	.w4(32'hbb1caf9a),
	.w5(32'hbb9dea3b),
	.w6(32'hbbc7c2da),
	.w7(32'hba999665),
	.w8(32'hbc0d5ff1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2272a3),
	.w1(32'h3b879f1f),
	.w2(32'h3af64ad7),
	.w3(32'hbb96659b),
	.w4(32'hbc10cc14),
	.w5(32'h3c4292b6),
	.w6(32'hbb54eedd),
	.w7(32'hbc235d2e),
	.w8(32'hba9da918),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c9508),
	.w1(32'hba832bfd),
	.w2(32'hbb9245fd),
	.w3(32'h3c05fa20),
	.w4(32'h3afcf772),
	.w5(32'h3984dacb),
	.w6(32'hbb18c8c3),
	.w7(32'h39c0c363),
	.w8(32'hbb40b9c2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf26e24),
	.w1(32'h3b7bb425),
	.w2(32'h3a8b4914),
	.w3(32'h3c708cc8),
	.w4(32'hbb0f6954),
	.w5(32'hbc122bdc),
	.w6(32'h3c255117),
	.w7(32'h3a9ee91e),
	.w8(32'hbb3ef36d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c44daf),
	.w1(32'h3bc3ed9a),
	.w2(32'h3a521618),
	.w3(32'hbb69cb59),
	.w4(32'h3aa6cf98),
	.w5(32'hba6ec8f0),
	.w6(32'hbb626830),
	.w7(32'h3a077bf9),
	.w8(32'hbadcec0d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b6944),
	.w1(32'hba03d156),
	.w2(32'hb9944804),
	.w3(32'h3922bc54),
	.w4(32'hba50a9d7),
	.w5(32'h39c1c145),
	.w6(32'h3ac8bb77),
	.w7(32'h3b37e851),
	.w8(32'h3a87efef),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab86aae),
	.w1(32'h3b918a79),
	.w2(32'h3bd4b559),
	.w3(32'hbaddaa51),
	.w4(32'hba111146),
	.w5(32'h3bc68d8f),
	.w6(32'h39973616),
	.w7(32'h3b72037e),
	.w8(32'h3bc7ad91),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba111db),
	.w1(32'hbb4e170d),
	.w2(32'hbb863bc7),
	.w3(32'h3af5004b),
	.w4(32'hbaf3b519),
	.w5(32'h3b9b6062),
	.w6(32'h3a1c5953),
	.w7(32'hbbf0ded2),
	.w8(32'hbbc395ec),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18f04f),
	.w1(32'h3ae9e1f4),
	.w2(32'hbacedea0),
	.w3(32'hba999b10),
	.w4(32'hbb3aa051),
	.w5(32'h398b8002),
	.w6(32'hbafc8872),
	.w7(32'hbb8be6f6),
	.w8(32'hbb74a0a0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25fbc),
	.w1(32'h3b1bd1f9),
	.w2(32'hbbc76e5a),
	.w3(32'hbb7b35de),
	.w4(32'hba8a2bb4),
	.w5(32'h3c957919),
	.w6(32'hbbfaecd9),
	.w7(32'hbbb50735),
	.w8(32'hbbe905ab),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbcf1a),
	.w1(32'hbc0f6506),
	.w2(32'hbb73474e),
	.w3(32'hba4c778b),
	.w4(32'hbc4ed47c),
	.w5(32'hb8b14343),
	.w6(32'hbc5c8e1a),
	.w7(32'hbbb1dce0),
	.w8(32'h3aa1e18d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b3223),
	.w1(32'h3a4f63fd),
	.w2(32'hba21e7df),
	.w3(32'hba45b2c9),
	.w4(32'h3ac5aeda),
	.w5(32'hbb455622),
	.w6(32'h3b8ad1ab),
	.w7(32'h3b37c904),
	.w8(32'h3afdbc55),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8f7b5),
	.w1(32'h3940b787),
	.w2(32'hbaa72f80),
	.w3(32'hbb4f380a),
	.w4(32'hb98034bc),
	.w5(32'hbbbc9455),
	.w6(32'hbb9ce528),
	.w7(32'hba1b83a5),
	.w8(32'hbaaad4a4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae7065),
	.w1(32'hbb51583d),
	.w2(32'hbad7fc4a),
	.w3(32'h3b2a7223),
	.w4(32'hbb91d4cc),
	.w5(32'hb99e9be2),
	.w6(32'hba50ac61),
	.w7(32'hbae0c515),
	.w8(32'hbb68828b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63ea3b),
	.w1(32'h3a7fa4b6),
	.w2(32'hba0bb662),
	.w3(32'hbb7610ed),
	.w4(32'h3b73d4bd),
	.w5(32'h3aa3b848),
	.w6(32'h394c539f),
	.w7(32'h3b2b4ab0),
	.w8(32'h3acf6483),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa45cf3),
	.w1(32'hbb2ef8e9),
	.w2(32'hbb8f4ef5),
	.w3(32'hbb673789),
	.w4(32'hbaff8952),
	.w5(32'hbb1aa9c8),
	.w6(32'hbb2f7a82),
	.w7(32'hbb304fe1),
	.w8(32'hbb046e86),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2054f4),
	.w1(32'hbb83eef3),
	.w2(32'hbb172b01),
	.w3(32'hbaa60080),
	.w4(32'hb9aad161),
	.w5(32'hbaceae0c),
	.w6(32'hbb144084),
	.w7(32'h3b1752e5),
	.w8(32'h3adbfe9c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5453e2),
	.w1(32'hba6da3e6),
	.w2(32'hb96a0a84),
	.w3(32'hbb86a2c0),
	.w4(32'hbb0a99db),
	.w5(32'hb8285daa),
	.w6(32'hbadfbea3),
	.w7(32'hbbe132d9),
	.w8(32'hbac7d2fc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb602ff8),
	.w1(32'h3a475bb6),
	.w2(32'h3ab242c4),
	.w3(32'hbb60f3c5),
	.w4(32'h3b05d4fb),
	.w5(32'h3a1521bc),
	.w6(32'h39fa1eff),
	.w7(32'h387b706d),
	.w8(32'h3ad2a86c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b236954),
	.w1(32'hbb0dc595),
	.w2(32'hbb2a46e2),
	.w3(32'h3b000fb9),
	.w4(32'hbb6bf5d2),
	.w5(32'hbb8cc9a2),
	.w6(32'h3a194a08),
	.w7(32'hbab4faa7),
	.w8(32'h3afa1262),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306292),
	.w1(32'h3ab83567),
	.w2(32'h3afe2e53),
	.w3(32'h3adf4ebe),
	.w4(32'h3af282fb),
	.w5(32'hba1f72fe),
	.w6(32'h38a231c5),
	.w7(32'hba212048),
	.w8(32'hba87850e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b698d94),
	.w1(32'hbb117dc7),
	.w2(32'hbb9cde45),
	.w3(32'h3b11d517),
	.w4(32'hbafbf979),
	.w5(32'h3b69a121),
	.w6(32'h3b0b3cfa),
	.w7(32'hbad74340),
	.w8(32'hbbb08111),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab192e3),
	.w1(32'h3b203350),
	.w2(32'h3c1a1318),
	.w3(32'h38a761e3),
	.w4(32'h3a8e1df4),
	.w5(32'hba888315),
	.w6(32'hbae4c0ba),
	.w7(32'hbb5c2003),
	.w8(32'hb9a49a9f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56aad8),
	.w1(32'hbc1ffa25),
	.w2(32'hbbde27c6),
	.w3(32'hbc456af6),
	.w4(32'hbc6c3e8b),
	.w5(32'h3aa3b562),
	.w6(32'hbc6a5841),
	.w7(32'hbbe231fe),
	.w8(32'hbb33fda9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb864d72),
	.w1(32'h3babf387),
	.w2(32'h3ad09d79),
	.w3(32'h3bb3789e),
	.w4(32'h3bb3269e),
	.w5(32'hbb397955),
	.w6(32'h3ac8f198),
	.w7(32'h3bd19f7f),
	.w8(32'h3a6e6f0e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af149bb),
	.w1(32'hbb033ec6),
	.w2(32'hbb96787e),
	.w3(32'hb93824a8),
	.w4(32'h3b566c01),
	.w5(32'h3b993040),
	.w6(32'h3a7b5d02),
	.w7(32'hbb19b7c9),
	.w8(32'hba625ad4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbd7ad),
	.w1(32'h3b099ab1),
	.w2(32'hbb717e0e),
	.w3(32'h399cffc8),
	.w4(32'h3b678248),
	.w5(32'h3b426404),
	.w6(32'hbb887d65),
	.w7(32'h3b1816ef),
	.w8(32'h3ac91651),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb2fe1),
	.w1(32'h3bc6d1ee),
	.w2(32'h3bc42b39),
	.w3(32'hbba49c21),
	.w4(32'h3a372def),
	.w5(32'h3b46eb86),
	.w6(32'hbb3c66fe),
	.w7(32'hbbb47c87),
	.w8(32'hbb78c39e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba83456),
	.w1(32'h3ad92fd5),
	.w2(32'hbaca03b5),
	.w3(32'h3ba075ca),
	.w4(32'h3b475e92),
	.w5(32'h3b5e710e),
	.w6(32'h3a5501ac),
	.w7(32'hb9d294c5),
	.w8(32'hb8fe2297),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57f38a),
	.w1(32'hbb63321d),
	.w2(32'hbb75a1ff),
	.w3(32'h3bbfbc64),
	.w4(32'h3a724adc),
	.w5(32'hbbd34a93),
	.w6(32'h3b49acc4),
	.w7(32'h3a01e13c),
	.w8(32'hbb2081c1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f2db2),
	.w1(32'hbb15f814),
	.w2(32'hbacbada9),
	.w3(32'h3a81dcb5),
	.w4(32'hb9f90558),
	.w5(32'hb9d2c920),
	.w6(32'h3b9a8806),
	.w7(32'hbac20087),
	.w8(32'hbb24bd03),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc7d47),
	.w1(32'h3b89d501),
	.w2(32'hba80754c),
	.w3(32'hbab800b8),
	.w4(32'hbaa3eed1),
	.w5(32'h39f5b38b),
	.w6(32'hbb520243),
	.w7(32'hba4a8b41),
	.w8(32'hbb89958b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb871457),
	.w1(32'hbbb05e1a),
	.w2(32'h3ab0a2a7),
	.w3(32'h3b7a18cc),
	.w4(32'hbb7c8681),
	.w5(32'hbb6120df),
	.w6(32'h3c1d721e),
	.w7(32'hbb343aba),
	.w8(32'hbba07e47),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10055e),
	.w1(32'hbc62ee93),
	.w2(32'hbc46965c),
	.w3(32'hbc950fae),
	.w4(32'hbc69c8e4),
	.w5(32'hbaa32d0a),
	.w6(32'hbc295f88),
	.w7(32'hbc362ef2),
	.w8(32'hbb2e4127),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc577dc9),
	.w1(32'h3b2a719a),
	.w2(32'h3a8afbf5),
	.w3(32'h3a436380),
	.w4(32'h3c013c32),
	.w5(32'h3c7d2776),
	.w6(32'h3abe9ee9),
	.w7(32'hbb157949),
	.w8(32'hbac4517d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2b6e7),
	.w1(32'h3a79e222),
	.w2(32'hba02128c),
	.w3(32'h3bfc16ab),
	.w4(32'h3a55b4cf),
	.w5(32'hbbbc4269),
	.w6(32'hbb089a38),
	.w7(32'hba8f1317),
	.w8(32'hbadab4f8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41084b),
	.w1(32'hbb85933e),
	.w2(32'hbb5d6c9e),
	.w3(32'h3ad04001),
	.w4(32'hba71cb21),
	.w5(32'hba960a1d),
	.w6(32'hba2d5e34),
	.w7(32'hbb089820),
	.w8(32'hbb87c83f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2bc40),
	.w1(32'hbb8afa5b),
	.w2(32'hbb709461),
	.w3(32'hbb848801),
	.w4(32'hba7e5f4c),
	.w5(32'hbb28670d),
	.w6(32'hbb5b5226),
	.w7(32'h39f1954c),
	.w8(32'h3a017808),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb347cbf),
	.w1(32'hbc87ef38),
	.w2(32'hbc46384e),
	.w3(32'hbc42f76a),
	.w4(32'hbc473314),
	.w5(32'hba9ac3bd),
	.w6(32'hbc3de51d),
	.w7(32'hbc0c3505),
	.w8(32'hbc03424c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dcee3),
	.w1(32'hba16a8b6),
	.w2(32'hba37d957),
	.w3(32'h3b89a35a),
	.w4(32'hba99d154),
	.w5(32'hba9c50da),
	.w6(32'h3b4f1b68),
	.w7(32'h3b3f0e82),
	.w8(32'h3b3a5465),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d3014),
	.w1(32'hbb7fe6c4),
	.w2(32'hbb9769dd),
	.w3(32'h3a12f87f),
	.w4(32'h3a07a2e6),
	.w5(32'hb7d0dc3a),
	.w6(32'h3a6cefbe),
	.w7(32'h3aa6c209),
	.w8(32'h3a72e5d9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74c88f),
	.w1(32'h3a71d2d9),
	.w2(32'h3b0e21a4),
	.w3(32'h39917338),
	.w4(32'hba19cd9f),
	.w5(32'hbb5c3ab4),
	.w6(32'h3b296812),
	.w7(32'hba8104ed),
	.w8(32'h393e3d2d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7954dc),
	.w1(32'h3b95f751),
	.w2(32'h3a80a369),
	.w3(32'h38842f3c),
	.w4(32'h3ade7a88),
	.w5(32'h3c15ce90),
	.w6(32'hbb63e8bd),
	.w7(32'h3ac0670c),
	.w8(32'h39af659e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0d471),
	.w1(32'hbac2f356),
	.w2(32'hbb64657b),
	.w3(32'h3bb93be7),
	.w4(32'h3bb7f062),
	.w5(32'h3c0920e7),
	.w6(32'h3b36ad99),
	.w7(32'hba52c978),
	.w8(32'hbac7a697),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0869b5),
	.w1(32'hbafabbab),
	.w2(32'hbb9c8d1e),
	.w3(32'h3be1513e),
	.w4(32'hbbb6fcc9),
	.w5(32'hbbbb40ba),
	.w6(32'h3ba24fca),
	.w7(32'h3a651445),
	.w8(32'h3a4067be),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10d644),
	.w1(32'hb835941e),
	.w2(32'hb980d82b),
	.w3(32'hbafb21fd),
	.w4(32'hbb76ab64),
	.w5(32'hb9b8bf35),
	.w6(32'hbb9e7043),
	.w7(32'hbb88238d),
	.w8(32'hbbba37aa),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1c37a),
	.w1(32'h3a5f15d6),
	.w2(32'h3b4a6789),
	.w3(32'hba6fd198),
	.w4(32'hbba95bab),
	.w5(32'h39375632),
	.w6(32'hbb13b2f0),
	.w7(32'hbb9769b6),
	.w8(32'hbafd9f90),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7e3b2),
	.w1(32'hbbfce9f2),
	.w2(32'hbc4a5253),
	.w3(32'hbc03759a),
	.w4(32'h3c12589a),
	.w5(32'h3c66eb24),
	.w6(32'hbbbeeb86),
	.w7(32'hbb897acc),
	.w8(32'hbc036471),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19cac1),
	.w1(32'h3b22f6d3),
	.w2(32'hbb163ea3),
	.w3(32'h3bef78de),
	.w4(32'h3ae5447b),
	.w5(32'h3a4baf8d),
	.w6(32'h3b024fba),
	.w7(32'h3a574992),
	.w8(32'h3ae8c09e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f36bf),
	.w1(32'hbb6683be),
	.w2(32'hbb164b9d),
	.w3(32'hba8df9eb),
	.w4(32'hbbcbe799),
	.w5(32'hbbb46ba5),
	.w6(32'h3aa13cd9),
	.w7(32'hbb9523a3),
	.w8(32'hbb143f8b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4af841),
	.w1(32'hbac65c65),
	.w2(32'hbba94738),
	.w3(32'hbb9510ba),
	.w4(32'hba867584),
	.w5(32'h3b6245fa),
	.w6(32'hbbafafa4),
	.w7(32'hba35acdc),
	.w8(32'hbb140880),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd16e8c),
	.w1(32'h3bd53d96),
	.w2(32'h3bb4bdc8),
	.w3(32'hbaf30b8e),
	.w4(32'hbacd2327),
	.w5(32'hbac29555),
	.w6(32'hbb00c0bb),
	.w7(32'hbb24e1bb),
	.w8(32'hbb83594a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f23b),
	.w1(32'h3a0839f4),
	.w2(32'hb982ef62),
	.w3(32'hb9a6113d),
	.w4(32'h3ae497a9),
	.w5(32'h3b7b3f3d),
	.w6(32'hba2239a6),
	.w7(32'h3a7fb559),
	.w8(32'hb9d9f5c0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9690e39),
	.w1(32'h3c17b2d3),
	.w2(32'h3b4902d0),
	.w3(32'h39b449d4),
	.w4(32'hbb8d5d1a),
	.w5(32'hbbbe282a),
	.w6(32'hba74f8cb),
	.w7(32'hbb7a45dd),
	.w8(32'hbbfc3e6e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb140c91),
	.w1(32'hb9ff0d64),
	.w2(32'h3b866651),
	.w3(32'hbb27e81f),
	.w4(32'h3ac26843),
	.w5(32'h3ad22476),
	.w6(32'hbb95c684),
	.w7(32'h399b0fbf),
	.w8(32'h3b7385de),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adde40b),
	.w1(32'hb9fab6bc),
	.w2(32'hbb1a9af5),
	.w3(32'hb9c14a1b),
	.w4(32'h3bbd9cc2),
	.w5(32'h3b864423),
	.w6(32'h392ac5b1),
	.w7(32'h3b314c56),
	.w8(32'hba8ccd7f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cc921),
	.w1(32'h3afe503a),
	.w2(32'h3a4392e1),
	.w3(32'h3c1c0bfb),
	.w4(32'hba1a80e8),
	.w5(32'hbbad8a05),
	.w6(32'h3ae1cf4f),
	.w7(32'h3a1fe975),
	.w8(32'hbb2db97a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4461a),
	.w1(32'h3b0d3f10),
	.w2(32'h3a8e4d6a),
	.w3(32'hbb42515c),
	.w4(32'h3b5f93b9),
	.w5(32'h3bbe6285),
	.w6(32'hbb285f2b),
	.w7(32'hba54f391),
	.w8(32'h3afc1269),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37d062),
	.w1(32'h3bdbdbfc),
	.w2(32'hb9cf6b26),
	.w3(32'h3baee5f9),
	.w4(32'h3b343818),
	.w5(32'h3c381fdd),
	.w6(32'h3b181adf),
	.w7(32'hb998865a),
	.w8(32'hbb19c926),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7be23a),
	.w1(32'hb9f8289a),
	.w2(32'hbbb4f0db),
	.w3(32'h3bb8274a),
	.w4(32'hbb1dde2f),
	.w5(32'h3a62baa1),
	.w6(32'hba581bc9),
	.w7(32'hbb862731),
	.w8(32'hbb47c823),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40fc8d),
	.w1(32'h3b7bcdc8),
	.w2(32'h3b06188f),
	.w3(32'h3a781d39),
	.w4(32'h3a11c7a9),
	.w5(32'hbae4b7dd),
	.w6(32'hbae35356),
	.w7(32'h3b2d22ee),
	.w8(32'h3b94947e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc6ff1),
	.w1(32'h3bc5c21f),
	.w2(32'h3be2574e),
	.w3(32'hb8da9352),
	.w4(32'h3981fc50),
	.w5(32'hbb6191e4),
	.w6(32'h39fa5833),
	.w7(32'hbb836be7),
	.w8(32'hbb351f96),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32c5de),
	.w1(32'hbad7e54d),
	.w2(32'hbb16bc47),
	.w3(32'hbba88e66),
	.w4(32'hbae0a785),
	.w5(32'h38a231a8),
	.w6(32'hbbe28278),
	.w7(32'hba9ff03d),
	.w8(32'hba588b4f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fefaa3),
	.w1(32'hbb65f1a9),
	.w2(32'hb9af3097),
	.w3(32'hb973d344),
	.w4(32'h3a9d0110),
	.w5(32'hbb3035e3),
	.w6(32'hbabc0e3e),
	.w7(32'h3b4c9292),
	.w8(32'h38648a09),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8681c0),
	.w1(32'h3bbd5440),
	.w2(32'hbb5733bb),
	.w3(32'h3ac9eca8),
	.w4(32'h3b9cd9f7),
	.w5(32'h3ceeffdc),
	.w6(32'h3aa1964f),
	.w7(32'hbc3ebdb2),
	.w8(32'hbc139d84),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d3375),
	.w1(32'h39e416c0),
	.w2(32'h37d74eef),
	.w3(32'h3c2e9f75),
	.w4(32'hb9077bdd),
	.w5(32'hbb88dbbd),
	.w6(32'h3a639911),
	.w7(32'h3aadca3b),
	.w8(32'hba86a858),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34893a),
	.w1(32'hbb343ceb),
	.w2(32'hbb199c85),
	.w3(32'hbb22d74c),
	.w4(32'h3970e208),
	.w5(32'h3ad2b20a),
	.w6(32'hbb52573b),
	.w7(32'hb78e24ee),
	.w8(32'h3ac239b7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb696009),
	.w1(32'hba5ec591),
	.w2(32'h3ad277e5),
	.w3(32'h3b15ae07),
	.w4(32'h39c2f279),
	.w5(32'h3b3948c1),
	.w6(32'h3b87d89d),
	.w7(32'hba3c5877),
	.w8(32'h3b4b8071),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5e4ec),
	.w1(32'hbb2e4cd7),
	.w2(32'hbb8b5072),
	.w3(32'hbc1972df),
	.w4(32'hbb0d84fc),
	.w5(32'h3b6fb60a),
	.w6(32'hbc15e49c),
	.w7(32'hbbed7308),
	.w8(32'hbc1c2808),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22ab06),
	.w1(32'h3be8b3c6),
	.w2(32'h3c0a9575),
	.w3(32'h3a938032),
	.w4(32'h3a9e6fb0),
	.w5(32'hbb2b5bdd),
	.w6(32'hbb0b03da),
	.w7(32'hbb91c84e),
	.w8(32'hbb9c4c05),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9568d9),
	.w1(32'hbb49a08f),
	.w2(32'hbae2906e),
	.w3(32'hbb2bee7d),
	.w4(32'hbb95bea9),
	.w5(32'hbc33da6c),
	.w6(32'hbbaec6f8),
	.w7(32'hbc18656a),
	.w8(32'hbc19fe0d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5923d7),
	.w1(32'hbc1b1c08),
	.w2(32'hbc438b5b),
	.w3(32'hbba8263b),
	.w4(32'hbb9bd08d),
	.w5(32'hb966d5a3),
	.w6(32'hbc0b9413),
	.w7(32'hbb81370c),
	.w8(32'hbb3e9c89),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb340da),
	.w1(32'h3b942c6c),
	.w2(32'h3bcd88c3),
	.w3(32'hbb73936d),
	.w4(32'hbb025d7a),
	.w5(32'h3b0b43da),
	.w6(32'h382bca01),
	.w7(32'hbacbf497),
	.w8(32'hba70fa13),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18d46a),
	.w1(32'h3b7b3758),
	.w2(32'h3adea58e),
	.w3(32'hb8894946),
	.w4(32'h39afa598),
	.w5(32'h3b689895),
	.w6(32'hba4d08ba),
	.w7(32'hba958f6f),
	.w8(32'h3a921382),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5d7e5),
	.w1(32'hba98aa4b),
	.w2(32'hb9af558c),
	.w3(32'h3b053cfe),
	.w4(32'hba3dcaca),
	.w5(32'hbb809880),
	.w6(32'h3b86aa72),
	.w7(32'h3938db77),
	.w8(32'h3b7520a8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87c048),
	.w1(32'h3a1bbd5b),
	.w2(32'h3aa756ed),
	.w3(32'h3a156983),
	.w4(32'h39f4603f),
	.w5(32'hbb80c2ee),
	.w6(32'h3bb9fb48),
	.w7(32'h3ba1951a),
	.w8(32'h3a63face),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e2279),
	.w1(32'h3b81f0bf),
	.w2(32'h3a1dcc8c),
	.w3(32'hbb6d6a10),
	.w4(32'hbb57e37f),
	.w5(32'h3a8e5d26),
	.w6(32'hb9ef41e7),
	.w7(32'hbb267dff),
	.w8(32'hbbaca8f4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4dd6a),
	.w1(32'hba702c49),
	.w2(32'hbae288d5),
	.w3(32'h3b32664b),
	.w4(32'hbb4a3098),
	.w5(32'hbb22fdfe),
	.w6(32'hbb013de3),
	.w7(32'hba8307ce),
	.w8(32'hbab6713b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a403f18),
	.w1(32'h3a8ab0bc),
	.w2(32'h39845917),
	.w3(32'h3aeb4e3a),
	.w4(32'hb9b119c0),
	.w5(32'h3ae7bed2),
	.w6(32'h3966bd1c),
	.w7(32'hbb4c3478),
	.w8(32'hba5d8162),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0661),
	.w1(32'h3b184d91),
	.w2(32'h38c2132c),
	.w3(32'hba9264bf),
	.w4(32'hbb54081e),
	.w5(32'hbb1ed777),
	.w6(32'hbaabdc9f),
	.w7(32'hb9d2ecaf),
	.w8(32'hbb1f52c6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83195e),
	.w1(32'h39dcef38),
	.w2(32'hbb7cf0a7),
	.w3(32'h3b4d6a6f),
	.w4(32'h398da91d),
	.w5(32'hbb15d2a2),
	.w6(32'h3afaa814),
	.w7(32'hbaa9f43d),
	.w8(32'hbb232d3b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59044b),
	.w1(32'hba70a305),
	.w2(32'h3ac69f99),
	.w3(32'hb9d6209b),
	.w4(32'h39198f79),
	.w5(32'h3aa2c97f),
	.w6(32'h3a6dfc17),
	.w7(32'hbae15270),
	.w8(32'h3b2e8f18),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb360e05),
	.w1(32'hbb7cf902),
	.w2(32'hbbbe2514),
	.w3(32'hba9acc5e),
	.w4(32'h3a9a03a7),
	.w5(32'hba415b78),
	.w6(32'h3a4b5b83),
	.w7(32'h38fa542c),
	.w8(32'h3bb8ad4f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6f5f0),
	.w1(32'h3b51c188),
	.w2(32'h3a2930e4),
	.w3(32'hba5ef7dd),
	.w4(32'h3ac80c89),
	.w5(32'hbb94e7f9),
	.w6(32'h3b7d8353),
	.w7(32'h3b621754),
	.w8(32'hba317fc2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8342d0),
	.w1(32'h3a1c0883),
	.w2(32'hbb9e8462),
	.w3(32'h3af1dc0d),
	.w4(32'h3a4326f1),
	.w5(32'hbae770c5),
	.w6(32'h3a80a99f),
	.w7(32'hbb170cd4),
	.w8(32'hbb6622bf),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f35d2),
	.w1(32'hbc14f111),
	.w2(32'hbc2c7de2),
	.w3(32'hbc029e25),
	.w4(32'h39cba868),
	.w5(32'hba3a6cd5),
	.w6(32'hbb8deed8),
	.w7(32'h3b113085),
	.w8(32'h3aeeb9f1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b01ec),
	.w1(32'h3bf94297),
	.w2(32'hb8af74a8),
	.w3(32'h3bb91bd4),
	.w4(32'h3c0ac161),
	.w5(32'hbb28c7bb),
	.w6(32'h3c29cef0),
	.w7(32'h3c0efa5d),
	.w8(32'h3a40e5a0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc764db),
	.w1(32'hbbaf1d2b),
	.w2(32'hbbde921c),
	.w3(32'h3b22cc2c),
	.w4(32'h3acc8afe),
	.w5(32'h3aa67b26),
	.w6(32'h3bd0e01e),
	.w7(32'h3ac8d1cd),
	.w8(32'h3b5d13ec),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf792a8),
	.w1(32'hba944388),
	.w2(32'h3b4d3c7d),
	.w3(32'hba00a50d),
	.w4(32'h3b3f6122),
	.w5(32'h3ba596d9),
	.w6(32'h393c9cb9),
	.w7(32'h3b63a0eb),
	.w8(32'h3b6c8e15),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15cdb0),
	.w1(32'h3bb20c12),
	.w2(32'h3b002eee),
	.w3(32'hba95c640),
	.w4(32'h3b6cd2af),
	.w5(32'hbae086e5),
	.w6(32'hbb345520),
	.w7(32'h3b370bb3),
	.w8(32'hbaf85532),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dc2b7),
	.w1(32'hbae423d0),
	.w2(32'h3b3c65ae),
	.w3(32'h3a0fae66),
	.w4(32'h3b7a3bb8),
	.w5(32'h3a84ec46),
	.w6(32'hb96f7bcb),
	.w7(32'hbaa82939),
	.w8(32'hb9125ba9),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb77229),
	.w1(32'h3bb88666),
	.w2(32'h3b4b6be2),
	.w3(32'h39cb8d9b),
	.w4(32'h3b58937a),
	.w5(32'h3ae6a254),
	.w6(32'h3adc046c),
	.w7(32'h3a3b76a2),
	.w8(32'h3b228828),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1738d6),
	.w1(32'hba32bf79),
	.w2(32'hbb623801),
	.w3(32'h3a257107),
	.w4(32'hb9ee49c3),
	.w5(32'h3a8bbf64),
	.w6(32'h3a06d09e),
	.w7(32'h3b1c3f3e),
	.w8(32'h3bd925c2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae00ba6),
	.w1(32'h3c022d31),
	.w2(32'h3b4b8c5b),
	.w3(32'h3aa09c02),
	.w4(32'h3b44bb7b),
	.w5(32'h3ba3ad6f),
	.w6(32'h3b9e8afb),
	.w7(32'hbaf72216),
	.w8(32'hbb2fa2b9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb053792),
	.w1(32'h3acaa63f),
	.w2(32'h3a8440fb),
	.w3(32'h3a299a8a),
	.w4(32'h399a7157),
	.w5(32'h3c0027b7),
	.w6(32'hbb6fdb86),
	.w7(32'hbbbac9c8),
	.w8(32'hbbc71b9a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e660e),
	.w1(32'hbb4b8313),
	.w2(32'hbadd9925),
	.w3(32'h3b54243a),
	.w4(32'h3a942247),
	.w5(32'h3b0a75f8),
	.w6(32'hba4d9271),
	.w7(32'hbaa35968),
	.w8(32'hbb0687ab),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb117ec3),
	.w1(32'hbbeda064),
	.w2(32'hbb9fb47a),
	.w3(32'hba723488),
	.w4(32'hbb4dd849),
	.w5(32'hbbede0fd),
	.w6(32'hbac58869),
	.w7(32'h3bda36a0),
	.w8(32'h3bbee081),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6c348),
	.w1(32'h3b164255),
	.w2(32'h3b088105),
	.w3(32'hbb989067),
	.w4(32'h3b151805),
	.w5(32'h39b6a409),
	.w6(32'h3a909d1c),
	.w7(32'h3a9ecb68),
	.w8(32'h39e16186),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c319410),
	.w1(32'hb81c4c8e),
	.w2(32'hbac2e73f),
	.w3(32'h3c166b90),
	.w4(32'h3b2f5d37),
	.w5(32'hba842fab),
	.w6(32'h3ba7d89c),
	.w7(32'hb97cddb7),
	.w8(32'hbb8b6fa8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ddcee),
	.w1(32'h3b82359a),
	.w2(32'h3bc11bf9),
	.w3(32'hbab843d5),
	.w4(32'h3a84ac97),
	.w5(32'h392ab89c),
	.w6(32'hbb3685e8),
	.w7(32'h3a766491),
	.w8(32'hba15aaa9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c12f8),
	.w1(32'hbb87d9df),
	.w2(32'hbb6ca19d),
	.w3(32'h3b695e47),
	.w4(32'hba930bd8),
	.w5(32'hba8ff6a9),
	.w6(32'h39a8f0de),
	.w7(32'hbaee7770),
	.w8(32'h38964e49),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb381fd1),
	.w1(32'hba6f7615),
	.w2(32'hbad53129),
	.w3(32'h3b92b7ac),
	.w4(32'hb8a21803),
	.w5(32'hbba42141),
	.w6(32'h3b028ef0),
	.w7(32'h3b0fbbbb),
	.w8(32'h3ae3e21e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b3535),
	.w1(32'h3a3aabbe),
	.w2(32'h3c0833ca),
	.w3(32'hbc0b44d2),
	.w4(32'hbc74a9aa),
	.w5(32'hbc42197a),
	.w6(32'hbc3effc8),
	.w7(32'hbc664fac),
	.w8(32'hbc3af112),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e53e4),
	.w1(32'h3b71e6a9),
	.w2(32'h3b16ffaa),
	.w3(32'hbb85ada2),
	.w4(32'h3a15c8d0),
	.w5(32'hbbb12e91),
	.w6(32'hbbd4876d),
	.w7(32'hb9c1a4c7),
	.w8(32'hbb87bcfa),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8acfcb),
	.w1(32'h38a8f4e3),
	.w2(32'hbb4e138c),
	.w3(32'h38fe02d9),
	.w4(32'hba01680a),
	.w5(32'hbbc085a4),
	.w6(32'hbac0d0df),
	.w7(32'h3ab66a7a),
	.w8(32'hbb6583e3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42b6d2),
	.w1(32'hbb066646),
	.w2(32'hbaa87d42),
	.w3(32'hba82e5b5),
	.w4(32'hb9aff94c),
	.w5(32'hbb2c0c94),
	.w6(32'h38eb5727),
	.w7(32'h3a5ae238),
	.w8(32'h3b335bcb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb579d83),
	.w1(32'h3a857b74),
	.w2(32'hbac34a94),
	.w3(32'hbb2ff300),
	.w4(32'h3a27a708),
	.w5(32'hba840285),
	.w6(32'hbae48eb0),
	.w7(32'hba2f0f2c),
	.w8(32'hbb45909f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b188cf8),
	.w1(32'hbb503fcf),
	.w2(32'hbb8013f8),
	.w3(32'hba1f7e1b),
	.w4(32'hbb0f9d16),
	.w5(32'hbac56347),
	.w6(32'hbb5662db),
	.w7(32'hbb1607db),
	.w8(32'hbad89479),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae83eb),
	.w1(32'hb73cacfd),
	.w2(32'hbb915ea1),
	.w3(32'hbb684d3a),
	.w4(32'hbaf6ec18),
	.w5(32'h3b12d0f8),
	.w6(32'hbbaaa667),
	.w7(32'hbb49f826),
	.w8(32'hb7c9e28f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46348b),
	.w1(32'h3b0fe83a),
	.w2(32'h3b972ce7),
	.w3(32'hbaf1c126),
	.w4(32'h37d6b7bc),
	.w5(32'hbb2c5043),
	.w6(32'h3ac7047c),
	.w7(32'hb9a2590c),
	.w8(32'hbb03b0f9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0b0e),
	.w1(32'hba21bb51),
	.w2(32'hbb80fd19),
	.w3(32'hb9d5985f),
	.w4(32'hba96a193),
	.w5(32'hbb2c315e),
	.w6(32'hbb5519aa),
	.w7(32'h3a5edf92),
	.w8(32'h3a4eff75),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d3ae3),
	.w1(32'h3b9a4a8b),
	.w2(32'h3a7316af),
	.w3(32'h39a20bfe),
	.w4(32'h3b375ea3),
	.w5(32'h3a8c0e4e),
	.w6(32'h3b4c3050),
	.w7(32'hbacf7b7e),
	.w8(32'hba5882a5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d120d3),
	.w1(32'hbbac243d),
	.w2(32'hb8b7b34e),
	.w3(32'h3a685930),
	.w4(32'hbb6254e7),
	.w5(32'hbbc59095),
	.w6(32'hb8f85292),
	.w7(32'h39be3007),
	.w8(32'hb8ab912d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb317f37),
	.w1(32'h3ac6785d),
	.w2(32'h3b6fc738),
	.w3(32'hbbace285),
	.w4(32'hb87a5f6c),
	.w5(32'h39f92aad),
	.w6(32'hba9bdc7f),
	.w7(32'hbb09cb19),
	.w8(32'hbb918fd6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a1346),
	.w1(32'hbaace4f1),
	.w2(32'hbb617a59),
	.w3(32'h399e432e),
	.w4(32'hba6fa8b0),
	.w5(32'hbb915a03),
	.w6(32'h3a9b1d56),
	.w7(32'hba4ae107),
	.w8(32'hbaea9484),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf0781),
	.w1(32'hbbd834bb),
	.w2(32'hbbfc5656),
	.w3(32'hbb754443),
	.w4(32'hbb68df57),
	.w5(32'hbc13adc4),
	.w6(32'hba999505),
	.w7(32'hba4b5a04),
	.w8(32'hba9b64fa),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7614d),
	.w1(32'h3b283a44),
	.w2(32'h3b1728e3),
	.w3(32'hbb6f47d2),
	.w4(32'hbb66fb79),
	.w5(32'hbac057a5),
	.w6(32'hbaa2fa1e),
	.w7(32'hbaab1d43),
	.w8(32'h3b12d6e5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdcdca),
	.w1(32'hba7aed95),
	.w2(32'hbace557b),
	.w3(32'h3b9c4840),
	.w4(32'hb9dde222),
	.w5(32'hbb4692ad),
	.w6(32'h3b019a4c),
	.w7(32'hbb7a20d3),
	.w8(32'hbb982deb),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24eb51),
	.w1(32'hbbf20f2a),
	.w2(32'hbba00f7d),
	.w3(32'h3b8d7c1a),
	.w4(32'hba693b64),
	.w5(32'h3a9fac2f),
	.w6(32'h3b35fccf),
	.w7(32'hbb37a8b4),
	.w8(32'hbb5248e0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc80226),
	.w1(32'hbb90ed85),
	.w2(32'hba43eb4f),
	.w3(32'hbafab799),
	.w4(32'hbb26bb2a),
	.w5(32'h3b23642d),
	.w6(32'hbbbbcb73),
	.w7(32'hbb91f75c),
	.w8(32'hba859d73),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08c4c1),
	.w1(32'hbb973d37),
	.w2(32'hbb744357),
	.w3(32'hbbab62e7),
	.w4(32'hbad83a1d),
	.w5(32'hbb68dbe1),
	.w6(32'hbadf29a5),
	.w7(32'hbb042f5e),
	.w8(32'hbb00d8d8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2419f8),
	.w1(32'hbb6b34e3),
	.w2(32'hbbd0f0af),
	.w3(32'hbc3169be),
	.w4(32'hbbe6257a),
	.w5(32'hbbe34968),
	.w6(32'hbc2b4718),
	.w7(32'h3ac9a5dd),
	.w8(32'hbb187f56),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20bc82),
	.w1(32'h3ac7ce3a),
	.w2(32'hb9badb3a),
	.w3(32'h3c1a6888),
	.w4(32'h3a7c3f1f),
	.w5(32'hbb9bdd1e),
	.w6(32'h3bb904a2),
	.w7(32'hb8f7ce28),
	.w8(32'hbaf363de),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb052902),
	.w1(32'h3b103751),
	.w2(32'h3b88eca7),
	.w3(32'hbb7cf54e),
	.w4(32'hba693829),
	.w5(32'h3b7a4875),
	.w6(32'hbb5934c3),
	.w7(32'hbb252f1d),
	.w8(32'hbb5a94e2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab76672),
	.w1(32'hbb019a6c),
	.w2(32'hbb00c099),
	.w3(32'h39cedf82),
	.w4(32'hbb99328d),
	.w5(32'hbc02ff2d),
	.w6(32'hbb77a08f),
	.w7(32'h3a55f6aa),
	.w8(32'hbb069bcf),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88151d),
	.w1(32'hbb938f7c),
	.w2(32'hbb62e61f),
	.w3(32'hbbc0236d),
	.w4(32'hbb9f69d9),
	.w5(32'hba2a0d8b),
	.w6(32'h3a93bad0),
	.w7(32'hbac67340),
	.w8(32'h3885d027),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74644d),
	.w1(32'h39620dc0),
	.w2(32'h38c6699d),
	.w3(32'hb88d6900),
	.w4(32'h3b30bf73),
	.w5(32'h3b6165a5),
	.w6(32'hb9cb622b),
	.w7(32'hba03c766),
	.w8(32'hb995cf94),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b134fce),
	.w1(32'h3aeb2bcb),
	.w2(32'hbac98351),
	.w3(32'h3b0287db),
	.w4(32'h3b81231a),
	.w5(32'h3b2b0b6a),
	.w6(32'hbb209ac3),
	.w7(32'h3aa056a4),
	.w8(32'hb974949c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b55b7),
	.w1(32'hbb979cd3),
	.w2(32'hbb08061b),
	.w3(32'h3b74b032),
	.w4(32'hbba5ac3b),
	.w5(32'hba079f00),
	.w6(32'h3ab3a248),
	.w7(32'hbb8b636d),
	.w8(32'hbadf5fc0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50c418),
	.w1(32'hbadc7b1c),
	.w2(32'h3aeb2ac4),
	.w3(32'h3a1f22b4),
	.w4(32'hbb8a1b98),
	.w5(32'hbbab9a00),
	.w6(32'hbb0ba80f),
	.w7(32'hbb14c98b),
	.w8(32'hbb8f0e9b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cd1f2),
	.w1(32'hbb7630dd),
	.w2(32'h3aafcaee),
	.w3(32'hbb7f01c8),
	.w4(32'hbbaf31ed),
	.w5(32'hbb05722a),
	.w6(32'h37f58a90),
	.w7(32'hbb9729bb),
	.w8(32'h3a3f77ab),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7b2a1),
	.w1(32'hbb4a32af),
	.w2(32'hbc115b69),
	.w3(32'hba9e4228),
	.w4(32'hba3f9aa9),
	.w5(32'h3b93c868),
	.w6(32'h3acd312e),
	.w7(32'hbb35cfb6),
	.w8(32'h3af850cb),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07c2e1),
	.w1(32'h3ad4934b),
	.w2(32'hbb5db24d),
	.w3(32'hbbfb3649),
	.w4(32'hbba2f158),
	.w5(32'h3bfc7224),
	.w6(32'hbc3a93c1),
	.w7(32'hbbdfcff2),
	.w8(32'hbb986cb7),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5715fe),
	.w1(32'hbc3f356d),
	.w2(32'h3aa6d898),
	.w3(32'hbb1fad7a),
	.w4(32'h3b4eb3e7),
	.w5(32'h3d0356ec),
	.w6(32'hbb68cd34),
	.w7(32'h39821585),
	.w8(32'hbbd09b8f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb4cda),
	.w1(32'hbbc60127),
	.w2(32'hbb4cf784),
	.w3(32'hbb5872b4),
	.w4(32'hbb484bd1),
	.w5(32'hbb03d175),
	.w6(32'hbc80e8ad),
	.w7(32'hbbbb0254),
	.w8(32'hbb479647),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32f057),
	.w1(32'h3b5affad),
	.w2(32'h3b80b5d4),
	.w3(32'hbb67978a),
	.w4(32'h3b83f225),
	.w5(32'h3c1227e5),
	.w6(32'hb9ab6d59),
	.w7(32'h3ba56ba8),
	.w8(32'h3b66e107),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00caf1),
	.w1(32'hbb0a0033),
	.w2(32'h3ae4fa74),
	.w3(32'hba939fd5),
	.w4(32'hbb3e465d),
	.w5(32'hbb728b59),
	.w6(32'h3ace050a),
	.w7(32'hbb965284),
	.w8(32'hb9f245d7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc975ee),
	.w1(32'hbb05533e),
	.w2(32'hbb3d3e9d),
	.w3(32'hbace3070),
	.w4(32'hbb22a50f),
	.w5(32'h3b559207),
	.w6(32'h39a75ddb),
	.w7(32'h3b1146f7),
	.w8(32'h3af9a2cb),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb795476),
	.w1(32'h3bfcc181),
	.w2(32'h3cb23a86),
	.w3(32'h3b8b6adb),
	.w4(32'h3ca120de),
	.w5(32'h3c705026),
	.w6(32'h3b272f51),
	.w7(32'h3bc2bc02),
	.w8(32'hba1994c9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c340764),
	.w1(32'hba02985a),
	.w2(32'hbba063d7),
	.w3(32'hbb237d64),
	.w4(32'hbb948acf),
	.w5(32'hbc4db13e),
	.w6(32'hbb03ec63),
	.w7(32'h3b3f4f60),
	.w8(32'hbbf43d71),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd7e99),
	.w1(32'h3b4011e1),
	.w2(32'hbbce3f31),
	.w3(32'h3a8c38fd),
	.w4(32'h3b4b983b),
	.w5(32'hbbfcd416),
	.w6(32'hbb079e10),
	.w7(32'h3ba955b2),
	.w8(32'h3b476ba3),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922e8bc),
	.w1(32'h3c3eca06),
	.w2(32'h3c858768),
	.w3(32'hba7a6132),
	.w4(32'hbaa94f27),
	.w5(32'h3c18a242),
	.w6(32'h3a25064e),
	.w7(32'h3b9a2044),
	.w8(32'h3c289a3c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8deeba),
	.w1(32'h3bfc571a),
	.w2(32'h3b3bacc2),
	.w3(32'hbbb39cd3),
	.w4(32'h3a893d40),
	.w5(32'hbc8fd189),
	.w6(32'hbc18d28d),
	.w7(32'h39f2434d),
	.w8(32'h3ba61548),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07839),
	.w1(32'h3b1a1bf2),
	.w2(32'h3bc4c0cc),
	.w3(32'h3b968cfe),
	.w4(32'hbb032404),
	.w5(32'hbbedfc14),
	.w6(32'h3bc01107),
	.w7(32'h3a11fafb),
	.w8(32'hb9f138cc),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a510e94),
	.w1(32'h3a875465),
	.w2(32'hbb25a808),
	.w3(32'hbbb63991),
	.w4(32'hbb8fdbc9),
	.w5(32'hbba25c4b),
	.w6(32'h3bab0c98),
	.w7(32'h3b16cfd2),
	.w8(32'hb88a6e64),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73b24e),
	.w1(32'hbbb41ff9),
	.w2(32'h3a861f0f),
	.w3(32'h3b669211),
	.w4(32'hbc072030),
	.w5(32'h3b22031d),
	.w6(32'hba06e659),
	.w7(32'hbbd747df),
	.w8(32'hbb89afdf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d1b77),
	.w1(32'hbbfd78f0),
	.w2(32'hbb8b8e9d),
	.w3(32'hbc1ccabb),
	.w4(32'hb9b1dc74),
	.w5(32'hbbf4e325),
	.w6(32'hbb9749ea),
	.w7(32'hbc1c77fa),
	.w8(32'hbc35f69f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b48ed),
	.w1(32'hbc3a9048),
	.w2(32'hbc6b8609),
	.w3(32'hbc0683a5),
	.w4(32'hbc8d2e42),
	.w5(32'hbbb85719),
	.w6(32'hbbef124b),
	.w7(32'hbb8aa712),
	.w8(32'h3b76e534),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb93df2),
	.w1(32'h3bd0238d),
	.w2(32'hbb0084c2),
	.w3(32'h3b885ba7),
	.w4(32'h39f3add6),
	.w5(32'hbba2a94d),
	.w6(32'h3c02b7c7),
	.w7(32'hbb549250),
	.w8(32'hbc0b13d0),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efb7c4),
	.w1(32'h3a3cde6a),
	.w2(32'h3a94a475),
	.w3(32'hbb9ea15b),
	.w4(32'hbb126cef),
	.w5(32'hbc22f3af),
	.w6(32'hbc28ff33),
	.w7(32'hba8f7424),
	.w8(32'hbadac2b7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f0c93d),
	.w1(32'hbb28a8bc),
	.w2(32'h3be6dbd8),
	.w3(32'hbc189d46),
	.w4(32'h3b7a4968),
	.w5(32'h3b0f25f5),
	.w6(32'h3c27ff89),
	.w7(32'hbb2c94a9),
	.w8(32'h3a8700d2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56859d),
	.w1(32'h38d2e16b),
	.w2(32'h3a998aa1),
	.w3(32'hbb314597),
	.w4(32'h3b605b03),
	.w5(32'hbbeafe55),
	.w6(32'hbbcfaae9),
	.w7(32'hba27425d),
	.w8(32'hbb06e4bd),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe58fa0),
	.w1(32'hbb9485e0),
	.w2(32'h39fa74ca),
	.w3(32'hbb687820),
	.w4(32'hbbc561f2),
	.w5(32'hb9bdaf7d),
	.w6(32'hba9ca132),
	.w7(32'hbc1b6580),
	.w8(32'hbb0aea3d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4c098),
	.w1(32'hbbd45e04),
	.w2(32'hbbee86d5),
	.w3(32'hbb99f77d),
	.w4(32'hbaf3f52e),
	.w5(32'hba570e5b),
	.w6(32'hbc50bcee),
	.w7(32'hbc4a2ea3),
	.w8(32'hbbd49f59),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30185f),
	.w1(32'hbb1429de),
	.w2(32'hbb63a6e5),
	.w3(32'hba84613b),
	.w4(32'hbb2a56ef),
	.w5(32'hbc087783),
	.w6(32'h3b84fe61),
	.w7(32'h3b2f223e),
	.w8(32'h3bb5ef78),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab650a0),
	.w1(32'hbb7b8ecd),
	.w2(32'hbc03d4b2),
	.w3(32'h3c33e1de),
	.w4(32'hbb6212d2),
	.w5(32'hbc2a12bd),
	.w6(32'h3b963266),
	.w7(32'hba9b74ae),
	.w8(32'h3b6e4c38),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a66df),
	.w1(32'h3bba8e96),
	.w2(32'hbadfaa57),
	.w3(32'h3b81258c),
	.w4(32'hba830af5),
	.w5(32'hbb6c3e2d),
	.w6(32'h3c6f45f9),
	.w7(32'hbbe70a03),
	.w8(32'hbc37391a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50c10a),
	.w1(32'hb95ccc8b),
	.w2(32'hbbcc2fa5),
	.w3(32'hbba62067),
	.w4(32'hbb6f50cb),
	.w5(32'h3cb668ac),
	.w6(32'hbbc7f454),
	.w7(32'hbafc43fd),
	.w8(32'hb9bb5035),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a8203),
	.w1(32'h3ada2e7d),
	.w2(32'hba83195c),
	.w3(32'h3bb61653),
	.w4(32'hbaa863ef),
	.w5(32'hbbe4c3e3),
	.w6(32'h3b320abe),
	.w7(32'hbc093539),
	.w8(32'hbbf1d9d9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac2225),
	.w1(32'hbbf93b3a),
	.w2(32'h3bfa3168),
	.w3(32'hbc3c59b9),
	.w4(32'hbace6189),
	.w5(32'h3be68dd2),
	.w6(32'h3b31f18a),
	.w7(32'h3aa738ac),
	.w8(32'h3b9ac2b1),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fb738),
	.w1(32'h3ad045ae),
	.w2(32'hbb02f839),
	.w3(32'h3c061895),
	.w4(32'h3b30298a),
	.w5(32'hbb45ecd3),
	.w6(32'h3adb60e1),
	.w7(32'hbb5a8384),
	.w8(32'hbc2fa859),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6a0f8),
	.w1(32'hbb5896b2),
	.w2(32'hbafb60bc),
	.w3(32'hba8c59a7),
	.w4(32'h3b8a30d1),
	.w5(32'h3c22e970),
	.w6(32'hbc3b15ff),
	.w7(32'hbbb4f5a6),
	.w8(32'hbc490219),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb455f38),
	.w1(32'h3bdb89cd),
	.w2(32'hbb924be6),
	.w3(32'h3c818300),
	.w4(32'hbb165c82),
	.w5(32'hbbc4c820),
	.w6(32'hbc5fc657),
	.w7(32'hbc03847c),
	.w8(32'hbbe06cd7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcdf7b),
	.w1(32'hbab1911f),
	.w2(32'hbb9f3da4),
	.w3(32'hbb350e70),
	.w4(32'hbaf7f606),
	.w5(32'hbc3ed3e9),
	.w6(32'h3ac3f878),
	.w7(32'h39594b53),
	.w8(32'hbb30f3db),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07c8c0),
	.w1(32'hbbb8ef6a),
	.w2(32'hbc1fb4fa),
	.w3(32'hbc2c5429),
	.w4(32'hbb17f769),
	.w5(32'h3bade19e),
	.w6(32'hbb3abeae),
	.w7(32'hb9bde44b),
	.w8(32'h3b304aca),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba201bbd),
	.w1(32'hbada5b77),
	.w2(32'hbb94709c),
	.w3(32'h3bcf0827),
	.w4(32'hba61d10e),
	.w5(32'hbc41ae95),
	.w6(32'hbb9725a1),
	.w7(32'hba7fcc28),
	.w8(32'hbbd1c7c4),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4133b9),
	.w1(32'h39db4bf2),
	.w2(32'h3b720917),
	.w3(32'hbba6292e),
	.w4(32'hba3e7d1c),
	.w5(32'hb9631b2d),
	.w6(32'hbb23d7b6),
	.w7(32'h3bb87434),
	.w8(32'hbaf5f58d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab21e31),
	.w1(32'hbc063c2e),
	.w2(32'hbb93b91a),
	.w3(32'h3a42b266),
	.w4(32'hbc00f6b5),
	.w5(32'hbbf664c4),
	.w6(32'hbaecf655),
	.w7(32'hbb97cb43),
	.w8(32'hb95a7c89),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb209e5e),
	.w1(32'h3b003a24),
	.w2(32'hbb77b6ab),
	.w3(32'hbacdd747),
	.w4(32'hbb8ba9b9),
	.w5(32'hbc06a811),
	.w6(32'h3bc02576),
	.w7(32'h3a3ca5a9),
	.w8(32'hbacc1891),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc021de6),
	.w1(32'hbb179170),
	.w2(32'hbbe2945c),
	.w3(32'hbb5adc57),
	.w4(32'hb9894e6d),
	.w5(32'hbc2137de),
	.w6(32'h3b921f0c),
	.w7(32'hbaa4e6d9),
	.w8(32'hb9957239),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ecc47),
	.w1(32'hbb4c85bb),
	.w2(32'hbaa95a6f),
	.w3(32'hba9f3bbf),
	.w4(32'hbb6bd2c6),
	.w5(32'hbb0e1af7),
	.w6(32'h3b22c36c),
	.w7(32'h3b080759),
	.w8(32'h3c31db57),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c9f07),
	.w1(32'h3abae475),
	.w2(32'hbb1ed6dd),
	.w3(32'h3c6cd36f),
	.w4(32'h3b4aba84),
	.w5(32'hbc507aab),
	.w6(32'h3b074e58),
	.w7(32'hba7ca1c3),
	.w8(32'hbc1bd299),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c20c7),
	.w1(32'h3a14ab0f),
	.w2(32'hba3d5918),
	.w3(32'hbb8a8173),
	.w4(32'hbbd4f468),
	.w5(32'hbb98125c),
	.w6(32'h3b4d4523),
	.w7(32'hbae89668),
	.w8(32'hbb189c34),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f8950),
	.w1(32'hbb290c5c),
	.w2(32'hbbcb02f0),
	.w3(32'hbc0e8914),
	.w4(32'hbbbaff9f),
	.w5(32'hbc27632d),
	.w6(32'h3a55b715),
	.w7(32'hbbf864a5),
	.w8(32'hbc3abe13),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6d80f),
	.w1(32'hbc0f016f),
	.w2(32'hbbc677a9),
	.w3(32'hbb262e42),
	.w4(32'hbb420cbb),
	.w5(32'h3a089efc),
	.w6(32'hbbab4264),
	.w7(32'h3af75fef),
	.w8(32'h3bb43900),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a64b1),
	.w1(32'hbb9674bf),
	.w2(32'hbb365417),
	.w3(32'hbaea6a86),
	.w4(32'hb9eed381),
	.w5(32'hbbff3687),
	.w6(32'hbac7308a),
	.w7(32'h3bc47263),
	.w8(32'hbb5c71ca),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1798fe),
	.w1(32'hbbacbebf),
	.w2(32'hbba863c3),
	.w3(32'hbbaf1ba8),
	.w4(32'hbb6daa57),
	.w5(32'h3bd5e2e1),
	.w6(32'hbb0b15dd),
	.w7(32'h3b1df944),
	.w8(32'hba996bc6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce3bc7),
	.w1(32'hbb5a2207),
	.w2(32'hbbfafa75),
	.w3(32'h3b89016d),
	.w4(32'hbbc884fe),
	.w5(32'hbb698cc5),
	.w6(32'h38dd6171),
	.w7(32'hba9473dd),
	.w8(32'h3a947cb5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b518ae6),
	.w1(32'hbb34b9f7),
	.w2(32'hbb09c836),
	.w3(32'hb917fca9),
	.w4(32'h3a482572),
	.w5(32'h3bd5fb0d),
	.w6(32'hba0f71f8),
	.w7(32'h3b68f9bf),
	.w8(32'h3baba351),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87222e),
	.w1(32'h3b8479b5),
	.w2(32'h3b8e74f1),
	.w3(32'h3b377835),
	.w4(32'h3bac5088),
	.w5(32'h3bcd6c44),
	.w6(32'hb90f806f),
	.w7(32'hbabfd59f),
	.w8(32'h3b6f0053),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb903457e),
	.w1(32'h3900593a),
	.w2(32'hbb2996ab),
	.w3(32'h3b5be6e9),
	.w4(32'hbb92211a),
	.w5(32'h3adf2f4e),
	.w6(32'hbadc9f10),
	.w7(32'h3ab030cc),
	.w8(32'h3b09b33d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c7bf0),
	.w1(32'hbbcc4a24),
	.w2(32'hbbbba29c),
	.w3(32'hbb713002),
	.w4(32'hbb91d301),
	.w5(32'h395c2d40),
	.w6(32'h3ba2a13f),
	.w7(32'h399cda8c),
	.w8(32'h3b8a2c2e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae01574),
	.w1(32'h3b20f1e1),
	.w2(32'h3c287ec7),
	.w3(32'hbaeeebed),
	.w4(32'h3c200ce8),
	.w5(32'h3b2cca11),
	.w6(32'hbbcc06cc),
	.w7(32'h3b92b763),
	.w8(32'hbb083f21),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33fe8390),
	.w1(32'hbbf1b0ac),
	.w2(32'hbbdb9999),
	.w3(32'hbc36d662),
	.w4(32'hbb64cbf3),
	.w5(32'hbbd50c8f),
	.w6(32'hba1ba3eb),
	.w7(32'hbb1ddcb8),
	.w8(32'h3ccf04a5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1031c2),
	.w1(32'h3b761c62),
	.w2(32'h3acfdd4d),
	.w3(32'h3ccdf036),
	.w4(32'hbb513f45),
	.w5(32'hbace8ab3),
	.w6(32'hbc0f3631),
	.w7(32'hbb90da1a),
	.w8(32'hbb3d5520),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7927ea),
	.w1(32'hba984c90),
	.w2(32'hbb6eb4a9),
	.w3(32'hbc05226c),
	.w4(32'hbbe8f872),
	.w5(32'hbc35e589),
	.w6(32'h3b893b68),
	.w7(32'hbad7fdc5),
	.w8(32'h3c0c9479),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f0414),
	.w1(32'hbbdc9eac),
	.w2(32'hbbb721d9),
	.w3(32'hbb9c5ac4),
	.w4(32'h3bcef498),
	.w5(32'h3b570d3c),
	.w6(32'h3b31ad0c),
	.w7(32'hbbab81ae),
	.w8(32'hbad7ee3b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995d550),
	.w1(32'hbb08e04a),
	.w2(32'h3bb7195d),
	.w3(32'hbb270112),
	.w4(32'h3c1626dc),
	.w5(32'h3c480502),
	.w6(32'hbc554aac),
	.w7(32'hb9c27afa),
	.w8(32'hbb5ac421),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbda9a3),
	.w1(32'h3ac00348),
	.w2(32'hbb3d1c3d),
	.w3(32'hbab31e71),
	.w4(32'hb9d35a5e),
	.w5(32'h3c7ea357),
	.w6(32'hbb09a82b),
	.w7(32'h39feca1a),
	.w8(32'hbaf0f992),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb59bb5),
	.w1(32'hbc171215),
	.w2(32'hbbaedde1),
	.w3(32'hbab8864b),
	.w4(32'hbbe86ab4),
	.w5(32'hba4a8cd6),
	.w6(32'hbc4695e5),
	.w7(32'hbbaac9bd),
	.w8(32'hbc04069c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule