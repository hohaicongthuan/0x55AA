module layer_8_featuremap_55(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad8ad4),
	.w1(32'hb9820bf1),
	.w2(32'h3a2cb9bd),
	.w3(32'hb90698c7),
	.w4(32'hb9d29735),
	.w5(32'hba0234b0),
	.w6(32'hb8ba3e0a),
	.w7(32'hb85e15a9),
	.w8(32'hb941fb92),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a5eef),
	.w1(32'h3a45b91b),
	.w2(32'h3a51eb06),
	.w3(32'h39d5e00c),
	.w4(32'h3a018aee),
	.w5(32'h3a0c82e9),
	.w6(32'h39c872bb),
	.w7(32'h39d77117),
	.w8(32'hb9c059ae),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9930e8c),
	.w1(32'hb92111d0),
	.w2(32'h391af3d9),
	.w3(32'hb93a81cd),
	.w4(32'hb97472a8),
	.w5(32'h398c2879),
	.w6(32'hb9e27c71),
	.w7(32'hb98fee7d),
	.w8(32'hb9984100),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ed7af),
	.w1(32'hbb40f771),
	.w2(32'hbad9ce32),
	.w3(32'hb9e9a2bb),
	.w4(32'hb9d8e2c8),
	.w5(32'hba282a45),
	.w6(32'hba857a54),
	.w7(32'hbad2465b),
	.w8(32'h39b41b1c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398046b4),
	.w1(32'h392158c4),
	.w2(32'h3a06ce04),
	.w3(32'hb8104db0),
	.w4(32'hb8a50631),
	.w5(32'hb8d5c55f),
	.w6(32'hb65fec77),
	.w7(32'h392d0c70),
	.w8(32'h3b5e95cd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a962b),
	.w1(32'h3b4e48c8),
	.w2(32'h3b1ad821),
	.w3(32'h3b907b46),
	.w4(32'h3b1f3d2b),
	.w5(32'h3a4cc640),
	.w6(32'h3b842f81),
	.w7(32'h3b4fe4fa),
	.w8(32'h3a767322),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08b5b3),
	.w1(32'h3a33d4a2),
	.w2(32'h3a21bd07),
	.w3(32'h3a26cb2c),
	.w4(32'h3a0ec9b0),
	.w5(32'h398b2201),
	.w6(32'h3a0c40b9),
	.w7(32'h3a652fbe),
	.w8(32'hba0e3f9c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f39a7),
	.w1(32'hb6e0c6f5),
	.w2(32'h3a2ce420),
	.w3(32'hbab99e36),
	.w4(32'hba26d0df),
	.w5(32'hb862112d),
	.w6(32'hba76a140),
	.w7(32'hb9ebe272),
	.w8(32'h39564451),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e27921),
	.w1(32'h392e1f4a),
	.w2(32'h3a41459b),
	.w3(32'hb98dc17a),
	.w4(32'h39918ecf),
	.w5(32'h3a5fad71),
	.w6(32'hb988b59d),
	.w7(32'h3a97ea99),
	.w8(32'h3a6a091d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2803bd),
	.w1(32'hbb8316cf),
	.w2(32'hbb33bb06),
	.w3(32'hbb5be4a6),
	.w4(32'hbb541eb4),
	.w5(32'hbb332e5e),
	.w6(32'hb9e472b0),
	.w7(32'hbb249f56),
	.w8(32'hbb187fa7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00390e),
	.w1(32'hbb254d8c),
	.w2(32'hbaaeadf0),
	.w3(32'hbb02b32c),
	.w4(32'hbb11fd32),
	.w5(32'hbae56870),
	.w6(32'hbb0b3dac),
	.w7(32'hbb15b909),
	.w8(32'hba2e040e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b1c28),
	.w1(32'h3992e6f5),
	.w2(32'h39be0562),
	.w3(32'h388072dc),
	.w4(32'hb84c89a5),
	.w5(32'hba2cf2d3),
	.w6(32'h3a19af74),
	.w7(32'h39808294),
	.w8(32'hba0b003b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39839128),
	.w1(32'h3a488642),
	.w2(32'h3a99f22b),
	.w3(32'hb972ae8a),
	.w4(32'hb9b151f6),
	.w5(32'h39046aab),
	.w6(32'h39906209),
	.w7(32'h3a09f545),
	.w8(32'h3ba541ea),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b785374),
	.w1(32'h3b263018),
	.w2(32'h3b041ec4),
	.w3(32'h3b61ac7b),
	.w4(32'h3b10e3e5),
	.w5(32'h3a418b6f),
	.w6(32'h3b3c226c),
	.w7(32'h3b291060),
	.w8(32'h3ae08360),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01036d),
	.w1(32'h3acb02c0),
	.w2(32'h3a94c310),
	.w3(32'h3aeaf830),
	.w4(32'h3ab5f58e),
	.w5(32'h39da7d90),
	.w6(32'h3ac150e4),
	.w7(32'h3a9eec94),
	.w8(32'hba0c13f6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13c8b0),
	.w1(32'hb9cb95c0),
	.w2(32'hb89ab31b),
	.w3(32'hb95ffceb),
	.w4(32'hb98eb4b6),
	.w5(32'hb690bfc3),
	.w6(32'hb9ad092f),
	.w7(32'hb933a57c),
	.w8(32'h3a44c3cf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad04926),
	.w1(32'hbb386070),
	.w2(32'hbb368163),
	.w3(32'hba57354c),
	.w4(32'hb9d39934),
	.w5(32'h38aaf2d0),
	.w6(32'hb9f92ad2),
	.w7(32'hb9ad0fef),
	.w8(32'hba861599),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba282bfe),
	.w1(32'hba207f5c),
	.w2(32'hb8bd76b3),
	.w3(32'hba326fc7),
	.w4(32'hba911e05),
	.w5(32'hba52a08f),
	.w6(32'hb99d8bc4),
	.w7(32'hba3bccf2),
	.w8(32'hbafaaee9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d4e18),
	.w1(32'hbb811114),
	.w2(32'hb972d482),
	.w3(32'hbb88916e),
	.w4(32'hbb567a7b),
	.w5(32'hbb5050c8),
	.w6(32'hbb9f56c4),
	.w7(32'hbb839a82),
	.w8(32'h3af3e770),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec26a0),
	.w1(32'h3ac2db47),
	.w2(32'hbaddc9c6),
	.w3(32'h39dbb200),
	.w4(32'hbb017ff2),
	.w5(32'hba768d10),
	.w6(32'h3a4d2b8c),
	.w7(32'hba6c23fe),
	.w8(32'hbae26896),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a398824),
	.w1(32'h37f0940c),
	.w2(32'hb90b95d3),
	.w3(32'h3a4dd216),
	.w4(32'hb91d2476),
	.w5(32'hb8eec611),
	.w6(32'hb987030c),
	.w7(32'h3877c8a4),
	.w8(32'h39e35bf7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a085e3b),
	.w1(32'h3a4cf82a),
	.w2(32'h3a71232f),
	.w3(32'h39064022),
	.w4(32'h38b7903b),
	.w5(32'h35ae18c9),
	.w6(32'h39b16a10),
	.w7(32'h3a12c3ce),
	.w8(32'h3a9344db),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e1083),
	.w1(32'hbb86196a),
	.w2(32'hba2943ce),
	.w3(32'hbae87861),
	.w4(32'hbb5b6628),
	.w5(32'hbabe99e5),
	.w6(32'hbb09277d),
	.w7(32'hbb105d12),
	.w8(32'hbad87927),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7316b1),
	.w1(32'hba509340),
	.w2(32'h39c57a82),
	.w3(32'hbabaa2d2),
	.w4(32'hba99dc36),
	.w5(32'h38e56a5d),
	.w6(32'hba59382b),
	.w7(32'hb9dbd77e),
	.w8(32'h39ceeae0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a89e78),
	.w1(32'h3a5be97f),
	.w2(32'h39c43bd3),
	.w3(32'hb9a8013c),
	.w4(32'hb8174278),
	.w5(32'h3a171422),
	.w6(32'hb94173de),
	.w7(32'hb9aa5e8a),
	.w8(32'h3a65a691),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92cc823),
	.w1(32'hbb07ff94),
	.w2(32'hb8ccfa10),
	.w3(32'h39e401fd),
	.w4(32'hbacc29f4),
	.w5(32'h38f04fdf),
	.w6(32'hba4f5975),
	.w7(32'hba34dca5),
	.w8(32'h3a2e21ce),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb7cc7),
	.w1(32'hbad8f2ed),
	.w2(32'hba53097a),
	.w3(32'hb8fa2cef),
	.w4(32'hba8b9f00),
	.w5(32'hb8816cd8),
	.w6(32'hba102c0b),
	.w7(32'hb93493be),
	.w8(32'h39cd9bd6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67d19f),
	.w1(32'hbb7d1293),
	.w2(32'h38afc7ec),
	.w3(32'hbaf7d9ee),
	.w4(32'hbb82d167),
	.w5(32'hbb5e6c08),
	.w6(32'hbbac72dc),
	.w7(32'hbbdee659),
	.w8(32'hbbc798e5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb281004),
	.w1(32'hbb70edfd),
	.w2(32'hb96d71d1),
	.w3(32'hbae63723),
	.w4(32'hbb6ecada),
	.w5(32'hbaedb52c),
	.w6(32'hb9da866a),
	.w7(32'hba8e25ec),
	.w8(32'hba37f742),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e804cd),
	.w1(32'hb96a29cb),
	.w2(32'hb93264de),
	.w3(32'hb9050fdb),
	.w4(32'hb98c376c),
	.w5(32'hb9a22172),
	.w6(32'hb9401687),
	.w7(32'hb936c536),
	.w8(32'hba472a14),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4c2d4),
	.w1(32'hbb088af7),
	.w2(32'hbb51eb5d),
	.w3(32'hbae1aa1c),
	.w4(32'hba848c16),
	.w5(32'hba3aacbe),
	.w6(32'hbaf69f55),
	.w7(32'hbb339d60),
	.w8(32'h3a744214),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea4a79),
	.w1(32'h3a4d5674),
	.w2(32'h3a746e90),
	.w3(32'h3af2f058),
	.w4(32'h3780bb7d),
	.w5(32'h3a7ae125),
	.w6(32'h39e1fcc3),
	.w7(32'h3a7ea440),
	.w8(32'h3ac82780),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38d933),
	.w1(32'hba489b52),
	.w2(32'hba31f4ec),
	.w3(32'h3a19d7cd),
	.w4(32'h3997e375),
	.w5(32'h38121418),
	.w6(32'h3a6c2783),
	.w7(32'hb9c60cde),
	.w8(32'hba1ebf72),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36769a),
	.w1(32'hba73d489),
	.w2(32'hbb211050),
	.w3(32'hbab25429),
	.w4(32'hbabd3dd2),
	.w5(32'hb983ebf2),
	.w6(32'hba997d52),
	.w7(32'hbb5486c5),
	.w8(32'h3b6a86c6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838d4a),
	.w1(32'h3b25e055),
	.w2(32'h3afeb5cf),
	.w3(32'h3b541acb),
	.w4(32'h3ac1c0b9),
	.w5(32'h39ba8371),
	.w6(32'h3b59f676),
	.w7(32'h3b14469b),
	.w8(32'hb8d37412),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba433502),
	.w1(32'hba378b9c),
	.w2(32'h39e76471),
	.w3(32'hba5fb724),
	.w4(32'hba5de8c4),
	.w5(32'hb9a12887),
	.w6(32'hba7bfcc1),
	.w7(32'hba11c931),
	.w8(32'hbad597c5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba550be5),
	.w1(32'hba8ebbf0),
	.w2(32'hbac1d28f),
	.w3(32'hba79179b),
	.w4(32'hbabf059f),
	.w5(32'hba1274ad),
	.w6(32'hbb066cb4),
	.w7(32'hbadbdf9b),
	.w8(32'hba895e1a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12ccea),
	.w1(32'hb9c4275e),
	.w2(32'hb9bd9da8),
	.w3(32'hba15d37e),
	.w4(32'hba03eddb),
	.w5(32'hba03c822),
	.w6(32'hb9d1e85d),
	.w7(32'hb95cf4f4),
	.w8(32'h3b4a1e72),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6139cb),
	.w1(32'h3b232190),
	.w2(32'h3af171ea),
	.w3(32'h3b3e28fd),
	.w4(32'h3b19a1cd),
	.w5(32'h3a07f610),
	.w6(32'h3b13e4be),
	.w7(32'h3adb3f7d),
	.w8(32'h39b07e34),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a092600),
	.w1(32'h39a0b65c),
	.w2(32'h3910d19e),
	.w3(32'h3a1760d6),
	.w4(32'hb97a09e8),
	.w5(32'h3993cdd7),
	.w6(32'h3716c0e0),
	.w7(32'h3968197e),
	.w8(32'h396d425a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b105029),
	.w1(32'h383439f2),
	.w2(32'h39af7e06),
	.w3(32'h3b132e5c),
	.w4(32'hb9b77f6f),
	.w5(32'hb9a32e23),
	.w6(32'h3b29c7df),
	.w7(32'h3a7e705a),
	.w8(32'h39c10da9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a480b4),
	.w1(32'hb9a961a3),
	.w2(32'hb9b868aa),
	.w3(32'hbabb5ba2),
	.w4(32'hba9139af),
	.w5(32'hba52fb15),
	.w6(32'hbab85423),
	.w7(32'hb99faee9),
	.w8(32'h3ac580ce),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad451c4),
	.w1(32'hbbafe9a3),
	.w2(32'h3a35e783),
	.w3(32'hb9826a16),
	.w4(32'hbba3630e),
	.w5(32'hbae9c523),
	.w6(32'h3b18b8ef),
	.w7(32'h3a51d599),
	.w8(32'hba59cb36),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba014411),
	.w1(32'hba3f3402),
	.w2(32'hb986f3af),
	.w3(32'hb96cbdeb),
	.w4(32'hb96c8bca),
	.w5(32'hba3045fa),
	.w6(32'hba42a9d1),
	.w7(32'hb9a0350f),
	.w8(32'h3a02f737),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9174b),
	.w1(32'hba08d2fb),
	.w2(32'h3aa3a2ab),
	.w3(32'h39b88ba2),
	.w4(32'hb9d6fd7e),
	.w5(32'hb9acce92),
	.w6(32'h39a2be98),
	.w7(32'h3a6d6cb9),
	.w8(32'h39a6fe33),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af658bb),
	.w1(32'h39fffafa),
	.w2(32'h3ae9716f),
	.w3(32'h3a059cfb),
	.w4(32'hba3c1407),
	.w5(32'h397b0a1e),
	.w6(32'h39118ab0),
	.w7(32'h3ab1c659),
	.w8(32'hbbd13cfb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccba51),
	.w1(32'h3bb4558a),
	.w2(32'h3b5d6fd3),
	.w3(32'hbb16ca6d),
	.w4(32'h3ae4e767),
	.w5(32'hbaedf578),
	.w6(32'hbbd7a761),
	.w7(32'hba61330c),
	.w8(32'h3abbe41c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98c0dd),
	.w1(32'hbb2f78a1),
	.w2(32'hbaae1c45),
	.w3(32'hba6fce4d),
	.w4(32'hba22eb29),
	.w5(32'h3a5358fd),
	.w6(32'hba51e0f1),
	.w7(32'hbb24d5c8),
	.w8(32'hba1a84cb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25f994),
	.w1(32'h398168df),
	.w2(32'h3aa51bf1),
	.w3(32'h3a3b3d23),
	.w4(32'h3a04c71d),
	.w5(32'h3ad892b7),
	.w6(32'hb972bf11),
	.w7(32'hba0827a5),
	.w8(32'h3a3096a2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf7ddf),
	.w1(32'hba05c832),
	.w2(32'h3a9d15cb),
	.w3(32'h3a934376),
	.w4(32'h398cf21a),
	.w5(32'h3a044757),
	.w6(32'h3a825200),
	.w7(32'h3b0eb430),
	.w8(32'h3a07ee96),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae8e3c),
	.w1(32'h3b2420e9),
	.w2(32'h3b092818),
	.w3(32'h3a520661),
	.w4(32'h3b066373),
	.w5(32'h3ad5e840),
	.w6(32'h3a9df159),
	.w7(32'h3b244ded),
	.w8(32'h3b07bf96),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d884e),
	.w1(32'hbad1ff1c),
	.w2(32'h39c45681),
	.w3(32'hb9c78d08),
	.w4(32'hb94d9566),
	.w5(32'hb9499d37),
	.w6(32'hbaba89d6),
	.w7(32'hba556b46),
	.w8(32'h3b05c964),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24fe09),
	.w1(32'hbc1930ac),
	.w2(32'hbbc2648f),
	.w3(32'hb9dc8e21),
	.w4(32'hbc1e6539),
	.w5(32'hbb831a68),
	.w6(32'hbb5f452d),
	.w7(32'hbb1174e0),
	.w8(32'hbb0b49a5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8af9b6),
	.w1(32'hbaef56d3),
	.w2(32'h38fb182e),
	.w3(32'hba32ac89),
	.w4(32'hbab73d34),
	.w5(32'hba41a22a),
	.w6(32'hbb0d7562),
	.w7(32'hbaad9fda),
	.w8(32'hba461d5c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2051e0),
	.w1(32'h3adef614),
	.w2(32'hbad74283),
	.w3(32'hbb2a84e5),
	.w4(32'h3b6ceec9),
	.w5(32'h375a11a0),
	.w6(32'h3b93fee1),
	.w7(32'hbaea5a73),
	.w8(32'h3a92181a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b559c92),
	.w1(32'hbaae6706),
	.w2(32'h399c9d08),
	.w3(32'h3b85f668),
	.w4(32'h3b808796),
	.w5(32'h3b07c662),
	.w6(32'hbadba8ce),
	.w7(32'h3b234d7e),
	.w8(32'hbb872583),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb380d3b),
	.w1(32'hbb16eee2),
	.w2(32'hbb00379a),
	.w3(32'hba990627),
	.w4(32'hbb11cdb7),
	.w5(32'hbb4897af),
	.w6(32'hbaf34e30),
	.w7(32'hbaa88a72),
	.w8(32'h3b8b83e3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1f132),
	.w1(32'hbb959c8e),
	.w2(32'hbb9a549c),
	.w3(32'h3ad3e3b2),
	.w4(32'h3a808858),
	.w5(32'hb9e01c87),
	.w6(32'h3af0f070),
	.w7(32'hbb9dad43),
	.w8(32'hb97d2531),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11cde2),
	.w1(32'hb9d7e89b),
	.w2(32'h388790b2),
	.w3(32'hba8f59f4),
	.w4(32'hba2df239),
	.w5(32'hba880524),
	.w6(32'hb9675a00),
	.w7(32'hb8520bd3),
	.w8(32'h3b2e5443),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52d2dc),
	.w1(32'h3b1b712a),
	.w2(32'h3b2e0d99),
	.w3(32'h3b3315b0),
	.w4(32'h3990b91b),
	.w5(32'h3b027401),
	.w6(32'h3b545310),
	.w7(32'h3b438967),
	.w8(32'hba920b6c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc247087),
	.w1(32'hbc04cb67),
	.w2(32'hbb5ac2a0),
	.w3(32'hbb6e48bd),
	.w4(32'hbac1590f),
	.w5(32'hbb7b9120),
	.w6(32'hbbe5ffcd),
	.w7(32'hbac5208d),
	.w8(32'h39cf1c7e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9574eef),
	.w1(32'hbb397e22),
	.w2(32'h392b9009),
	.w3(32'h3af722c9),
	.w4(32'h3b129171),
	.w5(32'h3b571b09),
	.w6(32'hba7bdc83),
	.w7(32'h3ad18330),
	.w8(32'h39f9dab7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f18fe),
	.w1(32'h3acfe87f),
	.w2(32'h3ae86f1f),
	.w3(32'h3acbcce6),
	.w4(32'h3a71c457),
	.w5(32'hb980aefe),
	.w6(32'h3a9a6190),
	.w7(32'h3b2072eb),
	.w8(32'h3a876fbd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d995c),
	.w1(32'hbbcba69d),
	.w2(32'hbb200a14),
	.w3(32'hbb0246e3),
	.w4(32'hbb86d234),
	.w5(32'hbb779fba),
	.w6(32'h3ab57075),
	.w7(32'hba95f7f3),
	.w8(32'hba9958d0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9291778),
	.w1(32'h3868f370),
	.w2(32'h38c375eb),
	.w3(32'hb7dcec36),
	.w4(32'h3851dd58),
	.w5(32'hb9c3f51b),
	.w6(32'h34f869c7),
	.w7(32'h3a5d65e4),
	.w8(32'h389cd2c9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4899b),
	.w1(32'hb9ae8aa0),
	.w2(32'hb936215e),
	.w3(32'hba31820b),
	.w4(32'hba0435ea),
	.w5(32'hb9f2dd0e),
	.w6(32'hb9ed4065),
	.w7(32'hb96b42ba),
	.w8(32'h3735ebad),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a536af1),
	.w1(32'h398e0259),
	.w2(32'h39f02da1),
	.w3(32'h3a7b1cb8),
	.w4(32'h39e20ff2),
	.w5(32'h39eeb24a),
	.w6(32'h3a1945e1),
	.w7(32'h3a757786),
	.w8(32'hbaa81061),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2b643),
	.w1(32'hbaa6e5ab),
	.w2(32'h3a2a435e),
	.w3(32'hbb6b695e),
	.w4(32'hbadce81c),
	.w5(32'hbae37bd8),
	.w6(32'hbb147b3d),
	.w7(32'hbafe8130),
	.w8(32'h3aa2b52c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51378b),
	.w1(32'hb89a2709),
	.w2(32'h3a2a8cbc),
	.w3(32'h3a144c11),
	.w4(32'hb8cfb4af),
	.w5(32'h38e2ff4f),
	.w6(32'h3a02aac0),
	.w7(32'h3ac369b9),
	.w8(32'h39b62d84),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39550c2f),
	.w1(32'hbb09da3a),
	.w2(32'hbb214f36),
	.w3(32'hba68108a),
	.w4(32'hbb308ec2),
	.w5(32'hbb94dc48),
	.w6(32'h3a3587da),
	.w7(32'hba7ce85e),
	.w8(32'hbadaa89c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b6336),
	.w1(32'h382478f6),
	.w2(32'hb991179d),
	.w3(32'hb95ff5de),
	.w4(32'hb9ef3fa0),
	.w5(32'hba47d49d),
	.w6(32'hb9b8bf5e),
	.w7(32'h3974336e),
	.w8(32'h3a40ca57),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d1cc0),
	.w1(32'hb9c46471),
	.w2(32'h3a7ae69c),
	.w3(32'h3a3f1947),
	.w4(32'hb9a3b28e),
	.w5(32'h39cd40b7),
	.w6(32'h3a26588d),
	.w7(32'h3ab24d35),
	.w8(32'hb97c094e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b7eef),
	.w1(32'hb91a456d),
	.w2(32'hb981c1c9),
	.w3(32'hb99190f8),
	.w4(32'hba64fa0c),
	.w5(32'hba8d6b12),
	.w6(32'hb9b450c1),
	.w7(32'h3a104c69),
	.w8(32'h3a03fc49),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b304d71),
	.w1(32'h399a0713),
	.w2(32'hbaea44b7),
	.w3(32'hbbb9b187),
	.w4(32'hbbc02f67),
	.w5(32'hbbd24833),
	.w6(32'hbb1ff9db),
	.w7(32'hbb64627c),
	.w8(32'h3a1e51f9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae864d7),
	.w1(32'h3a971b06),
	.w2(32'h3ad5cc07),
	.w3(32'h3a8f7e9d),
	.w4(32'h3a4ffe39),
	.w5(32'h3a56d6c4),
	.w6(32'h3a991c9b),
	.w7(32'h3ad82537),
	.w8(32'hba10d1cf),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e7729),
	.w1(32'hb9a065c0),
	.w2(32'hb9a08bc9),
	.w3(32'h383cfd6d),
	.w4(32'hb990e868),
	.w5(32'hba2664ef),
	.w6(32'hb95e916c),
	.w7(32'hb88cb4c4),
	.w8(32'hb945f12d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c075b),
	.w1(32'hb9088b88),
	.w2(32'h39452b2a),
	.w3(32'h38b08a52),
	.w4(32'h3960cf40),
	.w5(32'h39b63fcc),
	.w6(32'h392e86fe),
	.w7(32'h3a56e4b8),
	.w8(32'h39c45945),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba633994),
	.w1(32'hba801974),
	.w2(32'hba9ac428),
	.w3(32'hbb3a661e),
	.w4(32'hbb2f4c54),
	.w5(32'hbba2b419),
	.w6(32'h38b9a43d),
	.w7(32'h39c7d7a9),
	.w8(32'hb9cd0f5d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e2d7e),
	.w1(32'h3a02838a),
	.w2(32'hb9e562ec),
	.w3(32'hbaeb52fc),
	.w4(32'hba888cc4),
	.w5(32'hbb268dce),
	.w6(32'hb9bf10d4),
	.w7(32'hb938f6a3),
	.w8(32'hb822ccc4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6a268),
	.w1(32'hb8a56221),
	.w2(32'h399f6172),
	.w3(32'hb9edf24c),
	.w4(32'h3910c03b),
	.w5(32'h39650fcb),
	.w6(32'h3a17433e),
	.w7(32'h3932b836),
	.w8(32'hbadcb6f5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0ef7f),
	.w1(32'hba8cb6eb),
	.w2(32'hbaf0c748),
	.w3(32'hba8733d9),
	.w4(32'h3b38bab8),
	.w5(32'h3a2cbeba),
	.w6(32'hbb216625),
	.w7(32'hbafd5450),
	.w8(32'hb996a75c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa07f35),
	.w1(32'h39fcb5db),
	.w2(32'h3a4d6ad6),
	.w3(32'h3b15f684),
	.w4(32'h3ae08745),
	.w5(32'h3ad0078e),
	.w6(32'h3aaf2147),
	.w7(32'h3ad9043e),
	.w8(32'h3af65467),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0d76d),
	.w1(32'hb8ecced3),
	.w2(32'h3b16db2e),
	.w3(32'h3a41e38f),
	.w4(32'hba34a47e),
	.w5(32'h3a230ec4),
	.w6(32'h3aff5c9c),
	.w7(32'h3b44e71f),
	.w8(32'hbb162b92),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d8a78),
	.w1(32'hbb69ee9b),
	.w2(32'hba65739d),
	.w3(32'hb96d3b57),
	.w4(32'hbaa25e71),
	.w5(32'h3b02b9e5),
	.w6(32'hbb2c48a9),
	.w7(32'h3a9de93c),
	.w8(32'h3a84b2a6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10be4e),
	.w1(32'hbaf9397d),
	.w2(32'h39f9bc47),
	.w3(32'hb8509386),
	.w4(32'hbaf47d39),
	.w5(32'hbab9454a),
	.w6(32'hbab2b2a0),
	.w7(32'hbb026327),
	.w8(32'h39a31e13),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16bd23),
	.w1(32'hb9e71888),
	.w2(32'h3a3df68d),
	.w3(32'h3aa85362),
	.w4(32'h3880cd22),
	.w5(32'h3a140dec),
	.w6(32'h3a08c2cb),
	.w7(32'h3ad4a840),
	.w8(32'hba4ba3fe),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04d680),
	.w1(32'h39a500ba),
	.w2(32'h3ac25e7a),
	.w3(32'h3a5374d1),
	.w4(32'h3a6592e1),
	.w5(32'h3b1adf26),
	.w6(32'hba31b8e8),
	.w7(32'hba32ea36),
	.w8(32'hba3b53ee),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8b7d0),
	.w1(32'hb9d19865),
	.w2(32'hba12217d),
	.w3(32'h374a9e48),
	.w4(32'hb7bdc755),
	.w5(32'hb8e86fd3),
	.w6(32'h3978fb7c),
	.w7(32'h39825578),
	.w8(32'h3b2f899e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30f8ed),
	.w1(32'h3b1bd7b9),
	.w2(32'h3b03460d),
	.w3(32'h3a80f561),
	.w4(32'hb91d5e1e),
	.w5(32'h3b04a6c0),
	.w6(32'h3b4508b0),
	.w7(32'h3b277f26),
	.w8(32'hb9d39e97),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e0182),
	.w1(32'h399b437d),
	.w2(32'h3acfc320),
	.w3(32'h3a275542),
	.w4(32'h3a32c638),
	.w5(32'h3b12e956),
	.w6(32'hba1b32bf),
	.w7(32'hba442e0b),
	.w8(32'hb9ea6bdd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa75bff),
	.w1(32'h3a2db0de),
	.w2(32'h3abd9d7c),
	.w3(32'h3ab7cad2),
	.w4(32'h3a4381d4),
	.w5(32'h3b08c303),
	.w6(32'h39f36e13),
	.w7(32'hb974b188),
	.w8(32'hba19de29),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac3ae8),
	.w1(32'hb9fe98c2),
	.w2(32'h3989aedd),
	.w3(32'hb96389d6),
	.w4(32'hba82ef11),
	.w5(32'hb5138ede),
	.w6(32'hba837fd7),
	.w7(32'h380f0cdc),
	.w8(32'hb8e010ba),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3f0ac),
	.w1(32'hbaabb10e),
	.w2(32'hbba75e76),
	.w3(32'hbb0080f3),
	.w4(32'hbb6ec34d),
	.w5(32'hbbedf9c9),
	.w6(32'h3b8e87e9),
	.w7(32'hbb636f14),
	.w8(32'hb78d7024),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394933d3),
	.w1(32'h392e34e5),
	.w2(32'h39c55ae1),
	.w3(32'hb6bf5c62),
	.w4(32'hb8019d80),
	.w5(32'hb9479688),
	.w6(32'hb95981b2),
	.w7(32'hb90a03d4),
	.w8(32'h3a70c9a9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa14cf),
	.w1(32'hbb889687),
	.w2(32'hbb92387e),
	.w3(32'hbaf8ed27),
	.w4(32'h3aa72f23),
	.w5(32'hba3a4ab9),
	.w6(32'h37451c73),
	.w7(32'h3ae07f71),
	.w8(32'hbaf386aa),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a50fd),
	.w1(32'hba286521),
	.w2(32'hba01ceb7),
	.w3(32'hba4c06ab),
	.w4(32'hbb46c38c),
	.w5(32'hbb03d6d8),
	.w6(32'hbb1546fa),
	.w7(32'hbadab260),
	.w8(32'hbb201aa3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0028e7),
	.w1(32'h3b0ba4fd),
	.w2(32'h39932d7b),
	.w3(32'hb9e34504),
	.w4(32'h3aa71f3c),
	.w5(32'h3b00ba41),
	.w6(32'hba24cb4e),
	.w7(32'hbaa7114f),
	.w8(32'h3a7b5505),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfbb1e),
	.w1(32'hba2a3e76),
	.w2(32'hba675a7f),
	.w3(32'hbb37cff8),
	.w4(32'hbaadeee1),
	.w5(32'hbaf3c76f),
	.w6(32'hbacad9e7),
	.w7(32'h390e862f),
	.w8(32'h39aa4eba),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0590d1),
	.w1(32'hb8f66d25),
	.w2(32'hba84fa46),
	.w3(32'hbb096ac1),
	.w4(32'hbad799be),
	.w5(32'hbb80ae47),
	.w6(32'h3a766f3f),
	.w7(32'h3a945bbc),
	.w8(32'hb9be6ac2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e1508c),
	.w1(32'hb9c94351),
	.w2(32'hb9718ed1),
	.w3(32'hb7b74aab),
	.w4(32'hb9a18b2c),
	.w5(32'hb9566711),
	.w6(32'h395e4efd),
	.w7(32'h3a808285),
	.w8(32'h3acd0d40),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5c9c7),
	.w1(32'h3a633a87),
	.w2(32'h3a8213b1),
	.w3(32'h3aa2f1ca),
	.w4(32'h399db6e4),
	.w5(32'h3a5ab138),
	.w6(32'h3a9ab4a7),
	.w7(32'h3a54342c),
	.w8(32'hb99477f5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7ce63),
	.w1(32'h393fdcc3),
	.w2(32'h39f94af0),
	.w3(32'h39b6c616),
	.w4(32'h39786899),
	.w5(32'hb7a02491),
	.w6(32'hb97b4f50),
	.w7(32'h3a017eb7),
	.w8(32'hb9b4c036),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ac9f2c),
	.w1(32'h3ab02762),
	.w2(32'hbadcc7ac),
	.w3(32'hbac0469f),
	.w4(32'hba303b46),
	.w5(32'hbb71f04d),
	.w6(32'h3a161880),
	.w7(32'h3a05f65c),
	.w8(32'h38c7f251),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9521d),
	.w1(32'h3a70cf1d),
	.w2(32'h3a4d9ce6),
	.w3(32'h39f22c81),
	.w4(32'hba764583),
	.w5(32'h38750306),
	.w6(32'h3a6e15a0),
	.w7(32'h39dc6de8),
	.w8(32'hb9034a71),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1202a7),
	.w1(32'h398916c7),
	.w2(32'h3a3e9ba1),
	.w3(32'h3a0dfaab),
	.w4(32'h3985c594),
	.w5(32'h3a6fb4be),
	.w6(32'h390c90d2),
	.w7(32'hb93867cd),
	.w8(32'h391e02b7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91101c9),
	.w1(32'hba4a0406),
	.w2(32'h39095c3f),
	.w3(32'h392b68be),
	.w4(32'hba0ffd1b),
	.w5(32'hb99cd352),
	.w6(32'hba39502a),
	.w7(32'hbaadf952),
	.w8(32'hba50db95),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9874836),
	.w1(32'hb85c8988),
	.w2(32'h3750e0ee),
	.w3(32'hb959ceb7),
	.w4(32'hb9489c5f),
	.w5(32'hb92436bf),
	.w6(32'hb9d1a4ef),
	.w7(32'hb99cda7e),
	.w8(32'hb99cfc2f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e05b9e),
	.w1(32'hb87eb424),
	.w2(32'h3904cb6d),
	.w3(32'h391658a9),
	.w4(32'hb9bdbca2),
	.w5(32'hb9349b96),
	.w6(32'h39a8e2b9),
	.w7(32'hb8f7fc83),
	.w8(32'hb584d9db),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15ead2),
	.w1(32'h399c5abe),
	.w2(32'h36a87fe9),
	.w3(32'h39f0e0ed),
	.w4(32'h394e8a97),
	.w5(32'hb80b0df2),
	.w6(32'h3a181895),
	.w7(32'h39b21f9b),
	.w8(32'h398b7cce),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89724a5),
	.w1(32'hb85c324e),
	.w2(32'h36137f20),
	.w3(32'hb9b64f1e),
	.w4(32'hb99d5569),
	.w5(32'hb828f85f),
	.w6(32'hb98be0ad),
	.w7(32'hb8820cc8),
	.w8(32'h39369a24),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5576b6),
	.w1(32'h3a046955),
	.w2(32'h3a177e5a),
	.w3(32'hb881a8f8),
	.w4(32'hb99a103a),
	.w5(32'hb9b4ab8f),
	.w6(32'h3a06e2cb),
	.w7(32'h399ff28f),
	.w8(32'h3923c36d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86812b),
	.w1(32'h3a290bdd),
	.w2(32'h3a248747),
	.w3(32'h39cecb3b),
	.w4(32'h38c56d01),
	.w5(32'hb8d2453c),
	.w6(32'h3a799692),
	.w7(32'h3a42eb4c),
	.w8(32'h3a125156),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25c6a0),
	.w1(32'hb7c65ef4),
	.w2(32'h391f5e71),
	.w3(32'h3a0b3cf7),
	.w4(32'hb8a348da),
	.w5(32'hb9120eb6),
	.w6(32'h3a54c77b),
	.w7(32'h399d50ef),
	.w8(32'h39754668),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8600f54),
	.w1(32'hb868aac1),
	.w2(32'hb78b9c9f),
	.w3(32'hb7c959a4),
	.w4(32'hb795d5fe),
	.w5(32'h366f0dc2),
	.w6(32'hb8a07c53),
	.w7(32'hb8703980),
	.w8(32'hb803d235),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912e1b2),
	.w1(32'hb9871dff),
	.w2(32'hb8855a41),
	.w3(32'hb8b7304b),
	.w4(32'hb936922e),
	.w5(32'hb810ad65),
	.w6(32'hb90e8d9e),
	.w7(32'hb9264ef4),
	.w8(32'hb8c0174a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38592845),
	.w1(32'h38d52111),
	.w2(32'h38f1adf1),
	.w3(32'hb6edaf4a),
	.w4(32'hb8977610),
	.w5(32'hb8cf1fbd),
	.w6(32'h3798b596),
	.w7(32'h37929cc8),
	.w8(32'h372c513b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ef066),
	.w1(32'h39462d87),
	.w2(32'h38802582),
	.w3(32'h39ac47a6),
	.w4(32'h37ad5280),
	.w5(32'hb8ba9f54),
	.w6(32'h3a1a4cb8),
	.w7(32'h39896be6),
	.w8(32'h3962e4b3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d20e48),
	.w1(32'hb98f33d2),
	.w2(32'hb8e2f34f),
	.w3(32'h39bbed20),
	.w4(32'hb8e996d5),
	.w5(32'hb9c549ae),
	.w6(32'h39ac8ea9),
	.w7(32'hb7f2623e),
	.w8(32'h38726276),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d2ef14),
	.w1(32'hb70dd555),
	.w2(32'hb6bfe52d),
	.w3(32'hb69d5b9c),
	.w4(32'hb669100a),
	.w5(32'hb481d011),
	.w6(32'hb71c9153),
	.w7(32'hb6c5923e),
	.w8(32'hb6a65cf0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d7dc37),
	.w1(32'h37f2b727),
	.w2(32'h388e9409),
	.w3(32'hb7e574eb),
	.w4(32'h375a5497),
	.w5(32'hb7876847),
	.w6(32'hb7e31ef9),
	.w7(32'hb889b795),
	.w8(32'hb7bcd33e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03602b),
	.w1(32'h39907afe),
	.w2(32'h39731f67),
	.w3(32'h39de9c30),
	.w4(32'hb8e28859),
	.w5(32'hb88e9a5a),
	.w6(32'h3a7a027b),
	.w7(32'h399002dc),
	.w8(32'h3995d9dc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96615b5),
	.w1(32'hb95999ad),
	.w2(32'h35e181ee),
	.w3(32'hb8f996ca),
	.w4(32'hb9503be1),
	.w5(32'hb8e28dd0),
	.w6(32'hb99ea725),
	.w7(32'hb9721cfa),
	.w8(32'hb835c8ae),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379f7c5c),
	.w1(32'hb8853842),
	.w2(32'hb8dc277a),
	.w3(32'hb794f572),
	.w4(32'hb8c00ef7),
	.w5(32'hb9077dab),
	.w6(32'hb8a84b54),
	.w7(32'hb8eb5a18),
	.w8(32'h36b84f4d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2a440),
	.w1(32'h38f28afb),
	.w2(32'hb915c7c5),
	.w3(32'h38e30e05),
	.w4(32'h38e992c8),
	.w5(32'hb8cbf5d6),
	.w6(32'h3943475b),
	.w7(32'h398f4e9a),
	.w8(32'h39544a9d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc7488),
	.w1(32'h39ebca03),
	.w2(32'h396624cc),
	.w3(32'h399ee6cb),
	.w4(32'h39bb14ae),
	.w5(32'h39567ffa),
	.w6(32'h39f9bc05),
	.w7(32'h39cea187),
	.w8(32'h39b39e7d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992bbc3),
	.w1(32'hb3cc5ce0),
	.w2(32'h398e1438),
	.w3(32'hba3c6f1f),
	.w4(32'hb9b8ba24),
	.w5(32'h38fdace6),
	.w6(32'hba2b9f58),
	.w7(32'hb9a4fb2d),
	.w8(32'hb993d229),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384aa569),
	.w1(32'h38b22dd6),
	.w2(32'h39446401),
	.w3(32'hb8f0bcbd),
	.w4(32'hb9631ee7),
	.w5(32'hb8ce16b8),
	.w6(32'h379cc58f),
	.w7(32'hb8c70611),
	.w8(32'h3907e279),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9581444),
	.w1(32'hb94c346d),
	.w2(32'h3977bff1),
	.w3(32'hb9ada8ae),
	.w4(32'hb957c3de),
	.w5(32'h3903d2cd),
	.w6(32'hb9eba23a),
	.w7(32'hb98a4bf6),
	.w8(32'h38285c07),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule