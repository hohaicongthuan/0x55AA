module layer_10_featuremap_356(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4291d7),
	.w1(32'h39ef20ca),
	.w2(32'hba7a39e1),
	.w3(32'h3a51f612),
	.w4(32'hbb41d75d),
	.w5(32'hbb3430a1),
	.w6(32'hbba820a5),
	.w7(32'hbbd4928d),
	.w8(32'hba42a482),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1274a6),
	.w1(32'hba019f74),
	.w2(32'hb9e8af04),
	.w3(32'hbae46689),
	.w4(32'hb99125ef),
	.w5(32'h3a35ce77),
	.w6(32'hb8f27a80),
	.w7(32'h3a9143d7),
	.w8(32'hbac6deee),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c4d99),
	.w1(32'hbba6a03b),
	.w2(32'hbb1472ab),
	.w3(32'h3985332d),
	.w4(32'hb9852921),
	.w5(32'hb9c6d2e5),
	.w6(32'hbaa0094b),
	.w7(32'hbb177ac6),
	.w8(32'h3a46dcc7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc0193),
	.w1(32'hbaa46c80),
	.w2(32'hbae64876),
	.w3(32'hbadaecfc),
	.w4(32'hbace2262),
	.w5(32'hba3659d3),
	.w6(32'hbb413f8f),
	.w7(32'hbaea9f4d),
	.w8(32'hbbaf64ed),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd528e),
	.w1(32'h3b22237a),
	.w2(32'hbb866d2f),
	.w3(32'hbb6d0471),
	.w4(32'hbbb25d94),
	.w5(32'h3b733c5d),
	.w6(32'hbbedbec5),
	.w7(32'hbc454aa9),
	.w8(32'h3b69e4b6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44425a),
	.w1(32'hbb19e8be),
	.w2(32'h3aa1e2db),
	.w3(32'hb8f60caa),
	.w4(32'h3adbdca0),
	.w5(32'h3ae1e6fb),
	.w6(32'hbbd6530b),
	.w7(32'hbae91729),
	.w8(32'h3b9cfa20),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad65b03),
	.w1(32'hbb1f195e),
	.w2(32'hbb9132e3),
	.w3(32'hbb1a7edd),
	.w4(32'hbb8bbf5e),
	.w5(32'h3b428301),
	.w6(32'hbafabd6c),
	.w7(32'hbbd32ba6),
	.w8(32'h3a885b69),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a01a6f),
	.w1(32'hb96a0199),
	.w2(32'h3bb8f6bf),
	.w3(32'h3b7a242e),
	.w4(32'h3a322910),
	.w5(32'h3b654568),
	.w6(32'hba2be0b0),
	.w7(32'h39877b2a),
	.w8(32'h3b47d353),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b403df8),
	.w1(32'h3adc45d2),
	.w2(32'h3929f657),
	.w3(32'h3b8497b2),
	.w4(32'h39b11d68),
	.w5(32'h3b54a152),
	.w6(32'h3aaa64fc),
	.w7(32'hbb06a29f),
	.w8(32'h3b805b8a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b829e9a),
	.w1(32'hbac6c8b2),
	.w2(32'hb9e2cbe6),
	.w3(32'hba8443cc),
	.w4(32'h3b3c6c3b),
	.w5(32'h3b80da3b),
	.w6(32'hbbbd8124),
	.w7(32'hbb0dbba9),
	.w8(32'h3b9d1b25),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fc601),
	.w1(32'hbbac7c05),
	.w2(32'hbb12b22d),
	.w3(32'hbaa78572),
	.w4(32'hbb339a0b),
	.w5(32'h3aefad91),
	.w6(32'hbbb9b839),
	.w7(32'hbbbad8c2),
	.w8(32'h3b791843),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6e682),
	.w1(32'h384c303b),
	.w2(32'h3b52070e),
	.w3(32'h3b117d9b),
	.w4(32'hbb4a74f0),
	.w5(32'h3b5b7ec5),
	.w6(32'hba0d7a45),
	.w7(32'h3a58876d),
	.w8(32'h39da5e2b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900930),
	.w1(32'hb9332d57),
	.w2(32'hba8e9286),
	.w3(32'h3af08d5a),
	.w4(32'hba73e3ac),
	.w5(32'h3a5f917c),
	.w6(32'hbadff11e),
	.w7(32'hba19bd16),
	.w8(32'hba950d47),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a9576),
	.w1(32'h3af93245),
	.w2(32'h3ab2d406),
	.w3(32'h3a8b03df),
	.w4(32'hbb0d36bd),
	.w5(32'hb9fb96c7),
	.w6(32'h3ba0e0af),
	.w7(32'hbb008b30),
	.w8(32'h3a7372ff),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf77de),
	.w1(32'hba096b2b),
	.w2(32'h392665eb),
	.w3(32'h3a0ddaa6),
	.w4(32'hba142975),
	.w5(32'hbb368d38),
	.w6(32'hbab3c15d),
	.w7(32'hbac419b3),
	.w8(32'hbb726549),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba662f1),
	.w1(32'hbbad1af5),
	.w2(32'hbb3c666d),
	.w3(32'hbba8de17),
	.w4(32'hbb2d141b),
	.w5(32'h3a7044c2),
	.w6(32'hbb1ff8b8),
	.w7(32'hbb7401bc),
	.w8(32'h39135e48),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b454ae1),
	.w1(32'h3adeda10),
	.w2(32'h3bbac41b),
	.w3(32'h3a86c750),
	.w4(32'h3b49237e),
	.w5(32'h3b2f5962),
	.w6(32'hbb9dca44),
	.w7(32'h3aaf4ecf),
	.w8(32'h3b70aea8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ecd3a),
	.w1(32'hbabb6534),
	.w2(32'hbb01b953),
	.w3(32'h3a4eea30),
	.w4(32'hbac1d98e),
	.w5(32'h3a661c4a),
	.w6(32'hbac19b5d),
	.w7(32'hbb241573),
	.w8(32'hba33958a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18ab12),
	.w1(32'hbadb6c79),
	.w2(32'hbad6972e),
	.w3(32'h3a9ee0fa),
	.w4(32'h3a58b6bf),
	.w5(32'h3a8eb86c),
	.w6(32'hb9afe068),
	.w7(32'h39ad9cf9),
	.w8(32'hba665978),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88f4ee),
	.w1(32'hbb30ae05),
	.w2(32'hbb3fe065),
	.w3(32'hbb00550d),
	.w4(32'hbb723e55),
	.w5(32'hbb898eb4),
	.w6(32'h3b1165f9),
	.w7(32'hbb570d94),
	.w8(32'hbbbffdbe),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97bd4c),
	.w1(32'hba537ca6),
	.w2(32'hbbb0b2f5),
	.w3(32'hbb8af5f5),
	.w4(32'hbb142ba8),
	.w5(32'hbaa38b06),
	.w6(32'h397daae8),
	.w7(32'hbba0d7fe),
	.w8(32'h36b50a7c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16e7ca),
	.w1(32'h3bb8ed82),
	.w2(32'h3b6236ee),
	.w3(32'h3b408998),
	.w4(32'h3b852ad3),
	.w5(32'hbb213ec2),
	.w6(32'h3b57f9b9),
	.w7(32'h3b682d9b),
	.w8(32'hbb19f251),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f8280),
	.w1(32'hbada8bb0),
	.w2(32'hba8a592b),
	.w3(32'hbb3ff2c7),
	.w4(32'hbb115469),
	.w5(32'hbafe30bf),
	.w6(32'hbb1f96ee),
	.w7(32'hbb14773d),
	.w8(32'h3a6467f7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bd39e),
	.w1(32'hbc0d4efd),
	.w2(32'hbb226ca1),
	.w3(32'hbc11719d),
	.w4(32'hbbae7734),
	.w5(32'hba6a0d78),
	.w6(32'hbc26673b),
	.w7(32'hbbfdfb10),
	.w8(32'hbae25e82),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42e2ca),
	.w1(32'h3a0f691a),
	.w2(32'hbac3b6bb),
	.w3(32'hba93c7a8),
	.w4(32'h3886dd98),
	.w5(32'hbb02053c),
	.w6(32'hbaedd81d),
	.w7(32'hbaba34a4),
	.w8(32'hbb63fcff),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bc97f),
	.w1(32'hbb54bf7c),
	.w2(32'hb9058316),
	.w3(32'h39264fd8),
	.w4(32'hba16ea31),
	.w5(32'hba975031),
	.w6(32'hbb217834),
	.w7(32'hbaf2500b),
	.w8(32'hba2d0184),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9c1a3),
	.w1(32'hba9c1a05),
	.w2(32'h3b233ffc),
	.w3(32'h39768ae3),
	.w4(32'h3afd457e),
	.w5(32'h3bb043b3),
	.w6(32'h3a9377d7),
	.w7(32'h3b5cfc8c),
	.w8(32'h39522a3d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78ec18),
	.w1(32'h3af773c8),
	.w2(32'hb9bf53b0),
	.w3(32'h3b45f451),
	.w4(32'h3b449502),
	.w5(32'hba92e29c),
	.w6(32'hbbc4660e),
	.w7(32'hbb9b85eb),
	.w8(32'h3a83ab50),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af209c8),
	.w1(32'hbb24338f),
	.w2(32'hbacf73b0),
	.w3(32'hbb614df1),
	.w4(32'hbb5465da),
	.w5(32'h3c1266df),
	.w6(32'h3a9faf2b),
	.w7(32'hbaf28be7),
	.w8(32'h3c219cea),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21cf84),
	.w1(32'hbbea529a),
	.w2(32'h3a3931a0),
	.w3(32'hbbf2c5fe),
	.w4(32'hba9921c7),
	.w5(32'h3b0f4e44),
	.w6(32'hbb817057),
	.w7(32'h3aad8398),
	.w8(32'h3a03afc7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae003),
	.w1(32'hba8d296e),
	.w2(32'hbbcfbc0b),
	.w3(32'h3b59a83f),
	.w4(32'hba50081b),
	.w5(32'hbb62aff2),
	.w6(32'h3b09ae7b),
	.w7(32'hb8d8407e),
	.w8(32'hbaeb4063),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace6252),
	.w1(32'h3ab1b1aa),
	.w2(32'h3aba9fee),
	.w3(32'h3a369a65),
	.w4(32'h3a19b1b0),
	.w5(32'hbb302887),
	.w6(32'h3b84196b),
	.w7(32'h3aec4156),
	.w8(32'hba735fda),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0ce82),
	.w1(32'hbb10a05e),
	.w2(32'h3b056430),
	.w3(32'hbb651a52),
	.w4(32'hba8bf9d8),
	.w5(32'h3b233bf9),
	.w6(32'h3a807733),
	.w7(32'h3aecc29d),
	.w8(32'h3bc90a84),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e1284),
	.w1(32'hbb5b98e4),
	.w2(32'hbb8b1ee1),
	.w3(32'hbb482830),
	.w4(32'hbb8a47dc),
	.w5(32'hbadde63d),
	.w6(32'hbbcc29d0),
	.w7(32'hbbdf512d),
	.w8(32'hba489156),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b273940),
	.w1(32'hbb078dd3),
	.w2(32'hbb43e93d),
	.w3(32'hba5734cf),
	.w4(32'h3a3743d3),
	.w5(32'hbab3b41d),
	.w6(32'hb9f001e0),
	.w7(32'hba958a65),
	.w8(32'hbb0d5491),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb730a983),
	.w1(32'hbaff5a9b),
	.w2(32'hbaf98d2f),
	.w3(32'hbbbe302b),
	.w4(32'hbb662d47),
	.w5(32'hbb09b91e),
	.w6(32'hbbdf41ab),
	.w7(32'hbbc866e5),
	.w8(32'hbb4c4868),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae26038),
	.w1(32'hba7da614),
	.w2(32'hbbafcdd7),
	.w3(32'h3a2c9d04),
	.w4(32'h3a2e254d),
	.w5(32'hbab8e6b4),
	.w6(32'h3a3f625e),
	.w7(32'h3aca5cb1),
	.w8(32'h3a900f62),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90b375),
	.w1(32'hba58cfda),
	.w2(32'hbb34b9a1),
	.w3(32'h3b53252c),
	.w4(32'hb90d332c),
	.w5(32'hbb37a1f5),
	.w6(32'h3ba6ed30),
	.w7(32'hbae28000),
	.w8(32'h3b309a91),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87b41),
	.w1(32'h3b8d1a89),
	.w2(32'hbab5b6f7),
	.w3(32'hba725c64),
	.w4(32'h39402b17),
	.w5(32'h3b73cca9),
	.w6(32'hba2f5b44),
	.w7(32'hbb29bec9),
	.w8(32'h3b8265be),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb233b3),
	.w1(32'h3b9cd2af),
	.w2(32'hbb1bebb3),
	.w3(32'h3ba17a4a),
	.w4(32'hb850c265),
	.w5(32'h3bdd99e1),
	.w6(32'h3b7ef4c5),
	.w7(32'hbb90f7ef),
	.w8(32'h3b5a23b0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d255c),
	.w1(32'h3a4e7d9d),
	.w2(32'h3b28a161),
	.w3(32'h39f11ab8),
	.w4(32'h3a8c2130),
	.w5(32'hbba817d9),
	.w6(32'h3972f0ee),
	.w7(32'h3a316639),
	.w8(32'hbbbfe59b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e6cbf),
	.w1(32'hbbab381a),
	.w2(32'hbb07b481),
	.w3(32'hbb769a7f),
	.w4(32'hbac8a7cf),
	.w5(32'hb98a3b46),
	.w6(32'hbc140627),
	.w7(32'hbb93f68f),
	.w8(32'hb99b37e6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7e820),
	.w1(32'hb9a93a12),
	.w2(32'hbb7688c3),
	.w3(32'h3a82cbc5),
	.w4(32'hbade6d18),
	.w5(32'h3a063223),
	.w6(32'h3b7445d2),
	.w7(32'hbad78fdc),
	.w8(32'h3aa09b2d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68092e),
	.w1(32'hbb919795),
	.w2(32'hba588509),
	.w3(32'hb9f00585),
	.w4(32'h3af82d03),
	.w5(32'h3ac0fff1),
	.w6(32'hbb6a490c),
	.w7(32'hbab2eff8),
	.w8(32'h3ab214ed),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980c1d8),
	.w1(32'hbb801658),
	.w2(32'hba5ddbc2),
	.w3(32'hb8f003a4),
	.w4(32'h39b6d1c2),
	.w5(32'h3b4b73d7),
	.w6(32'hbb690202),
	.w7(32'hba686905),
	.w8(32'hba8003c2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b856c49),
	.w1(32'h3b814640),
	.w2(32'h3bc80305),
	.w3(32'h3a9caeed),
	.w4(32'h3bb2d177),
	.w5(32'h3a5906d2),
	.w6(32'hbbf38f82),
	.w7(32'hba80786b),
	.w8(32'hbae9309f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8daae6),
	.w1(32'hba9eebf0),
	.w2(32'h3b8ddde6),
	.w3(32'h39f625f0),
	.w4(32'h3b8e0b61),
	.w5(32'h39dceffb),
	.w6(32'hbb3ef110),
	.w7(32'h3b769c38),
	.w8(32'h3ab160b2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27e880),
	.w1(32'h3b7992f2),
	.w2(32'h3b0c294c),
	.w3(32'h3b389366),
	.w4(32'h3af77439),
	.w5(32'h3b0208ff),
	.w6(32'h3b6b8bfd),
	.w7(32'h3b362be0),
	.w8(32'h3b306c27),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b067dd7),
	.w1(32'hbb16152d),
	.w2(32'hbb37faad),
	.w3(32'hba309721),
	.w4(32'hbb0b5fed),
	.w5(32'h3a23f98b),
	.w6(32'hbb06b223),
	.w7(32'hbb30f736),
	.w8(32'hb8a06538),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f15a),
	.w1(32'h3b6a39e3),
	.w2(32'h3b08b29a),
	.w3(32'h3b013a80),
	.w4(32'h3afc4c4a),
	.w5(32'hbb381491),
	.w6(32'h3aea0f08),
	.w7(32'h3a35887f),
	.w8(32'hbbcdf932),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93ae6b),
	.w1(32'hbb59b9a9),
	.w2(32'hbb29608e),
	.w3(32'hbb876652),
	.w4(32'hba62bc14),
	.w5(32'hb9f7afa7),
	.w6(32'h38a5986f),
	.w7(32'hba11341d),
	.w8(32'hba6a1222),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5c74a),
	.w1(32'hbb1f2711),
	.w2(32'hbb2846dc),
	.w3(32'h39eb85cd),
	.w4(32'hb9ee469d),
	.w5(32'h3c03a7b9),
	.w6(32'hbb207a68),
	.w7(32'hbaefc1eb),
	.w8(32'h3b630034),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b7e83),
	.w1(32'hbb92ccf3),
	.w2(32'h3a050f42),
	.w3(32'hbb837d46),
	.w4(32'hbb167477),
	.w5(32'h3c19d4b3),
	.w6(32'hb97b94b9),
	.w7(32'h3b0322e6),
	.w8(32'h3c2696eb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e6672),
	.w1(32'hbb435a8c),
	.w2(32'hba89e86b),
	.w3(32'hbb6e4955),
	.w4(32'hbadef07f),
	.w5(32'h3a91f314),
	.w6(32'hbae03d2b),
	.w7(32'hbb05f0a0),
	.w8(32'h3a96b07e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba906769),
	.w1(32'hba80893c),
	.w2(32'hb9b76a3c),
	.w3(32'hbae1a96c),
	.w4(32'h3a2d69e4),
	.w5(32'hbb89d8ae),
	.w6(32'hb90469fb),
	.w7(32'hb88f92d2),
	.w8(32'hbb40652a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34183d),
	.w1(32'hbb1872bd),
	.w2(32'h399a73d3),
	.w3(32'hbb479343),
	.w4(32'hba934e57),
	.w5(32'hbb03d00c),
	.w6(32'hbaf01e56),
	.w7(32'hba8840cd),
	.w8(32'hbadcc912),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a162bb7),
	.w1(32'h3b0b636c),
	.w2(32'h3833e8f3),
	.w3(32'h39b02808),
	.w4(32'h3afa9427),
	.w5(32'h3a473e2b),
	.w6(32'h39114aef),
	.w7(32'hba69a099),
	.w8(32'hb9e8add1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeef60c),
	.w1(32'hbba660d5),
	.w2(32'hbb0c6242),
	.w3(32'hbbad1252),
	.w4(32'hbb39f528),
	.w5(32'hbac0c73e),
	.w6(32'hbb015dd2),
	.w7(32'hbab67d16),
	.w8(32'hbae6f4fd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c87a9a),
	.w1(32'h398fd864),
	.w2(32'hbb3a85e2),
	.w3(32'h367eb16e),
	.w4(32'hbb3b254a),
	.w5(32'hbbb3d53b),
	.w6(32'hb90c390b),
	.w7(32'hbba6e7d3),
	.w8(32'hbbea2195),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d7743),
	.w1(32'h3a43a336),
	.w2(32'hbb42409f),
	.w3(32'h3a0da583),
	.w4(32'h3b410a85),
	.w5(32'hbb0529f0),
	.w6(32'h3b528ae5),
	.w7(32'hba9bfbfc),
	.w8(32'h3bc504a5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbd06a),
	.w1(32'h3b6e3af0),
	.w2(32'hbae29b14),
	.w3(32'hbabcbaff),
	.w4(32'h3b3c4b73),
	.w5(32'h3b4a1e25),
	.w6(32'h3a7822fc),
	.w7(32'hbae544c4),
	.w8(32'hba8f2ba2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49a775),
	.w1(32'hbaf953cf),
	.w2(32'h3b1406ff),
	.w3(32'hbadfdb73),
	.w4(32'h396305a8),
	.w5(32'hbb349c18),
	.w6(32'hbbf03911),
	.w7(32'hb9f590cb),
	.w8(32'hbbd804bc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915e8cc),
	.w1(32'h39bba28a),
	.w2(32'hb8a9f696),
	.w3(32'h3a807b7f),
	.w4(32'h3b27c33d),
	.w5(32'hba2c0c4b),
	.w6(32'hbb26708d),
	.w7(32'hbb444c6d),
	.w8(32'hbad0d990),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f6fe9),
	.w1(32'h3aa17b6e),
	.w2(32'h3ae74e05),
	.w3(32'h3aa7b3ff),
	.w4(32'h3aaa22f9),
	.w5(32'hbb98cb33),
	.w6(32'h3a74e2c2),
	.w7(32'h389c4bc8),
	.w8(32'hbb268fc6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab93cc9),
	.w1(32'hbba52d47),
	.w2(32'hbab389a7),
	.w3(32'hbb8cf9d3),
	.w4(32'h3b14f638),
	.w5(32'h3b8e1d5b),
	.w6(32'hbad7e917),
	.w7(32'h3a7eb1ea),
	.w8(32'h3951382a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf781c1),
	.w1(32'hbb72ce80),
	.w2(32'hbb1a7f9c),
	.w3(32'h3aa3b78a),
	.w4(32'hba05e33e),
	.w5(32'h3bad6a8a),
	.w6(32'hbaa28164),
	.w7(32'hba3772fd),
	.w8(32'h3b12516b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b713a97),
	.w1(32'hb9f095c3),
	.w2(32'h3bb7379b),
	.w3(32'h3b5da9b8),
	.w4(32'h391cd986),
	.w5(32'hbb650315),
	.w6(32'hbb843ade),
	.w7(32'h3acdb31b),
	.w8(32'hbbb02a59),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0e403),
	.w1(32'hbbb25006),
	.w2(32'hbb8a4a10),
	.w3(32'hbb1173c0),
	.w4(32'hbb37e462),
	.w5(32'hbbb61ecb),
	.w6(32'hbb95d717),
	.w7(32'hbb884b26),
	.w8(32'hbbbb7db7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc04a9e),
	.w1(32'hbbbf8348),
	.w2(32'hbb941884),
	.w3(32'hbbcaecbd),
	.w4(32'hbb84939a),
	.w5(32'h3b903c31),
	.w6(32'hbb28af32),
	.w7(32'hbbba08e7),
	.w8(32'h3bb9d55c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38897f),
	.w1(32'hb98c8f94),
	.w2(32'h39b2a54d),
	.w3(32'h3ba3a157),
	.w4(32'h3b590065),
	.w5(32'hbb11148b),
	.w6(32'hbb4aba8b),
	.w7(32'hba95d7d3),
	.w8(32'hbb17fe69),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bd0e0),
	.w1(32'hb6dc9a47),
	.w2(32'hb9b7e563),
	.w3(32'hb5a1285d),
	.w4(32'hba4f6b75),
	.w5(32'hbbe605d0),
	.w6(32'h3afdbf63),
	.w7(32'h3aa264b4),
	.w8(32'hbb660ea1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77aac8),
	.w1(32'h3c039d9d),
	.w2(32'hbb1246c4),
	.w3(32'hbab28e24),
	.w4(32'h3b372705),
	.w5(32'hbb761066),
	.w6(32'h3b4d3e99),
	.w7(32'hbb67c34e),
	.w8(32'hbab2536a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a4efa),
	.w1(32'hbb12f778),
	.w2(32'hbb1f8560),
	.w3(32'hbb2a23ae),
	.w4(32'hbb08211d),
	.w5(32'h3b2ca79c),
	.w6(32'hb8b5c427),
	.w7(32'hb926a936),
	.w8(32'h3b920c33),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d5074),
	.w1(32'h3b148c94),
	.w2(32'hbb11b72d),
	.w3(32'hbadaeb4a),
	.w4(32'hba16b98c),
	.w5(32'h3c1c1a5d),
	.w6(32'h3a6b16ec),
	.w7(32'hbb5c92b2),
	.w8(32'h3c14a3a8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce91e0),
	.w1(32'hb8d5e8b4),
	.w2(32'h3af65ccf),
	.w3(32'h3b1fc27e),
	.w4(32'hbaebebc9),
	.w5(32'h3a8df1f8),
	.w6(32'hbad442ee),
	.w7(32'hbad29638),
	.w8(32'h3abf057b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7cfd1),
	.w1(32'h3a6b3784),
	.w2(32'hbb25e0b3),
	.w3(32'h39af5c9b),
	.w4(32'hba778001),
	.w5(32'h3b5c0118),
	.w6(32'hba515adc),
	.w7(32'hbb1916a6),
	.w8(32'h3a5754d3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2db01),
	.w1(32'hba1d5303),
	.w2(32'hb9dab91f),
	.w3(32'h3731a41d),
	.w4(32'hba9ae3bb),
	.w5(32'h3b17c6a9),
	.w6(32'hb714987f),
	.w7(32'hbacb0e92),
	.w8(32'h3b210b20),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa052b0),
	.w1(32'hba00d9fe),
	.w2(32'hba3faefe),
	.w3(32'h3aaa0bfd),
	.w4(32'hba50e251),
	.w5(32'h3b5dee59),
	.w6(32'hbadc10be),
	.w7(32'hbaafb4c2),
	.w8(32'h3b8b781c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43da84),
	.w1(32'h3af6bd75),
	.w2(32'hbad5639f),
	.w3(32'h3b15af49),
	.w4(32'hb9eed4ad),
	.w5(32'h3bb8735c),
	.w6(32'h3a90abf2),
	.w7(32'hbadc7046),
	.w8(32'h3b96821a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb83825),
	.w1(32'h3a759183),
	.w2(32'h3b43aba9),
	.w3(32'h3b3f7946),
	.w4(32'h3b5cf7d6),
	.w5(32'hbb389126),
	.w6(32'hbbc7238c),
	.w7(32'hbaa40e21),
	.w8(32'h3981e4ef),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20f7cd),
	.w1(32'h3ae1012d),
	.w2(32'h3a406627),
	.w3(32'hbb081f1f),
	.w4(32'hba8390d9),
	.w5(32'h3b3d7984),
	.w6(32'h3b8195a0),
	.w7(32'h3b338b67),
	.w8(32'h3b694c21),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad33619),
	.w1(32'h3a312b86),
	.w2(32'hbb3ebb9c),
	.w3(32'hba572a56),
	.w4(32'hbaff5dad),
	.w5(32'h3a24d3cb),
	.w6(32'hb9b59ef0),
	.w7(32'hbb89dfdf),
	.w8(32'hbb804d0c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51eee5),
	.w1(32'hbb33193e),
	.w2(32'hb9ca4f75),
	.w3(32'hbb54d7c9),
	.w4(32'h3a21148f),
	.w5(32'hbabff20b),
	.w6(32'h3aad61fb),
	.w7(32'h3a7d73eb),
	.w8(32'hba69a71f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05f11c),
	.w1(32'hbbcc3418),
	.w2(32'hbbe07726),
	.w3(32'hbbb127d2),
	.w4(32'hbc035684),
	.w5(32'h3a6acb76),
	.w6(32'hbbaf6934),
	.w7(32'hbbc4bcd5),
	.w8(32'hbadb031a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba968f11),
	.w1(32'h3a15109a),
	.w2(32'h3b2f68f3),
	.w3(32'hba4e59ef),
	.w4(32'h3b3d67c3),
	.w5(32'h3b89c119),
	.w6(32'h3a1a1dd8),
	.w7(32'h3b364e54),
	.w8(32'h3aba4ccc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66f775),
	.w1(32'hbb3234b9),
	.w2(32'h3a8b05a2),
	.w3(32'h3a835e12),
	.w4(32'hb9519893),
	.w5(32'hbb1178e5),
	.w6(32'hbba1a8a2),
	.w7(32'hbb6c5342),
	.w8(32'hbb05c9c3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9904d5),
	.w1(32'hbba66b11),
	.w2(32'h385e99ef),
	.w3(32'hbb4ed580),
	.w4(32'hba924833),
	.w5(32'hb9afee34),
	.w6(32'hbb3d1ca9),
	.w7(32'hba5fa649),
	.w8(32'hbb68b012),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb4f6c),
	.w1(32'hbb5a9842),
	.w2(32'hba837e0b),
	.w3(32'hb8cc59d8),
	.w4(32'hba1b7204),
	.w5(32'h3b84b366),
	.w6(32'hba155c39),
	.w7(32'hbaaaf4d3),
	.w8(32'h3b29f76e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58b176),
	.w1(32'h3acb3574),
	.w2(32'h3b57bf4a),
	.w3(32'h3b6ac577),
	.w4(32'h3b5e6902),
	.w5(32'h3c8da02e),
	.w6(32'hba26803c),
	.w7(32'h3a6c69b7),
	.w8(32'h3c24f482),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba73f59),
	.w1(32'hbab20ff2),
	.w2(32'h3c167912),
	.w3(32'h3aeb00f6),
	.w4(32'h3bc18bdb),
	.w5(32'h3a96089c),
	.w6(32'hbb4da769),
	.w7(32'h3c191d2f),
	.w8(32'h3ba45de1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb200e3),
	.w1(32'hbb31e19e),
	.w2(32'hbb9886bd),
	.w3(32'hbb0b52c8),
	.w4(32'hbbc8de63),
	.w5(32'hba5075b3),
	.w6(32'hbbf08e3c),
	.w7(32'hbc2c305a),
	.w8(32'hbb4b71b8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb734007),
	.w1(32'hbc45707c),
	.w2(32'hba0864b2),
	.w3(32'hbc39d5b4),
	.w4(32'hbb8c3b91),
	.w5(32'hbba71081),
	.w6(32'hbbdbe4ce),
	.w7(32'hb972b31a),
	.w8(32'hbb92ba4e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb666110),
	.w1(32'hbb7ea73a),
	.w2(32'hbb3f2a05),
	.w3(32'hbb487495),
	.w4(32'hbb43fec9),
	.w5(32'h3ac94f20),
	.w6(32'hbb1d2d95),
	.w7(32'hbba39731),
	.w8(32'hbac0ab75),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb266573),
	.w1(32'hbb9f723d),
	.w2(32'h3b0b1229),
	.w3(32'hbab2d6e3),
	.w4(32'h3b725b4c),
	.w5(32'h3abe48f5),
	.w6(32'hbb5711ca),
	.w7(32'h3ae73218),
	.w8(32'hbaa6cf08),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba444cd1),
	.w1(32'h3bc50a40),
	.w2(32'h3afe9b1e),
	.w3(32'h3b2f26f8),
	.w4(32'h3b58d3f8),
	.w5(32'hb945d696),
	.w6(32'h3bb7aef7),
	.w7(32'h3b31851a),
	.w8(32'hba9670ff),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba14f48),
	.w1(32'hbad3f933),
	.w2(32'hbb671714),
	.w3(32'h3bc672e6),
	.w4(32'hb8772330),
	.w5(32'hbb053772),
	.w6(32'h3bc95b70),
	.w7(32'h37fde808),
	.w8(32'hbaa29012),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44fae8),
	.w1(32'hb84dbbce),
	.w2(32'hbb9f6821),
	.w3(32'hbb31b75c),
	.w4(32'hbb9e7c52),
	.w5(32'hb975c1ea),
	.w6(32'hbafcad6c),
	.w7(32'hbb887758),
	.w8(32'hbb2d19ab),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44050),
	.w1(32'hbb20839a),
	.w2(32'h3a947b21),
	.w3(32'hbb26e768),
	.w4(32'hba90c6c7),
	.w5(32'hba153c29),
	.w6(32'hb9ca1ed9),
	.w7(32'h3aed7d87),
	.w8(32'h3a3dea87),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0924c3),
	.w1(32'hbb202794),
	.w2(32'hbae25382),
	.w3(32'hbb11fffd),
	.w4(32'hba3250c2),
	.w5(32'h3b0ac22b),
	.w6(32'hbb0cee2a),
	.w7(32'hbabe260e),
	.w8(32'h3b021f4e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cbd9b),
	.w1(32'h3b4aa83c),
	.w2(32'h3aef3030),
	.w3(32'h3b3e0f69),
	.w4(32'h3ab7c7d2),
	.w5(32'hb8b850f9),
	.w6(32'h3bc8ed81),
	.w7(32'h3b451496),
	.w8(32'hba0e4333),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6127d1),
	.w1(32'h3a6d82bf),
	.w2(32'hbbacf275),
	.w3(32'hb9a728eb),
	.w4(32'hbb8b6407),
	.w5(32'h38ff390c),
	.w6(32'h39821c99),
	.w7(32'hbbddd488),
	.w8(32'h3b883d0a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8c1a9),
	.w1(32'hbaca150a),
	.w2(32'hbab3373b),
	.w3(32'hb9b97ca1),
	.w4(32'h3b3b8778),
	.w5(32'hb9806235),
	.w6(32'h3b0d4c1e),
	.w7(32'hb93528ed),
	.w8(32'hba06f154),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac583a4),
	.w1(32'hb94fad13),
	.w2(32'hbb599d1a),
	.w3(32'hba94f7dd),
	.w4(32'h39157054),
	.w5(32'hbbd25b5c),
	.w6(32'hb94cd30b),
	.w7(32'hbab79007),
	.w8(32'hbbf7b22a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb73589),
	.w1(32'hbb3744c7),
	.w2(32'h3a6ff00d),
	.w3(32'hbb986b8e),
	.w4(32'hba0074ef),
	.w5(32'h3bd44c94),
	.w6(32'hbb673ef4),
	.w7(32'h3b618c80),
	.w8(32'h3bd2c613),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30b884),
	.w1(32'hbb0756dc),
	.w2(32'hbbb12e65),
	.w3(32'hb68f84e4),
	.w4(32'hbb991578),
	.w5(32'hba62f0b5),
	.w6(32'hba6d1586),
	.w7(32'hbba10b8e),
	.w8(32'h3b10ef4f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956404d),
	.w1(32'hbb3c38fd),
	.w2(32'hbaa5aec0),
	.w3(32'hbaddd207),
	.w4(32'hbadff31b),
	.w5(32'h3ae8d1e7),
	.w6(32'hb96ffbec),
	.w7(32'hbb214cc9),
	.w8(32'h3bd0a723),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28922e),
	.w1(32'h3b82fe1b),
	.w2(32'hb9a26048),
	.w3(32'h3ab7bfc2),
	.w4(32'hbb8e2a3b),
	.w5(32'hb9aff9d7),
	.w6(32'h3b33b9b0),
	.w7(32'hbb936883),
	.w8(32'hbacbc5d7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98f31c),
	.w1(32'hba83b0ad),
	.w2(32'h3ac9a1c5),
	.w3(32'h39e90602),
	.w4(32'h3aa3e22a),
	.w5(32'hbc36c597),
	.w6(32'hbab3e375),
	.w7(32'h38f191c6),
	.w8(32'hbc1c267c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc202644),
	.w1(32'hbc01be68),
	.w2(32'hbb9c8897),
	.w3(32'hbc283f95),
	.w4(32'hbb8fd898),
	.w5(32'hbb966f93),
	.w6(32'hbc1b3326),
	.w7(32'hbb999720),
	.w8(32'hbb8692c2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c9e35),
	.w1(32'hbb90f5c9),
	.w2(32'hbb0b8607),
	.w3(32'hbbb2552c),
	.w4(32'hbae987ac),
	.w5(32'h3a6f4ade),
	.w6(32'hbbcbb6ab),
	.w7(32'hbb571af8),
	.w8(32'h3b9536c8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23ffc9),
	.w1(32'hbabc6451),
	.w2(32'hbaa5dd22),
	.w3(32'h3ab1c83b),
	.w4(32'hbb9bb650),
	.w5(32'h3b3edd58),
	.w6(32'h36b496d7),
	.w7(32'hbb57d4bb),
	.w8(32'h3a9af2d6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3e6a6),
	.w1(32'hba00c147),
	.w2(32'hbbb5540c),
	.w3(32'hbae47e21),
	.w4(32'hbb29faa2),
	.w5(32'h39c0abbf),
	.w6(32'hbb72242a),
	.w7(32'hbb5e719b),
	.w8(32'h3a74bfc8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39703a5d),
	.w1(32'hbad01d01),
	.w2(32'hb9886079),
	.w3(32'h3a3452e5),
	.w4(32'hba1db0e9),
	.w5(32'h3a9d27ec),
	.w6(32'hbaea4228),
	.w7(32'hbb76777b),
	.w8(32'h3b5259df),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af68063),
	.w1(32'hbad19778),
	.w2(32'hbb2803b7),
	.w3(32'hbb1ca3c0),
	.w4(32'hbb175ee1),
	.w5(32'hba51e6fd),
	.w6(32'hba95a9d5),
	.w7(32'hbb0c0207),
	.w8(32'h39896f16),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6930f5),
	.w1(32'h3bb8a2ef),
	.w2(32'h3bb09392),
	.w3(32'hba06ea4d),
	.w4(32'hba6b2fe1),
	.w5(32'h3adc2a78),
	.w6(32'h3bfde973),
	.w7(32'h3b823cd4),
	.w8(32'h3b44d21a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba590a0),
	.w1(32'h3b21bb1c),
	.w2(32'h398f8c7a),
	.w3(32'h391815f8),
	.w4(32'h3b103403),
	.w5(32'h3b929470),
	.w6(32'hba8eb46b),
	.w7(32'h3ae14b17),
	.w8(32'h3b8a7d1f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51697c),
	.w1(32'h3a5915c8),
	.w2(32'hbb3b1918),
	.w3(32'h3b40801e),
	.w4(32'h3a875d64),
	.w5(32'h3a6d1f8d),
	.w6(32'h3ae58dfd),
	.w7(32'hba9274b1),
	.w8(32'h3b2cdf97),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a5ce8),
	.w1(32'h3a06f404),
	.w2(32'hba2c0858),
	.w3(32'h3a4380cb),
	.w4(32'h3b751d11),
	.w5(32'h3bc459ba),
	.w6(32'h3b8a0b0e),
	.w7(32'h3a9a09c1),
	.w8(32'h3bba64ae),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87533c),
	.w1(32'hbac6d798),
	.w2(32'hbaac49f8),
	.w3(32'h3accea3e),
	.w4(32'h3ad5e1e8),
	.w5(32'hbbef817c),
	.w6(32'h3ac81632),
	.w7(32'h390e7580),
	.w8(32'hbc1379d7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd7613),
	.w1(32'hbc11f7ca),
	.w2(32'hbbcbdb62),
	.w3(32'hbc054461),
	.w4(32'hbb92c3ef),
	.w5(32'h3b1ee881),
	.w6(32'hbbfc2f4e),
	.w7(32'hbbe7e17d),
	.w8(32'h3b3e4954),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c611c),
	.w1(32'h39492942),
	.w2(32'h3a0f59bf),
	.w3(32'hbab6473b),
	.w4(32'h393f61f6),
	.w5(32'hbab474b0),
	.w6(32'hbb4fe23f),
	.w7(32'h39e8e5dd),
	.w8(32'hbb995948),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88595f),
	.w1(32'h3b9cd313),
	.w2(32'h3c556b02),
	.w3(32'h3b831325),
	.w4(32'h3c1a134b),
	.w5(32'hbc171305),
	.w6(32'h3b530033),
	.w7(32'h3bfb345e),
	.w8(32'h3992d103),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c262e52),
	.w1(32'h3c15b22e),
	.w2(32'h3c0ecb01),
	.w3(32'hbc019825),
	.w4(32'hbabff386),
	.w5(32'h3b85c919),
	.w6(32'h3b69a875),
	.w7(32'h3bcc2f77),
	.w8(32'hb9e662a4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ca5cf),
	.w1(32'h3b912388),
	.w2(32'h3b99cdac),
	.w3(32'h3bb6dbcd),
	.w4(32'h3bb8fd1f),
	.w5(32'hbbfc2dc6),
	.w6(32'h3b9d4041),
	.w7(32'h3b747433),
	.w8(32'hbb030629),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa5b58),
	.w1(32'h3bc6a1a3),
	.w2(32'h3c049a82),
	.w3(32'hbbc8872b),
	.w4(32'hbabd7671),
	.w5(32'hbb130a6f),
	.w6(32'hb8aaf1fb),
	.w7(32'h3bc2ea84),
	.w8(32'h3a62f5f3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfc18a),
	.w1(32'hbb2b25c7),
	.w2(32'hbb41785d),
	.w3(32'hbb653067),
	.w4(32'hbbc51df0),
	.w5(32'hba6fd887),
	.w6(32'hb95e7689),
	.w7(32'hbb8de969),
	.w8(32'h3912faba),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2c19c),
	.w1(32'hbaea489f),
	.w2(32'hbb0e90b5),
	.w3(32'hbb2b6be9),
	.w4(32'hbaed1ad8),
	.w5(32'h3a5d57e8),
	.w6(32'hbb384bd5),
	.w7(32'hbb0045c3),
	.w8(32'h3a42056f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad60537),
	.w1(32'h3c064832),
	.w2(32'h3b57f2e1),
	.w3(32'h3afd80e8),
	.w4(32'hb9fe253a),
	.w5(32'hbbeca5a2),
	.w6(32'h3bbe964a),
	.w7(32'h37deb769),
	.w8(32'hbc0645e7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cc419),
	.w1(32'hbc27ce0a),
	.w2(32'hbbfa2120),
	.w3(32'hbbd8281a),
	.w4(32'hbbef5f6b),
	.w5(32'hb9adfc0b),
	.w6(32'hbbeccf30),
	.w7(32'hbc10948d),
	.w8(32'hb99a3e45),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb086935),
	.w1(32'hba873443),
	.w2(32'h3b1e8a65),
	.w3(32'hbaa1c998),
	.w4(32'hb8c76161),
	.w5(32'h3aef6490),
	.w6(32'hb8d0c55a),
	.w7(32'hba61f95b),
	.w8(32'h3b6a09ef),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d37bc),
	.w1(32'h3a10f43b),
	.w2(32'h395eca47),
	.w3(32'hbb0566bf),
	.w4(32'hbb42815a),
	.w5(32'hba262155),
	.w6(32'hbb4bcf83),
	.w7(32'hbb06818e),
	.w8(32'hbabc58d9),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c5890),
	.w1(32'h3a502c68),
	.w2(32'h3b33a6ec),
	.w3(32'hb789e905),
	.w4(32'h3ae75394),
	.w5(32'h3bccf306),
	.w6(32'hba84071c),
	.w7(32'h3b29d36b),
	.w8(32'h3b8cc5d5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd442ac),
	.w1(32'h3c2d519b),
	.w2(32'h3c36f2be),
	.w3(32'h3b997a53),
	.w4(32'h3c2fa89a),
	.w5(32'h3a53eca7),
	.w6(32'h3c545b70),
	.w7(32'h3c4fdeed),
	.w8(32'h3b56186d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b392385),
	.w1(32'h3a2aebad),
	.w2(32'h3b06ff0a),
	.w3(32'hba0e60b1),
	.w4(32'h39c56603),
	.w5(32'h3b50006e),
	.w6(32'hba1e2097),
	.w7(32'h3935fbcb),
	.w8(32'h3b850424),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26830c),
	.w1(32'hba181751),
	.w2(32'h371823f7),
	.w3(32'h39a20419),
	.w4(32'h393a79a4),
	.w5(32'h3b86f315),
	.w6(32'hba6f750b),
	.w7(32'hba731619),
	.w8(32'h3b41e0ec),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05523e),
	.w1(32'hbbaa0797),
	.w2(32'hbb225463),
	.w3(32'h3b67cf20),
	.w4(32'hbb16a41d),
	.w5(32'h38d5332b),
	.w6(32'h3a84f9af),
	.w7(32'hbb0a87b4),
	.w8(32'h3a3ea76e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2ee02),
	.w1(32'hbb2b0ed7),
	.w2(32'hb9ab5ad4),
	.w3(32'hbaa11e05),
	.w4(32'h3a498288),
	.w5(32'h3a9f1eaa),
	.w6(32'hbb3ca048),
	.w7(32'hbb043a82),
	.w8(32'h3b2dc8c5),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2db96a),
	.w1(32'hb951d11e),
	.w2(32'h39f77668),
	.w3(32'hb9bece8d),
	.w4(32'h3a08cc36),
	.w5(32'h3affedc0),
	.w6(32'hbabda5fa),
	.w7(32'hb91351d9),
	.w8(32'h3b805334),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9167d9),
	.w1(32'h3b838b9b),
	.w2(32'h3bc2a6e9),
	.w3(32'h3ab8f964),
	.w4(32'h3a8cc0b7),
	.w5(32'hba3916ae),
	.w6(32'h3acf4c57),
	.w7(32'h3b19f982),
	.w8(32'h3ae35477),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79c7d9),
	.w1(32'hbb2cc35d),
	.w2(32'hbb559d9e),
	.w3(32'hba5acfb7),
	.w4(32'hbac63b76),
	.w5(32'hbb190787),
	.w6(32'hb859cc1b),
	.w7(32'hba9953be),
	.w8(32'hbb1e3fe0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68eb3d),
	.w1(32'h3b1089ec),
	.w2(32'h3a7da910),
	.w3(32'h38817600),
	.w4(32'hb8e434cf),
	.w5(32'hbb508824),
	.w6(32'hba050c64),
	.w7(32'h3ad09f87),
	.w8(32'hbbc1cd0b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb483af9),
	.w1(32'h3a2a9166),
	.w2(32'hba0f2e62),
	.w3(32'h3a1db84a),
	.w4(32'hba89fd77),
	.w5(32'h3b6ed78b),
	.w6(32'h3a055e77),
	.w7(32'h39d75055),
	.w8(32'h3bb2ddad),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f5c6d),
	.w1(32'h3b3aae54),
	.w2(32'h3b7ccf46),
	.w3(32'h3b690a81),
	.w4(32'h39f58a53),
	.w5(32'h39668289),
	.w6(32'h3aca1532),
	.w7(32'h3aa2b987),
	.w8(32'h3a9712fa),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b852c),
	.w1(32'hbb9942e3),
	.w2(32'hba923f00),
	.w3(32'hbb501d3c),
	.w4(32'hbae62244),
	.w5(32'h3af7126b),
	.w6(32'hbbc8a97d),
	.w7(32'hbb803c42),
	.w8(32'h3ac68d9b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37304aa6),
	.w1(32'hbac5a525),
	.w2(32'h3a663ae8),
	.w3(32'hb9825979),
	.w4(32'hb9cccc4e),
	.w5(32'hbb28fd88),
	.w6(32'hbb195845),
	.w7(32'hbaeb446a),
	.w8(32'hb9673ee8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa38489),
	.w1(32'h3ab777b9),
	.w2(32'h3b55e849),
	.w3(32'hbaac9a9d),
	.w4(32'h3a1c78d9),
	.w5(32'h3a81e2ec),
	.w6(32'h3a885e17),
	.w7(32'h3b0908f7),
	.w8(32'h3b4a4c58),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac837e9),
	.w1(32'hb8b9c979),
	.w2(32'h3a5be5a2),
	.w3(32'hb9c7d785),
	.w4(32'hbacd2abf),
	.w5(32'h3b4aa1e8),
	.w6(32'h3a633463),
	.w7(32'hbb02b221),
	.w8(32'h3b41b6f1),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0b20c),
	.w1(32'hbada7bf3),
	.w2(32'hba835a4d),
	.w3(32'h3a2227cd),
	.w4(32'hbb72d836),
	.w5(32'h3aab2510),
	.w6(32'h3a945e2b),
	.w7(32'hba4863b3),
	.w8(32'h3b40971e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0df687),
	.w1(32'hbb82a9fd),
	.w2(32'hba917dd1),
	.w3(32'hbba603bc),
	.w4(32'hbb82fac3),
	.w5(32'h3b269d0a),
	.w6(32'hbc03ec44),
	.w7(32'hbb974f9e),
	.w8(32'h3b25ae3a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42bc54),
	.w1(32'hb84f5989),
	.w2(32'hbb37b047),
	.w3(32'h3aa39f9f),
	.w4(32'h398f0bcf),
	.w5(32'h3aa62e45),
	.w6(32'hb9fd626e),
	.w7(32'hbb2ef14d),
	.w8(32'h3b09f7f6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba203d4c),
	.w1(32'h399e20ee),
	.w2(32'h3966fd5a),
	.w3(32'hb989e486),
	.w4(32'hba9942d4),
	.w5(32'h3b6dfe8b),
	.w6(32'hba81f2e7),
	.w7(32'hba02eb66),
	.w8(32'hbb1b74a6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac22426),
	.w1(32'hbba66805),
	.w2(32'h3b97f16a),
	.w3(32'hbbaf846d),
	.w4(32'hb7acb732),
	.w5(32'hbb08a95e),
	.w6(32'hbc273143),
	.w7(32'h3b5a9adc),
	.w8(32'hbac4b5eb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb382734),
	.w1(32'hbbb2b7d8),
	.w2(32'hbb8d1db5),
	.w3(32'hbb6b00a5),
	.w4(32'hba81cc0f),
	.w5(32'h3b795fe9),
	.w6(32'hbb748906),
	.w7(32'hbba3be07),
	.w8(32'h3bc2c965),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6f64f),
	.w1(32'h3b17d1e6),
	.w2(32'hbb6b71cb),
	.w3(32'h3b8c4cfe),
	.w4(32'hbb3c9c09),
	.w5(32'hbbe6ca8c),
	.w6(32'h3b47f5f3),
	.w7(32'hbb929b94),
	.w8(32'hbc17a8d0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe35c49),
	.w1(32'hbbc23dfc),
	.w2(32'hbbe2f5f1),
	.w3(32'hbbf8bc48),
	.w4(32'hbbf91fb5),
	.w5(32'hbbf568e0),
	.w6(32'hbc192a5c),
	.w7(32'hbc07fca3),
	.w8(32'hbbd12d60),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd27eae),
	.w1(32'hbbf7f66f),
	.w2(32'hbba3ad1c),
	.w3(32'hbc05c69f),
	.w4(32'hbb893230),
	.w5(32'hbafb817b),
	.w6(32'hbc0107db),
	.w7(32'hbbd3aad4),
	.w8(32'hbb26c710),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8093e7),
	.w1(32'hba97ddf3),
	.w2(32'h39923ccc),
	.w3(32'hba400911),
	.w4(32'hbac51923),
	.w5(32'h3b2863ad),
	.w6(32'h3b09ad61),
	.w7(32'hbb2e50aa),
	.w8(32'hb9311617),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b33dde),
	.w1(32'h3c06144f),
	.w2(32'h3bf88c40),
	.w3(32'h3c01a024),
	.w4(32'h3c04ec81),
	.w5(32'h3ba8d487),
	.w6(32'h3c17d0dc),
	.w7(32'h3bfb1089),
	.w8(32'h3b270674),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92c8e0c),
	.w1(32'hbaf99248),
	.w2(32'hba5c3e5b),
	.w3(32'hbabbf8be),
	.w4(32'h3b971044),
	.w5(32'h3b0bd04d),
	.w6(32'h3b635acd),
	.w7(32'h3b444846),
	.w8(32'h3bc0c0cb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3634f),
	.w1(32'hba2d882c),
	.w2(32'hbb1cbe2a),
	.w3(32'hbb3ebfdd),
	.w4(32'hbbc27c54),
	.w5(32'h3b19c8f5),
	.w6(32'h3ad4b6f9),
	.w7(32'hbb64f885),
	.w8(32'h3a86f922),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82ca20),
	.w1(32'h3b99267e),
	.w2(32'hbb47a85f),
	.w3(32'h3b5c9116),
	.w4(32'hb7c0041d),
	.w5(32'hbb123a7b),
	.w6(32'h3bbc5c9b),
	.w7(32'hbaa2d691),
	.w8(32'hba378099),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eae7a),
	.w1(32'hba1ad208),
	.w2(32'h3b3a3359),
	.w3(32'hbafd25f1),
	.w4(32'hba2bb391),
	.w5(32'hbb363563),
	.w6(32'h394c54f4),
	.w7(32'h38638e13),
	.w8(32'hbad456eb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2012b3),
	.w1(32'hbba0651c),
	.w2(32'hbb58858c),
	.w3(32'hbb23de2f),
	.w4(32'hbb6bf598),
	.w5(32'h3ba67dd3),
	.w6(32'hbb08b7f9),
	.w7(32'hbb8fb69b),
	.w8(32'h3be87a29),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82ce23),
	.w1(32'hb99986ea),
	.w2(32'h3bd11c0e),
	.w3(32'h3a45cfb9),
	.w4(32'h3b8e273d),
	.w5(32'h3b310000),
	.w6(32'h389a3538),
	.w7(32'h3b2f28eb),
	.w8(32'h3b9a0819),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af77a15),
	.w1(32'hba9acc84),
	.w2(32'h3a3f44ac),
	.w3(32'h3afe7934),
	.w4(32'h3b4cfb66),
	.w5(32'hbb5b684f),
	.w6(32'h3b8bb10a),
	.w7(32'hba83021e),
	.w8(32'hbb009b22),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab052c5),
	.w1(32'h3aa1e488),
	.w2(32'hbb01155b),
	.w3(32'hbae9de10),
	.w4(32'hbb5a3809),
	.w5(32'h3b562181),
	.w6(32'hb9e2048d),
	.w7(32'hbb26a7e6),
	.w8(32'hbb9b223d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffa173),
	.w1(32'hbb85d9d6),
	.w2(32'h3a3940bd),
	.w3(32'h3bb28887),
	.w4(32'h3a8d0a06),
	.w5(32'hbb8228bd),
	.w6(32'hba7d1ee5),
	.w7(32'h3af00986),
	.w8(32'hbb52f5d5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949fd65),
	.w1(32'hbb27a9ca),
	.w2(32'hbb30069f),
	.w3(32'hbb271231),
	.w4(32'h3a99c990),
	.w5(32'hbb66bea8),
	.w6(32'hbb624dce),
	.w7(32'hba32672d),
	.w8(32'hbb6a363b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b75b3),
	.w1(32'hbbbd28dc),
	.w2(32'hbbf29e33),
	.w3(32'hbb82b1a9),
	.w4(32'hbb69d6b2),
	.w5(32'h3a7d680d),
	.w6(32'hbb4ebb80),
	.w7(32'hbb9cebf3),
	.w8(32'h3b069eba),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ee8ce),
	.w1(32'hbb1b230d),
	.w2(32'hbb9e2cd1),
	.w3(32'hba339b91),
	.w4(32'hbb63e7d1),
	.w5(32'hbaada234),
	.w6(32'hbb5322e2),
	.w7(32'hbbc4b6a2),
	.w8(32'hba9f1c43),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aea37f),
	.w1(32'hbb3ea709),
	.w2(32'hbba63246),
	.w3(32'hbb3bbb45),
	.w4(32'hbb6c6e5e),
	.w5(32'h39918d61),
	.w6(32'hbb095747),
	.w7(32'hbbd6fcf6),
	.w8(32'hbaf297b7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20ca7c),
	.w1(32'hbb38345a),
	.w2(32'h3a06e196),
	.w3(32'hbb9fb36b),
	.w4(32'hbbd540de),
	.w5(32'hb9a33525),
	.w6(32'hbb2378f7),
	.w7(32'hbbbe57c4),
	.w8(32'hba952115),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e402a4),
	.w1(32'hba9a2fa7),
	.w2(32'hbb93e709),
	.w3(32'hbaddcb89),
	.w4(32'hbb434906),
	.w5(32'hbb866e28),
	.w6(32'hbb2a6d6c),
	.w7(32'hbbe27d6c),
	.w8(32'hbbad2922),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce0729),
	.w1(32'hbbbed39b),
	.w2(32'hbbfbae1a),
	.w3(32'hbb4e6c65),
	.w4(32'hbb7b3966),
	.w5(32'hbbb2f210),
	.w6(32'hbb80d994),
	.w7(32'hbb5dc193),
	.w8(32'hbbe09444),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc42cab),
	.w1(32'hbbb23116),
	.w2(32'hbbe23ea5),
	.w3(32'hbba1375f),
	.w4(32'hbba3fcc3),
	.w5(32'h3b92f85a),
	.w6(32'hbbc0abb1),
	.w7(32'hbbdaa906),
	.w8(32'h3b614543),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b741fbe),
	.w1(32'h3ae539ad),
	.w2(32'hbacb338f),
	.w3(32'h3b213bbc),
	.w4(32'h3a996ff2),
	.w5(32'hbb3b7d41),
	.w6(32'hba036feb),
	.w7(32'hbb45c888),
	.w8(32'hbb8814a8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ba113),
	.w1(32'hbada3e93),
	.w2(32'h38faf8b0),
	.w3(32'hbb658ab1),
	.w4(32'hbb1f888f),
	.w5(32'h3a72a9d2),
	.w6(32'hbb7a9366),
	.w7(32'hba761f8f),
	.w8(32'h3a8e5659),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5843d),
	.w1(32'hba30ce93),
	.w2(32'hbb81abb0),
	.w3(32'h3a00f39b),
	.w4(32'hbab94b5a),
	.w5(32'h3aa00fa1),
	.w6(32'hbb03c069),
	.w7(32'hbb7a1ca0),
	.w8(32'hbadbae20),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05873b),
	.w1(32'hba0e2b7d),
	.w2(32'h3ae844f0),
	.w3(32'hbb2d80ed),
	.w4(32'h3b11ce00),
	.w5(32'h3ad66776),
	.w6(32'hbb6c337e),
	.w7(32'h3b88a36e),
	.w8(32'h3acf119d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac35529),
	.w1(32'hba695fa4),
	.w2(32'hbb1265f2),
	.w3(32'hb98aac68),
	.w4(32'hb96aea13),
	.w5(32'hba8f6792),
	.w6(32'h3b6d3d43),
	.w7(32'hba2f3ae6),
	.w8(32'hbaa3e36a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4db2c),
	.w1(32'hbb444ec5),
	.w2(32'h3a0829bf),
	.w3(32'hbb850133),
	.w4(32'hbb5ae5ed),
	.w5(32'h3a05c62a),
	.w6(32'hbb91ef7a),
	.w7(32'hba559448),
	.w8(32'h3af2a92c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b357698),
	.w1(32'h3b034ce2),
	.w2(32'h3a9193a7),
	.w3(32'h3ae27d7e),
	.w4(32'h3b160307),
	.w5(32'hba142eec),
	.w6(32'h3b3da848),
	.w7(32'h3ad41cf3),
	.w8(32'hb9bb9909),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86b332),
	.w1(32'hbb337bd8),
	.w2(32'hbac6d442),
	.w3(32'hbb179144),
	.w4(32'hbba070be),
	.w5(32'hba54cd1f),
	.w6(32'hbb2bceb8),
	.w7(32'hbb309fbf),
	.w8(32'h3a026479),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396eb30f),
	.w1(32'h397e926b),
	.w2(32'hba4157d8),
	.w3(32'hba2ee75d),
	.w4(32'hba8b8fbd),
	.w5(32'hbb03bdfa),
	.w6(32'h3b3892a5),
	.w7(32'hbaeb0c26),
	.w8(32'hbab4a32b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae44721),
	.w1(32'hbb308f66),
	.w2(32'hbb24c83b),
	.w3(32'hba7cd51d),
	.w4(32'hb9ca1932),
	.w5(32'h39e459ed),
	.w6(32'hba441e95),
	.w7(32'hbb0f07b6),
	.w8(32'hba0b8460),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf918eb),
	.w1(32'hbaa313c8),
	.w2(32'hbaf4d8d4),
	.w3(32'h3908bee0),
	.w4(32'hbad27f97),
	.w5(32'h3b24a9be),
	.w6(32'hbb0cd394),
	.w7(32'hbb167e40),
	.w8(32'h3b5414ec),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d22a3),
	.w1(32'hba1e9e9b),
	.w2(32'hbb58e8b4),
	.w3(32'h3ae258db),
	.w4(32'hb9f3a3a2),
	.w5(32'h3bbba876),
	.w6(32'hbaa05f7a),
	.w7(32'hbb6cf500),
	.w8(32'h3bf972da),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5d9d5),
	.w1(32'h3acfcb1c),
	.w2(32'hbad680e4),
	.w3(32'h3b6329f9),
	.w4(32'h3a864d30),
	.w5(32'h3b1fc6e1),
	.w6(32'h3b7d661e),
	.w7(32'h3a91b87e),
	.w8(32'hbaa45e0d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1f47),
	.w1(32'hba665958),
	.w2(32'h3ac84a70),
	.w3(32'h3bbeb664),
	.w4(32'h3a954647),
	.w5(32'h3b256017),
	.w6(32'h3b365acc),
	.w7(32'h3ac9861d),
	.w8(32'h3b67b364),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989647d),
	.w1(32'hba694a07),
	.w2(32'hbb46aa09),
	.w3(32'h3ac17219),
	.w4(32'hbb202dde),
	.w5(32'hbb0a3330),
	.w6(32'h3a69bb3d),
	.w7(32'hbb442d65),
	.w8(32'hbb680613),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43e802),
	.w1(32'hb91919f3),
	.w2(32'hb8b5cca8),
	.w3(32'hbb2d3a9e),
	.w4(32'hbb60d866),
	.w5(32'hbac897f0),
	.w6(32'hbacb1179),
	.w7(32'hba4fc01b),
	.w8(32'hbb2a8558),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafc7b5),
	.w1(32'hbaf96119),
	.w2(32'hbb074e2a),
	.w3(32'hba9c34fa),
	.w4(32'hb9b8e8a7),
	.w5(32'hbb0827ab),
	.w6(32'hba8c155a),
	.w7(32'hbb536ad7),
	.w8(32'hbba2480e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7e6ac),
	.w1(32'hbb06168a),
	.w2(32'hbbbe9a7a),
	.w3(32'hb7a5b7ac),
	.w4(32'hbbd86a83),
	.w5(32'hbb65de6c),
	.w6(32'h3a93410f),
	.w7(32'hbb692a9d),
	.w8(32'hbadcda4c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e6907),
	.w1(32'hbb279bb6),
	.w2(32'hbb1fbd8e),
	.w3(32'hbbb9dbbb),
	.w4(32'hbbaf72a2),
	.w5(32'h3a1e167a),
	.w6(32'hbaae89b5),
	.w7(32'hbab8b61b),
	.w8(32'h39d8ef93),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39853cae),
	.w1(32'hbb44671d),
	.w2(32'h3a720309),
	.w3(32'h399714b1),
	.w4(32'hbb208927),
	.w5(32'h3ba67fe6),
	.w6(32'hbaa079ca),
	.w7(32'hba133378),
	.w8(32'h3ac4ae12),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f70b1),
	.w1(32'h3c0cf835),
	.w2(32'h3bfc6e30),
	.w3(32'h3b88fc6e),
	.w4(32'h3bdad4f9),
	.w5(32'hba3ef8e2),
	.w6(32'h3b39902f),
	.w7(32'h3b62377c),
	.w8(32'hb926bbb1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4e68d),
	.w1(32'h3ba14039),
	.w2(32'h3a19a69f),
	.w3(32'h3b0fa944),
	.w4(32'hba4c2287),
	.w5(32'h3bc8859e),
	.w6(32'h3aeca4c3),
	.w7(32'h3a38b855),
	.w8(32'h3bd173a4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beadd1e),
	.w1(32'h3bae025b),
	.w2(32'h3b6e303b),
	.w3(32'h3baa7ca3),
	.w4(32'h3b4344d6),
	.w5(32'h3ac4c766),
	.w6(32'h3ba478ed),
	.w7(32'hba1e3f35),
	.w8(32'h3a950533),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc4a72),
	.w1(32'hba5b112c),
	.w2(32'hbb334049),
	.w3(32'hba961cf2),
	.w4(32'hbb1b696d),
	.w5(32'h3acdf290),
	.w6(32'hbabe2066),
	.w7(32'hbb8bd8b6),
	.w8(32'h3983924f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39196ee3),
	.w1(32'hbbe50e2a),
	.w2(32'hbabbb1e4),
	.w3(32'h3ae80c13),
	.w4(32'hbb0bbd9f),
	.w5(32'h3b1385c3),
	.w6(32'hbbbb162b),
	.w7(32'hbb43daae),
	.w8(32'hbac67685),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2383ee),
	.w1(32'hbbfdafd3),
	.w2(32'hbabe9008),
	.w3(32'h3b309b50),
	.w4(32'h3a25781a),
	.w5(32'hb9080eba),
	.w6(32'hba4c8a79),
	.w7(32'h3a507d36),
	.w8(32'hbb083c9f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e73dc),
	.w1(32'hbac58f0d),
	.w2(32'hbb377c70),
	.w3(32'hb92a383b),
	.w4(32'hbaaa1b93),
	.w5(32'hbb1e1853),
	.w6(32'h3b212e8b),
	.w7(32'hba3323f9),
	.w8(32'hbb28651b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c7075),
	.w1(32'hbb54d5e3),
	.w2(32'h3aa2a065),
	.w3(32'hbb3a1777),
	.w4(32'hbb05d1d9),
	.w5(32'hbb411238),
	.w6(32'hbb325473),
	.w7(32'hbb132fa5),
	.w8(32'hbb3bd7ec),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16a463),
	.w1(32'hba88ca3f),
	.w2(32'h39eefc01),
	.w3(32'hbb13774d),
	.w4(32'hba7d296a),
	.w5(32'hbaf32133),
	.w6(32'hbaa175b8),
	.w7(32'h3a9f434b),
	.w8(32'hbb240cc7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb200de8),
	.w1(32'hbb5df969),
	.w2(32'hbbb74933),
	.w3(32'hbb88c55f),
	.w4(32'hbb34e98c),
	.w5(32'h3b0e8e6a),
	.w6(32'hbb2616d3),
	.w7(32'hbb6109eb),
	.w8(32'h3a248c2e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa95dda),
	.w1(32'h3ae79611),
	.w2(32'h3ac876a4),
	.w3(32'h3af1519b),
	.w4(32'h3b2e6201),
	.w5(32'hbbb121cf),
	.w6(32'h3b64df2a),
	.w7(32'h3b045588),
	.w8(32'hbb4e75e3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c025a),
	.w1(32'hbada763c),
	.w2(32'h3adc98d8),
	.w3(32'hbaad73a0),
	.w4(32'hba938b04),
	.w5(32'h3812ed90),
	.w6(32'h3a21f4ba),
	.w7(32'h3b45a6ee),
	.w8(32'h3a4f7b29),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9b7d0),
	.w1(32'hba55cdea),
	.w2(32'h3b1872ae),
	.w3(32'hba55f369),
	.w4(32'hba038a50),
	.w5(32'h3b8004af),
	.w6(32'hbb131729),
	.w7(32'hb9a0a8f9),
	.w8(32'h3ac94b56),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a832d),
	.w1(32'hbb25823a),
	.w2(32'hbb5ec3ac),
	.w3(32'h3aa8b7d5),
	.w4(32'hbb46c46c),
	.w5(32'hbb169de4),
	.w6(32'hba3874f4),
	.w7(32'hbb94d8e3),
	.w8(32'hbaafccb0),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbcde5),
	.w1(32'hbb3c3169),
	.w2(32'hbb03fee5),
	.w3(32'hbb003c03),
	.w4(32'hbae051e4),
	.w5(32'hbb90fa71),
	.w6(32'hb93ecb8a),
	.w7(32'hbb1a915b),
	.w8(32'hbb3f9c77),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ad406),
	.w1(32'hbae7b55a),
	.w2(32'hbb1c9e4c),
	.w3(32'hbb510876),
	.w4(32'hba60e8fc),
	.w5(32'hbba1694f),
	.w6(32'hbb308c9b),
	.w7(32'h3998244e),
	.w8(32'hbc36e4be),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb899e4f),
	.w1(32'h3c07f19f),
	.w2(32'h3c7d6bf6),
	.w3(32'h3ac3ea94),
	.w4(32'h3c06ae9c),
	.w5(32'hbbd4a860),
	.w6(32'hbaff5b8d),
	.w7(32'h3c3952c7),
	.w8(32'hbb472824),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0158ee),
	.w1(32'h3864a5c6),
	.w2(32'hb8bc059f),
	.w3(32'hbbc94fc0),
	.w4(32'hbaf0f0bb),
	.w5(32'h3abffdd3),
	.w6(32'hbb696f49),
	.w7(32'h3a4a3226),
	.w8(32'h3a4e5488),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74a255),
	.w1(32'hba6c86cd),
	.w2(32'hba632a18),
	.w3(32'hbb15f173),
	.w4(32'hbb8b5471),
	.w5(32'h3b42db08),
	.w6(32'h3a877d25),
	.w7(32'h3a62bf0c),
	.w8(32'h3b4391b4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00120e),
	.w1(32'hbb858d5c),
	.w2(32'hbb8f0d71),
	.w3(32'hbac4bfe3),
	.w4(32'hbb9c9136),
	.w5(32'h3a6fc21a),
	.w6(32'hbb867076),
	.w7(32'hbbcef3ad),
	.w8(32'h3b0197fd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8db964),
	.w1(32'hbb622c72),
	.w2(32'hbb92a1be),
	.w3(32'hba71e512),
	.w4(32'hbb3a3ce5),
	.w5(32'hbaa89c02),
	.w6(32'h3ad8f23b),
	.w7(32'hbb0f1d36),
	.w8(32'hb9da7274),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0690c9),
	.w1(32'hbba87551),
	.w2(32'hbb345806),
	.w3(32'hbb78ed58),
	.w4(32'hbb6a6594),
	.w5(32'hbb7e5936),
	.w6(32'hbbbf594e),
	.w7(32'hbb99efd0),
	.w8(32'hbb418f8c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac58ae8),
	.w1(32'h3c0673f3),
	.w2(32'h3c171dfa),
	.w3(32'h3ba583b6),
	.w4(32'h3c0c2408),
	.w5(32'hbbada11b),
	.w6(32'h3c38f839),
	.w7(32'h3c14598a),
	.w8(32'hbbecbe0b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbb371),
	.w1(32'hbb8e7189),
	.w2(32'h3b90dbb6),
	.w3(32'hbb93cd9a),
	.w4(32'h3a3c1d95),
	.w5(32'h3b369d06),
	.w6(32'hbc1fc0a7),
	.w7(32'h3afb65b1),
	.w8(32'h39a61cbd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393aa2d7),
	.w1(32'h3c8d292d),
	.w2(32'h3b848bf4),
	.w3(32'h3c74939f),
	.w4(32'h3bac25f9),
	.w5(32'hba70844c),
	.w6(32'h3ccb6877),
	.w7(32'h3c185d73),
	.w8(32'hbaa40244),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba303c7c),
	.w1(32'h3bb942a5),
	.w2(32'h3b960c26),
	.w3(32'h3a9a9d1e),
	.w4(32'hba8f3013),
	.w5(32'h3acac5b5),
	.w6(32'h3b3f8424),
	.w7(32'hb8f1844d),
	.w8(32'h3acbd940),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b7567),
	.w1(32'h3a7e7b45),
	.w2(32'hbb2d3244),
	.w3(32'h3ad0519a),
	.w4(32'hb9ac704a),
	.w5(32'hbb168948),
	.w6(32'h3b0ee734),
	.w7(32'hbab25adf),
	.w8(32'hbad67967),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf27495),
	.w1(32'h3a897b8a),
	.w2(32'hba996a50),
	.w3(32'h3b130ef2),
	.w4(32'hba043137),
	.w5(32'hb926ac8d),
	.w6(32'h3b1ada60),
	.w7(32'hbaa1b173),
	.w8(32'h3b615b38),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2ba8c),
	.w1(32'hbad9a904),
	.w2(32'hbb17f4db),
	.w3(32'hbb3885f5),
	.w4(32'hbbd2c050),
	.w5(32'hbb816d18),
	.w6(32'hb837edf7),
	.w7(32'hbb9f4b61),
	.w8(32'hbb6e7a6a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb188719),
	.w1(32'h3a1eb711),
	.w2(32'h3a92e285),
	.w3(32'hbb0b5101),
	.w4(32'h3b424dfb),
	.w5(32'h3ab9e47e),
	.w6(32'hba485bb3),
	.w7(32'h3ba773b5),
	.w8(32'hbabb8e88),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac060e4),
	.w1(32'h3bbfc3b3),
	.w2(32'hbabf8e24),
	.w3(32'h3a5adbd8),
	.w4(32'h3b3dec32),
	.w5(32'h39fb6cf5),
	.w6(32'h3bc33a38),
	.w7(32'h3b04cbbc),
	.w8(32'h3a97edf4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22f771),
	.w1(32'h3a8f291c),
	.w2(32'h3a397165),
	.w3(32'h39f27f52),
	.w4(32'h39982100),
	.w5(32'hba033297),
	.w6(32'h3afc133f),
	.w7(32'h3a4e08bc),
	.w8(32'h398129df),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9b587),
	.w1(32'hbb371f9c),
	.w2(32'h3a83a8da),
	.w3(32'h3b597e37),
	.w4(32'hba8782c6),
	.w5(32'hb80f5622),
	.w6(32'h39d6a5ad),
	.w7(32'h3a20e417),
	.w8(32'h392378ec),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c87640),
	.w1(32'h3a919b39),
	.w2(32'h3a23e5b2),
	.w3(32'h3acb6250),
	.w4(32'h3aace4e7),
	.w5(32'hba52d2a1),
	.w6(32'h38b1a44b),
	.w7(32'h3a5ce0d7),
	.w8(32'hb96865d2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92c840),
	.w1(32'hb99e9560),
	.w2(32'h3a2a7820),
	.w3(32'hba66ddff),
	.w4(32'hb97d1f2a),
	.w5(32'h3a75a012),
	.w6(32'h3ab6c702),
	.w7(32'hb8944630),
	.w8(32'h3a3e9087),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa65738),
	.w1(32'h3a26f4d9),
	.w2(32'h3a856096),
	.w3(32'hb95aa7b3),
	.w4(32'h390acf4c),
	.w5(32'hbad2231a),
	.w6(32'hb9adc7f3),
	.w7(32'hba74dc28),
	.w8(32'hbaa7218f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27d94d),
	.w1(32'hbb7f1169),
	.w2(32'hbb2bd7d8),
	.w3(32'hba5a5fa0),
	.w4(32'hbb14583e),
	.w5(32'hba685f9f),
	.w6(32'h3a1a6fe7),
	.w7(32'hbad37ba6),
	.w8(32'h3a7cca69),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba17ac),
	.w1(32'h3a6f70eb),
	.w2(32'h3ac088d0),
	.w3(32'hbb6fa85b),
	.w4(32'hbb1be7fb),
	.w5(32'h39b84bdf),
	.w6(32'h3b21f05d),
	.w7(32'h39bdbe2a),
	.w8(32'h375f3afb),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67dc44),
	.w1(32'hbb8ff540),
	.w2(32'hb9ffa983),
	.w3(32'h3b9258f4),
	.w4(32'h3b24b42f),
	.w5(32'hbb0ff949),
	.w6(32'hb981b9c0),
	.w7(32'h3b2afeaf),
	.w8(32'hba35672b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c60765),
	.w1(32'hbb459c66),
	.w2(32'h3af9ca12),
	.w3(32'hbb875920),
	.w4(32'hba99fe4c),
	.w5(32'hb8971e0a),
	.w6(32'hbaf42330),
	.w7(32'h38eea128),
	.w8(32'h3a02e71c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842e814),
	.w1(32'hba8bce56),
	.w2(32'hba4096fc),
	.w3(32'hb9e23e26),
	.w4(32'hba3cbef3),
	.w5(32'hba4e8324),
	.w6(32'h3a137121),
	.w7(32'hb8d7ef8f),
	.w8(32'h39def2ad),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6af55),
	.w1(32'h39f850d0),
	.w2(32'h39553348),
	.w3(32'hba79ba45),
	.w4(32'hba9f08e6),
	.w5(32'hb9f2ec07),
	.w6(32'h3ac38345),
	.w7(32'h3a25d4ec),
	.w8(32'h3a8673b4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b915e8),
	.w1(32'hb9964581),
	.w2(32'hbadc7e5f),
	.w3(32'h3830ae11),
	.w4(32'h38f1be0c),
	.w5(32'hb902f984),
	.w6(32'h39c6cd2d),
	.w7(32'hb9c1bdaf),
	.w8(32'hba024957),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b9d73),
	.w1(32'h3a2a92fd),
	.w2(32'h3a09f4e0),
	.w3(32'h39037e6f),
	.w4(32'h3a119800),
	.w5(32'hbad203d4),
	.w6(32'h39bfbdca),
	.w7(32'hb8a5a48c),
	.w8(32'hba6760f8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba841468),
	.w1(32'hba40ad61),
	.w2(32'h3a471b57),
	.w3(32'hbaa89155),
	.w4(32'h394b59a8),
	.w5(32'h399641a3),
	.w6(32'hba12a7f0),
	.w7(32'h3984e22c),
	.w8(32'hb91e1be3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa53716),
	.w1(32'h3a83fd5b),
	.w2(32'h3a14b87a),
	.w3(32'hb9fc7ab6),
	.w4(32'h3a7fdae9),
	.w5(32'h3a72f535),
	.w6(32'h392116f3),
	.w7(32'h3a87db2a),
	.w8(32'hba3b7869),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba386b64),
	.w1(32'hba75a4de),
	.w2(32'h3a1fdd1c),
	.w3(32'h3a3cdb38),
	.w4(32'h3ab3a9e6),
	.w5(32'h399b0dd2),
	.w6(32'hb938851f),
	.w7(32'h3a4d3dd9),
	.w8(32'hba4fe5bb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb148df0),
	.w1(32'hbb5ccb7e),
	.w2(32'hb994c8f2),
	.w3(32'hba37b4b5),
	.w4(32'hba8a2a23),
	.w5(32'hba90860e),
	.w6(32'hb9e457b9),
	.w7(32'hba358457),
	.w8(32'hbaa40baa),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba819809),
	.w1(32'hba97f703),
	.w2(32'hb9ad5963),
	.w3(32'hbafd2828),
	.w4(32'h3a2a4369),
	.w5(32'h3a6869d1),
	.w6(32'hb9fbce37),
	.w7(32'h39a77593),
	.w8(32'h3acb2fb4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9edf7b),
	.w1(32'h3aa6a389),
	.w2(32'h3aaae277),
	.w3(32'h3989ac4d),
	.w4(32'h3a9a49e7),
	.w5(32'h3a59fc86),
	.w6(32'h3a373e05),
	.w7(32'h3aa9d324),
	.w8(32'h3b169008),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0350f9),
	.w1(32'h3aa059c0),
	.w2(32'h391f9c90),
	.w3(32'h3aa7aad7),
	.w4(32'hbab53e1f),
	.w5(32'hb7b3ff61),
	.w6(32'h3b56f8ba),
	.w7(32'h3b0b92ee),
	.w8(32'h3b0181c6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac613c1),
	.w1(32'h39fad581),
	.w2(32'hb922c832),
	.w3(32'hba753c51),
	.w4(32'hba605b7f),
	.w5(32'hbac3fc21),
	.w6(32'h3a55bd01),
	.w7(32'h39c44bac),
	.w8(32'hb9f5667e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5f84d),
	.w1(32'hba6d958c),
	.w2(32'hbaa98a4b),
	.w3(32'h3b079a07),
	.w4(32'hbaa09bdf),
	.w5(32'hbaaf6b6c),
	.w6(32'h3b62cc7f),
	.w7(32'h3a1dca50),
	.w8(32'hbaa2108c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a23ad),
	.w1(32'hbae2c93f),
	.w2(32'hbabdb93d),
	.w3(32'hbb316540),
	.w4(32'hb978ffed),
	.w5(32'h3aa3a771),
	.w6(32'hbaff36f4),
	.w7(32'hb9a229a0),
	.w8(32'h3ade0061),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76b69e),
	.w1(32'h3a0becba),
	.w2(32'h3a049ab8),
	.w3(32'hba61c3df),
	.w4(32'hb8a9e568),
	.w5(32'h3a0a96ca),
	.w6(32'h3b12d516),
	.w7(32'hb87e63ee),
	.w8(32'hba11b2c2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba5044),
	.w1(32'hb9a53973),
	.w2(32'h3a34babb),
	.w3(32'hbaa65222),
	.w4(32'h3aae3fe3),
	.w5(32'hbafac705),
	.w6(32'h3aa43773),
	.w7(32'h39a8e672),
	.w8(32'hba1b0ba3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba866bb6),
	.w1(32'hb7d4c697),
	.w2(32'hbaa32289),
	.w3(32'hb888009a),
	.w4(32'h3a741263),
	.w5(32'h3a311dd6),
	.w6(32'hbabaa712),
	.w7(32'hba00c0df),
	.w8(32'h3aaab68b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39819e38),
	.w1(32'h3a6623f6),
	.w2(32'h3a9d6582),
	.w3(32'hba9266bd),
	.w4(32'h3ac05b98),
	.w5(32'hb99f61ac),
	.w6(32'h3ae3a907),
	.w7(32'h3a8b95c5),
	.w8(32'h39cc88d9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b8daa),
	.w1(32'h39704a45),
	.w2(32'h3a1047dd),
	.w3(32'h390a53eb),
	.w4(32'hb9d614f0),
	.w5(32'hb9162d94),
	.w6(32'h3ade5a42),
	.w7(32'h3ae982e6),
	.w8(32'h3a9a6d99),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b7c16e),
	.w1(32'h3a372297),
	.w2(32'hbae5209c),
	.w3(32'hbadbb54b),
	.w4(32'h39ae824e),
	.w5(32'h3a122e16),
	.w6(32'hba0b243b),
	.w7(32'hba7116da),
	.w8(32'hba842a5c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0075b2),
	.w1(32'hbb42cf40),
	.w2(32'hbaa99c13),
	.w3(32'h3a3e32de),
	.w4(32'hbad50922),
	.w5(32'hba7e1b5e),
	.w6(32'hb99f5ab6),
	.w7(32'hba14553e),
	.w8(32'hba83fc1d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule