module layer_10_featuremap_429(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89df8a),
	.w1(32'hbb3ebdc1),
	.w2(32'hbb912ac5),
	.w3(32'hbb120ea1),
	.w4(32'h3b126b80),
	.w5(32'h3b88662e),
	.w6(32'hbc318754),
	.w7(32'hb9fa01e5),
	.w8(32'h3b596bf9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7c11c),
	.w1(32'hbb4b16cb),
	.w2(32'hbc07ce5c),
	.w3(32'h3c1128fe),
	.w4(32'hbba8c261),
	.w5(32'hba7cb21b),
	.w6(32'h3c19926c),
	.w7(32'hbc121fc5),
	.w8(32'hbc251f49),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a68c6),
	.w1(32'hbc3129e7),
	.w2(32'h3c5c0b1f),
	.w3(32'hbc351b21),
	.w4(32'h3cefa704),
	.w5(32'hbc2618db),
	.w6(32'hbc219d82),
	.w7(32'h3b12c60b),
	.w8(32'h3aefe608),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199823),
	.w1(32'hbb665086),
	.w2(32'h3c66f351),
	.w3(32'hbb4242fe),
	.w4(32'h3c8d6153),
	.w5(32'h3c96526f),
	.w6(32'hbb9397e0),
	.w7(32'h3bec6b1b),
	.w8(32'hbc491427),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb184b08),
	.w1(32'h3b35bbbf),
	.w2(32'hbc12ab70),
	.w3(32'hbb81897f),
	.w4(32'h3bdd1181),
	.w5(32'hbc2fcd5b),
	.w6(32'h3cb0d74a),
	.w7(32'hbb42763b),
	.w8(32'h3bf0d13f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e5fb4),
	.w1(32'h3a24d011),
	.w2(32'hbb6b6435),
	.w3(32'hba569a65),
	.w4(32'hbb68695a),
	.w5(32'h3bd4944a),
	.w6(32'h3ac3e81e),
	.w7(32'h3b177fc0),
	.w8(32'hbbbfbca4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec913),
	.w1(32'hbbc11f6e),
	.w2(32'hb9938040),
	.w3(32'hbc094a7d),
	.w4(32'hbc6c630f),
	.w5(32'h3ad30ad6),
	.w6(32'hba7de61d),
	.w7(32'hbb97848c),
	.w8(32'h39b9afe1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91e109),
	.w1(32'hbc2dd6a6),
	.w2(32'h3bc5d8ef),
	.w3(32'hbc1eae59),
	.w4(32'h3c3ae119),
	.w5(32'hbbd56120),
	.w6(32'hbb4ccf36),
	.w7(32'h3c424b02),
	.w8(32'h3bf8ff6f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23d08b),
	.w1(32'hbc2fbeda),
	.w2(32'h3c915dad),
	.w3(32'hbc60925b),
	.w4(32'hbc3cb1d4),
	.w5(32'h3c58f764),
	.w6(32'hbb2aacf1),
	.w7(32'h38d60dda),
	.w8(32'hbcf30408),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fe7b2),
	.w1(32'h3b9d0769),
	.w2(32'h3b918885),
	.w3(32'hbc110b00),
	.w4(32'hbad86bee),
	.w5(32'h3b447f36),
	.w6(32'h3c6153b0),
	.w7(32'hbc108983),
	.w8(32'h3ac76d01),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae65ba),
	.w1(32'hbb023d47),
	.w2(32'h3a2705a6),
	.w3(32'hbbbae1cc),
	.w4(32'hbbd6ac23),
	.w5(32'hbc74e06c),
	.w6(32'hba542585),
	.w7(32'hbc536e49),
	.w8(32'hbc165142),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1475c2),
	.w1(32'hbb1aeb5f),
	.w2(32'h3aa3b6e5),
	.w3(32'hbb959135),
	.w4(32'hbb9468c9),
	.w5(32'hbae3f369),
	.w6(32'hbc8f40d7),
	.w7(32'hba68ca1d),
	.w8(32'h3bd301b4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd79eac),
	.w1(32'hbb08fe15),
	.w2(32'h3c28c9eb),
	.w3(32'hbb0f5a37),
	.w4(32'h3b4349b8),
	.w5(32'h3cbc7445),
	.w6(32'h3b626f82),
	.w7(32'h3bc58bb6),
	.w8(32'hbb8fed57),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b287bf9),
	.w1(32'h3c3e0cc5),
	.w2(32'hbbc8a9ae),
	.w3(32'hbb65c4e1),
	.w4(32'hbc1508e5),
	.w5(32'h3adb1842),
	.w6(32'h3beec938),
	.w7(32'hbbc7bd51),
	.w8(32'hbb083f68),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc369874),
	.w1(32'h3bd22ef3),
	.w2(32'h3c0fb9ca),
	.w3(32'h3bbdc8ac),
	.w4(32'h3c05407e),
	.w5(32'hbca4e5a2),
	.w6(32'h3aa06811),
	.w7(32'hbb8eaddd),
	.w8(32'h3c85dcbb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bf85c),
	.w1(32'hbb822a76),
	.w2(32'h3b278892),
	.w3(32'h3c22e3a0),
	.w4(32'hbb47e466),
	.w5(32'hbbad039b),
	.w6(32'hbc0a0813),
	.w7(32'hba57f985),
	.w8(32'h3b182c9c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f1140),
	.w1(32'h3ac5d222),
	.w2(32'hbba6d991),
	.w3(32'hbb62a502),
	.w4(32'h3b57f195),
	.w5(32'hbae8672f),
	.w6(32'hbb799cdc),
	.w7(32'h3bc69431),
	.w8(32'h3a64d76f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e13fd),
	.w1(32'hbbc17d83),
	.w2(32'h3b4555dd),
	.w3(32'hbc7d58a3),
	.w4(32'hbb3615a0),
	.w5(32'h3b892583),
	.w6(32'hbbca139e),
	.w7(32'h3bd563b4),
	.w8(32'h3b284ac7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997eff0),
	.w1(32'hbb3c04e5),
	.w2(32'h3c5121c8),
	.w3(32'hbb4e782f),
	.w4(32'hbb7ad3a3),
	.w5(32'h3b94cf68),
	.w6(32'hbb55ced9),
	.w7(32'h3ba89a15),
	.w8(32'h3bbb4e44),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c2dd0),
	.w1(32'h3a776633),
	.w2(32'hbaf5d3d2),
	.w3(32'h3abd9c6a),
	.w4(32'hbc2676e2),
	.w5(32'h3b0d944e),
	.w6(32'h3b96b356),
	.w7(32'hbb8a9c61),
	.w8(32'hbbbf733a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1941),
	.w1(32'hb9b8e706),
	.w2(32'h3bc79916),
	.w3(32'hbc14b7c6),
	.w4(32'hbadc1022),
	.w5(32'h3bb0db99),
	.w6(32'hbb237eba),
	.w7(32'h39917169),
	.w8(32'hbba3c0a3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc967e1),
	.w1(32'h3b88d83e),
	.w2(32'hbb6e0477),
	.w3(32'hbada7c7c),
	.w4(32'h3c2ea59c),
	.w5(32'h3b1f8788),
	.w6(32'h3b9f3b4c),
	.w7(32'h3c0a1a86),
	.w8(32'h3a79d9f4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9afade),
	.w1(32'hbc0e63dc),
	.w2(32'h39f74016),
	.w3(32'hbc24ecc5),
	.w4(32'h3b545315),
	.w5(32'h3beefa06),
	.w6(32'hba89c59e),
	.w7(32'h3b87d761),
	.w8(32'h3b9cf2b2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aa991),
	.w1(32'h3bafc4d1),
	.w2(32'h3c73b704),
	.w3(32'hbba2f11f),
	.w4(32'hbb201470),
	.w5(32'h3b9f497b),
	.w6(32'hbb8f6665),
	.w7(32'hbc26513d),
	.w8(32'h3bc2ba5a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3812b5),
	.w1(32'hba8b507c),
	.w2(32'h3b936699),
	.w3(32'h39eca678),
	.w4(32'hba973eb6),
	.w5(32'h39a97933),
	.w6(32'h3b55d431),
	.w7(32'hbc0191c4),
	.w8(32'hbbce8ade),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1067e),
	.w1(32'h3b8f562e),
	.w2(32'h3bf72e7a),
	.w3(32'h3b223308),
	.w4(32'h3bbf7561),
	.w5(32'h3a9f3a9e),
	.w6(32'h3ab46582),
	.w7(32'h389a9dc1),
	.w8(32'hbaea7a56),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3931ab4a),
	.w1(32'h3b9f25c6),
	.w2(32'h3bec0363),
	.w3(32'h3b6d2526),
	.w4(32'h3a0f5568),
	.w5(32'hbbf1cfc6),
	.w6(32'hb901d901),
	.w7(32'h3a84a38a),
	.w8(32'hbba650d3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaec91b),
	.w1(32'hbbd1a664),
	.w2(32'hbb6cc61a),
	.w3(32'hbc3f106b),
	.w4(32'hbbdd50b6),
	.w5(32'hbbbe9e6c),
	.w6(32'h3ad9414b),
	.w7(32'hbbb2d540),
	.w8(32'hbbc408f5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd88a05),
	.w1(32'hbbcbc474),
	.w2(32'h390903a2),
	.w3(32'hbb9f9c55),
	.w4(32'hba06ae9f),
	.w5(32'hbbf69388),
	.w6(32'hbbf26919),
	.w7(32'hbb33a209),
	.w8(32'hbb71f73e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b376972),
	.w1(32'h39034297),
	.w2(32'h3c65854d),
	.w3(32'h3bbb0b39),
	.w4(32'hbb8c82e8),
	.w5(32'h3c64cda9),
	.w6(32'h3a4c3f2e),
	.w7(32'hbbab1671),
	.w8(32'hbb1ab017),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01d0db),
	.w1(32'h3c039a5f),
	.w2(32'hbbb95f4f),
	.w3(32'h3b1c178b),
	.w4(32'hbb3efd78),
	.w5(32'hbb764b94),
	.w6(32'h3b8d10cf),
	.w7(32'h3b6255c1),
	.w8(32'h3b44dd9b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f60f7),
	.w1(32'hbabca56b),
	.w2(32'hbc5cf689),
	.w3(32'h3b75da12),
	.w4(32'h3c0d78c8),
	.w5(32'hbc927994),
	.w6(32'h3b0b97ca),
	.w7(32'h3c016912),
	.w8(32'h3c1ff497),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3da2ae),
	.w1(32'h3c043796),
	.w2(32'h3bbf280b),
	.w3(32'h3b72d0e2),
	.w4(32'hbc60dbd0),
	.w5(32'h3c849c59),
	.w6(32'hbc585ef5),
	.w7(32'hbb0c951a),
	.w8(32'hbb1f6059),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3e1ce),
	.w1(32'h3c0d3b9a),
	.w2(32'h3b1f2140),
	.w3(32'h3bc88ce7),
	.w4(32'hbb3c1059),
	.w5(32'h3c846260),
	.w6(32'hbb9e4bd4),
	.w7(32'h3bdbc449),
	.w8(32'h3c9a2614),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bda37),
	.w1(32'h3c45b61d),
	.w2(32'hbc28fff4),
	.w3(32'h3cae0492),
	.w4(32'hbce64f26),
	.w5(32'h3ce7f30e),
	.w6(32'h3a96c188),
	.w7(32'hbc325873),
	.w8(32'hbb5d26df),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34054b),
	.w1(32'hbc07dfd8),
	.w2(32'h3c90cd9c),
	.w3(32'h3cbd9f80),
	.w4(32'h3b19ef64),
	.w5(32'h3cb622a8),
	.w6(32'hbb269f64),
	.w7(32'h3b069304),
	.w8(32'hbcab3b39),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17665a),
	.w1(32'hbc3fe5c7),
	.w2(32'hba817769),
	.w3(32'hbc891a90),
	.w4(32'hbc29dd0d),
	.w5(32'hbbcf1456),
	.w6(32'h3bb51bb9),
	.w7(32'hb9ff8db3),
	.w8(32'hbc1b5ac3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18f8e6),
	.w1(32'h3c354f3a),
	.w2(32'h3a3f67aa),
	.w3(32'hba8613b2),
	.w4(32'hbaa932bc),
	.w5(32'h3c01599a),
	.w6(32'hbadb8a8d),
	.w7(32'hbb63eb2f),
	.w8(32'hbc9f269d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7297c7),
	.w1(32'h3bd66b09),
	.w2(32'hbc3f4d35),
	.w3(32'h3b5486fe),
	.w4(32'h3c162698),
	.w5(32'hbcd5a5bf),
	.w6(32'h3ba6cbb1),
	.w7(32'hbbd7c084),
	.w8(32'h3ca129e2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6379f0),
	.w1(32'h3b1e2a72),
	.w2(32'hbb9ee842),
	.w3(32'h3c939f26),
	.w4(32'hbbed9031),
	.w5(32'h3c2e3485),
	.w6(32'h3aa059be),
	.w7(32'hbae2cab7),
	.w8(32'hbca1625e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57b3b4),
	.w1(32'h3caede2f),
	.w2(32'hbc85d43e),
	.w3(32'hbb92e57f),
	.w4(32'h3c222afd),
	.w5(32'hbb2eef07),
	.w6(32'h3b5ad2da),
	.w7(32'hbca860f1),
	.w8(32'h3cec8970),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abab198),
	.w1(32'h3bb7afdf),
	.w2(32'hbaa0dda2),
	.w3(32'h3c823999),
	.w4(32'h3a1cf422),
	.w5(32'hbc0688ee),
	.w6(32'hbb17775d),
	.w7(32'hbb437d55),
	.w8(32'h3c91bf0c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3325ad),
	.w1(32'hbac49920),
	.w2(32'h3c293f89),
	.w3(32'h3c3bb23c),
	.w4(32'h3ba4a97c),
	.w5(32'h3caa3a56),
	.w6(32'hbbe78510),
	.w7(32'h3ac3bd9b),
	.w8(32'hbc463b51),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95897a),
	.w1(32'h3ba89ba8),
	.w2(32'h3b5f02e7),
	.w3(32'hbb6d9adc),
	.w4(32'h3b9b1b54),
	.w5(32'h3be79472),
	.w6(32'h3ba7a22d),
	.w7(32'hba810789),
	.w8(32'h3c2272f2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc09e11),
	.w1(32'h3bc2d0ec),
	.w2(32'h3c3f4f7e),
	.w3(32'h3bd19f06),
	.w4(32'h3aa49bcd),
	.w5(32'hb9c9d5c1),
	.w6(32'h3bc780f9),
	.w7(32'h3a911a13),
	.w8(32'h3bd0ca57),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03558e),
	.w1(32'h3bb03881),
	.w2(32'h3c0f07fd),
	.w3(32'h3abd19cd),
	.w4(32'hbb22710d),
	.w5(32'h3abd3039),
	.w6(32'h3b0db0a9),
	.w7(32'hbb9c70eb),
	.w8(32'hbb0add5f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbdc1c),
	.w1(32'h3b40f62e),
	.w2(32'h3c20c387),
	.w3(32'hbba783d3),
	.w4(32'h3c2780a7),
	.w5(32'h3ae18033),
	.w6(32'hbaa30182),
	.w7(32'h3b104e62),
	.w8(32'h3bf87a39),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb535f8),
	.w1(32'hbbc01af2),
	.w2(32'hbab107a2),
	.w3(32'hbc30a286),
	.w4(32'hbb0376c8),
	.w5(32'hba7e52ff),
	.w6(32'h3b50fef7),
	.w7(32'hbac104d6),
	.w8(32'h3c65f24a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb864c5b),
	.w1(32'h3b7bb262),
	.w2(32'h3c83f902),
	.w3(32'hbaf65695),
	.w4(32'hbb996966),
	.w5(32'h3c2f5501),
	.w6(32'hbaceeb80),
	.w7(32'hbb4e49fc),
	.w8(32'hbc81b8c4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46e564),
	.w1(32'hba577334),
	.w2(32'hbca46c27),
	.w3(32'hbbf7e882),
	.w4(32'h3ad91346),
	.w5(32'hbc90e930),
	.w6(32'h3c21f90b),
	.w7(32'h3aa5cbd6),
	.w8(32'h3cba62a2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca63fca),
	.w1(32'h3a6e83af),
	.w2(32'h3a839ee5),
	.w3(32'h3c48cd4d),
	.w4(32'h3b294d45),
	.w5(32'h3ba6d547),
	.w6(32'hbc5a1ca5),
	.w7(32'hb8f660b0),
	.w8(32'h3b7e3a5c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bc92f),
	.w1(32'h3b08bacc),
	.w2(32'h3b034b2c),
	.w3(32'hb88b1b6a),
	.w4(32'hbb1a4c68),
	.w5(32'hbb7a64a7),
	.w6(32'hbac10c19),
	.w7(32'hbb08f8f1),
	.w8(32'h3ad51ffe),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1c44d),
	.w1(32'h3b7575ca),
	.w2(32'hbbecacce),
	.w3(32'hbbe33422),
	.w4(32'hbc408c34),
	.w5(32'h3c33241f),
	.w6(32'hbafb2ec5),
	.w7(32'h3a600a56),
	.w8(32'h3bbb95a3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75a7fb),
	.w1(32'h3bf65077),
	.w2(32'h39938d14),
	.w3(32'hbaabe6c2),
	.w4(32'hbceb909b),
	.w5(32'h3d229274),
	.w6(32'hbc26c266),
	.w7(32'hbb854930),
	.w8(32'hbc5c6839),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc45681),
	.w1(32'h3afcec2e),
	.w2(32'hbc5ccb3d),
	.w3(32'h3c9eddac),
	.w4(32'hbbf2c7f5),
	.w5(32'hb9dbcfd2),
	.w6(32'h3b49bf90),
	.w7(32'hbc1aa47f),
	.w8(32'hbc89ef70),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b61a0),
	.w1(32'hbb76a93b),
	.w2(32'h3c8f9334),
	.w3(32'hbc2ad769),
	.w4(32'hbc89c664),
	.w5(32'h3d4d6684),
	.w6(32'hbb147318),
	.w7(32'h3b4374ff),
	.w8(32'hbd01591e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a161833),
	.w1(32'h3bac2adc),
	.w2(32'hbb8156ef),
	.w3(32'hb990403e),
	.w4(32'h3b80dd3e),
	.w5(32'h3b13660c),
	.w6(32'h3b4c021c),
	.w7(32'h3b937ef6),
	.w8(32'h3b9f4877),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b468cec),
	.w1(32'h39a44b4c),
	.w2(32'h3ba15492),
	.w3(32'h3b4ceb78),
	.w4(32'h39e7187d),
	.w5(32'hbaad5ebf),
	.w6(32'h3b4191be),
	.w7(32'hb9f31eba),
	.w8(32'hbb61f27b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2cf99),
	.w1(32'h3b006786),
	.w2(32'h3bcf94cb),
	.w3(32'hbb5c05d2),
	.w4(32'h3b90a75a),
	.w5(32'h3c178992),
	.w6(32'hbc05642b),
	.w7(32'h3a8de9df),
	.w8(32'h3b828c14),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c575ee),
	.w1(32'h3b140721),
	.w2(32'hba972409),
	.w3(32'h3a6bc735),
	.w4(32'hbc36fe68),
	.w5(32'hbba0f22b),
	.w6(32'hbb05cf5e),
	.w7(32'hbb4258fe),
	.w8(32'hbc3fd22e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9c9f1),
	.w1(32'h3b85b557),
	.w2(32'h3bec1c1e),
	.w3(32'hbc30a565),
	.w4(32'h3bf2bca3),
	.w5(32'h3bdaae76),
	.w6(32'hbbcac10a),
	.w7(32'h3b54fa5b),
	.w8(32'h3bf368be),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b431842),
	.w1(32'hba0d69ef),
	.w2(32'hbba183f5),
	.w3(32'hbb295ba7),
	.w4(32'h3c2ef59c),
	.w5(32'hbc75b570),
	.w6(32'h3aaa1f21),
	.w7(32'h3b03496a),
	.w8(32'h3cb79e23),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb33370),
	.w1(32'h3a3799b5),
	.w2(32'hbb8f18b9),
	.w3(32'h3c133016),
	.w4(32'h3a8528f2),
	.w5(32'h3bdbbf4d),
	.w6(32'hbc5110a1),
	.w7(32'hbc0dd995),
	.w8(32'hbc6c0c1d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2e560),
	.w1(32'h3c101aad),
	.w2(32'hb96ffc3c),
	.w3(32'hba8f933b),
	.w4(32'h3bcee712),
	.w5(32'h3b63154f),
	.w6(32'h3b04bbd1),
	.w7(32'h3b3f4a52),
	.w8(32'h3b6e7cf2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a7806),
	.w1(32'h38cc6c6a),
	.w2(32'h3b080dbd),
	.w3(32'h3b0ed573),
	.w4(32'h3ac069e1),
	.w5(32'h3c14c65c),
	.w6(32'h3ba122ef),
	.w7(32'h3bd5f311),
	.w8(32'hbb2cf426),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39010593),
	.w1(32'h37e0a5b1),
	.w2(32'hbb062324),
	.w3(32'hbaa112de),
	.w4(32'hbb975fde),
	.w5(32'hbc4cd34b),
	.w6(32'h3c3e21cc),
	.w7(32'hbba9ad9b),
	.w8(32'h3bd5457a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd98f44),
	.w1(32'h3af4e5ad),
	.w2(32'h3bf67c74),
	.w3(32'h3a98663c),
	.w4(32'h3a05a7b9),
	.w5(32'hbac71a0a),
	.w6(32'hbb9797ff),
	.w7(32'hbaeb0bd7),
	.w8(32'h3b8ae529),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69bb9c),
	.w1(32'hbc5af7a6),
	.w2(32'h3b283f1e),
	.w3(32'hbba31649),
	.w4(32'hbc764494),
	.w5(32'h3c1e657c),
	.w6(32'hbbc01786),
	.w7(32'hbc047158),
	.w8(32'hbc104e25),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91cac1),
	.w1(32'hb80def5f),
	.w2(32'hba838630),
	.w3(32'hbaf75fb0),
	.w4(32'h3ad49f85),
	.w5(32'hb992a9f6),
	.w6(32'hbbcfe974),
	.w7(32'hbb87a4d7),
	.w8(32'h3ad7e87a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8af2f3),
	.w1(32'h3b8d6e96),
	.w2(32'h3ba535aa),
	.w3(32'h3c16377f),
	.w4(32'hbb4ad538),
	.w5(32'hb9ac50bf),
	.w6(32'hb8c133d2),
	.w7(32'hbb92b4b3),
	.w8(32'hbbee3920),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbe336),
	.w1(32'hbba5fc1a),
	.w2(32'h3b937f9d),
	.w3(32'hbc35b049),
	.w4(32'hbb7decc8),
	.w5(32'h3c2a3fd3),
	.w6(32'hbb76a2cb),
	.w7(32'hbc02e444),
	.w8(32'h3b47d510),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaef667),
	.w1(32'h3c3d3792),
	.w2(32'h3bb472a6),
	.w3(32'hbbbc26fd),
	.w4(32'h3c1f6d50),
	.w5(32'hba8bf7ac),
	.w6(32'hbc4211dd),
	.w7(32'h3be8e5d0),
	.w8(32'hbac81a1e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c79c7),
	.w1(32'h39bb8691),
	.w2(32'h3c72a11c),
	.w3(32'h3b801c4e),
	.w4(32'h3bb4b492),
	.w5(32'h3c255ead),
	.w6(32'h3b66cb30),
	.w7(32'h3b1683fd),
	.w8(32'h3b1e6284),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20771b),
	.w1(32'h3a8b1beb),
	.w2(32'hbb624101),
	.w3(32'h3ba20f72),
	.w4(32'h3a512232),
	.w5(32'hbb85a1ff),
	.w6(32'h3c134201),
	.w7(32'h3b1c7be7),
	.w8(32'hbb281cb6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393300d4),
	.w1(32'h3a91ad32),
	.w2(32'hbb9ce52d),
	.w3(32'h3abe527f),
	.w4(32'hbb8c2d82),
	.w5(32'hbc17f523),
	.w6(32'h3b4e3a4d),
	.w7(32'hbba47cb8),
	.w8(32'h3b864463),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc531619),
	.w1(32'hbb9a00a0),
	.w2(32'h3acf7313),
	.w3(32'hbbaea08a),
	.w4(32'hbb8c9c1d),
	.w5(32'hbb3fc7e8),
	.w6(32'h39d0b597),
	.w7(32'h3b099945),
	.w8(32'h393b734c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc428945),
	.w1(32'h3bc96e67),
	.w2(32'hbab41104),
	.w3(32'hbbf503e3),
	.w4(32'h3bac771c),
	.w5(32'hbb1461b0),
	.w6(32'hbbc960b2),
	.w7(32'h3c17538a),
	.w8(32'h3b3c5173),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada1b82),
	.w1(32'hbb5251b6),
	.w2(32'h3b29c27a),
	.w3(32'h399f2a08),
	.w4(32'hbbb0e61b),
	.w5(32'hbb6087b8),
	.w6(32'h3a11bb10),
	.w7(32'hbae09714),
	.w8(32'h3c4d30db),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba354dbd),
	.w1(32'h3bd2a314),
	.w2(32'h394f4240),
	.w3(32'hbbaa6662),
	.w4(32'h3b7f20ac),
	.w5(32'hbb8dca16),
	.w6(32'h3b87e682),
	.w7(32'h3b4e265d),
	.w8(32'h3ab99e80),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd90c0b),
	.w1(32'h3bfa3db6),
	.w2(32'h3b8c8e5b),
	.w3(32'hbb60850f),
	.w4(32'h3c38d57f),
	.w5(32'h3a9d4be1),
	.w6(32'hbb2f2e35),
	.w7(32'h3c307bc0),
	.w8(32'hbbc1ebe5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fca29),
	.w1(32'h3c80aae6),
	.w2(32'h3b9c54ad),
	.w3(32'h3c1e9d19),
	.w4(32'h3c5d8762),
	.w5(32'hbc155c41),
	.w6(32'h3b05e409),
	.w7(32'h3c311878),
	.w8(32'hbafaf121),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fa86f),
	.w1(32'hbc361e4f),
	.w2(32'h3b305751),
	.w3(32'hbbaea66b),
	.w4(32'hbbe69544),
	.w5(32'h3c2e47fb),
	.w6(32'hbbcb99db),
	.w7(32'hbb50e11a),
	.w8(32'h3c0cf303),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad9f4a),
	.w1(32'hbab3961a),
	.w2(32'h39a59726),
	.w3(32'h3a43bef6),
	.w4(32'hbb0b8cc5),
	.w5(32'h38340edc),
	.w6(32'hba6de47c),
	.w7(32'hb9f7ffaa),
	.w8(32'h3977eb2e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e33dc),
	.w1(32'h39f1fdad),
	.w2(32'hbba50ac5),
	.w3(32'hb94be00c),
	.w4(32'hbb192194),
	.w5(32'h3c8bb676),
	.w6(32'hb964f69e),
	.w7(32'hbb56531b),
	.w8(32'h3c1f2cc1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0233b6),
	.w1(32'hbbb7257c),
	.w2(32'h3acdd66a),
	.w3(32'h3c5d268b),
	.w4(32'hbbb81c4f),
	.w5(32'h3b90aa15),
	.w6(32'hbbfa0752),
	.w7(32'hbbc4da0f),
	.w8(32'hb941a825),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b945e06),
	.w1(32'hbc65d0a6),
	.w2(32'h3c9ca11f),
	.w3(32'hba0d7a9c),
	.w4(32'hbc3dddeb),
	.w5(32'h3d51b0fe),
	.w6(32'h3a6930b0),
	.w7(32'h3becb5dc),
	.w8(32'hbaf33bd7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fc592),
	.w1(32'h3c8f8416),
	.w2(32'h3b0691f9),
	.w3(32'h3bc60386),
	.w4(32'h3c6080da),
	.w5(32'hbbd96ff2),
	.w6(32'hbaee9b4b),
	.w7(32'h3a6cee0e),
	.w8(32'hbc3fae2b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c1ef9),
	.w1(32'h3b292f45),
	.w2(32'h3ab38a4c),
	.w3(32'h3b981266),
	.w4(32'hbad12f70),
	.w5(32'h3b512d4f),
	.w6(32'h39f1cd76),
	.w7(32'hbbceb370),
	.w8(32'hb8ecd4c3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2528f0),
	.w1(32'h3c23603f),
	.w2(32'h3aa3db7c),
	.w3(32'h38eb9dd2),
	.w4(32'h3b9d09f7),
	.w5(32'hbc319502),
	.w6(32'hbae5956f),
	.w7(32'hbb8f74a8),
	.w8(32'h3c1d9a2f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeb8f7),
	.w1(32'hb9912d54),
	.w2(32'h3b7a397d),
	.w3(32'h3c0d979f),
	.w4(32'h3bafecb1),
	.w5(32'h3ad4af2c),
	.w6(32'h3b480337),
	.w7(32'h3bdbd4d1),
	.w8(32'h3c120960),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb62cf5),
	.w1(32'hbbfcbb47),
	.w2(32'hbc5aeb74),
	.w3(32'hbb8c9f48),
	.w4(32'hbb82457a),
	.w5(32'hbc178986),
	.w6(32'h3983b62e),
	.w7(32'hbb52bb08),
	.w8(32'hbbe845a9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa84d82),
	.w1(32'hbacd6cf9),
	.w2(32'hbb7ed2f9),
	.w3(32'hbc2a49f6),
	.w4(32'hbbc222f6),
	.w5(32'h3c786b32),
	.w6(32'hbc3b07f3),
	.w7(32'h3b39bf16),
	.w8(32'hbb1777aa),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3701f8),
	.w1(32'h3994d215),
	.w2(32'h3b72a762),
	.w3(32'h3c3f8b4e),
	.w4(32'hbb407ec6),
	.w5(32'h39f9c4b5),
	.w6(32'h3a454930),
	.w7(32'h3b1b4592),
	.w8(32'hbb80d913),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b988de2),
	.w1(32'h3bf2c318),
	.w2(32'h3c197154),
	.w3(32'hbabd71f5),
	.w4(32'h3b2e50bf),
	.w5(32'h3bea465e),
	.w6(32'h3a6c8f86),
	.w7(32'h3b33ee50),
	.w8(32'h3a534841),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c010475),
	.w1(32'h3b2a73ed),
	.w2(32'h3c409b48),
	.w3(32'hba5701fc),
	.w4(32'h3b197a7e),
	.w5(32'h3be9e60e),
	.w6(32'hbadf3c11),
	.w7(32'h3c2e0bfe),
	.w8(32'h3b499af8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f02b4),
	.w1(32'h3b5733b9),
	.w2(32'hbc03d32e),
	.w3(32'h3c272fc2),
	.w4(32'h3ba0748d),
	.w5(32'hbbccbb98),
	.w6(32'h3a4021f4),
	.w7(32'hba208c25),
	.w8(32'hbbbeb0ec),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394474fb),
	.w1(32'hbbdcf483),
	.w2(32'h3beb0914),
	.w3(32'h3bbf0362),
	.w4(32'hbbdda6ef),
	.w5(32'h3cbc87ab),
	.w6(32'hba3c51ad),
	.w7(32'hbbe85f4d),
	.w8(32'h3bf86007),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1f662),
	.w1(32'hbb3576f9),
	.w2(32'h3bff1d3a),
	.w3(32'h3b3b0555),
	.w4(32'hbc205dd2),
	.w5(32'h3b9f9869),
	.w6(32'hbb5ebbe9),
	.w7(32'hbbc7c59a),
	.w8(32'h3c24a977),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12575c),
	.w1(32'hbb4cf1b7),
	.w2(32'h3bd36c25),
	.w3(32'hbb3888a4),
	.w4(32'hbbdc4608),
	.w5(32'h3be13eff),
	.w6(32'hbb0a00e5),
	.w7(32'hbbe64b7a),
	.w8(32'h3af87e7b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d8ace),
	.w1(32'hbbbb1a3b),
	.w2(32'h3a67d2d3),
	.w3(32'hbc20c06c),
	.w4(32'hbbac96d5),
	.w5(32'h3bb3d94e),
	.w6(32'h3abf93f8),
	.w7(32'h3b860ecf),
	.w8(32'h3c791c68),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4598f1),
	.w1(32'h3c12fb3f),
	.w2(32'hbbc5a786),
	.w3(32'h3a94af18),
	.w4(32'hbaadd222),
	.w5(32'hbc15e7e8),
	.w6(32'h3bee1fd4),
	.w7(32'hbc5f5d5c),
	.w8(32'hbc68116c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08e2d5),
	.w1(32'hbb85ee24),
	.w2(32'h3be0917c),
	.w3(32'h3bdb8c85),
	.w4(32'hbbba1b84),
	.w5(32'h3c2f74a3),
	.w6(32'h399e627a),
	.w7(32'hbb146a87),
	.w8(32'h3c2d1f32),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa81cc9),
	.w1(32'h3b0c5b38),
	.w2(32'h3b1f7227),
	.w3(32'hbae3f2d9),
	.w4(32'h3a6604a8),
	.w5(32'h3bf75cc4),
	.w6(32'hbb6e9481),
	.w7(32'h39eceed2),
	.w8(32'h3bbec2f2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a067b15),
	.w1(32'h3acec613),
	.w2(32'h3b34d02e),
	.w3(32'h3b9ab689),
	.w4(32'h3b26e564),
	.w5(32'h3c15c4da),
	.w6(32'h3a85e32e),
	.w7(32'hba5fd6cb),
	.w8(32'h3ba132b1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13baef),
	.w1(32'hbc2b1247),
	.w2(32'hbb889a37),
	.w3(32'hbc55bcee),
	.w4(32'hba66b178),
	.w5(32'h3be7a6a2),
	.w6(32'hbbe72e91),
	.w7(32'h3c64ccb6),
	.w8(32'h3c871f14),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96adb2),
	.w1(32'hbba10a8e),
	.w2(32'h3a801dbf),
	.w3(32'h3a4bb97c),
	.w4(32'hbbe72674),
	.w5(32'h3bbc6a51),
	.w6(32'h3ba41445),
	.w7(32'hbb8db32f),
	.w8(32'hbbb30337),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96adf7),
	.w1(32'hbbdcfac1),
	.w2(32'h3ba01cda),
	.w3(32'h3ae6582d),
	.w4(32'hbb320f1f),
	.w5(32'h3c20ddcc),
	.w6(32'h3ae67ad4),
	.w7(32'h38db6dcc),
	.w8(32'h3b92ca3c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66714c),
	.w1(32'h3b2808a4),
	.w2(32'hbb3ab942),
	.w3(32'hbbe647d0),
	.w4(32'hbb8bdab2),
	.w5(32'hbb3e3536),
	.w6(32'hbc06983d),
	.w7(32'hbb867baf),
	.w8(32'hbb1d32f8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0df1d),
	.w1(32'h3aea67f5),
	.w2(32'h3bf1d404),
	.w3(32'hbb754cc0),
	.w4(32'hbbfa895c),
	.w5(32'hbba13118),
	.w6(32'h39be150f),
	.w7(32'hbb73a51d),
	.w8(32'hbb417bda),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1036d),
	.w1(32'hba911922),
	.w2(32'h3b2dd3af),
	.w3(32'hbb44f68a),
	.w4(32'h3b73322d),
	.w5(32'hbab4ffa2),
	.w6(32'hbb35b18b),
	.w7(32'h3b694d58),
	.w8(32'h3abae26a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ae183),
	.w1(32'hbb9cf241),
	.w2(32'h3bbd6f1d),
	.w3(32'h3bebe4c2),
	.w4(32'h3bb353ea),
	.w5(32'h3c0fa2bb),
	.w6(32'h3b87cdcb),
	.w7(32'hbb85dd52),
	.w8(32'hbba0c3f1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b756c0f),
	.w1(32'hbb7720ef),
	.w2(32'h3b11f76b),
	.w3(32'h3b97ecb7),
	.w4(32'hb5a3e3cf),
	.w5(32'h3bdafe34),
	.w6(32'h3b42fe6f),
	.w7(32'h3bb4f236),
	.w8(32'h3bef52ec),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb290f86),
	.w1(32'hba1777b6),
	.w2(32'hbbbf7c49),
	.w3(32'hbbb021a3),
	.w4(32'hbbc66e5b),
	.w5(32'h3b8ab0d8),
	.w6(32'hbb94570e),
	.w7(32'hbbbc7262),
	.w8(32'hbb5925a5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5049d),
	.w1(32'hba92a550),
	.w2(32'h3b574d97),
	.w3(32'hb98480df),
	.w4(32'hbb938c9f),
	.w5(32'hbb8115a9),
	.w6(32'hbb1cffc6),
	.w7(32'h3b123369),
	.w8(32'h39f3c57b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63b1e1),
	.w1(32'h3c2f35e1),
	.w2(32'hbbcaf0c7),
	.w3(32'h3c071961),
	.w4(32'h3a296ef8),
	.w5(32'hbbcc7824),
	.w6(32'h3b798001),
	.w7(32'hba7e599f),
	.w8(32'hbc25fcde),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813e8f),
	.w1(32'h3b95ecf3),
	.w2(32'hbac498df),
	.w3(32'hbade0d7c),
	.w4(32'h3b87753b),
	.w5(32'hbc153782),
	.w6(32'h3bdbd1eb),
	.w7(32'hba305e88),
	.w8(32'hbbc1fd4d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37a863),
	.w1(32'h3b9336d5),
	.w2(32'hbbaa1c8b),
	.w3(32'hbb389c1f),
	.w4(32'h3b7417d2),
	.w5(32'hbb6d6336),
	.w6(32'h3ab60dff),
	.w7(32'h3b4852e9),
	.w8(32'h3a65d484),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b860138),
	.w1(32'h3b004cd1),
	.w2(32'h3b19911e),
	.w3(32'h3a12b234),
	.w4(32'h3a3dd242),
	.w5(32'hbb03ace1),
	.w6(32'h3b6ea934),
	.w7(32'h3b446cdd),
	.w8(32'hbb811678),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3666a5),
	.w1(32'h3b1b72e6),
	.w2(32'hbb2bf5e9),
	.w3(32'hba57d6b3),
	.w4(32'hbaa15d69),
	.w5(32'hbc042bcd),
	.w6(32'h3b438a60),
	.w7(32'h3a205801),
	.w8(32'hbb1ffd20),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f1807),
	.w1(32'h3c6d1a09),
	.w2(32'h3bd8a078),
	.w3(32'h3ae06100),
	.w4(32'h3c144880),
	.w5(32'h3b480bff),
	.w6(32'h3b26c185),
	.w7(32'h3ae0d0fe),
	.w8(32'h37af35e9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb976f44),
	.w1(32'h3bc9eb31),
	.w2(32'hbc016256),
	.w3(32'hbb74c2bd),
	.w4(32'h3b52b460),
	.w5(32'hbc62fa51),
	.w6(32'hbbe1fbad),
	.w7(32'h3a8dea3d),
	.w8(32'hbb9a12cc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a615bb4),
	.w1(32'hbbf67880),
	.w2(32'hbc072cbf),
	.w3(32'h3aaee779),
	.w4(32'hbc0edbe3),
	.w5(32'hbb228e2a),
	.w6(32'hbb19cf77),
	.w7(32'hbb01580a),
	.w8(32'h3abd78c6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01759e),
	.w1(32'hbb2a2f8f),
	.w2(32'h3b88af2f),
	.w3(32'hbb918851),
	.w4(32'hbbaf7f25),
	.w5(32'h3c399513),
	.w6(32'hbc0fe15a),
	.w7(32'hbc2a047a),
	.w8(32'hbb025e51),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb1a6a),
	.w1(32'hbbb4a7af),
	.w2(32'hbb111363),
	.w3(32'hb9769534),
	.w4(32'hbb8081bc),
	.w5(32'hb99b37b5),
	.w6(32'h3a428f90),
	.w7(32'h3b02bdfe),
	.w8(32'h3b3f0816),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe869fa),
	.w1(32'h3a9adc54),
	.w2(32'h3b916ef9),
	.w3(32'hbbd10c74),
	.w4(32'hbae41e83),
	.w5(32'hbc011de6),
	.w6(32'hba4247b8),
	.w7(32'h3b7792c2),
	.w8(32'h3ab6ca78),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12c00c),
	.w1(32'hba50fb0f),
	.w2(32'hbb0559cc),
	.w3(32'h3a3e4cf5),
	.w4(32'hbb41abfb),
	.w5(32'h3afb806e),
	.w6(32'h3b109aa3),
	.w7(32'h3a34fd33),
	.w8(32'hbbaf2d7e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6ba3),
	.w1(32'hbc494553),
	.w2(32'hbc2dcaf2),
	.w3(32'hbb197c9b),
	.w4(32'hbc190655),
	.w5(32'h3ba5db96),
	.w6(32'h3b1b7ce5),
	.w7(32'hbc319f84),
	.w8(32'hbadf7a0f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31df87),
	.w1(32'h3a18b9b2),
	.w2(32'hbb61030c),
	.w3(32'h3b83140e),
	.w4(32'hbbb19311),
	.w5(32'h3c439676),
	.w6(32'h3b02fd68),
	.w7(32'hbb88b859),
	.w8(32'h3b152af2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8636a),
	.w1(32'h3c1da9c4),
	.w2(32'h3ba4c4be),
	.w3(32'h3b1b4845),
	.w4(32'h3bad3d42),
	.w5(32'hbb9a3e01),
	.w6(32'hbba226b5),
	.w7(32'h3bb76cb0),
	.w8(32'hbb27354d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d7afb),
	.w1(32'hbb0cf333),
	.w2(32'hbb19ece1),
	.w3(32'hbaf8a1d4),
	.w4(32'hba588f5e),
	.w5(32'h3b65446a),
	.w6(32'hb994efd1),
	.w7(32'hbaa6835e),
	.w8(32'hb9a67a7b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30ee6a),
	.w1(32'h3be39da1),
	.w2(32'h3be61ef1),
	.w3(32'hbade1935),
	.w4(32'h3b82d790),
	.w5(32'h3bd9c2b4),
	.w6(32'h3b12a1c0),
	.w7(32'h3ba528ad),
	.w8(32'h3c0d0763),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3520c8),
	.w1(32'h3bf176a2),
	.w2(32'h3ab1daba),
	.w3(32'h393014e7),
	.w4(32'h3c071d26),
	.w5(32'hbb97a986),
	.w6(32'h3b7dfee6),
	.w7(32'h3b05e002),
	.w8(32'hbbc4addc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f11fa8),
	.w1(32'hbaeb0a0f),
	.w2(32'h39f4e9bb),
	.w3(32'h3a069431),
	.w4(32'hba059761),
	.w5(32'hbb9c1db1),
	.w6(32'h3b6ccb3c),
	.w7(32'hbaafebd1),
	.w8(32'h39cbd39a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3194d9),
	.w1(32'h3bda9a33),
	.w2(32'hbb767c32),
	.w3(32'hbb3b096a),
	.w4(32'hbbe34ebe),
	.w5(32'h3b9ef9c3),
	.w6(32'hbaf8b10b),
	.w7(32'h3b801729),
	.w8(32'h3c55a541),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35a2bf),
	.w1(32'hba098b95),
	.w2(32'h3aa9c63c),
	.w3(32'hbc5fa340),
	.w4(32'hbae69fe2),
	.w5(32'hb9f62bb8),
	.w6(32'hba69ea5a),
	.w7(32'h3a97d9fa),
	.w8(32'h3b01c2cb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18d2c0),
	.w1(32'hb89c4099),
	.w2(32'h3c1b3292),
	.w3(32'h3ba15350),
	.w4(32'hbbd1385b),
	.w5(32'h398280e5),
	.w6(32'h3aa2a2c3),
	.w7(32'hbb690622),
	.w8(32'hbbae0bad),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcfb9e),
	.w1(32'h3bfc10ed),
	.w2(32'hbae6dd1f),
	.w3(32'hbb6162cc),
	.w4(32'h3bda4a85),
	.w5(32'h3b62bfc4),
	.w6(32'hbbbd05a0),
	.w7(32'h3ab081f2),
	.w8(32'hbbe093f7),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4ae30),
	.w1(32'hba87a1c5),
	.w2(32'h3aa13d07),
	.w3(32'hbb7a2e48),
	.w4(32'hbb4862e2),
	.w5(32'h3a10ad93),
	.w6(32'hbb8b0586),
	.w7(32'hbbbc2856),
	.w8(32'hbb1ee843),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973eb3),
	.w1(32'h3b3ff8e8),
	.w2(32'h3ae029df),
	.w3(32'hbbb969bd),
	.w4(32'h39cc8044),
	.w5(32'hb9adf6fe),
	.w6(32'hbb135be1),
	.w7(32'hba4e64b5),
	.w8(32'h3b9f95ac),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a47af),
	.w1(32'hbb7ebf4b),
	.w2(32'h3b19ac97),
	.w3(32'h3afdba08),
	.w4(32'hbb73493d),
	.w5(32'h3be541f1),
	.w6(32'h3bfd3f82),
	.w7(32'h3824cbf7),
	.w8(32'h3bac9c93),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32c045),
	.w1(32'hbc0b5066),
	.w2(32'hbb782442),
	.w3(32'hba83ce66),
	.w4(32'hbc029bd6),
	.w5(32'h3cab4601),
	.w6(32'hbb5bb384),
	.w7(32'hbb21bf78),
	.w8(32'h3c355f72),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c610d10),
	.w1(32'h3bdd1e08),
	.w2(32'h3bc1afa5),
	.w3(32'h3bc320a2),
	.w4(32'hbbe144ce),
	.w5(32'hbb36ec65),
	.w6(32'hbba3baad),
	.w7(32'hbc0bb68d),
	.w8(32'h3b1456ab),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1e618),
	.w1(32'hbbf6f1e6),
	.w2(32'h3bd9e019),
	.w3(32'hbaade279),
	.w4(32'hbb251215),
	.w5(32'h3c15111c),
	.w6(32'h3bbc377c),
	.w7(32'h3b013dd7),
	.w8(32'h3c29ad51),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbc861),
	.w1(32'hbabccc48),
	.w2(32'h3c0561a7),
	.w3(32'hbb2d9cf1),
	.w4(32'h3b894f10),
	.w5(32'h3c4512ab),
	.w6(32'hbb00d465),
	.w7(32'h3b66a83c),
	.w8(32'hba38506f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bbd68),
	.w1(32'h3b3065e3),
	.w2(32'hbb0ba035),
	.w3(32'h3bb6f960),
	.w4(32'h3b707552),
	.w5(32'hb9f8d39e),
	.w6(32'h3afc6e31),
	.w7(32'h3c031707),
	.w8(32'h3bc96ced),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e2099),
	.w1(32'h3b685580),
	.w2(32'hbb8db6ca),
	.w3(32'hb9ad9d34),
	.w4(32'h3a04e145),
	.w5(32'hbc24f799),
	.w6(32'h3b44e835),
	.w7(32'h3b0b9afa),
	.w8(32'hbc2babb6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf347e),
	.w1(32'hbaf07518),
	.w2(32'hbabaa547),
	.w3(32'hbaaae50f),
	.w4(32'hbb547ab1),
	.w5(32'hba2aa89c),
	.w6(32'h3b46240b),
	.w7(32'hbbfe06e2),
	.w8(32'h3acdf586),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb99b77),
	.w1(32'hbbef704b),
	.w2(32'h3bb90212),
	.w3(32'h3b63928e),
	.w4(32'hbaf85143),
	.w5(32'hbbb85a4b),
	.w6(32'h3a4c2e4a),
	.w7(32'hbb038088),
	.w8(32'hbb8d1c97),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc12c5),
	.w1(32'hbba87175),
	.w2(32'hbb350011),
	.w3(32'hbc3e8d7d),
	.w4(32'hbc0b8ce3),
	.w5(32'h3c26e454),
	.w6(32'h3b9a6540),
	.w7(32'hbb8d66aa),
	.w8(32'h3c09dcaa),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ae664),
	.w1(32'hbb65c51e),
	.w2(32'h3c2106d0),
	.w3(32'hbb8ad800),
	.w4(32'hbc0174b5),
	.w5(32'h3cabfb10),
	.w6(32'hbc29ed45),
	.w7(32'hbac14712),
	.w8(32'h3c9f08de),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c482391),
	.w1(32'hba5e7651),
	.w2(32'hbb3ba4cb),
	.w3(32'h3b800c9a),
	.w4(32'hbb19b320),
	.w5(32'hbbde6e9f),
	.w6(32'hb6043a41),
	.w7(32'hbb86605b),
	.w8(32'hbb78687b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe16c6e),
	.w1(32'hbbceab29),
	.w2(32'h388cb888),
	.w3(32'hbc31cdd0),
	.w4(32'hbc053224),
	.w5(32'hbb4a56ce),
	.w6(32'h3b7f63de),
	.w7(32'hbc28911b),
	.w8(32'hbb4ed0a0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b012305),
	.w1(32'hbb9757fe),
	.w2(32'hbbd068e4),
	.w3(32'h3a87885b),
	.w4(32'h3b2a971a),
	.w5(32'hbbf3c642),
	.w6(32'h3abcfce2),
	.w7(32'hbb24cd14),
	.w8(32'hbbf0e650),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab01495),
	.w1(32'h398021b3),
	.w2(32'h3b442ee0),
	.w3(32'hbb61cb61),
	.w4(32'hbaf4e2c4),
	.w5(32'hbba43e97),
	.w6(32'hbb870852),
	.w7(32'hbadc6f15),
	.w8(32'hbb6cca76),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8c4b1),
	.w1(32'hbba931b7),
	.w2(32'hbc0e5533),
	.w3(32'hbbe16ca6),
	.w4(32'hbbf141fd),
	.w5(32'hb98a0f96),
	.w6(32'h3b055dbb),
	.w7(32'hbb9e98d2),
	.w8(32'h3af24aeb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c175cfd),
	.w1(32'hbbb64743),
	.w2(32'hbb0b7e15),
	.w3(32'h3c3adbcc),
	.w4(32'hbb6f870f),
	.w5(32'h39421567),
	.w6(32'hbabe3115),
	.w7(32'hbb3f5a97),
	.w8(32'hbb7c00b3),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054204),
	.w1(32'h3ba9a495),
	.w2(32'hbbb89e14),
	.w3(32'hbbbbd288),
	.w4(32'h3af45412),
	.w5(32'hbb8e234a),
	.w6(32'hba6117bb),
	.w7(32'h39e9fe43),
	.w8(32'hbc001ac0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6440d5),
	.w1(32'hbbeae3f7),
	.w2(32'h3beea3f9),
	.w3(32'hbaa64331),
	.w4(32'hbb89df7b),
	.w5(32'h3bf2aca0),
	.w6(32'h3b36b50e),
	.w7(32'h391c5334),
	.w8(32'h3bdae23a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4637c),
	.w1(32'h3c0f159e),
	.w2(32'h3b8cabcc),
	.w3(32'hbbcb00cb),
	.w4(32'h3b7cf339),
	.w5(32'hba285eb5),
	.w6(32'hbbe99d0d),
	.w7(32'h3ab54c0b),
	.w8(32'hbb814cff),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeee64d),
	.w1(32'h3ba1f1be),
	.w2(32'h3ab101e9),
	.w3(32'h3b92c9d7),
	.w4(32'h3b07d88b),
	.w5(32'h3b8d4820),
	.w6(32'h3ba715a7),
	.w7(32'h3a2761a1),
	.w8(32'h3b98cb1e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947c41),
	.w1(32'h3a2172ce),
	.w2(32'h3be159d5),
	.w3(32'hbbddac18),
	.w4(32'hba568593),
	.w5(32'h3ab70d8a),
	.w6(32'hbbd2f23f),
	.w7(32'h3ac54dee),
	.w8(32'h3bc98ff6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386f52ad),
	.w1(32'h3bc668f9),
	.w2(32'h3b12ac4f),
	.w3(32'h3b0639b3),
	.w4(32'h3b805170),
	.w5(32'h3b0ca729),
	.w6(32'h3b7efe46),
	.w7(32'hb99c8fdb),
	.w8(32'hba3cdc23),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25967b),
	.w1(32'h3be07788),
	.w2(32'h3c3962a7),
	.w3(32'h3b27a341),
	.w4(32'h3bb41d54),
	.w5(32'h3b6bfeb9),
	.w6(32'h3be47889),
	.w7(32'h3aa57e62),
	.w8(32'h3a9f8828),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf4fdf),
	.w1(32'h3c2f5632),
	.w2(32'hbc154877),
	.w3(32'hba6e0f70),
	.w4(32'h3c2fb3bd),
	.w5(32'hbc31711c),
	.w6(32'h3b8d5058),
	.w7(32'h3bea7336),
	.w8(32'hbc215e1e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd2e2f),
	.w1(32'hba95b5cf),
	.w2(32'hbb038725),
	.w3(32'hbbd5a0fc),
	.w4(32'h3b09fb3e),
	.w5(32'h3b1f71c5),
	.w6(32'hbad09f10),
	.w7(32'hbb39712b),
	.w8(32'h3a4a64ff),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2f3e9),
	.w1(32'hbb764ac2),
	.w2(32'hbc483203),
	.w3(32'h3b1ca8e9),
	.w4(32'hbacde85e),
	.w5(32'hbbde4a6a),
	.w6(32'h3ae6af7f),
	.w7(32'hbafecf9c),
	.w8(32'h3a82e9b4),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb107b71),
	.w1(32'h3c04912a),
	.w2(32'hbba71542),
	.w3(32'hbb61738e),
	.w4(32'h3c2efe5c),
	.w5(32'hbbab4b47),
	.w6(32'hbaaa8a7a),
	.w7(32'h3c02da95),
	.w8(32'hbbd6719d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b837e83),
	.w1(32'h3ab088a4),
	.w2(32'hbbc55fd1),
	.w3(32'h3bb1f813),
	.w4(32'hb8a01426),
	.w5(32'hbc1459e0),
	.w6(32'h3a671511),
	.w7(32'hbb3445ff),
	.w8(32'hbc12a19f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c4bd3),
	.w1(32'hbb168508),
	.w2(32'h3c2116ea),
	.w3(32'hbc18c763),
	.w4(32'hb9cacf8c),
	.w5(32'hb9d49743),
	.w6(32'hbc08d090),
	.w7(32'hb9b35c0b),
	.w8(32'h3be28192),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0ea2c),
	.w1(32'hbbdb4eab),
	.w2(32'h3b214ca5),
	.w3(32'hba16187d),
	.w4(32'hbb864157),
	.w5(32'h3c9415b7),
	.w6(32'hbb86a7ba),
	.w7(32'hbb2b7eee),
	.w8(32'h3c1eddb4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebdca5),
	.w1(32'h3beb6685),
	.w2(32'h3c0b2e2d),
	.w3(32'h3bd3031f),
	.w4(32'h3bc728c1),
	.w5(32'h39c96c05),
	.w6(32'hba523ab0),
	.w7(32'h3bba6693),
	.w8(32'hb999ddc0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc99f52),
	.w1(32'h3a7e2462),
	.w2(32'hb836bea6),
	.w3(32'h3b07365b),
	.w4(32'h3b5672ad),
	.w5(32'hbb65929f),
	.w6(32'h3c2e0b3d),
	.w7(32'h3aef9060),
	.w8(32'hba986d65),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c76ad),
	.w1(32'hbae5f5c7),
	.w2(32'hba413251),
	.w3(32'hbbe76d0b),
	.w4(32'hb9863aac),
	.w5(32'h3ac98d18),
	.w6(32'hbbf0b092),
	.w7(32'hbbac3198),
	.w8(32'h3b176151),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23542e),
	.w1(32'h3abe03d5),
	.w2(32'h3c2846c0),
	.w3(32'hbb996580),
	.w4(32'h3b230e22),
	.w5(32'h3c9bf932),
	.w6(32'hbbadcf7b),
	.w7(32'h3a6bdef7),
	.w8(32'h3b769af4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2abf1f),
	.w1(32'hbb8bb9c3),
	.w2(32'h3c26f638),
	.w3(32'hbbadff70),
	.w4(32'hbb7fe9e0),
	.w5(32'h3ca80e57),
	.w6(32'hbb6fb205),
	.w7(32'h3afbafa0),
	.w8(32'h3bab0548),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca5fb1),
	.w1(32'h3b25f7e4),
	.w2(32'h3a32dbae),
	.w3(32'h3b0e2730),
	.w4(32'hba96950b),
	.w5(32'h3b1dcae9),
	.w6(32'h3a56e06b),
	.w7(32'h39ecb9a5),
	.w8(32'hbae15c94),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f78ea),
	.w1(32'hbb1480dd),
	.w2(32'h3aca8d6b),
	.w3(32'hbac2baf2),
	.w4(32'hbb1d6a42),
	.w5(32'h3b0150ae),
	.w6(32'hbb7bac33),
	.w7(32'h3b78aa2f),
	.w8(32'h3b5f1413),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b559ff4),
	.w1(32'h3bc7ba0d),
	.w2(32'hba35bb5e),
	.w3(32'hbaf6b513),
	.w4(32'h3ba93d25),
	.w5(32'hbba2074b),
	.w6(32'hb9adcd6c),
	.w7(32'h3c1b24c5),
	.w8(32'hb9b4e527),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b0f5b),
	.w1(32'h3bab9e2c),
	.w2(32'hbc0b1a2a),
	.w3(32'hbc3592ff),
	.w4(32'hbb8ac8b5),
	.w5(32'hbbe46089),
	.w6(32'hbc30e4cc),
	.w7(32'hbb4e3000),
	.w8(32'hbc6637e1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89299),
	.w1(32'h3c011395),
	.w2(32'h3ab9b934),
	.w3(32'hbb673ac6),
	.w4(32'h3b833e70),
	.w5(32'hbad23e80),
	.w6(32'hbb28d8ae),
	.w7(32'h3a768f6a),
	.w8(32'hbb84912a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6946c),
	.w1(32'h3bf61dfd),
	.w2(32'h3b640016),
	.w3(32'h3b43f88a),
	.w4(32'h3aef95d3),
	.w5(32'hbb8a38ae),
	.w6(32'h3b051d91),
	.w7(32'h3b24dd9f),
	.w8(32'hbb82d1f4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407242),
	.w1(32'h3c092cec),
	.w2(32'h3c2c52f0),
	.w3(32'hba70df5a),
	.w4(32'h3b4536fc),
	.w5(32'h3b189eb3),
	.w6(32'h3abf343c),
	.w7(32'hbb6ae464),
	.w8(32'hbb075eea),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be717a2),
	.w1(32'hb8e55361),
	.w2(32'hbbcaa626),
	.w3(32'h3967a289),
	.w4(32'h3b428ffc),
	.w5(32'hbba08400),
	.w6(32'hba3d690a),
	.w7(32'hbac1b49b),
	.w8(32'hbbe28a62),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f4a09),
	.w1(32'h39b6b868),
	.w2(32'hbb3d9060),
	.w3(32'h3b67d701),
	.w4(32'h38cfd44c),
	.w5(32'hba8ad79e),
	.w6(32'h3ada04f5),
	.w7(32'hba03a9a4),
	.w8(32'hbaca25ec),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c85b1),
	.w1(32'hbace9387),
	.w2(32'hbb395656),
	.w3(32'hbb0be193),
	.w4(32'h3aaecd3c),
	.w5(32'hbb37f1a4),
	.w6(32'hbaa18890),
	.w7(32'hb99db3ea),
	.w8(32'hbb57e6df),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc78d2),
	.w1(32'hbbcc2edc),
	.w2(32'h3c19474a),
	.w3(32'hbba97598),
	.w4(32'hbc0bc57e),
	.w5(32'h3c9f503c),
	.w6(32'hba093386),
	.w7(32'hbb6df83b),
	.w8(32'h3cb29c13),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabecff),
	.w1(32'hbb613a81),
	.w2(32'hbb10bc63),
	.w3(32'hba170cdb),
	.w4(32'hba276f40),
	.w5(32'hbc252378),
	.w6(32'h3b6fbcce),
	.w7(32'h3b2fbee9),
	.w8(32'hbc281c8e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f5839),
	.w1(32'h3bec083d),
	.w2(32'h3725a0d6),
	.w3(32'hbc35584b),
	.w4(32'h3c02b73f),
	.w5(32'h3b86e70b),
	.w6(32'hbbf6aaf3),
	.w7(32'hbb4676e0),
	.w8(32'h3b4628a1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c013d),
	.w1(32'h3b464345),
	.w2(32'hbb7c1182),
	.w3(32'h3b444d10),
	.w4(32'hba32055a),
	.w5(32'h3c376f89),
	.w6(32'h3b95f57e),
	.w7(32'hb9d3fc6e),
	.w8(32'h3ac4921f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17da3c),
	.w1(32'hbb8f9518),
	.w2(32'hbb31497c),
	.w3(32'h3a928af1),
	.w4(32'hbba39a84),
	.w5(32'hbb041150),
	.w6(32'h395e663f),
	.w7(32'hbabf7d91),
	.w8(32'h3a924b3a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fbcb0),
	.w1(32'hbb7e59ca),
	.w2(32'hbb7df930),
	.w3(32'h3a21e674),
	.w4(32'hbb052dbf),
	.w5(32'h39eff20b),
	.w6(32'h3ab9efe6),
	.w7(32'hbc09f917),
	.w8(32'hbb59a1ab),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcef5e),
	.w1(32'h39051083),
	.w2(32'hbb4a8237),
	.w3(32'h3bad444f),
	.w4(32'h3aa2c830),
	.w5(32'hbc33170b),
	.w6(32'h3ad2200e),
	.w7(32'hbb066aa3),
	.w8(32'hbb92347e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb937291),
	.w1(32'h3bf9070d),
	.w2(32'h3b210d8f),
	.w3(32'hbbaab947),
	.w4(32'h3be67612),
	.w5(32'hbb4b16de),
	.w6(32'h3ae73940),
	.w7(32'h3ba743a8),
	.w8(32'h3b0fcdbf),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba439ae4),
	.w1(32'h3b57911a),
	.w2(32'hbb447cbe),
	.w3(32'hba6a16f2),
	.w4(32'h3b829b5e),
	.w5(32'hbb5fa395),
	.w6(32'hbaa5f0cf),
	.w7(32'h3a249b23),
	.w8(32'hbb0ee280),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2ef47),
	.w1(32'hbb1bd36d),
	.w2(32'hbb01d19c),
	.w3(32'hbaad4850),
	.w4(32'hb9a253f1),
	.w5(32'h3ba07f81),
	.w6(32'hb94a61c7),
	.w7(32'h3aff6ce2),
	.w8(32'h3a8fdccb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a88e85),
	.w1(32'hbb6df0bf),
	.w2(32'h3ad8248f),
	.w3(32'hbb3f67c2),
	.w4(32'hbc539a16),
	.w5(32'h3c021dab),
	.w6(32'hbb3d6fb5),
	.w7(32'hbb1b897e),
	.w8(32'h3b8c8b27),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2ecca),
	.w1(32'h3c4415af),
	.w2(32'h3b795a63),
	.w3(32'hbbb4440f),
	.w4(32'h3b80a5c8),
	.w5(32'h3bb19e0d),
	.w6(32'hbaec70bd),
	.w7(32'hbbd51b06),
	.w8(32'hbb4efae7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9886bc3),
	.w1(32'h3c1c4aad),
	.w2(32'h3bc0efe9),
	.w3(32'h39f2b895),
	.w4(32'h3c4b0ce3),
	.w5(32'hba838425),
	.w6(32'hbb8f7ae8),
	.w7(32'h3bfdd956),
	.w8(32'h3b0562a9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923d2d3),
	.w1(32'hbc378ac3),
	.w2(32'hbbd58169),
	.w3(32'hbb2172cc),
	.w4(32'hbc134957),
	.w5(32'hbbcf0a1c),
	.w6(32'h390deffc),
	.w7(32'hbbcd79d5),
	.w8(32'hbbbdba21),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0107b9),
	.w1(32'h3b2c4bfc),
	.w2(32'h3aed3cb3),
	.w3(32'hbba559e0),
	.w4(32'h398e297f),
	.w5(32'h3b04b442),
	.w6(32'hbad5acbd),
	.w7(32'hbb3f9249),
	.w8(32'hbb5412e4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1dbb9),
	.w1(32'h3a9a6fc4),
	.w2(32'h3b2175b7),
	.w3(32'h39d4361c),
	.w4(32'h3bd4e075),
	.w5(32'h3c1fb984),
	.w6(32'hbb5ef644),
	.w7(32'h398f77ee),
	.w8(32'h3b3ace8e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab09c79),
	.w1(32'h3b4fee7e),
	.w2(32'h3b3668c3),
	.w3(32'h3b14b223),
	.w4(32'h3bab8609),
	.w5(32'h3bab5577),
	.w6(32'h3b2fb1f6),
	.w7(32'h3b7f6b07),
	.w8(32'h3b88c046),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27e68b),
	.w1(32'h3b096e54),
	.w2(32'h3afb2cb3),
	.w3(32'hb8d40194),
	.w4(32'h3b17163b),
	.w5(32'h3b43c661),
	.w6(32'h3a89f66d),
	.w7(32'h3bd345e5),
	.w8(32'h3b963cdf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a606c38),
	.w1(32'h3b8f3b68),
	.w2(32'h3b513bbc),
	.w3(32'h3be10e76),
	.w4(32'hbb9cb986),
	.w5(32'hbb9d7501),
	.w6(32'h3b8eca62),
	.w7(32'hbba1aed8),
	.w8(32'hbc03ce0f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dc14a),
	.w1(32'h3c1b99d7),
	.w2(32'h3c16396b),
	.w3(32'hbb6d0eb2),
	.w4(32'h3b808068),
	.w5(32'h3c620d03),
	.w6(32'hbb57a573),
	.w7(32'h3a6b81b0),
	.w8(32'h3bedd5ae),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c1d96),
	.w1(32'h3bd1d077),
	.w2(32'hb9bc5a8f),
	.w3(32'h3bf4cc5b),
	.w4(32'h3c1b1307),
	.w5(32'h3b26fbac),
	.w6(32'h3b62a799),
	.w7(32'h3b6cae19),
	.w8(32'hbb27bb39),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc14ac8),
	.w1(32'h3bb3d7cb),
	.w2(32'h3bb2b735),
	.w3(32'h3acc86be),
	.w4(32'h3c0ca38c),
	.w5(32'h3c00e469),
	.w6(32'hbb811688),
	.w7(32'h3babff98),
	.w8(32'h3bcec684),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5589d),
	.w1(32'h3b1f4423),
	.w2(32'hb94a40ad),
	.w3(32'hbbaaefcc),
	.w4(32'h3c09ad50),
	.w5(32'h3b66869e),
	.w6(32'hbb9671e4),
	.w7(32'h3c5fde36),
	.w8(32'h3c15ccbc),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88684),
	.w1(32'hbb9c4d62),
	.w2(32'h3b954adc),
	.w3(32'hbb943f6f),
	.w4(32'hbb6bba40),
	.w5(32'h3c332d0e),
	.w6(32'hbae06fcb),
	.w7(32'hbbde29b5),
	.w8(32'h3b856da3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba72f6d),
	.w1(32'hbc13271d),
	.w2(32'hbba1c8b1),
	.w3(32'hbbf2a49a),
	.w4(32'hbc1b2de2),
	.w5(32'hbbe8d22c),
	.w6(32'hbc07d088),
	.w7(32'hbc0955c5),
	.w8(32'hbb96eedc),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3b8af),
	.w1(32'hbb873f6c),
	.w2(32'h3af765a6),
	.w3(32'hba82547e),
	.w4(32'hba371a10),
	.w5(32'h3b2c7cc9),
	.w6(32'h3a343325),
	.w7(32'hba4d78a9),
	.w8(32'h3b0bc8df),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bed28),
	.w1(32'hbbc09bcd),
	.w2(32'h3b64a7aa),
	.w3(32'hba0dd192),
	.w4(32'h3b2d3ca9),
	.w5(32'h3b148b19),
	.w6(32'hbacf8577),
	.w7(32'hbb95659a),
	.w8(32'hbb1aa286),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71679b),
	.w1(32'hbbae0ca2),
	.w2(32'h3bbfc6b9),
	.w3(32'hba1238de),
	.w4(32'hbb517962),
	.w5(32'h3c058678),
	.w6(32'hbb9d5b17),
	.w7(32'hbbdceb66),
	.w8(32'h3b5f53a6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5beaa1),
	.w1(32'h3a51c4c2),
	.w2(32'hbb4e381b),
	.w3(32'h3a691a80),
	.w4(32'hbb924df9),
	.w5(32'hbb6171f6),
	.w6(32'h3af7f341),
	.w7(32'hbb2b146b),
	.w8(32'hbb8c50f7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba994864),
	.w1(32'h3b1e1372),
	.w2(32'hbb430ccb),
	.w3(32'h3a79bf44),
	.w4(32'h3ae3114e),
	.w5(32'hbbe979a5),
	.w6(32'hb8d1cca4),
	.w7(32'h3a7048a5),
	.w8(32'hbb510ff3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16743f),
	.w1(32'hbb3a7e64),
	.w2(32'hbc08cc27),
	.w3(32'hbc1227bd),
	.w4(32'hbbb14351),
	.w5(32'hbc4ebf21),
	.w6(32'hbbf35a4e),
	.w7(32'hbbb9566f),
	.w8(32'hbbd8ffd6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5dc5),
	.w1(32'hbc132dd2),
	.w2(32'hbb621672),
	.w3(32'hbc2bdf16),
	.w4(32'hbbbc8a7b),
	.w5(32'h3b3fde78),
	.w6(32'hbbf50799),
	.w7(32'hbb5473bf),
	.w8(32'h39e091d6),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7087b9),
	.w1(32'hbbe32790),
	.w2(32'hbbab6feb),
	.w3(32'hbb9e441f),
	.w4(32'hbb7e1e0d),
	.w5(32'hbad13b1c),
	.w6(32'hbb99e069),
	.w7(32'h3b24639a),
	.w8(32'hb92ee7e0),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb979ed2),
	.w1(32'hbc6d704f),
	.w2(32'h3b89c22c),
	.w3(32'hbbe905ee),
	.w4(32'hbc400912),
	.w5(32'h3bcbe722),
	.w6(32'hbb71bdee),
	.w7(32'hbc349609),
	.w8(32'h3b5f710b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba50f32),
	.w1(32'hbaf26728),
	.w2(32'h3b8c0891),
	.w3(32'hbb87b46e),
	.w4(32'hbb9296d2),
	.w5(32'h3b19afd2),
	.w6(32'hbbcd7ae0),
	.w7(32'h3ad4ebc8),
	.w8(32'h3af6cc28),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c041151),
	.w1(32'h3b9929a2),
	.w2(32'h3b8c14b9),
	.w3(32'h3be1f59d),
	.w4(32'h3c06dc8f),
	.w5(32'h3b2fba43),
	.w6(32'hbae8e8bc),
	.w7(32'h3b8d8031),
	.w8(32'h3a24cd01),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae3908),
	.w1(32'h3ba8fb41),
	.w2(32'h39bdbf88),
	.w3(32'h3b70e14e),
	.w4(32'h3b452b0b),
	.w5(32'h3b32b2f3),
	.w6(32'h3bacfeb3),
	.w7(32'hb9c10be4),
	.w8(32'hbb4f942c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6642b8),
	.w1(32'hbbddb23d),
	.w2(32'hbbdd2752),
	.w3(32'hba141920),
	.w4(32'h3a24779f),
	.w5(32'hba60a4c0),
	.w6(32'h3a32fac9),
	.w7(32'h3c439546),
	.w8(32'h3badde92),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fe10f),
	.w1(32'h3b9838c3),
	.w2(32'h3c0420ab),
	.w3(32'hba0c3008),
	.w4(32'h3b9d9630),
	.w5(32'h3c68c0a0),
	.w6(32'h3ab8cee5),
	.w7(32'h3becbe9c),
	.w8(32'h3c3a1a36),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6aa22),
	.w1(32'hba43903c),
	.w2(32'h3a916dd5),
	.w3(32'h3bef766b),
	.w4(32'hbb81e8c2),
	.w5(32'hbb462e48),
	.w6(32'h3ba47e4a),
	.w7(32'hbaf915dd),
	.w8(32'hbabe7f02),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c70b7),
	.w1(32'h3b80aa7e),
	.w2(32'h39a3107e),
	.w3(32'h3a3aafb6),
	.w4(32'hb9eed054),
	.w5(32'h3b5266f7),
	.w6(32'h3a7e4ff8),
	.w7(32'h3b2e05bb),
	.w8(32'h39a42781),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae68257),
	.w1(32'hbb85cd17),
	.w2(32'hbaee35fb),
	.w3(32'hba84dcc4),
	.w4(32'hbbf2b6b9),
	.w5(32'hbb7b2c2c),
	.w6(32'hbaf3b32e),
	.w7(32'h39fb66a3),
	.w8(32'h3a81e2fe),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcff17e),
	.w1(32'h3c05a50e),
	.w2(32'h3c74307e),
	.w3(32'h3bc71b20),
	.w4(32'hbb76a77f),
	.w5(32'hbb1df850),
	.w6(32'h3ba792e0),
	.w7(32'h3af5cdf2),
	.w8(32'h3abe4d6a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07cf34),
	.w1(32'hbb2911b6),
	.w2(32'hb7f9eb06),
	.w3(32'h3ab14205),
	.w4(32'hbb458bf4),
	.w5(32'h3b665227),
	.w6(32'h3b7a988e),
	.w7(32'h3a9c44d0),
	.w8(32'h3b9341d4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7a34),
	.w1(32'h3b7fe57e),
	.w2(32'h3b985744),
	.w3(32'h3b067e27),
	.w4(32'hba722df0),
	.w5(32'h3b037892),
	.w6(32'h3c04de34),
	.w7(32'hb9a1a7bc),
	.w8(32'h398a0332),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20266c),
	.w1(32'hbb6df398),
	.w2(32'h3c4bca5d),
	.w3(32'hbbdbea2d),
	.w4(32'h3a98328e),
	.w5(32'h3c7a4c5b),
	.w6(32'hbae6c62b),
	.w7(32'h3b96bba1),
	.w8(32'h3c3fb0ca),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22ae94),
	.w1(32'hbbaa1268),
	.w2(32'h3bb4de41),
	.w3(32'h3bd37850),
	.w4(32'h39d236b3),
	.w5(32'h3bb72e2d),
	.w6(32'hb9ef07a8),
	.w7(32'hbb43066b),
	.w8(32'h3b7a400b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30c4e1),
	.w1(32'hba2bd03f),
	.w2(32'h3af96701),
	.w3(32'h3a928553),
	.w4(32'h3872e28e),
	.w5(32'h3b0166de),
	.w6(32'hb9c6d8fe),
	.w7(32'h3a0142be),
	.w8(32'hba571c67),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36a885),
	.w1(32'hbbfb4528),
	.w2(32'hbaab564c),
	.w3(32'hbb03abf6),
	.w4(32'hbbb5b45a),
	.w5(32'h3ac2d349),
	.w6(32'hba2a20bc),
	.w7(32'hb92a95d4),
	.w8(32'h3bb14818),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd0255),
	.w1(32'h3c131bc0),
	.w2(32'h39fad87c),
	.w3(32'h3a9a9e37),
	.w4(32'h3c1cbad0),
	.w5(32'hbad21980),
	.w6(32'h3b0098f0),
	.w7(32'h3bc49d7c),
	.w8(32'hbb4c6f1e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb939a6c),
	.w1(32'h3b468644),
	.w2(32'h3b687d0c),
	.w3(32'hbc0c102c),
	.w4(32'h3b27fb47),
	.w5(32'hbad49d9c),
	.w6(32'hbbdc2469),
	.w7(32'h3b1ec4e8),
	.w8(32'h39e0b5d1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c951c4),
	.w1(32'h3bcd519b),
	.w2(32'h3ba4fbf8),
	.w3(32'h3b78f8f2),
	.w4(32'h3b162a24),
	.w5(32'h39a24c80),
	.w6(32'h3beb2d51),
	.w7(32'h3b47054b),
	.w8(32'hbb0fd613),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c4780),
	.w1(32'h3bf668b7),
	.w2(32'h3c12b236),
	.w3(32'hbaa83dd8),
	.w4(32'h3bc5fda4),
	.w5(32'h3c8cd012),
	.w6(32'hbb84087c),
	.w7(32'hba14a3d7),
	.w8(32'h3c23a123),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ed067),
	.w1(32'hba1c1d6c),
	.w2(32'hbb9bed0c),
	.w3(32'h3c632f93),
	.w4(32'hbbf5e462),
	.w5(32'hbbdaa313),
	.w6(32'h3c71ac69),
	.w7(32'hbb69ba53),
	.w8(32'hba98923d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c50eb0),
	.w1(32'h3c001f01),
	.w2(32'h3c6de554),
	.w3(32'hbb87422a),
	.w4(32'hbb99394e),
	.w5(32'h3c142ab9),
	.w6(32'h38feba0d),
	.w7(32'hbb97ff00),
	.w8(32'h3aaafdc1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52a47),
	.w1(32'h3b8852bf),
	.w2(32'h3be2eb3b),
	.w3(32'h3ac277d5),
	.w4(32'h3b23db6b),
	.w5(32'h3ae52eac),
	.w6(32'hba9bf363),
	.w7(32'h3b45ea49),
	.w8(32'h3b5b5333),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3871605a),
	.w1(32'hba9a6d57),
	.w2(32'h3c3f044f),
	.w3(32'hbb5f58ed),
	.w4(32'h3c0715b1),
	.w5(32'h3cc4a4c6),
	.w6(32'hbbd6b390),
	.w7(32'hba85f936),
	.w8(32'h3c210bc8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea5ab2),
	.w1(32'hbabff115),
	.w2(32'hb9d4a6af),
	.w3(32'h3b439015),
	.w4(32'h3b6a6b75),
	.w5(32'h3b5a8dfe),
	.w6(32'h3b060aca),
	.w7(32'h3a690af9),
	.w8(32'h3b4332fb),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ae553),
	.w1(32'h3b328b7e),
	.w2(32'h3b3a2fff),
	.w3(32'hbb5d469d),
	.w4(32'h395f463f),
	.w5(32'h3b015269),
	.w6(32'hbb9f2b52),
	.w7(32'hb9be782c),
	.w8(32'h3b47ae30),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03bcd1),
	.w1(32'h3b58c4ae),
	.w2(32'h3bfa1695),
	.w3(32'h3addfd5b),
	.w4(32'h3be647d6),
	.w5(32'h3c1674fc),
	.w6(32'h3ad934bd),
	.w7(32'h3b326d4a),
	.w8(32'h3c01396b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb1dbe),
	.w1(32'h3b89eb68),
	.w2(32'hb9b25e0c),
	.w3(32'h3bfb5ed6),
	.w4(32'hbb09171d),
	.w5(32'hbc013296),
	.w6(32'h3b79e777),
	.w7(32'hbbebc3a1),
	.w8(32'hbc3bb361),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c52e87),
	.w1(32'h3a6dfeca),
	.w2(32'h3bd0dfb7),
	.w3(32'hbc0b0908),
	.w4(32'h3be65814),
	.w5(32'h3c2cde00),
	.w6(32'hbc0e2b04),
	.w7(32'h3c2a54f6),
	.w8(32'h3c466913),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c3f09),
	.w1(32'hba16eafa),
	.w2(32'h3b9d60e8),
	.w3(32'h3bd47ea2),
	.w4(32'h3aa25d66),
	.w5(32'h3c515adc),
	.w6(32'h3b9f6f6f),
	.w7(32'h3b938746),
	.w8(32'h3c11e63f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc2bcf),
	.w1(32'hbb0a2af9),
	.w2(32'hbabea6ed),
	.w3(32'h3bed4a7c),
	.w4(32'h3aff67da),
	.w5(32'h3bec1313),
	.w6(32'h3b625ebe),
	.w7(32'hbb69bc85),
	.w8(32'hb9ec59bb),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd9db7),
	.w1(32'h3a871f18),
	.w2(32'h3bd79dea),
	.w3(32'hbb76674a),
	.w4(32'h3c041eae),
	.w5(32'hba4990ab),
	.w6(32'hbbd91795),
	.w7(32'h3c317d5d),
	.w8(32'h3a91d683),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb27024),
	.w1(32'hbc50d8c9),
	.w2(32'hbc04c5ac),
	.w3(32'hbb1aafc2),
	.w4(32'hbc68040c),
	.w5(32'hbc3336cb),
	.w6(32'hbb3db83a),
	.w7(32'hbc688ab4),
	.w8(32'hbbd427eb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc108858),
	.w1(32'hbb8314b4),
	.w2(32'h37b31f8e),
	.w3(32'hbbe2bc48),
	.w4(32'hbb26108b),
	.w5(32'hbb812f63),
	.w6(32'hbbe13ffc),
	.w7(32'hb9985dfa),
	.w8(32'hbaf16819),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24ff73),
	.w1(32'hbaf2c38c),
	.w2(32'h3a3e0abc),
	.w3(32'hbb57dfd1),
	.w4(32'hbc1adbc7),
	.w5(32'hbc4e15c0),
	.w6(32'hbb5a9058),
	.w7(32'hbc4dfe13),
	.w8(32'hbc89988a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b3e5f),
	.w1(32'h3c2b8f06),
	.w2(32'h3c7267dd),
	.w3(32'hbc53dd0c),
	.w4(32'h3c76c048),
	.w5(32'h3c971024),
	.w6(32'hbc8628c7),
	.w7(32'h3be47902),
	.w8(32'h3c46f8f6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b116880),
	.w1(32'hbbaaf125),
	.w2(32'hbb567eae),
	.w3(32'h3bc33301),
	.w4(32'hbc3168be),
	.w5(32'hbc066def),
	.w6(32'h3b9eaba9),
	.w7(32'hbbf272d3),
	.w8(32'hbbb6335c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9957328),
	.w1(32'hbb9c880d),
	.w2(32'hba8375a6),
	.w3(32'h3b94e69c),
	.w4(32'hbaac7506),
	.w5(32'h3bcc9b29),
	.w6(32'h3a1e9452),
	.w7(32'h3abc2177),
	.w8(32'h3c040426),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule