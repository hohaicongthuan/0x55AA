module layer_10_featuremap_52(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab6428),
	.w1(32'hbc709e21),
	.w2(32'hbb99613e),
	.w3(32'hbc7524dd),
	.w4(32'hbc4be99d),
	.w5(32'h3c7e54d9),
	.w6(32'hbbe050ee),
	.w7(32'hba2f2f4d),
	.w8(32'h3c4b1fcd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91d7f6),
	.w1(32'hbc513bf3),
	.w2(32'hbc735725),
	.w3(32'hbbe105d9),
	.w4(32'hbca89f3b),
	.w5(32'hbd368115),
	.w6(32'h3bd0ef6d),
	.w7(32'hbc453482),
	.w8(32'hbcb888a9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0dd820),
	.w1(32'hbc440e5a),
	.w2(32'h3bfa4468),
	.w3(32'hbd8310de),
	.w4(32'hbcbc36e0),
	.w5(32'h3befacc8),
	.w6(32'hbd038d6d),
	.w7(32'hbc692a38),
	.w8(32'h3bbde6af),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0905d0),
	.w1(32'h3bfaab6d),
	.w2(32'h3b30df93),
	.w3(32'h3cb817e6),
	.w4(32'h3c8f998b),
	.w5(32'h3a7f5e89),
	.w6(32'h3c1e470a),
	.w7(32'h3c5fb533),
	.w8(32'hbc1cc3f8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c1496),
	.w1(32'h38d3f844),
	.w2(32'hbc0ac7ae),
	.w3(32'hba4c387d),
	.w4(32'h3b88fcf1),
	.w5(32'hbc3e7331),
	.w6(32'hbc1d15a5),
	.w7(32'hbc0bf05d),
	.w8(32'hbbee6715),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98dec5),
	.w1(32'hbc2ae88d),
	.w2(32'h3ba03034),
	.w3(32'hbcfdf364),
	.w4(32'hbcd5236e),
	.w5(32'h3bd50b34),
	.w6(32'hbcd7a7cc),
	.w7(32'hbc91a006),
	.w8(32'h3c0d4e17),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49be10),
	.w1(32'h3c306308),
	.w2(32'hbc53d87d),
	.w3(32'h3c3f7e6f),
	.w4(32'h3c38e365),
	.w5(32'hbc3adb22),
	.w6(32'h3c40cc94),
	.w7(32'h3c42e74d),
	.w8(32'hbbd7117c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd01d0c),
	.w1(32'hbc0bf5dc),
	.w2(32'hbc74ac48),
	.w3(32'hbca70c95),
	.w4(32'hbb40df9c),
	.w5(32'hbc9bf540),
	.w6(32'hbc7cd6d0),
	.w7(32'hbaae083b),
	.w8(32'hbc9c9bc6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73e83c),
	.w1(32'hbbb66edb),
	.w2(32'h3c40eefb),
	.w3(32'hbb5bc425),
	.w4(32'hbc172c26),
	.w5(32'h3c63ff49),
	.w6(32'hbc07ba78),
	.w7(32'hbb9aeae1),
	.w8(32'h3c1d09a0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4465f6),
	.w1(32'h3b5abcc4),
	.w2(32'h3c196b37),
	.w3(32'h3c2dbf71),
	.w4(32'hb846bda6),
	.w5(32'h3b649dc2),
	.w6(32'h3b9d4ac2),
	.w7(32'hbb480e12),
	.w8(32'hbb6d2184),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3bf3a),
	.w1(32'h3b5ca084),
	.w2(32'hb883515a),
	.w3(32'h3be65a56),
	.w4(32'h3b9320a0),
	.w5(32'h3b86907e),
	.w6(32'h3b890bad),
	.w7(32'h3abdf52f),
	.w8(32'h3b5aa634),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36e45c),
	.w1(32'h3c7a5376),
	.w2(32'hbb8d1cc7),
	.w3(32'h3c84afd8),
	.w4(32'h3cb75bda),
	.w5(32'hbb3944bb),
	.w6(32'h3c8555b4),
	.w7(32'h3caeea1c),
	.w8(32'hbb593271),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2255b),
	.w1(32'h392efd48),
	.w2(32'h3bd94b37),
	.w3(32'hbc1bc744),
	.w4(32'hbbc8c223),
	.w5(32'h3b6fa6b0),
	.w6(32'hbb86e406),
	.w7(32'hb8388add),
	.w8(32'hbc373ec2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39b9d1),
	.w1(32'h3b4a102d),
	.w2(32'hbc6c7eb9),
	.w3(32'h3b395874),
	.w4(32'h3c2546dc),
	.w5(32'hbcb0762f),
	.w6(32'hbb1667a0),
	.w7(32'hbab94382),
	.w8(32'hbc372842),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07a422),
	.w1(32'hbb21bdca),
	.w2(32'h3b5c8aa2),
	.w3(32'hbc7d888f),
	.w4(32'hbc84acfd),
	.w5(32'h38fdc4e1),
	.w6(32'hbc262c28),
	.w7(32'hbbc425f3),
	.w8(32'h3b8b5fb7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9d209),
	.w1(32'hb9f51380),
	.w2(32'hba69bcfa),
	.w3(32'hbb6d05dc),
	.w4(32'hbc116b6a),
	.w5(32'h39c09436),
	.w6(32'h39758c24),
	.w7(32'hbb2c5a7a),
	.w8(32'hbbd9d16e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26b191),
	.w1(32'h38fdb064),
	.w2(32'hbc6663fb),
	.w3(32'hbb035413),
	.w4(32'h399eeb60),
	.w5(32'hbc9eb8d4),
	.w6(32'hba85dcc4),
	.w7(32'hb9650e88),
	.w8(32'hbaaa7394),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd2ce59),
	.w1(32'hbc8c78c3),
	.w2(32'hbcb7eeb3),
	.w3(32'hbd1b5e77),
	.w4(32'hbcb07983),
	.w5(32'hbbd71942),
	.w6(32'hbcab6a6a),
	.w7(32'hbc745bd6),
	.w8(32'hbbe69c97),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb930b223),
	.w1(32'h3b9beb5d),
	.w2(32'hbb9917fc),
	.w3(32'h3b11ba1a),
	.w4(32'h3bac50df),
	.w5(32'hbb569d96),
	.w6(32'h3abcc5d2),
	.w7(32'h3b24de33),
	.w8(32'hbc02f151),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa95106),
	.w1(32'h3b05ea45),
	.w2(32'h3af99ed6),
	.w3(32'h3b5c075f),
	.w4(32'h3b2f322a),
	.w5(32'h3735a8f0),
	.w6(32'h39d00d59),
	.w7(32'h3b0b650f),
	.w8(32'h3b379821),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a021baa),
	.w1(32'h3b3338c5),
	.w2(32'h3b71758d),
	.w3(32'h3addab2c),
	.w4(32'hba66ff83),
	.w5(32'h3c5c14f6),
	.w6(32'hba5b362f),
	.w7(32'hba968b8a),
	.w8(32'h3c2cd16c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7880aa),
	.w1(32'h3c11aa74),
	.w2(32'h396ba2f4),
	.w3(32'h3cba074d),
	.w4(32'h3c8642dc),
	.w5(32'h3aa9d7b8),
	.w6(32'h3c971dc5),
	.w7(32'h3c5f4199),
	.w8(32'h3b3812e2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9209c),
	.w1(32'hbc4852a8),
	.w2(32'hbcc092cb),
	.w3(32'hbbd746c8),
	.w4(32'h3b192c42),
	.w5(32'hbc39bbc6),
	.w6(32'hbb951914),
	.w7(32'hbac0f2f0),
	.w8(32'hbc3b9878),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c3c86),
	.w1(32'h3be60c6e),
	.w2(32'h3b070beb),
	.w3(32'h3c35e1b2),
	.w4(32'h3c0b1968),
	.w5(32'h3b831628),
	.w6(32'h3bc1a252),
	.w7(32'h3bb1c004),
	.w8(32'hba3afb22),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38666796),
	.w1(32'h3ba5a5b2),
	.w2(32'h3bbd9c86),
	.w3(32'h3c3b7783),
	.w4(32'h3c2e19d3),
	.w5(32'hbbacb7f2),
	.w6(32'hb9d3767d),
	.w7(32'hbb4b22a8),
	.w8(32'hbb98989d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900ccde),
	.w1(32'h3a11d416),
	.w2(32'h3b9340ad),
	.w3(32'h3b3d8ed0),
	.w4(32'h3bf991cf),
	.w5(32'h3c4bfc86),
	.w6(32'h3bc166b4),
	.w7(32'h3bfca0f3),
	.w8(32'hbb44447a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47bebd),
	.w1(32'h3c1de44e),
	.w2(32'h3b2f0203),
	.w3(32'h3cd213c1),
	.w4(32'h3c888916),
	.w5(32'h39e186ab),
	.w6(32'h3c2a589f),
	.w7(32'h3be4a3ae),
	.w8(32'h3a81c19f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf10554),
	.w1(32'h3ba40b8b),
	.w2(32'h399b0949),
	.w3(32'h3c4100f2),
	.w4(32'h3995eb35),
	.w5(32'h3c6065dc),
	.w6(32'h3ad14daf),
	.w7(32'hbb044ab9),
	.w8(32'h3a700d4d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3760b6),
	.w1(32'h3c1c2b0a),
	.w2(32'hbc15b106),
	.w3(32'h3cb2941e),
	.w4(32'h3ca7a352),
	.w5(32'hbbcab1b3),
	.w6(32'h3c2d793e),
	.w7(32'h3b052481),
	.w8(32'hbc2abd59),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41795f),
	.w1(32'h3a53ac9b),
	.w2(32'h3c1e72ed),
	.w3(32'h3c07011e),
	.w4(32'h3b38ead7),
	.w5(32'h38bc5a61),
	.w6(32'hbbd200a7),
	.w7(32'hbb2498be),
	.w8(32'hbbfa183c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b330443),
	.w1(32'h38d335ee),
	.w2(32'hbb813950),
	.w3(32'h3a80527e),
	.w4(32'hba52b829),
	.w5(32'hbc786900),
	.w6(32'hbbce59c2),
	.w7(32'hbbcfa135),
	.w8(32'hbc66f0d5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06e189),
	.w1(32'hbbdca191),
	.w2(32'h3720b84f),
	.w3(32'hbc325dcb),
	.w4(32'hbc368052),
	.w5(32'h3b8e883a),
	.w6(32'h3bb5af02),
	.w7(32'h3c95be1d),
	.w8(32'hbc66b8c7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf590f0),
	.w1(32'hba25dcbd),
	.w2(32'h3aa8f799),
	.w3(32'hbafec2a6),
	.w4(32'h3abc6cd5),
	.w5(32'h3b508729),
	.w6(32'hbbf81e4e),
	.w7(32'hbc72d100),
	.w8(32'hbaf352db),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ee82e),
	.w1(32'h3b830d51),
	.w2(32'h3c47cfcc),
	.w3(32'h3c457952),
	.w4(32'h3bee90ac),
	.w5(32'hbb19d2f7),
	.w6(32'h3b08a48b),
	.w7(32'hbbcf5ec6),
	.w8(32'h3b978d12),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51a896),
	.w1(32'hbb25ff8d),
	.w2(32'hba782f2c),
	.w3(32'hbb271407),
	.w4(32'hbb3dc589),
	.w5(32'h3a8a99cf),
	.w6(32'h38985ba4),
	.w7(32'hb8518870),
	.w8(32'h3b23c9c0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb774b06e),
	.w1(32'h3b6299be),
	.w2(32'hbbb3d2c1),
	.w3(32'h3b458c9d),
	.w4(32'h3b9f4d59),
	.w5(32'h3bc199d0),
	.w6(32'h3b659fc9),
	.w7(32'h3b6cc45a),
	.w8(32'h3bcf319f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16906d),
	.w1(32'hbad16e6f),
	.w2(32'hbb30f245),
	.w3(32'hbaf61655),
	.w4(32'h3bb888cd),
	.w5(32'h3c317ec2),
	.w6(32'h3b02a13f),
	.w7(32'h3c4ec3d2),
	.w8(32'hbace3089),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f8bea),
	.w1(32'h3c36713c),
	.w2(32'h3ba1b35f),
	.w3(32'h3cccc37f),
	.w4(32'h3c5651ae),
	.w5(32'h3ae1e7bb),
	.w6(32'hbbf13d36),
	.w7(32'hbc9762c3),
	.w8(32'hbc68cf2d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c729017),
	.w1(32'h3caac632),
	.w2(32'hb9d9be90),
	.w3(32'h3d5e4b83),
	.w4(32'h3d5970f8),
	.w5(32'hbbc4b6b5),
	.w6(32'h3c9742f7),
	.w7(32'h3c9cdb54),
	.w8(32'hbc323c41),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3b8e0),
	.w1(32'hbb2e6dcb),
	.w2(32'h3b4aa0ae),
	.w3(32'h3bb4a68c),
	.w4(32'h3a97f742),
	.w5(32'hba88463a),
	.w6(32'h3c1be42c),
	.w7(32'h3bdb0a6c),
	.w8(32'hbac9cff7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aba65),
	.w1(32'hbc42335b),
	.w2(32'hbc10dabd),
	.w3(32'hba984c41),
	.w4(32'hbb3ca597),
	.w5(32'h3aa85352),
	.w6(32'h3c37b7cb),
	.w7(32'h3c4b3751),
	.w8(32'hbb1b529a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf96236),
	.w1(32'h3b7af4b5),
	.w2(32'hbc1dd4eb),
	.w3(32'h3c35a86c),
	.w4(32'h3c5ee128),
	.w5(32'hbc1f5561),
	.w6(32'h3be9178f),
	.w7(32'h3c0e8915),
	.w8(32'hbbfa58b2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12d32e),
	.w1(32'h3a1691c4),
	.w2(32'h3b2e1a46),
	.w3(32'hbab42f86),
	.w4(32'h3c01f9f2),
	.w5(32'h3b57d86f),
	.w6(32'hbbb4c232),
	.w7(32'h3c65e45e),
	.w8(32'h3a7231d4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb922b88f),
	.w1(32'h3b83b533),
	.w2(32'hbc3c23c8),
	.w3(32'hbb8949af),
	.w4(32'hbaf36d96),
	.w5(32'hbc8e92fe),
	.w6(32'hbbc7eb82),
	.w7(32'hbc0602a4),
	.w8(32'hbc84d24a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3c48e),
	.w1(32'hbc347513),
	.w2(32'h3bfdda04),
	.w3(32'hbc75c059),
	.w4(32'hbc776214),
	.w5(32'h3ba5aba1),
	.w6(32'hbc5582ac),
	.w7(32'hbc0e7f27),
	.w8(32'h3a78a8cf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb543cb1),
	.w1(32'hbb869f0f),
	.w2(32'h3b2f92a3),
	.w3(32'h3b611c3c),
	.w4(32'h3ba927a4),
	.w5(32'hbbe47a02),
	.w6(32'h3c00da8b),
	.w7(32'h3ac25b7f),
	.w8(32'hbab0774b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc082b80),
	.w1(32'h3aec21db),
	.w2(32'hbbdf6376),
	.w3(32'hbc337011),
	.w4(32'h38e683ab),
	.w5(32'hbc4e46df),
	.w6(32'hba5b9c09),
	.w7(32'h3a524465),
	.w8(32'hbbd05754),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc642a34),
	.w1(32'hbc6755bd),
	.w2(32'hbccfd897),
	.w3(32'hbd0c7152),
	.w4(32'hbc24146b),
	.w5(32'hbbfa8693),
	.w6(32'hbbd6949e),
	.w7(32'h3a52004f),
	.w8(32'hbb6de61f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7a227),
	.w1(32'hbb006277),
	.w2(32'h3c3a0eb6),
	.w3(32'hbb1738f5),
	.w4(32'hba466031),
	.w5(32'hbbb16085),
	.w6(32'h3b8b965e),
	.w7(32'h3aa0e76c),
	.w8(32'h3be40a8b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c902f67),
	.w1(32'h3c007e7f),
	.w2(32'hbb6dc656),
	.w3(32'h3c44c66e),
	.w4(32'h3c2e5777),
	.w5(32'hbbe3c303),
	.w6(32'hbb756695),
	.w7(32'hbb7af330),
	.w8(32'hbbbcb980),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd458d1),
	.w1(32'hbc17b71c),
	.w2(32'hbca20753),
	.w3(32'hbb12d283),
	.w4(32'hbc560403),
	.w5(32'hbc825293),
	.w6(32'hbb9e2447),
	.w7(32'hbae05181),
	.w8(32'hbc39e4b4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca12fbd),
	.w1(32'hbc2dee41),
	.w2(32'hb9fa1f8b),
	.w3(32'hbca9f745),
	.w4(32'h39905d49),
	.w5(32'hbaa35088),
	.w6(32'hbab9b246),
	.w7(32'h3ca6727d),
	.w8(32'hbb98fdc9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9197e9),
	.w1(32'hbbfa892b),
	.w2(32'h39ff9e94),
	.w3(32'h3bf4fb74),
	.w4(32'h3bb86c7e),
	.w5(32'hbbb7ad03),
	.w6(32'h399e224c),
	.w7(32'h3c0d7515),
	.w8(32'hbc3425d3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab23fc),
	.w1(32'hbbb1902b),
	.w2(32'hbc2bfa09),
	.w3(32'hbd00210a),
	.w4(32'hbcb679dc),
	.w5(32'h3bd873f0),
	.w6(32'hbc87cf40),
	.w7(32'hbc495fb1),
	.w8(32'hbc2a13b2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199c2c),
	.w1(32'h3bf62cfc),
	.w2(32'h3bf654fc),
	.w3(32'h3c0dc46d),
	.w4(32'h3bcea12d),
	.w5(32'h3beb00f0),
	.w6(32'h3bd67e69),
	.w7(32'hbba22aa7),
	.w8(32'hbbb52008),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c337e32),
	.w1(32'h3bd3d01f),
	.w2(32'h3bc40fd2),
	.w3(32'h3c1eb9d5),
	.w4(32'h3b4aff52),
	.w5(32'hbbad8700),
	.w6(32'h3b3db7e1),
	.w7(32'hbaa185a9),
	.w8(32'hb93c158e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ac07a),
	.w1(32'h3ba7d5c5),
	.w2(32'hbc0760cd),
	.w3(32'hbb8fca86),
	.w4(32'hbadf90fc),
	.w5(32'hbbb01e77),
	.w6(32'hbb319ece),
	.w7(32'hbc4c6b29),
	.w8(32'hba2de3ca),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf27ab4),
	.w1(32'hbbce6ce0),
	.w2(32'hbadb0ae7),
	.w3(32'h3b94a353),
	.w4(32'h3b0c0c25),
	.w5(32'hbba444c7),
	.w6(32'h3c7ed5fd),
	.w7(32'h3c0d2778),
	.w8(32'hbc0ffd68),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e2d79),
	.w1(32'hba99f667),
	.w2(32'hbc32cb94),
	.w3(32'h3ac960c7),
	.w4(32'h3adc01ed),
	.w5(32'hbc1b870a),
	.w6(32'hbb23e28b),
	.w7(32'h3a9d724b),
	.w8(32'hbb8d3f5b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a57c),
	.w1(32'hbbe6eaa0),
	.w2(32'hba7ba082),
	.w3(32'hb8d058f5),
	.w4(32'h3b8a044a),
	.w5(32'hba309193),
	.w6(32'h3c324866),
	.w7(32'h3bd1fbbb),
	.w8(32'h3a937225),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f1eb1),
	.w1(32'h390c56a2),
	.w2(32'hbc497288),
	.w3(32'hbbd2591b),
	.w4(32'h3a1e00c0),
	.w5(32'hbbcf0c98),
	.w6(32'hba60905e),
	.w7(32'hbb0839b3),
	.w8(32'hbc1c980d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc40ded),
	.w1(32'hbc3f1a6f),
	.w2(32'hbc46bc7e),
	.w3(32'hbc241872),
	.w4(32'hbb2f805c),
	.w5(32'hbbdd8331),
	.w6(32'hb907de08),
	.w7(32'h3ba7d0bb),
	.w8(32'h3b4c830e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ffb77),
	.w1(32'hbb1da3c3),
	.w2(32'hbb20cd0a),
	.w3(32'h3afd96d1),
	.w4(32'hba0dcb81),
	.w5(32'h3c186020),
	.w6(32'h3b50809a),
	.w7(32'hb9eae84a),
	.w8(32'h3a30bacd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98687c),
	.w1(32'hb9048eae),
	.w2(32'hba2949d7),
	.w3(32'h3cbf20bf),
	.w4(32'h3c996800),
	.w5(32'hbc127988),
	.w6(32'h3c855da8),
	.w7(32'h3c94d722),
	.w8(32'hbb3e986f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb105af6),
	.w1(32'hbaf33ff4),
	.w2(32'h3bcb8aec),
	.w3(32'hbbdc3a95),
	.w4(32'hbbbc7b8e),
	.w5(32'h3b96c623),
	.w6(32'h3724dee4),
	.w7(32'hba8ec55e),
	.w8(32'h3b070e8e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42b128),
	.w1(32'hba9cc7d6),
	.w2(32'h3b940e0d),
	.w3(32'hba0e9418),
	.w4(32'hbbc83505),
	.w5(32'h3bc18159),
	.w6(32'hba06b2fe),
	.w7(32'hbbe54073),
	.w8(32'hbb94fad9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf889ed),
	.w1(32'hbba50148),
	.w2(32'hbb3aaf6c),
	.w3(32'h3b0735cc),
	.w4(32'hbbf5c396),
	.w5(32'hbbf39da4),
	.w6(32'hbc7d9824),
	.w7(32'hbc94abbc),
	.w8(32'hbbef6e67),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba802219),
	.w1(32'hbc6aac15),
	.w2(32'hbbade2ce),
	.w3(32'hbad76d33),
	.w4(32'hbb77926d),
	.w5(32'hbb1b4228),
	.w6(32'hbb46eef2),
	.w7(32'h3b97ae3e),
	.w8(32'hbbec2e93),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33737b),
	.w1(32'hbc2e38a8),
	.w2(32'hbbb313b4),
	.w3(32'hbba5501c),
	.w4(32'h3adb4cdc),
	.w5(32'h3a21c46e),
	.w6(32'h3a0bfe52),
	.w7(32'hbc1c66b7),
	.w8(32'hbc09ba94),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5720df),
	.w1(32'h3c394b9f),
	.w2(32'h3b2d8130),
	.w3(32'h3cc849d4),
	.w4(32'h3c26e8dd),
	.w5(32'hbb9a8801),
	.w6(32'h3c83d0db),
	.w7(32'hb89d5694),
	.w8(32'hbbf99e52),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a7d32),
	.w1(32'h3abc049c),
	.w2(32'hba152fa3),
	.w3(32'hbbe5b500),
	.w4(32'hb9c0b89a),
	.w5(32'hbb0f81df),
	.w6(32'hbb9bad9e),
	.w7(32'h3bb5ecdb),
	.w8(32'h3b3656c2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ed348),
	.w1(32'hbbdcf99c),
	.w2(32'hbbc67f40),
	.w3(32'hbc023091),
	.w4(32'hbbd41409),
	.w5(32'hbb90c227),
	.w6(32'h3b66f46e),
	.w7(32'h3b55c6b9),
	.w8(32'h3a72984a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dbbb3),
	.w1(32'hbc1aef6d),
	.w2(32'hbaebfa79),
	.w3(32'hbc1d779b),
	.w4(32'hbc08aa5e),
	.w5(32'hbb17119f),
	.w6(32'hbb87072d),
	.w7(32'hbb9fb60b),
	.w8(32'hbb03b5f6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab02dbc),
	.w1(32'hbb98c867),
	.w2(32'hbba01ab3),
	.w3(32'h3bb68ff4),
	.w4(32'h3b8cc389),
	.w5(32'hbad55ab6),
	.w6(32'h3b009c37),
	.w7(32'hb9c13c73),
	.w8(32'hb939526b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb318d25),
	.w1(32'h3b33e109),
	.w2(32'hbc6b6d6b),
	.w3(32'hba6276d5),
	.w4(32'h3b380c1e),
	.w5(32'hbc916a00),
	.w6(32'h39b9fd8f),
	.w7(32'h3aec0014),
	.w8(32'hbbe22871),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc929029),
	.w1(32'hbc928f8e),
	.w2(32'hbc7ff995),
	.w3(32'hbca5ff76),
	.w4(32'hbbcab59b),
	.w5(32'hbc4d7e91),
	.w6(32'h3ac72798),
	.w7(32'h3c1a53b3),
	.w8(32'hbbb22ae8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e1ede),
	.w1(32'hbc53ddd9),
	.w2(32'hbcfad34c),
	.w3(32'hbc9a7879),
	.w4(32'hbb75181a),
	.w5(32'hbc7f82eb),
	.w6(32'hbc3340b5),
	.w7(32'hbb702747),
	.w8(32'hbc303968),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3af79a),
	.w1(32'hbc31846f),
	.w2(32'h3b958ac6),
	.w3(32'hbba079d7),
	.w4(32'h3a846a2c),
	.w5(32'hbbcbc43b),
	.w6(32'h3bd23540),
	.w7(32'h3c235ac1),
	.w8(32'hbbca42aa),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a953848),
	.w1(32'h3c077cc0),
	.w2(32'h3a55dba7),
	.w3(32'hbbf57d0d),
	.w4(32'hbb555d53),
	.w5(32'hba03513b),
	.w6(32'h3b2b205e),
	.w7(32'h39730713),
	.w8(32'hbb1185c9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c077f79),
	.w1(32'h3a39062a),
	.w2(32'h3bf25b24),
	.w3(32'h3ba51348),
	.w4(32'hb99ba362),
	.w5(32'hb9bdd493),
	.w6(32'h3bce12c6),
	.w7(32'hb900eae9),
	.w8(32'hbc04869d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab849d),
	.w1(32'h3aad031a),
	.w2(32'h3c058d9b),
	.w3(32'hbb316c35),
	.w4(32'hbb68ae01),
	.w5(32'h3b6350e8),
	.w6(32'hbbd3fb63),
	.w7(32'hbb8e758e),
	.w8(32'hbbcabe89),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd93a66),
	.w1(32'h3a25a4d4),
	.w2(32'hbc2439ab),
	.w3(32'hbb5e6490),
	.w4(32'hbb9f8c04),
	.w5(32'h3b6a59e0),
	.w6(32'hbc4e02e1),
	.w7(32'hbc60bbc8),
	.w8(32'h3c09dc17),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec7fec),
	.w1(32'hbbc72b1b),
	.w2(32'hbbbf5ef5),
	.w3(32'h3b57fb25),
	.w4(32'hbbbcf592),
	.w5(32'h3b670ca6),
	.w6(32'h3b9de28c),
	.w7(32'hbbee7ba0),
	.w8(32'h3c19eb4d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc490f22),
	.w1(32'hbc55f46d),
	.w2(32'hbbef6b7f),
	.w3(32'h38ca7826),
	.w4(32'hbbc8e84a),
	.w5(32'hbb2ba2b8),
	.w6(32'h3c0bf325),
	.w7(32'h3c7c6ca4),
	.w8(32'h3bf767f9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7824b),
	.w1(32'h3bad4e5b),
	.w2(32'hbc42faec),
	.w3(32'hbb800a48),
	.w4(32'h3b83e885),
	.w5(32'h394fe24d),
	.w6(32'h3bce8de2),
	.w7(32'h3adc8454),
	.w8(32'h3c80be41),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb740a9),
	.w1(32'hbca2c6b9),
	.w2(32'h3bf23a16),
	.w3(32'h3caa276a),
	.w4(32'h3c093434),
	.w5(32'h3c493c46),
	.w6(32'h3d3308c5),
	.w7(32'h3bb8d243),
	.w8(32'h3c562f26),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f6a31),
	.w1(32'hbc287e46),
	.w2(32'h3bcf4bcc),
	.w3(32'h3c13287e),
	.w4(32'hbbead125),
	.w5(32'h39c4effc),
	.w6(32'h3c0236be),
	.w7(32'hbabacdb2),
	.w8(32'hbb5d16e1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1129fd),
	.w1(32'hbb2f0103),
	.w2(32'hbb87fdb9),
	.w3(32'hb94d821f),
	.w4(32'hba9394fc),
	.w5(32'hbbdcdb49),
	.w6(32'hbae9de75),
	.w7(32'h3a341cf4),
	.w8(32'hbbd57e53),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22b574),
	.w1(32'hbc19b4b3),
	.w2(32'h3be52330),
	.w3(32'hbc20c505),
	.w4(32'hbb107cc1),
	.w5(32'h3bd69ffc),
	.w6(32'h3c0b19f5),
	.w7(32'h3b5e8592),
	.w8(32'hbc077cc3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba4d0a),
	.w1(32'hbc04df50),
	.w2(32'hbc609c28),
	.w3(32'hbbf87b02),
	.w4(32'hba954a5b),
	.w5(32'hbc438229),
	.w6(32'hbca3b040),
	.w7(32'hbc88d728),
	.w8(32'hbcbfa8ee),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3405e1),
	.w1(32'h3bff0600),
	.w2(32'h3bb5c10b),
	.w3(32'hbcb2da59),
	.w4(32'hbcd76fc3),
	.w5(32'h3bd09b18),
	.w6(32'hbce48928),
	.w7(32'hbcc432ba),
	.w8(32'h3a037e96),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3154ef),
	.w1(32'h3c200d52),
	.w2(32'hbb2a8f1e),
	.w3(32'hbb98d4f2),
	.w4(32'h3b6f10bf),
	.w5(32'h3b3bda1f),
	.w6(32'hbb87f9bf),
	.w7(32'h3b510882),
	.w8(32'hbb4ac1e3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd41400),
	.w1(32'h3b99c05a),
	.w2(32'h3b47c061),
	.w3(32'h3c3e40f8),
	.w4(32'h3bad43d9),
	.w5(32'hbbc0edbe),
	.w6(32'h3bdf99bf),
	.w7(32'hb9f34ae0),
	.w8(32'hbbdb2af7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97e165),
	.w1(32'hbbcceab6),
	.w2(32'h3a1a94f4),
	.w3(32'hbc14006f),
	.w4(32'hbc128796),
	.w5(32'hbc136b12),
	.w6(32'hbba7b324),
	.w7(32'hbb43414b),
	.w8(32'hbc270930),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb6036),
	.w1(32'hbb0a0ef5),
	.w2(32'h3a99f5f5),
	.w3(32'h3bb231de),
	.w4(32'hbb41ad86),
	.w5(32'hbc1e71d3),
	.w6(32'h3b986e49),
	.w7(32'h3aa50958),
	.w8(32'hbb6b43f0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6eb56),
	.w1(32'hbbfc0993),
	.w2(32'h3bb4040a),
	.w3(32'hbc543158),
	.w4(32'hbc5f37dc),
	.w5(32'hbb855da2),
	.w6(32'hbbf9dd37),
	.w7(32'hbc95e981),
	.w8(32'h3a0b5647),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8de530),
	.w1(32'h3ba0f9be),
	.w2(32'hba703d8f),
	.w3(32'h393ca04f),
	.w4(32'h3c2fec61),
	.w5(32'h39aa5286),
	.w6(32'hb786747a),
	.w7(32'hbb8d510e),
	.w8(32'hbae413c5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814e71),
	.w1(32'h3b3d34f9),
	.w2(32'hbc8c88bb),
	.w3(32'hbbfa4729),
	.w4(32'h3bd55d0e),
	.w5(32'hbc5a117c),
	.w6(32'hbb0f4194),
	.w7(32'h3b04d86a),
	.w8(32'hbbb6c661),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71fbff),
	.w1(32'hbbcce66e),
	.w2(32'h3b4bd885),
	.w3(32'h3baf91ef),
	.w4(32'hbb0d80b6),
	.w5(32'h3babeafc),
	.w6(32'h3c5cf42b),
	.w7(32'hb997dada),
	.w8(32'hbbd7b01c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba982eb9),
	.w1(32'hbbdfc672),
	.w2(32'hbca37af5),
	.w3(32'hbcd31635),
	.w4(32'hbb88e541),
	.w5(32'h3b0600a5),
	.w6(32'hbd071aaf),
	.w7(32'hbc3444b8),
	.w8(32'h3b52e1e7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8007d9),
	.w1(32'h3c0efb76),
	.w2(32'h3b920133),
	.w3(32'h3bf0d57f),
	.w4(32'h3c5a6c72),
	.w5(32'hbc9d4e70),
	.w6(32'h3bca12f2),
	.w7(32'h3c0bb3e6),
	.w8(32'hbbba853c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0c6c4),
	.w1(32'h3b867357),
	.w2(32'h3bcea160),
	.w3(32'hba00145e),
	.w4(32'hbb7a9c3a),
	.w5(32'hbb904981),
	.w6(32'h3c79f77c),
	.w7(32'h3c36634c),
	.w8(32'hbbdce648),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb168616),
	.w1(32'h3a4017d4),
	.w2(32'h3bac1b99),
	.w3(32'hbb250eae),
	.w4(32'h3c927713),
	.w5(32'h3c15c96a),
	.w6(32'hbb982914),
	.w7(32'h3c5d6ae8),
	.w8(32'hbc025d4c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d80aa),
	.w1(32'hbb18227a),
	.w2(32'h3ade1638),
	.w3(32'hbcad0362),
	.w4(32'hbcb9542a),
	.w5(32'hbb9de4c3),
	.w6(32'hbcebd8ae),
	.w7(32'hbcc36813),
	.w8(32'h3b0e4db1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccab97b),
	.w1(32'hbc859e83),
	.w2(32'hbce9455e),
	.w3(32'hbc9b9b4a),
	.w4(32'hbca57b69),
	.w5(32'hbb6a43ad),
	.w6(32'hbbc95be0),
	.w7(32'hbbca5eeb),
	.w8(32'h3bc9306d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9739ac),
	.w1(32'hbbb530c8),
	.w2(32'h3bb3a48b),
	.w3(32'h3bd47177),
	.w4(32'h3bc4ee12),
	.w5(32'h3c060a6f),
	.w6(32'h3c82bc5e),
	.w7(32'h3c3a1b0b),
	.w8(32'h3c40db34),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb948a203),
	.w1(32'hb96f18f6),
	.w2(32'h3ac60c19),
	.w3(32'h3bba3400),
	.w4(32'h3ac99d22),
	.w5(32'hbbf404f9),
	.w6(32'h3c8a3615),
	.w7(32'h3c1b1964),
	.w8(32'hbbe97802),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2674b1),
	.w1(32'h3c0dc030),
	.w2(32'hbb464e23),
	.w3(32'hbab677eb),
	.w4(32'h3c8aa437),
	.w5(32'hb9b835b6),
	.w6(32'h3b1e4682),
	.w7(32'h3bf5dafc),
	.w8(32'h3b1d1101),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46d249),
	.w1(32'h3c2dfe80),
	.w2(32'hba10a0dd),
	.w3(32'hbabb9f4c),
	.w4(32'h3a7ae23e),
	.w5(32'h3a06dee2),
	.w6(32'h3b29053f),
	.w7(32'hbb5a0c91),
	.w8(32'hbbbd41e1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba84ec7),
	.w1(32'hbbc1be15),
	.w2(32'h3bbe8692),
	.w3(32'h3bd40fd2),
	.w4(32'h3bfbcc23),
	.w5(32'h3b3eca6c),
	.w6(32'h3bd2330e),
	.w7(32'h3ba04e92),
	.w8(32'h3b87d841),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00d950),
	.w1(32'hbbfb0805),
	.w2(32'hbc369082),
	.w3(32'h3994fc7d),
	.w4(32'hb9cc8326),
	.w5(32'hbc381381),
	.w6(32'h3b5da3ac),
	.w7(32'h3932885e),
	.w8(32'hbae9c6bd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b8416),
	.w1(32'hbc16e6bb),
	.w2(32'h3c33f819),
	.w3(32'hbc312ce8),
	.w4(32'hbbd9e59c),
	.w5(32'h3b9f7ebb),
	.w6(32'hb9762022),
	.w7(32'hbbea5b71),
	.w8(32'hbbd6e3d9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3d598),
	.w1(32'h3a08209b),
	.w2(32'h3ae40d71),
	.w3(32'hbb6f5e13),
	.w4(32'hb9d2e924),
	.w5(32'hbb9b80a0),
	.w6(32'hbc352443),
	.w7(32'h3b827304),
	.w8(32'h39c76a5d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dddd3),
	.w1(32'hbc3921ef),
	.w2(32'hbcaa8d8b),
	.w3(32'hbc131234),
	.w4(32'hbbb9d60f),
	.w5(32'hbc936a4a),
	.w6(32'h3a24e0d7),
	.w7(32'h3c1e2163),
	.w8(32'hbc2aab09),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc273dec),
	.w1(32'hbbd575e3),
	.w2(32'h3bdea04d),
	.w3(32'hbc68ef85),
	.w4(32'hbc6ee357),
	.w5(32'h3c0a4ea7),
	.w6(32'hbba0a541),
	.w7(32'hbbb6ae20),
	.w8(32'hbbb6f058),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18aac1),
	.w1(32'h3c98e50d),
	.w2(32'h3aeb2bf7),
	.w3(32'h3ca9c9fe),
	.w4(32'h3cd047c0),
	.w5(32'h3ba0eed9),
	.w6(32'h3aa79c9f),
	.w7(32'h3ba62094),
	.w8(32'hbb25b297),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f84e0f),
	.w1(32'hbb77572f),
	.w2(32'hba7284ea),
	.w3(32'hbb98d011),
	.w4(32'hbc15e562),
	.w5(32'h3bf67b94),
	.w6(32'hbbb7fd1c),
	.w7(32'hbbfa858d),
	.w8(32'hbbc32cdb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bec39),
	.w1(32'h3b9d2c79),
	.w2(32'hbbae5871),
	.w3(32'h3ca49281),
	.w4(32'h3caaab45),
	.w5(32'hbbec9319),
	.w6(32'h3c0d1278),
	.w7(32'h3c5f62ae),
	.w8(32'h3be9890a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf42917),
	.w1(32'hba2ac312),
	.w2(32'hbb26d127),
	.w3(32'h3c6c44bc),
	.w4(32'h3c9c7433),
	.w5(32'hbb65c927),
	.w6(32'h3c71e1bb),
	.w7(32'h3bcc4aa2),
	.w8(32'hbb9a1e33),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ffbb1),
	.w1(32'h3b79e36a),
	.w2(32'h3b8775fb),
	.w3(32'h3b266549),
	.w4(32'hbace9209),
	.w5(32'h3b692c9e),
	.w6(32'h3bfb897a),
	.w7(32'h3c441216),
	.w8(32'h3a971567),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d3d06),
	.w1(32'hbb880d42),
	.w2(32'hba4e8a4d),
	.w3(32'h3a9fd2a6),
	.w4(32'h3b4ccc65),
	.w5(32'hb9a0d210),
	.w6(32'h3a73fe06),
	.w7(32'hba166cea),
	.w8(32'hbb20b7c3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4370),
	.w1(32'hbb0ea36c),
	.w2(32'hbb28d246),
	.w3(32'hbb3b7826),
	.w4(32'hba9bb0c0),
	.w5(32'hbb3973d9),
	.w6(32'hbbf6b198),
	.w7(32'hbbbad034),
	.w8(32'hbb5757d9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2ed82),
	.w1(32'hba759df0),
	.w2(32'hbc0a0cca),
	.w3(32'h3a582c1b),
	.w4(32'hbb23e3c9),
	.w5(32'hbc46c6bf),
	.w6(32'h3b726936),
	.w7(32'hbaa06b28),
	.w8(32'hbbee192e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d947c),
	.w1(32'hbc1b2c79),
	.w2(32'hba45b92d),
	.w3(32'hb9a5d55a),
	.w4(32'hba6a2d52),
	.w5(32'h3c3dd0e2),
	.w6(32'h3b60fdf8),
	.w7(32'h3c3f39a1),
	.w8(32'h3c23a2d7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ea2d),
	.w1(32'hb9e46361),
	.w2(32'hbb6cd299),
	.w3(32'h3c9d16cb),
	.w4(32'h3c46c1a8),
	.w5(32'hbbb9101e),
	.w6(32'h3c9631f2),
	.w7(32'h3c455850),
	.w8(32'h3b8da04b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab965d4),
	.w1(32'hbc0a072b),
	.w2(32'hba3ce75b),
	.w3(32'h3bcc901a),
	.w4(32'h3bcec7bf),
	.w5(32'hbb64d7f8),
	.w6(32'h3c88bda3),
	.w7(32'h3c490c0c),
	.w8(32'hbb7ad4b7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe012a5),
	.w1(32'hbb107795),
	.w2(32'h3a03640a),
	.w3(32'hbb84d477),
	.w4(32'hbb32ce50),
	.w5(32'hbb42968f),
	.w6(32'h3981a9c7),
	.w7(32'h3b571a10),
	.w8(32'hbbe84bcd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b823f),
	.w1(32'hbc15ac47),
	.w2(32'hbc2d84ec),
	.w3(32'hbbf3a64f),
	.w4(32'hbbda6d60),
	.w5(32'hbd0a3353),
	.w6(32'h3b49b15e),
	.w7(32'hbb5edeb4),
	.w8(32'hbb4ac4b3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc963bc9),
	.w1(32'hbc01aec0),
	.w2(32'hbba5ac12),
	.w3(32'hbc9ff0dc),
	.w4(32'hbb9ffeaa),
	.w5(32'hbc2ca02a),
	.w6(32'h3c36ecc8),
	.w7(32'h3c490042),
	.w8(32'hbc324bf5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba10589),
	.w1(32'h3a0db010),
	.w2(32'h3b6cf429),
	.w3(32'hbc56e5c1),
	.w4(32'hbba01257),
	.w5(32'h3c2b6953),
	.w6(32'hbc03330d),
	.w7(32'hbc1292cf),
	.w8(32'hbb18bfd6),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e630),
	.w1(32'h3b029b1b),
	.w2(32'hbb2b7abd),
	.w3(32'h3b20f857),
	.w4(32'hbc3985ed),
	.w5(32'hba94ddcf),
	.w6(32'hbc512230),
	.w7(32'hbc40ea05),
	.w8(32'h3b0a37e5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb515774),
	.w1(32'h3bfb0fc4),
	.w2(32'hbb82a000),
	.w3(32'h398c9827),
	.w4(32'h3b61a6a4),
	.w5(32'h3c5ad164),
	.w6(32'h3b9d0ef5),
	.w7(32'h3b91d25a),
	.w8(32'h3b231700),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c29fb),
	.w1(32'h3bc337a4),
	.w2(32'h3bd684d1),
	.w3(32'h3d011986),
	.w4(32'h3caef300),
	.w5(32'h3973b16c),
	.w6(32'h3bd726d0),
	.w7(32'hbbffe8e6),
	.w8(32'hb6f0fbae),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc024c35),
	.w1(32'hbb08610f),
	.w2(32'h3c602d43),
	.w3(32'hbb99a9ee),
	.w4(32'hbb315be9),
	.w5(32'h3bf21380),
	.w6(32'h3ad381a8),
	.w7(32'hbabe9f15),
	.w8(32'h3bbc719b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84cd7d),
	.w1(32'h3b60ec84),
	.w2(32'hbca6692f),
	.w3(32'hbc08fa93),
	.w4(32'h3a44169c),
	.w5(32'h3a665de3),
	.w6(32'hbc0e2bde),
	.w7(32'hbbb5f52b),
	.w8(32'hbc3ae9dc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d90be),
	.w1(32'hbb18c2f5),
	.w2(32'h3c12200c),
	.w3(32'h3cbd7c97),
	.w4(32'h3c5d6f04),
	.w5(32'hbb6604a1),
	.w6(32'h3c5dbc21),
	.w7(32'h3a9291c0),
	.w8(32'hbbf00fa8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb241612),
	.w1(32'hbba5b017),
	.w2(32'hbc0869be),
	.w3(32'hbc70b390),
	.w4(32'hbc8bf8ab),
	.w5(32'hbab09e92),
	.w6(32'hbc3abd63),
	.w7(32'hbc3ecbfb),
	.w8(32'h3a8b8a03),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab24899),
	.w1(32'h3b89df4e),
	.w2(32'hbbc005c3),
	.w3(32'h3b5ee6a2),
	.w4(32'h3c30f485),
	.w5(32'hba931b77),
	.w6(32'h3c0d1e6e),
	.w7(32'h3c54bfb0),
	.w8(32'hbb88603e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafffcc6),
	.w1(32'h3afcc01e),
	.w2(32'h3b9660b8),
	.w3(32'hbabd2e40),
	.w4(32'h3a32dc97),
	.w5(32'hbbf66482),
	.w6(32'hbbb5741d),
	.w7(32'hbacd59c3),
	.w8(32'hbb388bfe),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb237b27),
	.w1(32'hba80b354),
	.w2(32'hbc353474),
	.w3(32'hbbe7c936),
	.w4(32'hbb1cead2),
	.w5(32'hbc162682),
	.w6(32'h3a5d6d7d),
	.w7(32'h3bde320d),
	.w8(32'hbb897fec),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11fc14),
	.w1(32'hbbde2f96),
	.w2(32'h3b03cbfd),
	.w3(32'hbbc48925),
	.w4(32'h39e48239),
	.w5(32'h3b84d43f),
	.w6(32'h3be06a16),
	.w7(32'h3c17650e),
	.w8(32'h398547cd),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed6edb),
	.w1(32'h3c1ba77c),
	.w2(32'hbbea388e),
	.w3(32'h3bb2c90f),
	.w4(32'h3c096b10),
	.w5(32'hbba81f4b),
	.w6(32'h3c1d0e16),
	.w7(32'h390f3310),
	.w8(32'h3be85bbc),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca8c4e),
	.w1(32'hbc9b36f7),
	.w2(32'h3a89dcdc),
	.w3(32'hbc632897),
	.w4(32'hbbe962e5),
	.w5(32'hbb32065c),
	.w6(32'h3bab8743),
	.w7(32'h3b8233d4),
	.w8(32'hbc238230),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b375e0c),
	.w1(32'h3ba231c8),
	.w2(32'h3b596f4e),
	.w3(32'h3be7e005),
	.w4(32'h3c173e1a),
	.w5(32'h39e6fcdd),
	.w6(32'h3a4a0c59),
	.w7(32'h3bc4f0bb),
	.w8(32'hbae5432a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26dd1a),
	.w1(32'h3b05af06),
	.w2(32'h3c77a3fe),
	.w3(32'h38b41e52),
	.w4(32'hba16c497),
	.w5(32'h3abe2e66),
	.w6(32'hbaa2d739),
	.w7(32'h3823db8e),
	.w8(32'h3a940cbe),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd99f0f),
	.w1(32'h3cb41c84),
	.w2(32'h3bc9a53b),
	.w3(32'hbbc3cccf),
	.w4(32'hbb5608bd),
	.w5(32'h3a8ff473),
	.w6(32'hbc38df0a),
	.w7(32'hbca93cb3),
	.w8(32'h3aa3380e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb874cf5),
	.w1(32'h3b2b9b88),
	.w2(32'h3b29963c),
	.w3(32'hbb47fab9),
	.w4(32'h3a90b1c7),
	.w5(32'h3c1187b1),
	.w6(32'hbb45af94),
	.w7(32'hba3576b7),
	.w8(32'h3b96363f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c234751),
	.w1(32'h3b7b10da),
	.w2(32'h3c88a639),
	.w3(32'h3c1db02b),
	.w4(32'h3c821745),
	.w5(32'h3c0a9d63),
	.w6(32'h3cbb8295),
	.w7(32'h3c2eb63e),
	.w8(32'hbb322610),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03306a),
	.w1(32'h3a518063),
	.w2(32'hbad6495f),
	.w3(32'hbb725cd9),
	.w4(32'hbc143420),
	.w5(32'h3aae89ce),
	.w6(32'hbc58d270),
	.w7(32'hbc40465c),
	.w8(32'hbb5bf333),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39748d0a),
	.w1(32'h3c676080),
	.w2(32'hbc1b8937),
	.w3(32'hbb8b75f9),
	.w4(32'hbb2d6920),
	.w5(32'hbc122057),
	.w6(32'h3b840361),
	.w7(32'h3bb1630d),
	.w8(32'hbc1f2f84),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0173dc),
	.w1(32'hbc0ad7b0),
	.w2(32'h38b681b1),
	.w3(32'hb88c8fe8),
	.w4(32'h3ad0ba09),
	.w5(32'hbb10e0fe),
	.w6(32'h3bc59d9d),
	.w7(32'h3b1868a6),
	.w8(32'hbb0818f3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61d200),
	.w1(32'hbac35c0d),
	.w2(32'hbbe1bdc8),
	.w3(32'h3a4f9a54),
	.w4(32'h3bc73899),
	.w5(32'h3ba843c6),
	.w6(32'h3aae9b49),
	.w7(32'h3ba1a43f),
	.w8(32'h39ce4c86),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0695b7),
	.w1(32'hbb6bbef3),
	.w2(32'hbc18a879),
	.w3(32'h3c2f768b),
	.w4(32'h3bcd34ff),
	.w5(32'hbc5c8447),
	.w6(32'h3c5c7927),
	.w7(32'h3b8f08b7),
	.w8(32'hba115f63),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aed4d),
	.w1(32'hbc52a06c),
	.w2(32'hbbb4be44),
	.w3(32'hbb99d670),
	.w4(32'h39de5c82),
	.w5(32'hbc89b196),
	.w6(32'hbbc37d59),
	.w7(32'hbb195af7),
	.w8(32'hbc1af19b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf23078),
	.w1(32'hbc0747a7),
	.w2(32'h3bba2222),
	.w3(32'hbb9c28d9),
	.w4(32'hbb3b8840),
	.w5(32'h3b8ef315),
	.w6(32'h3b28e48f),
	.w7(32'h3b40f119),
	.w8(32'h3bba5fbf),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbd791),
	.w1(32'h3bb55e06),
	.w2(32'h3bc9aa10),
	.w3(32'h3b9c8871),
	.w4(32'h3ba62808),
	.w5(32'h3bb3d2f8),
	.w6(32'h3b3a84e9),
	.w7(32'h3b8fc896),
	.w8(32'h3abe7d99),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb241031),
	.w1(32'hbae33591),
	.w2(32'h3bb6b20f),
	.w3(32'h3c0b52aa),
	.w4(32'h3bbae72a),
	.w5(32'h3bda9b25),
	.w6(32'h3beb199d),
	.w7(32'h3b78ebc8),
	.w8(32'h39c18d44),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9ca44),
	.w1(32'h3c030b8c),
	.w2(32'hbcd056c0),
	.w3(32'h3b2df323),
	.w4(32'h3b16ccc3),
	.w5(32'hbc13d995),
	.w6(32'h3b9bd228),
	.w7(32'h3bf09a37),
	.w8(32'hbc991095),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48686b),
	.w1(32'hbccebb15),
	.w2(32'hbb902745),
	.w3(32'h3c8f0fb8),
	.w4(32'h3b26e654),
	.w5(32'hbb32212d),
	.w6(32'h3b4f216e),
	.w7(32'hbc1822ad),
	.w8(32'h3ab74805),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03c46f),
	.w1(32'hbafad9ce),
	.w2(32'h3b809633),
	.w3(32'h3c1ecde9),
	.w4(32'h3b506d56),
	.w5(32'hba01a515),
	.w6(32'h3c1ea1be),
	.w7(32'h3b377b71),
	.w8(32'hbb2d59ff),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c52c8),
	.w1(32'h3c22350f),
	.w2(32'hbce0c879),
	.w3(32'h39476d58),
	.w4(32'h3acdf0d8),
	.w5(32'h3b89fc6d),
	.w6(32'h3b2d7b43),
	.w7(32'hbb223c4a),
	.w8(32'hbc556664),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb81bc2),
	.w1(32'hbce3177f),
	.w2(32'hbc0c137f),
	.w3(32'h3d251fb7),
	.w4(32'h3c1c0bd7),
	.w5(32'hbc9c7356),
	.w6(32'h3c95729b),
	.w7(32'hbc11911d),
	.w8(32'hbbdba2f4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc48b0),
	.w1(32'hbc073050),
	.w2(32'h3ac757a4),
	.w3(32'hbc386bb0),
	.w4(32'h3b10b89c),
	.w5(32'hbb948b16),
	.w6(32'hbbff3631),
	.w7(32'h3c220b4b),
	.w8(32'hbba92611),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda07cf),
	.w1(32'hbb22ba04),
	.w2(32'hbaec5b89),
	.w3(32'hbc8f64cc),
	.w4(32'hbc50c972),
	.w5(32'hbb9b5ac0),
	.w6(32'hbc5b665b),
	.w7(32'hbc02cfef),
	.w8(32'hbc4ee651),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87133a),
	.w1(32'h3b0f62ba),
	.w2(32'h3cc7104d),
	.w3(32'h3c332907),
	.w4(32'hba9aa11e),
	.w5(32'h3d817d1b),
	.w6(32'hbbf62c94),
	.w7(32'hbc29bf1f),
	.w8(32'h3d39b668),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3c43ec),
	.w1(32'h3ca96847),
	.w2(32'h3b5cfdf6),
	.w3(32'h3dcf4e5f),
	.w4(32'h3d866054),
	.w5(32'hbba13b0d),
	.w6(32'h3dacb0cd),
	.w7(32'h3d4a4ba7),
	.w8(32'h39e09c6c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8508e),
	.w1(32'h3c2cb73d),
	.w2(32'hbbb4d9b5),
	.w3(32'hb99ac588),
	.w4(32'h3bca5158),
	.w5(32'h3b2189fb),
	.w6(32'hbb5424ab),
	.w7(32'hba1f62c8),
	.w8(32'h3c90f61f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc809206),
	.w1(32'hbc7298a5),
	.w2(32'h3b730a3b),
	.w3(32'hbba3f1e8),
	.w4(32'hbc3d02a0),
	.w5(32'hbba98132),
	.w6(32'h3baba912),
	.w7(32'hbc112221),
	.w8(32'hba891587),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cebb8),
	.w1(32'h3be758a9),
	.w2(32'hbc18f2f4),
	.w3(32'hbc1f1208),
	.w4(32'hbb67b4ac),
	.w5(32'hbbb356ce),
	.w6(32'hbc4e6fab),
	.w7(32'hbbe3798e),
	.w8(32'hbc4407a7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b165201),
	.w1(32'h3bd510be),
	.w2(32'h3b3e9fed),
	.w3(32'h3bf0c81e),
	.w4(32'hb9c11456),
	.w5(32'h3b8966f9),
	.w6(32'hbc28a414),
	.w7(32'hbbf371ef),
	.w8(32'h3aa6e010),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8332a6),
	.w1(32'h3c69fb5e),
	.w2(32'h3ce7193f),
	.w3(32'h3c33ad2f),
	.w4(32'h3baa0522),
	.w5(32'h3c55308e),
	.w6(32'h3be67db7),
	.w7(32'h3a142cd7),
	.w8(32'h3c99f09f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b647a),
	.w1(32'h3ce9fd7c),
	.w2(32'hba533531),
	.w3(32'h3a75f51e),
	.w4(32'h3c7eb137),
	.w5(32'hbc484da2),
	.w6(32'h3c3e2243),
	.w7(32'h3cc6ed7f),
	.w8(32'hbc0bbc56),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db21d),
	.w1(32'h3c00c67b),
	.w2(32'hbb097041),
	.w3(32'hbbf50f22),
	.w4(32'h3b3e9d92),
	.w5(32'h3b351a3c),
	.w6(32'hba9f6689),
	.w7(32'h3b777db0),
	.w8(32'h3af57b7c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bdafd),
	.w1(32'hbb96575a),
	.w2(32'hbbf60e6e),
	.w3(32'hbb7b7b5d),
	.w4(32'hbc1225b4),
	.w5(32'hbc062e90),
	.w6(32'hbb1f0969),
	.w7(32'hbc093cdc),
	.w8(32'hbc48f870),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23e502),
	.w1(32'hbb27f398),
	.w2(32'hbc1c54b4),
	.w3(32'hbbb6eae3),
	.w4(32'h3b218f41),
	.w5(32'hbcc06aaf),
	.w6(32'h3ac0cf6c),
	.w7(32'hba172e23),
	.w8(32'hbca0ed95),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c78de),
	.w1(32'h3becb93d),
	.w2(32'h3c30e21d),
	.w3(32'hbc5b37b8),
	.w4(32'h3c3dc6d9),
	.w5(32'hbaca632c),
	.w6(32'hbc3e383c),
	.w7(32'h3bf78806),
	.w8(32'h3c0fad4f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d4488),
	.w1(32'h3be7a868),
	.w2(32'hbb711218),
	.w3(32'hbcb4ddb4),
	.w4(32'hbc10c4f6),
	.w5(32'h3b029b8e),
	.w6(32'hbbdae731),
	.w7(32'h3b9dbdc1),
	.w8(32'h3b33e2d0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03455),
	.w1(32'hbc1781d0),
	.w2(32'hbb798a89),
	.w3(32'h3ab8a941),
	.w4(32'hbc2215e8),
	.w5(32'hbb6d1875),
	.w6(32'h3c0f273a),
	.w7(32'h3ae633ae),
	.w8(32'hbb26e1b8),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17a293),
	.w1(32'hbb234e33),
	.w2(32'h3be26a08),
	.w3(32'h3c0397f0),
	.w4(32'h3903f769),
	.w5(32'h3bb445b8),
	.w6(32'h3afea10c),
	.w7(32'hbb86a382),
	.w8(32'hba6d9f7a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba11dc5),
	.w1(32'h3a3354b4),
	.w2(32'hbbed6bfb),
	.w3(32'h3af0f0f1),
	.w4(32'h3c16b28a),
	.w5(32'hbaf2e26a),
	.w6(32'h3b83acfa),
	.w7(32'h3b81a94d),
	.w8(32'hbb821c10),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54f713),
	.w1(32'hbbdf6aef),
	.w2(32'h3c982e66),
	.w3(32'h3b8736f5),
	.w4(32'hbc1eb552),
	.w5(32'h3c4c6f07),
	.w6(32'hbb6fb609),
	.w7(32'hbbfaec39),
	.w8(32'hbb04ef00),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca40113),
	.w1(32'h3c6e56ef),
	.w2(32'h39d69a2b),
	.w3(32'h3c8ef2a7),
	.w4(32'h3c467711),
	.w5(32'h3b5be297),
	.w6(32'h3ba198d8),
	.w7(32'h3bd6ccfd),
	.w8(32'hbc05833c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d2c68),
	.w1(32'hbbfaa6a4),
	.w2(32'h398814e8),
	.w3(32'h3c747d66),
	.w4(32'h3b283b78),
	.w5(32'hbb114a3b),
	.w6(32'hbbaf9376),
	.w7(32'hbc1ac5c4),
	.w8(32'h3bf936b8),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae40e39),
	.w1(32'hbae208d8),
	.w2(32'hbb8b923e),
	.w3(32'h3b1b031c),
	.w4(32'h3be8bd38),
	.w5(32'h3b732f5d),
	.w6(32'h3bedbc46),
	.w7(32'h3c7ad395),
	.w8(32'h3b67cf37),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4be045),
	.w1(32'h3bd24f10),
	.w2(32'hbcd6c77c),
	.w3(32'h3c29f1cb),
	.w4(32'h3b2c94d3),
	.w5(32'hbceeabb0),
	.w6(32'h3b7ddaf0),
	.w7(32'hba06c30d),
	.w8(32'hbcbc3a28),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31b847),
	.w1(32'h3c44d7c1),
	.w2(32'h3c367056),
	.w3(32'hbc1073b8),
	.w4(32'h3cd4b622),
	.w5(32'h3ca673b5),
	.w6(32'h3b572c63),
	.w7(32'h3d1d3f04),
	.w8(32'h3c2d3d77),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ebbfc),
	.w1(32'h3a9b5a32),
	.w2(32'hbc78fd02),
	.w3(32'h3d02a06f),
	.w4(32'h3c7d9bc1),
	.w5(32'hbbe7af6f),
	.w6(32'h3c9c5057),
	.w7(32'h3bd836ee),
	.w8(32'h3cafe772),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd06025),
	.w1(32'hbcd13c39),
	.w2(32'hbc82a91e),
	.w3(32'hbc15cf15),
	.w4(32'hbc05c777),
	.w5(32'hbcad3062),
	.w6(32'h3d05f4a9),
	.w7(32'h3ccff0ee),
	.w8(32'hbc5249fd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ce13f),
	.w1(32'h3bd1275f),
	.w2(32'h3c2e6ebe),
	.w3(32'h3be11f7b),
	.w4(32'h3be58a5b),
	.w5(32'h3c049d81),
	.w6(32'h3ba96eb6),
	.w7(32'h3c26ff1d),
	.w8(32'h3b12156e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88320e),
	.w1(32'h3c180f5e),
	.w2(32'h3b932cc4),
	.w3(32'h3c571432),
	.w4(32'h3c0f5dcf),
	.w5(32'h3b8d89f3),
	.w6(32'h3c07eeb6),
	.w7(32'h3808129c),
	.w8(32'hb73831fd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b943cb1),
	.w1(32'hbb78e2c6),
	.w2(32'h3b90251d),
	.w3(32'hb796c473),
	.w4(32'h3a8da08d),
	.w5(32'h3c9285e9),
	.w6(32'h3bb7eb7a),
	.w7(32'h3981a9aa),
	.w8(32'h39ff1dc4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11e1fc),
	.w1(32'hbc01f0ee),
	.w2(32'hbb12fd10),
	.w3(32'h3cb78723),
	.w4(32'h3c14d7fb),
	.w5(32'hbbd5e003),
	.w6(32'hbab332f3),
	.w7(32'hbbf588c3),
	.w8(32'hbb8228c8),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fa923),
	.w1(32'hbae09c72),
	.w2(32'hbb69e4ba),
	.w3(32'hbbd4ddac),
	.w4(32'hbb168c0a),
	.w5(32'hbba86508),
	.w6(32'hbb451c09),
	.w7(32'hbb934ce6),
	.w8(32'hbc36bff1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf63abc),
	.w1(32'h3c4ec893),
	.w2(32'h3b658924),
	.w3(32'h3b6310db),
	.w4(32'h3bdae4e8),
	.w5(32'h3c1ae17b),
	.w6(32'hbbcbb95b),
	.w7(32'hbae58ce4),
	.w8(32'h3aa62cde),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59826),
	.w1(32'h3b076002),
	.w2(32'hbc013482),
	.w3(32'h3c7cfd0f),
	.w4(32'h3c467231),
	.w5(32'h3aa2ff70),
	.w6(32'h3c137b3c),
	.w7(32'h3b816290),
	.w8(32'hbb24f738),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf5670),
	.w1(32'hbb0c8432),
	.w2(32'h3be6fa4c),
	.w3(32'h3a6435f9),
	.w4(32'h3b07f7e0),
	.w5(32'h3b2dd886),
	.w6(32'h3a6fbd79),
	.w7(32'hbb2baa3a),
	.w8(32'hbb059b17),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfc863),
	.w1(32'hba9b3be4),
	.w2(32'hbbd6e8b2),
	.w3(32'h3af2b852),
	.w4(32'hbb95489a),
	.w5(32'hbc0b8810),
	.w6(32'hbaffb8e6),
	.w7(32'h3b05126c),
	.w8(32'hbc28ac84),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc223cd0),
	.w1(32'hbc0e824f),
	.w2(32'h3c33b4b2),
	.w3(32'hbc272096),
	.w4(32'hbc1e5740),
	.w5(32'h3c5bf9b0),
	.w6(32'hbc3174d3),
	.w7(32'hbc32b8a7),
	.w8(32'h3c9517f9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9655f7),
	.w1(32'hbd00b52f),
	.w2(32'h3c107aeb),
	.w3(32'hbc580d3f),
	.w4(32'hbd257ce4),
	.w5(32'h3bdacf36),
	.w6(32'hbb80163d),
	.w7(32'hbce33fe0),
	.w8(32'h3bec0b8a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c207342),
	.w1(32'h3ca91393),
	.w2(32'h3b34e400),
	.w3(32'h3ba160e1),
	.w4(32'h3c80ad7e),
	.w5(32'h3aa2a60d),
	.w6(32'h3a38aeb3),
	.w7(32'h3c323816),
	.w8(32'h3b640a86),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc200442),
	.w1(32'hbbe41dc7),
	.w2(32'hbb0ad32f),
	.w3(32'hbb53d330),
	.w4(32'hbb6308f9),
	.w5(32'hba940afa),
	.w6(32'h38d6395f),
	.w7(32'h3b16b5e7),
	.w8(32'hbc12b12e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a996f0a),
	.w1(32'hba3da8dd),
	.w2(32'hbc5149e7),
	.w3(32'h3c03738b),
	.w4(32'hba8abe52),
	.w5(32'hbcaf86ba),
	.w6(32'hbbd52946),
	.w7(32'hbc798bcb),
	.w8(32'hbc934b58),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0dcb7),
	.w1(32'hbc7b970d),
	.w2(32'hbbcdbedd),
	.w3(32'hbd1a588d),
	.w4(32'hbceba4e2),
	.w5(32'h39018006),
	.w6(32'hbd096747),
	.w7(32'hbcce8781),
	.w8(32'hbb7ffa25),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb935456),
	.w1(32'hbb9288df),
	.w2(32'hbbc5fbb4),
	.w3(32'h3c87263a),
	.w4(32'h3b088f96),
	.w5(32'h3bc69a68),
	.w6(32'h3bf05dd9),
	.w7(32'hbb2a1265),
	.w8(32'hbc226f30),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23f1dd),
	.w1(32'h3b7e72c4),
	.w2(32'h3b005639),
	.w3(32'h3c2f130d),
	.w4(32'h3b4d38db),
	.w5(32'hbb2f2efe),
	.w6(32'h3bae6e97),
	.w7(32'hbb895986),
	.w8(32'hbb9d9480),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b7ff4),
	.w1(32'h3b0356b7),
	.w2(32'hb99ab4f5),
	.w3(32'h3c1fbf19),
	.w4(32'h3c302d05),
	.w5(32'h3af9896d),
	.w6(32'hbb083c09),
	.w7(32'hbac10336),
	.w8(32'hbc0158f4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4402d5),
	.w1(32'hbb450eeb),
	.w2(32'h3c190fce),
	.w3(32'h3c7fa8dc),
	.w4(32'h3b213497),
	.w5(32'hbb7949c9),
	.w6(32'h3a6dbeed),
	.w7(32'h3c3f308a),
	.w8(32'h3a9ad50c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982735a),
	.w1(32'h3b89413f),
	.w2(32'h3b643deb),
	.w3(32'hbc2f36ea),
	.w4(32'hbbbb889a),
	.w5(32'hbb67cbec),
	.w6(32'hbb8320be),
	.w7(32'h3a828b0c),
	.w8(32'hbb583e4b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a511eba),
	.w1(32'hbba51a4e),
	.w2(32'hbbe374c0),
	.w3(32'h3b88450c),
	.w4(32'hbc4179f0),
	.w5(32'h3a87e7d7),
	.w6(32'h3bf3b59d),
	.w7(32'hbb99311f),
	.w8(32'hbc3bb329),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab252ba),
	.w1(32'hbc222069),
	.w2(32'h3b70dd5d),
	.w3(32'h3ca34c5f),
	.w4(32'h3bc44692),
	.w5(32'h3b3581c9),
	.w6(32'h3b45bcdc),
	.w7(32'hbbca9941),
	.w8(32'hbb63c371),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc114042),
	.w1(32'hbac74108),
	.w2(32'h3bbcae12),
	.w3(32'hbaa4fd50),
	.w4(32'h3a635f0b),
	.w5(32'h3c2b8af6),
	.w6(32'hba47be16),
	.w7(32'hbb58676e),
	.w8(32'h3c40085a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34c1d6),
	.w1(32'h3c059c51),
	.w2(32'hbbd70dda),
	.w3(32'h3c92f39a),
	.w4(32'h3c205d15),
	.w5(32'h3a1c1283),
	.w6(32'h3c6ac1dd),
	.w7(32'h3c4d1f9a),
	.w8(32'hbb684a1f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000ec3),
	.w1(32'hbc14bfdf),
	.w2(32'hbba40e0b),
	.w3(32'h3b44513c),
	.w4(32'hbb9a6d89),
	.w5(32'hbc1b7883),
	.w6(32'hbc30c061),
	.w7(32'hbc81751b),
	.w8(32'hbca9f102),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b325be6),
	.w1(32'h370765de),
	.w2(32'h3b9f7168),
	.w3(32'hb904b104),
	.w4(32'hbacc4621),
	.w5(32'hbb0b1969),
	.w6(32'hbae951eb),
	.w7(32'h3ba5f5b4),
	.w8(32'hbb7dea70),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87f919),
	.w1(32'h3c2a9b4d),
	.w2(32'h3b99a266),
	.w3(32'h3ca01912),
	.w4(32'h3c80aa8e),
	.w5(32'h3b363e61),
	.w6(32'h3c9efba3),
	.w7(32'h3c56b406),
	.w8(32'hbb4ce69d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a392e7d),
	.w1(32'h3a0ba94a),
	.w2(32'hbc016c5a),
	.w3(32'hbc09f840),
	.w4(32'hbbf24a36),
	.w5(32'hbb33c235),
	.w6(32'hbbaa93e2),
	.w7(32'hbba31be7),
	.w8(32'hbb9f1b33),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31a0b8),
	.w1(32'hb9ef7499),
	.w2(32'hbb5761ae),
	.w3(32'h3c1d9c09),
	.w4(32'h3953462a),
	.w5(32'hbbcd9355),
	.w6(32'h3a709d5e),
	.w7(32'h3b35c49c),
	.w8(32'hbc2914cb),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce9264),
	.w1(32'h3aefdb78),
	.w2(32'hbb899e4b),
	.w3(32'hbc0494c8),
	.w4(32'h3bed5732),
	.w5(32'h3beec037),
	.w6(32'hbbd0a33a),
	.w7(32'h3c76290b),
	.w8(32'hbaa91676),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85662c),
	.w1(32'h3b28a17c),
	.w2(32'hbce83535),
	.w3(32'h3c18c33b),
	.w4(32'h3c2cbcee),
	.w5(32'hbd1e2fcc),
	.w6(32'h3b8c717c),
	.w7(32'hbab6e799),
	.w8(32'hbd1082e5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0f49e),
	.w1(32'hbc06ced2),
	.w2(32'hbb9f5d92),
	.w3(32'hbd512884),
	.w4(32'hbd04d2d1),
	.w5(32'h3abe6c6c),
	.w6(32'hbd4d4887),
	.w7(32'hbccbb46f),
	.w8(32'h3b173949),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d680a),
	.w1(32'h3a3b6088),
	.w2(32'h3c5e77b9),
	.w3(32'h3b2233b8),
	.w4(32'h3ad91700),
	.w5(32'h3bb38f69),
	.w6(32'h3a1de94c),
	.w7(32'hba7b12b6),
	.w8(32'h3c363b2e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15ae40),
	.w1(32'h3c92935d),
	.w2(32'hbb49cada),
	.w3(32'h3b3101a6),
	.w4(32'h3c2e7bbc),
	.w5(32'h39588ac2),
	.w6(32'h3c03699d),
	.w7(32'h3c655eca),
	.w8(32'hbb5c724c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b749c2c),
	.w1(32'h3b48a116),
	.w2(32'h3c0b1c57),
	.w3(32'h3b897927),
	.w4(32'h3b24fbf8),
	.w5(32'h3b828000),
	.w6(32'hbb3f2dcd),
	.w7(32'hbbdc7fb4),
	.w8(32'hbac4979d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b471c3d),
	.w1(32'h3b4eab55),
	.w2(32'h3bcc819d),
	.w3(32'h399293a6),
	.w4(32'h3bee79e3),
	.w5(32'h3c497211),
	.w6(32'hbb9c8bb3),
	.w7(32'h3b013961),
	.w8(32'h3b9670cb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2813c),
	.w1(32'hbb8ed283),
	.w2(32'h3a7db0a6),
	.w3(32'h3c9e8e37),
	.w4(32'h3afb04cf),
	.w5(32'h39daad79),
	.w6(32'h3c548023),
	.w7(32'h3b33fbe7),
	.w8(32'hbc01158d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cb7a3),
	.w1(32'hbb3c8e1e),
	.w2(32'h3be97387),
	.w3(32'h3bed3987),
	.w4(32'h3b3858e0),
	.w5(32'h3c5a48de),
	.w6(32'h3b6b648f),
	.w7(32'hbbd7124d),
	.w8(32'h3a909c97),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c245f83),
	.w1(32'h3b05ee18),
	.w2(32'hba4d2448),
	.w3(32'h3c9df02b),
	.w4(32'h3c974b54),
	.w5(32'h3b88598d),
	.w6(32'h3c847939),
	.w7(32'h3c49c90b),
	.w8(32'h3b5509ea),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6939a),
	.w1(32'hbb4d3d31),
	.w2(32'hbb4ed52e),
	.w3(32'h3c1ad9f8),
	.w4(32'hbaf2854a),
	.w5(32'hba01f8d8),
	.w6(32'h3c27a1ac),
	.w7(32'hbb5673c1),
	.w8(32'hbc4a18ff),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a990169),
	.w1(32'hbb28a3dc),
	.w2(32'hbbf233a7),
	.w3(32'h3b522ae9),
	.w4(32'h3b8d9dde),
	.w5(32'hba53aad6),
	.w6(32'hbb026274),
	.w7(32'hbb5469e1),
	.w8(32'hbbe223f1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cd588),
	.w1(32'hbbf788c3),
	.w2(32'h3afd1785),
	.w3(32'hba858724),
	.w4(32'hbb94e611),
	.w5(32'hba10fa7e),
	.w6(32'hba8ee1a4),
	.w7(32'hb9d4de7b),
	.w8(32'hbbfaf7b7),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0644b4),
	.w1(32'h3a232b7f),
	.w2(32'hbb92bb50),
	.w3(32'hbb67232b),
	.w4(32'h3a93b655),
	.w5(32'h3b68d843),
	.w6(32'hbb8ba629),
	.w7(32'h3badd1cb),
	.w8(32'hbb6abe64),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb532759),
	.w1(32'hbbf516c6),
	.w2(32'h3b0520ca),
	.w3(32'hbbe8975f),
	.w4(32'hbc059e44),
	.w5(32'h3b282c28),
	.w6(32'hbc08e741),
	.w7(32'hbc099524),
	.w8(32'h3a053373),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9301e7),
	.w1(32'hbbc9b093),
	.w2(32'h3c172457),
	.w3(32'h3aeadec9),
	.w4(32'h3aca49e8),
	.w5(32'h3b97f95e),
	.w6(32'h3c17ace9),
	.w7(32'h3b296be9),
	.w8(32'hbb077408),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f6b48),
	.w1(32'h3c034162),
	.w2(32'hb981f48d),
	.w3(32'h3b9fe9ce),
	.w4(32'h3c6ec0cd),
	.w5(32'h3b635ad9),
	.w6(32'h3b5a6ec2),
	.w7(32'h3c7c1d45),
	.w8(32'hb89ca622),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4de312),
	.w1(32'hbb00b071),
	.w2(32'h3a189888),
	.w3(32'h3c1c285d),
	.w4(32'h3b9c53fe),
	.w5(32'hbbada7ef),
	.w6(32'h3c24feda),
	.w7(32'h3c10d597),
	.w8(32'hbb8677d4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd0975),
	.w1(32'h3a0241ac),
	.w2(32'hbbad7240),
	.w3(32'h3c361145),
	.w4(32'h3b036f13),
	.w5(32'h3bbb4b0c),
	.w6(32'h3ba70059),
	.w7(32'h3b9d89ab),
	.w8(32'hb8683cf2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08ed0f),
	.w1(32'h3a0e3fd4),
	.w2(32'hbaa28a25),
	.w3(32'h3c0f431a),
	.w4(32'hba86774d),
	.w5(32'h3bfe44da),
	.w6(32'h3baaedf0),
	.w7(32'h3b4798aa),
	.w8(32'h3a207895),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f544d),
	.w1(32'h3b0b7086),
	.w2(32'h3adde00f),
	.w3(32'h3c1a5b3a),
	.w4(32'h3b810c91),
	.w5(32'hb9832ac1),
	.w6(32'h3bec350f),
	.w7(32'h3ba33491),
	.w8(32'hbb906855),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4a739),
	.w1(32'hbb031105),
	.w2(32'hbbbecec4),
	.w3(32'h3bb5af21),
	.w4(32'h3b879bdc),
	.w5(32'hbba244c2),
	.w6(32'hbb6425fc),
	.w7(32'hbb63e261),
	.w8(32'hbbd3c0f9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd5edb),
	.w1(32'hbb829979),
	.w2(32'h3a640b12),
	.w3(32'h3b2ea4e0),
	.w4(32'h3a497474),
	.w5(32'h3c26b477),
	.w6(32'h3bd9b547),
	.w7(32'h3a27bd07),
	.w8(32'hbbc69f45),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe04c2),
	.w1(32'hbb22cbc8),
	.w2(32'hbb85b6e2),
	.w3(32'h3c1aeeb1),
	.w4(32'hb9cc0f63),
	.w5(32'h3b04cb59),
	.w6(32'h3acbaeca),
	.w7(32'h3b28b729),
	.w8(32'h3a2d902c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23aca8),
	.w1(32'h3b5ffd8e),
	.w2(32'hbc02f6c7),
	.w3(32'h3c36aaf4),
	.w4(32'h3c20e177),
	.w5(32'hbbf131bf),
	.w6(32'h3c798e60),
	.w7(32'h3c1c3411),
	.w8(32'hbbc41d8b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb8aaa),
	.w1(32'h3b1e510d),
	.w2(32'hbc2b652b),
	.w3(32'h3b8d5d58),
	.w4(32'h3b476d36),
	.w5(32'hbbd0c687),
	.w6(32'h3c01fcd3),
	.w7(32'h3c2a3c2b),
	.w8(32'h3b3f5ee5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41df1e),
	.w1(32'hbc4b24b5),
	.w2(32'h3cb85946),
	.w3(32'hbbdf90a9),
	.w4(32'hbbd7ac66),
	.w5(32'h3b95e276),
	.w6(32'h3aa7127d),
	.w7(32'h3b91503a),
	.w8(32'hbcf78b26),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfe70b7),
	.w1(32'h3ce29657),
	.w2(32'hbc057cd8),
	.w3(32'h3c8d217a),
	.w4(32'h3c3fa4ed),
	.w5(32'h3b89e915),
	.w6(32'hbd04a431),
	.w7(32'hbcb88fd2),
	.w8(32'h3acc877c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeddfc7),
	.w1(32'hbc3e93d3),
	.w2(32'hbac8db64),
	.w3(32'h3c0ba45e),
	.w4(32'h3b6e430a),
	.w5(32'h3a070964),
	.w6(32'h3b868095),
	.w7(32'h3bb26410),
	.w8(32'hbacf77d3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99bd16),
	.w1(32'hbb3fe531),
	.w2(32'hbc4edc84),
	.w3(32'hbb3e16ff),
	.w4(32'h3b3b3f28),
	.w5(32'hbc076fad),
	.w6(32'h3b19336c),
	.w7(32'h3bfba4d4),
	.w8(32'hbc65afc1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea82a),
	.w1(32'hbbe90524),
	.w2(32'hbb2a08ec),
	.w3(32'hbbef8de4),
	.w4(32'hbbaaa928),
	.w5(32'hbb8b122b),
	.w6(32'hba9c59e6),
	.w7(32'hbbfa125e),
	.w8(32'h3b2d087f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fc08c),
	.w1(32'h3b7776a3),
	.w2(32'hbbf2b9b6),
	.w3(32'h3b3dcf64),
	.w4(32'h3b49ecaf),
	.w5(32'hbbcb83bb),
	.w6(32'h3b217adc),
	.w7(32'h398ff7ca),
	.w8(32'hbb991b17),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11ad46),
	.w1(32'hbbf24a09),
	.w2(32'hbc7708b7),
	.w3(32'hbac4523c),
	.w4(32'hbb39b9bc),
	.w5(32'hbc1fa33f),
	.w6(32'hb8a15617),
	.w7(32'hbb17510b),
	.w8(32'hbc37da82),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda5993),
	.w1(32'hbc3d900e),
	.w2(32'h3bcdb5d0),
	.w3(32'h3ba5d913),
	.w4(32'hbb8dbcf3),
	.w5(32'h3c23db9d),
	.w6(32'hbb330f61),
	.w7(32'hbc0a0a1a),
	.w8(32'h3bb02bc5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7396e9),
	.w1(32'hbb256097),
	.w2(32'hbb570809),
	.w3(32'h3cf7a88a),
	.w4(32'h3c47e562),
	.w5(32'hbbbb68f1),
	.w6(32'h3cb28d47),
	.w7(32'h3c6e4b65),
	.w8(32'hbb023992),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d218f),
	.w1(32'h3b14ac77),
	.w2(32'h3b2b875f),
	.w3(32'h39b2e87a),
	.w4(32'h3bf90886),
	.w5(32'h3ba35915),
	.w6(32'h3bbb69e5),
	.w7(32'h3c67723e),
	.w8(32'h3b900c43),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61fbdb),
	.w1(32'h3961d0b0),
	.w2(32'hbc7dad3c),
	.w3(32'h3c731511),
	.w4(32'h3c91c012),
	.w5(32'hbbc927bb),
	.w6(32'h3c23438b),
	.w7(32'h3c961c18),
	.w8(32'hbc51663e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39188e93),
	.w1(32'hbac577ca),
	.w2(32'hbbcc5c37),
	.w3(32'h3c090d4b),
	.w4(32'h3c0be94b),
	.w5(32'hbb96ad08),
	.w6(32'h3b1d4bf4),
	.w7(32'h3c0b2e06),
	.w8(32'hbbca056f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e2df6),
	.w1(32'hbbb78112),
	.w2(32'hbc0ab253),
	.w3(32'hbb0eb199),
	.w4(32'h39858d76),
	.w5(32'h3b722047),
	.w6(32'hbbd77e90),
	.w7(32'hbbf32fb8),
	.w8(32'h3b080305),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule