module layer_10_featuremap_104(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396af20b),
	.w1(32'hb85e0963),
	.w2(32'h38916bd9),
	.w3(32'h3991ec9c),
	.w4(32'h39a64f4a),
	.w5(32'h381ece41),
	.w6(32'hb8da27fc),
	.w7(32'h38d989a1),
	.w8(32'hb8cd875a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ad6d5),
	.w1(32'hb99f1dd8),
	.w2(32'hb9f597d6),
	.w3(32'hb8fe3687),
	.w4(32'hb82805e9),
	.w5(32'h371d47dc),
	.w6(32'h38c6cc13),
	.w7(32'h37d8f77d),
	.w8(32'h395ac995),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ebd5c),
	.w1(32'hb92b0d1a),
	.w2(32'hb9a8dbca),
	.w3(32'h3912ebdb),
	.w4(32'hb8b731d3),
	.w5(32'hb89f5412),
	.w6(32'h3814554a),
	.w7(32'hb8b51fcc),
	.w8(32'h3918c7e8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934eccb),
	.w1(32'hb9e71403),
	.w2(32'hb8206d1a),
	.w3(32'hb98d765f),
	.w4(32'hb9295b55),
	.w5(32'h37947279),
	.w6(32'hb949bdae),
	.w7(32'hb9c7b31c),
	.w8(32'hb99c8b9c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d858fd),
	.w1(32'h398afd82),
	.w2(32'hb918a546),
	.w3(32'h38796edb),
	.w4(32'h3880ccbd),
	.w5(32'hb9b931f6),
	.w6(32'hb9095ccc),
	.w7(32'hb803008a),
	.w8(32'hb90094b1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fd28bf),
	.w1(32'h39b452f6),
	.w2(32'h3684925e),
	.w3(32'h367b17d9),
	.w4(32'h39b018bf),
	.w5(32'h38f73533),
	.w6(32'h39c89a27),
	.w7(32'h39a41614),
	.w8(32'h3a106a3c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efa82c),
	.w1(32'h394cc80b),
	.w2(32'h3825d0f1),
	.w3(32'h3a2427de),
	.w4(32'h38c041c9),
	.w5(32'h39895bd9),
	.w6(32'h3900b3db),
	.w7(32'hb98114ec),
	.w8(32'h392c9a81),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a149e4),
	.w1(32'h39867813),
	.w2(32'h3997a7fc),
	.w3(32'hb90941d5),
	.w4(32'hb8b8bb1f),
	.w5(32'h3903d7a2),
	.w6(32'hb937f469),
	.w7(32'hb8937a54),
	.w8(32'h3980a085),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391dda04),
	.w1(32'h396e8148),
	.w2(32'h39474d79),
	.w3(32'h399b5d44),
	.w4(32'h39fd2ef2),
	.w5(32'h39ec03a3),
	.w6(32'h39de93e3),
	.w7(32'h39b2f2b9),
	.w8(32'h39bb2681),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cff1b),
	.w1(32'hbb1b2983),
	.w2(32'hbb5000cd),
	.w3(32'hbb430175),
	.w4(32'hbb3ef6a1),
	.w5(32'hbb6b2f8d),
	.w6(32'hbb5bea68),
	.w7(32'hbb4582f6),
	.w8(32'hbb4b578b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d2e602),
	.w1(32'hb98eb724),
	.w2(32'hb99e21c3),
	.w3(32'h3930d921),
	.w4(32'h383d3aa3),
	.w5(32'h391481b4),
	.w6(32'hb888c6a1),
	.w7(32'h37a18b42),
	.w8(32'hb7839445),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1dad5),
	.w1(32'h3a33bbf6),
	.w2(32'h3aa93f9e),
	.w3(32'h3a65559d),
	.w4(32'h3a40e647),
	.w5(32'h3ac332fc),
	.w6(32'h3a0e6b92),
	.w7(32'h3a35bb18),
	.w8(32'h3ab6f702),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb1da1),
	.w1(32'hba8d0d7f),
	.w2(32'hbb0eb7b0),
	.w3(32'hbb29db5d),
	.w4(32'hbae2d8eb),
	.w5(32'hbb30aabd),
	.w6(32'hbb2ff99c),
	.w7(32'hbb0307cc),
	.w8(32'hbb10413b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba512c34),
	.w1(32'hba406c9b),
	.w2(32'hb9fd4e60),
	.w3(32'hba1c53f6),
	.w4(32'hba1b83c5),
	.w5(32'hba035f83),
	.w6(32'hba6de09b),
	.w7(32'hba4de6fd),
	.w8(32'hba6836f4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385f47f7),
	.w1(32'h3897a7dc),
	.w2(32'h3809452d),
	.w3(32'hb844f43d),
	.w4(32'h38d48674),
	.w5(32'hb5144e16),
	.w6(32'hb97d08f8),
	.w7(32'h39379127),
	.w8(32'h37113ee1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9c91a),
	.w1(32'hba876bdd),
	.w2(32'hbaebde36),
	.w3(32'hbac26d21),
	.w4(32'hba9ae29f),
	.w5(32'hbadcbdfb),
	.w6(32'hbacb79ec),
	.w7(32'hba7aae36),
	.w8(32'hbab26fad),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8e453),
	.w1(32'h39bcd16e),
	.w2(32'h39aba8da),
	.w3(32'h397405f0),
	.w4(32'h38ddff87),
	.w5(32'h38ac976a),
	.w6(32'h38f57e21),
	.w7(32'h39450f27),
	.w8(32'h39ac9107),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba152258),
	.w1(32'h39d46455),
	.w2(32'h39934ee4),
	.w3(32'hba9232d2),
	.w4(32'h38104096),
	.w5(32'hb9f6d1b7),
	.w6(32'hbaae50fe),
	.w7(32'hb9ce0dc2),
	.w8(32'hba0fa1dc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2d9b6),
	.w1(32'hb98c48f1),
	.w2(32'hba8697c9),
	.w3(32'hba4f4bfc),
	.w4(32'hba2fef06),
	.w5(32'hba9964f2),
	.w6(32'hbab9c864),
	.w7(32'hba89796d),
	.w8(32'hba9d4c27),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380f5130),
	.w1(32'h391065ee),
	.w2(32'h384bc50a),
	.w3(32'h3695f4b1),
	.w4(32'h3962c0c0),
	.w5(32'h39a477bb),
	.w6(32'h395662d8),
	.w7(32'h38817f93),
	.w8(32'h394b0743),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3347a),
	.w1(32'h389142a3),
	.w2(32'hb9613dbc),
	.w3(32'h39b00768),
	.w4(32'h39bf075e),
	.w5(32'h399e0306),
	.w6(32'h3971db80),
	.w7(32'hb79d8b46),
	.w8(32'h3967f18f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a126dc6),
	.w1(32'h3a5fb5f9),
	.w2(32'h3a32b05b),
	.w3(32'h3a4276cd),
	.w4(32'h3a08f077),
	.w5(32'h3a2c920d),
	.w6(32'h3a0ded7c),
	.w7(32'h39e2744b),
	.w8(32'h3a1504bd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e57fa7),
	.w1(32'h3a65de86),
	.w2(32'h3a23149d),
	.w3(32'hbb03fdeb),
	.w4(32'h39ee2f7e),
	.w5(32'h3a27ba48),
	.w6(32'hbaf653ff),
	.w7(32'h39e3bade),
	.w8(32'hb7e1b5f3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099da8),
	.w1(32'hba9c830c),
	.w2(32'hbb188423),
	.w3(32'hbb08c776),
	.w4(32'hba95ca90),
	.w5(32'hbb05e339),
	.w6(32'hbaea3282),
	.w7(32'hba73bf85),
	.w8(32'hbac8cd6d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bcf7a),
	.w1(32'hba24495c),
	.w2(32'hbaace552),
	.w3(32'hba0d45b2),
	.w4(32'hb6a576f9),
	.w5(32'hb9e54743),
	.w6(32'hb9037778),
	.w7(32'h39c8f02b),
	.w8(32'hb8cc1601),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f09a9f),
	.w1(32'h38fc63b5),
	.w2(32'h38b052dc),
	.w3(32'hba44834a),
	.w4(32'hb86f3789),
	.w5(32'h39b9d57e),
	.w6(32'hb9d1ce9b),
	.w7(32'h3847baf3),
	.w8(32'h395dda42),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b3061),
	.w1(32'h3913b39c),
	.w2(32'h387ac8b0),
	.w3(32'h39fb272d),
	.w4(32'h398757cb),
	.w5(32'h39b2bfad),
	.w6(32'h396fcb59),
	.w7(32'h38b8e565),
	.w8(32'h397fa24d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d996f9),
	.w1(32'hb92d3963),
	.w2(32'hb8faa457),
	.w3(32'h397844f1),
	.w4(32'h3810247e),
	.w5(32'h397081a8),
	.w6(32'h39544825),
	.w7(32'h3783a034),
	.w8(32'h39a41597),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a194838),
	.w1(32'h39e5f6a7),
	.w2(32'h39859a55),
	.w3(32'h39a7f744),
	.w4(32'h39d4baad),
	.w5(32'h3a123295),
	.w6(32'h3a5fbdfb),
	.w7(32'h3a0a13cc),
	.w8(32'h39e6891a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23fadf),
	.w1(32'hbade0465),
	.w2(32'hbb2b8949),
	.w3(32'hbb3714fd),
	.w4(32'hbb055e03),
	.w5(32'hbb158c7b),
	.w6(32'hbb4390b4),
	.w7(32'hbae2ee7b),
	.w8(32'hbb108e6e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8499071),
	.w1(32'h38ce857e),
	.w2(32'hb8b7ea6f),
	.w3(32'hb8a19a2f),
	.w4(32'h3993c78c),
	.w5(32'h3941dd9b),
	.w6(32'h39429832),
	.w7(32'h38f2788c),
	.w8(32'h3940cef7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389889db),
	.w1(32'h39c28c12),
	.w2(32'h39310ba7),
	.w3(32'h397ce9be),
	.w4(32'h3a0138b1),
	.w5(32'h39b44234),
	.w6(32'h39d6a26a),
	.w7(32'h398bf8fd),
	.w8(32'h39b2d592),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba136fac),
	.w1(32'hb8f8a836),
	.w2(32'hba07eaae),
	.w3(32'hb9f18a74),
	.w4(32'h385a5903),
	.w5(32'hb9d36513),
	.w6(32'hba2e0b1a),
	.w7(32'hb9c682a0),
	.w8(32'hba42a8ac),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba062bd8),
	.w1(32'h3a676d37),
	.w2(32'h395c9c20),
	.w3(32'hb835f374),
	.w4(32'h3a3c088d),
	.w5(32'h397a31b3),
	.w6(32'h3a680b00),
	.w7(32'h3a234281),
	.w8(32'h3a15c299),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1df47c),
	.w1(32'hb8243b7f),
	.w2(32'hb7ea176f),
	.w3(32'h39c26b05),
	.w4(32'h392ce0b1),
	.w5(32'h39704f80),
	.w6(32'h3986d598),
	.w7(32'h38514235),
	.w8(32'h39effbcf),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b7f71),
	.w1(32'h39dfb258),
	.w2(32'h38fa6c7b),
	.w3(32'h3a0f7836),
	.w4(32'h3a05d45a),
	.w5(32'h39b00bf1),
	.w6(32'h39739396),
	.w7(32'h3920d158),
	.w8(32'h39325886),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957c99d),
	.w1(32'h38af972a),
	.w2(32'hb96a8474),
	.w3(32'hb9af1d92),
	.w4(32'hb8aebb65),
	.w5(32'h38a094cd),
	.w6(32'hba4a9a71),
	.w7(32'h3825f248),
	.w8(32'h3a19bdd6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7060f7),
	.w1(32'h3912ff7e),
	.w2(32'h38a5646d),
	.w3(32'h3952ecd1),
	.w4(32'h3aa33a20),
	.w5(32'h3ab6c0a3),
	.w6(32'h3a28508a),
	.w7(32'h3abe6165),
	.w8(32'h3b156aa6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66a993),
	.w1(32'h3a8bb6f6),
	.w2(32'h3a28095a),
	.w3(32'h3abb76f0),
	.w4(32'h3ab2a404),
	.w5(32'h3aed5a2f),
	.w6(32'h3adcf503),
	.w7(32'h3ada503b),
	.w8(32'h3b207569),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e42262),
	.w1(32'hb89044fc),
	.w2(32'hb9b4aa45),
	.w3(32'h391d8d89),
	.w4(32'hb86d57ec),
	.w5(32'hb7f3aeb2),
	.w6(32'hb9804f27),
	.w7(32'hb9567321),
	.w8(32'h37180b4f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38888585),
	.w1(32'h39a18433),
	.w2(32'h39d96d19),
	.w3(32'h381224df),
	.w4(32'h3983aca8),
	.w5(32'h39a7c431),
	.w6(32'h37b39bed),
	.w7(32'h39909f9a),
	.w8(32'hb8333104),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39003b01),
	.w1(32'hb85c9fcc),
	.w2(32'h391e7089),
	.w3(32'hb7ff1b00),
	.w4(32'hb7cb14f5),
	.w5(32'hb7572177),
	.w6(32'h3913e9d7),
	.w7(32'h3755dd1f),
	.w8(32'h39300947),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a8b42),
	.w1(32'h39d2b87e),
	.w2(32'h3a50e795),
	.w3(32'h38be3e08),
	.w4(32'h3a2e01b9),
	.w5(32'h3a370a7f),
	.w6(32'h39c2b45b),
	.w7(32'h39c35e53),
	.w8(32'h3a35a215),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb375c25),
	.w1(32'hbb3a7080),
	.w2(32'hbb745c28),
	.w3(32'hbb411ce8),
	.w4(32'hbb4ccc9c),
	.w5(32'hbb691b52),
	.w6(32'hbb7711bb),
	.w7(32'hbb335ae5),
	.w8(32'hbb54d78b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5920c),
	.w1(32'hbad838f7),
	.w2(32'hbb0733b0),
	.w3(32'hbac08f5a),
	.w4(32'hbab55a9c),
	.w5(32'hbada8e13),
	.w6(32'hbaf7ab90),
	.w7(32'hba797357),
	.w8(32'hba9cae33),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20664c),
	.w1(32'hbacd0c5a),
	.w2(32'hbb1ecdb0),
	.w3(32'hbb13a70e),
	.w4(32'hbab537ab),
	.w5(32'hbaeda770),
	.w6(32'hbb09475c),
	.w7(32'hbaa1b212),
	.w8(32'hbab0e499),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9859060),
	.w1(32'hba345c5f),
	.w2(32'h39d1c3cc),
	.w3(32'h39747346),
	.w4(32'hb942c5a3),
	.w5(32'hb7ab3b64),
	.w6(32'hb97e90bf),
	.w7(32'h395aaa10),
	.w8(32'h3814017c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de1261),
	.w1(32'h38abe365),
	.w2(32'hba13106f),
	.w3(32'hbafbdc05),
	.w4(32'hb9dfaec2),
	.w5(32'hba5d16de),
	.w6(32'hbb20a20c),
	.w7(32'hba9fb53d),
	.w8(32'hbae051a5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917913d),
	.w1(32'h3a01750f),
	.w2(32'h39c98354),
	.w3(32'h39b8877f),
	.w4(32'h39fcf9d8),
	.w5(32'h39f2abed),
	.w6(32'h39f4c76c),
	.w7(32'h39b87d3c),
	.w8(32'h39b95e79),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fec533),
	.w1(32'hb8ac89b4),
	.w2(32'hb997aac8),
	.w3(32'h395711ab),
	.w4(32'hb9998406),
	.w5(32'hb9a9a8aa),
	.w6(32'hb9824f72),
	.w7(32'hb7a0e48a),
	.w8(32'h35e64f22),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a44c21),
	.w1(32'hb960d425),
	.w2(32'hb980127b),
	.w3(32'h373b64a5),
	.w4(32'hb94cf4ed),
	.w5(32'hb8f45694),
	.w6(32'hb9412227),
	.w7(32'hb8f35212),
	.w8(32'h3981f864),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53e77a),
	.w1(32'hba8ecec5),
	.w2(32'hba81e195),
	.w3(32'hba9e81a2),
	.w4(32'hba829787),
	.w5(32'hba90d382),
	.w6(32'hbaa5d598),
	.w7(32'hbaa7ee62),
	.w8(32'hbaa34b0d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b25ba3),
	.w1(32'h38b140a1),
	.w2(32'hb8fa0d62),
	.w3(32'hb9accf6a),
	.w4(32'h380ad90a),
	.w5(32'hb7381831),
	.w6(32'h38aa2cae),
	.w7(32'h38bab139),
	.w8(32'h3920a259),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa77198),
	.w1(32'hb90c93a9),
	.w2(32'hbac37905),
	.w3(32'hbad4ff85),
	.w4(32'hb9e8a5b5),
	.w5(32'hbac80f13),
	.w6(32'hbafdcf9f),
	.w7(32'hba3e4db5),
	.w8(32'hbadb7d36),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eaeee2),
	.w1(32'h3a164995),
	.w2(32'h3a308238),
	.w3(32'h3a22cab5),
	.w4(32'h39da91aa),
	.w5(32'h3a16ee36),
	.w6(32'h3a458b0e),
	.w7(32'h3a4d8ea2),
	.w8(32'h3a3a3951),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39505838),
	.w1(32'h39aeaf5e),
	.w2(32'h39a4856f),
	.w3(32'hb787e5ec),
	.w4(32'h39b9a7a7),
	.w5(32'h36a6ee6a),
	.w6(32'hb9d577a9),
	.w7(32'hb7da4992),
	.w8(32'hb91da025),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89741e8),
	.w1(32'hb99b0748),
	.w2(32'hb98d8261),
	.w3(32'hba1f8b7b),
	.w4(32'hb965dc2f),
	.w5(32'hb82b7640),
	.w6(32'hb9246943),
	.w7(32'hb930bbee),
	.w8(32'h361d92a7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3818096f),
	.w1(32'h3a2c6553),
	.w2(32'h39c4fe7c),
	.w3(32'h38bc90b0),
	.w4(32'h3a010308),
	.w5(32'hb897dd71),
	.w6(32'h39556dae),
	.w7(32'h39b79cd8),
	.w8(32'h39b3b83e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a046a),
	.w1(32'h380f9ae9),
	.w2(32'h3990031e),
	.w3(32'h3a0e39c4),
	.w4(32'hb87ce5a4),
	.w5(32'h39613cf2),
	.w6(32'h38925090),
	.w7(32'hb8ae4d08),
	.w8(32'h39311e8d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b9592a),
	.w1(32'h399e57f8),
	.w2(32'h38a1e77b),
	.w3(32'h393c73f4),
	.w4(32'h39b50ecd),
	.w5(32'h3934a69d),
	.w6(32'h39aa5fca),
	.w7(32'h3920d641),
	.w8(32'h39956922),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384122fd),
	.w1(32'hb6c4d6fd),
	.w2(32'hb99a2cc1),
	.w3(32'hb87b4a2a),
	.w4(32'hb9804ee9),
	.w5(32'hba15a0b6),
	.w6(32'hba1ca483),
	.w7(32'hb9a4ff5d),
	.w8(32'hb9ec1c92),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be0a70),
	.w1(32'h38bc5b9b),
	.w2(32'hb8f0f41a),
	.w3(32'hba1c2f32),
	.w4(32'hb8814ad0),
	.w5(32'hb9971c2f),
	.w6(32'hba287378),
	.w7(32'hb8eb3fdc),
	.w8(32'hb66608e5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913359c),
	.w1(32'h39a8ba50),
	.w2(32'h39d50b62),
	.w3(32'h362e0021),
	.w4(32'h39bee8af),
	.w5(32'h39c65a11),
	.w6(32'hb8979f74),
	.w7(32'hb908bb51),
	.w8(32'hba2887c9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc5713),
	.w1(32'hb9813964),
	.w2(32'hb925fec4),
	.w3(32'hb75eba4c),
	.w4(32'hb93c2bd2),
	.w5(32'hb891f87a),
	.w6(32'hb8821481),
	.w7(32'hb96a580b),
	.w8(32'h38c5c1ef),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989d203),
	.w1(32'h38433ce6),
	.w2(32'h3851115e),
	.w3(32'h398e7bb5),
	.w4(32'h38163f8a),
	.w5(32'hb8b57c63),
	.w6(32'h38cfb539),
	.w7(32'hb86face7),
	.w8(32'h38f648fa),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c7bda),
	.w1(32'h3a470683),
	.w2(32'h3a04f4fa),
	.w3(32'h3947a839),
	.w4(32'h3a10e459),
	.w5(32'h38b745e7),
	.w6(32'h391f052d),
	.w7(32'h3a01a335),
	.w8(32'h39d364ff),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399395e0),
	.w1(32'h39a90cfc),
	.w2(32'h3a0c3614),
	.w3(32'h39c19e71),
	.w4(32'h396ab79b),
	.w5(32'h3a01f731),
	.w6(32'hb982f821),
	.w7(32'h38defd62),
	.w8(32'hb99397c5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3335c),
	.w1(32'hb9c02f9c),
	.w2(32'hba88402f),
	.w3(32'h387d3f54),
	.w4(32'h38c98a5a),
	.w5(32'hba333d58),
	.w6(32'h3992375a),
	.w7(32'h3a30642e),
	.w8(32'hb924e590),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9581b60),
	.w1(32'h3aaa4db1),
	.w2(32'h3acc9ec4),
	.w3(32'h38706603),
	.w4(32'h3ad330d9),
	.w5(32'h3af22e0c),
	.w6(32'h3ab7ff74),
	.w7(32'h3b03e537),
	.w8(32'h3b232f94),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c97c0),
	.w1(32'hb9fdbe59),
	.w2(32'hbb07068d),
	.w3(32'hb9ae3c46),
	.w4(32'h39036662),
	.w5(32'hba190bb0),
	.w6(32'hb753c077),
	.w7(32'h3a7942a2),
	.w8(32'h3a4e0adc),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c017ee),
	.w1(32'hb8e98538),
	.w2(32'hb8946e07),
	.w3(32'h39c91555),
	.w4(32'h3824535b),
	.w5(32'h38c3ca97),
	.w6(32'h34c83abc),
	.w7(32'hb92e7e2a),
	.w8(32'h38513ee3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0e0c2),
	.w1(32'h395d9e01),
	.w2(32'h38c06052),
	.w3(32'h3955f796),
	.w4(32'h39b80163),
	.w5(32'h3907cad4),
	.w6(32'h3919ab62),
	.w7(32'h3947f373),
	.w8(32'h39563732),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38daa08c),
	.w1(32'h3931682a),
	.w2(32'h3830e26a),
	.w3(32'h3929ade9),
	.w4(32'h3994f243),
	.w5(32'h3937f0b9),
	.w6(32'h392d4606),
	.w7(32'h38b419d4),
	.w8(32'h39735cdb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39230170),
	.w1(32'h39e9c25a),
	.w2(32'h395caab5),
	.w3(32'h3991827f),
	.w4(32'h3a49ca15),
	.w5(32'h3a1e1b51),
	.w6(32'h39f0c74b),
	.w7(32'h39670c46),
	.w8(32'h3986655c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d8c0a),
	.w1(32'hb91414b5),
	.w2(32'hb834f8e5),
	.w3(32'h3a14032a),
	.w4(32'hb93daf8c),
	.w5(32'hb914be7e),
	.w6(32'h38726fe9),
	.w7(32'h36cf6f15),
	.w8(32'h39088b00),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a98af1),
	.w1(32'hb6d04547),
	.w2(32'h3ac75f78),
	.w3(32'hb9c3b738),
	.w4(32'h3931d110),
	.w5(32'h3a21d776),
	.w6(32'hba20107d),
	.w7(32'h391acd53),
	.w8(32'h3a4342d5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ccbf1),
	.w1(32'hb91bec75),
	.w2(32'hb9ba7390),
	.w3(32'hba097772),
	.w4(32'hb988ded0),
	.w5(32'h387e9ee0),
	.w6(32'hb9835495),
	.w7(32'h37370955),
	.w8(32'hb709d8f1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8eeaa),
	.w1(32'hba739c10),
	.w2(32'hbab7fafd),
	.w3(32'hba967ddd),
	.w4(32'hba5648dd),
	.w5(32'hba95674e),
	.w6(32'hbabd76dd),
	.w7(32'hba3013df),
	.w8(32'hba52da30),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba934690),
	.w1(32'hb91aaea7),
	.w2(32'hb97e5aec),
	.w3(32'hba738cff),
	.w4(32'hb56d149c),
	.w5(32'hb90d7e9a),
	.w6(32'h39960045),
	.w7(32'h3a377a1f),
	.w8(32'h39a21aa5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d7f172),
	.w1(32'hb84bb945),
	.w2(32'hb9acdb01),
	.w3(32'hb9073fd9),
	.w4(32'h39875467),
	.w5(32'hb9653e2e),
	.w6(32'h3966af6c),
	.w7(32'h38a8b428),
	.w8(32'h39265bcf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48c0fe),
	.w1(32'hb9d8ec1b),
	.w2(32'hba6fe4f9),
	.w3(32'hba36c60f),
	.w4(32'hba04436d),
	.w5(32'hba452c91),
	.w6(32'hba771b49),
	.w7(32'hba02af32),
	.w8(32'hba84a192),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28b980),
	.w1(32'h39947526),
	.w2(32'h3903207a),
	.w3(32'hba693d12),
	.w4(32'hb9c835c1),
	.w5(32'hb9b21631),
	.w6(32'hba13fa51),
	.w7(32'hb90a43a0),
	.w8(32'hb9a06d69),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9ebb3),
	.w1(32'h37bdd491),
	.w2(32'hb8c08e71),
	.w3(32'h39853558),
	.w4(32'h38f88e3c),
	.w5(32'h38bc99c3),
	.w6(32'h38f8d1ce),
	.w7(32'h38a63d72),
	.w8(32'hb78f23ae),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93890e4),
	.w1(32'hb86808c4),
	.w2(32'hb76db9bd),
	.w3(32'hb7baaa09),
	.w4(32'hb8a62507),
	.w5(32'h38443a31),
	.w6(32'h38599a67),
	.w7(32'hb7c51c4c),
	.w8(32'hb8afd0fb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e8423d),
	.w1(32'h395763f4),
	.w2(32'h38b4bec9),
	.w3(32'h36f586bb),
	.w4(32'h3982c7bd),
	.w5(32'h39a38845),
	.w6(32'h3979c35c),
	.w7(32'h3a0c746c),
	.w8(32'h39d75a05),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce87d1),
	.w1(32'hb969c5b1),
	.w2(32'hb9027042),
	.w3(32'h3982e619),
	.w4(32'hb968e0a3),
	.w5(32'hb7fe80cc),
	.w6(32'hb98f7618),
	.w7(32'hb986fe38),
	.w8(32'hb98fe5f0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa16ce),
	.w1(32'h3a92253d),
	.w2(32'h3a618760),
	.w3(32'h397d4dbe),
	.w4(32'h3ac5bd51),
	.w5(32'h3ac4d4ec),
	.w6(32'h3a129898),
	.w7(32'h3ace840e),
	.w8(32'h3b1243b3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9b545),
	.w1(32'h39584b72),
	.w2(32'h39919907),
	.w3(32'h3984bdee),
	.w4(32'h39fbf491),
	.w5(32'h3a2b770a),
	.w6(32'h39a07b57),
	.w7(32'h397a1ba1),
	.w8(32'h3a0b6b54),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba335a4e),
	.w1(32'hb9f86c0a),
	.w2(32'hba8fd334),
	.w3(32'hba45ba2e),
	.w4(32'hba6782dd),
	.w5(32'hba89c6ad),
	.w6(32'hb9c60a4b),
	.w7(32'hb9adee49),
	.w8(32'hba15e223),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c365b),
	.w1(32'hba492680),
	.w2(32'hb88adf4c),
	.w3(32'hba959a48),
	.w4(32'hb8455bd2),
	.w5(32'hb8298f22),
	.w6(32'hba176460),
	.w7(32'hb9c40d58),
	.w8(32'h394368f7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e6712),
	.w1(32'h3a622976),
	.w2(32'h3a122714),
	.w3(32'h3a79965d),
	.w4(32'h3aa990e1),
	.w5(32'h3aa57baf),
	.w6(32'h3a7cd53d),
	.w7(32'h3abeaadc),
	.w8(32'h3ad7d91e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1618b),
	.w1(32'hb9f38528),
	.w2(32'h38ada2b6),
	.w3(32'hb9603d23),
	.w4(32'hb9bfa2a8),
	.w5(32'hb9bbb1cc),
	.w6(32'hba12845b),
	.w7(32'hb9860307),
	.w8(32'h39816fc9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01b6c0),
	.w1(32'hb95eec1b),
	.w2(32'h39980ca7),
	.w3(32'hb99960a1),
	.w4(32'hb998e1db),
	.w5(32'h37eec4bd),
	.w6(32'hb7dd7542),
	.w7(32'h39cdf4cd),
	.w8(32'h3a62c454),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba45a4),
	.w1(32'hba8100e5),
	.w2(32'hbaa8b353),
	.w3(32'hba87907c),
	.w4(32'hb7d7c699),
	.w5(32'h3824fd40),
	.w6(32'hb895228d),
	.w7(32'h3a2279a0),
	.w8(32'h39e55c0c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba710e7c),
	.w1(32'hb9ef4074),
	.w2(32'hba4c8e2b),
	.w3(32'hba5e86de),
	.w4(32'hba069237),
	.w5(32'hba1952dd),
	.w6(32'hba30cd1b),
	.w7(32'hb85df199),
	.w8(32'hb8fa774c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba572b98),
	.w1(32'h39149081),
	.w2(32'hba1bc80d),
	.w3(32'hb99a4893),
	.w4(32'h39908450),
	.w5(32'hb971277e),
	.w6(32'hb8b9ff4a),
	.w7(32'h3a25c041),
	.w8(32'h3994b2b2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b66e05),
	.w1(32'h398c227e),
	.w2(32'h39cc82ef),
	.w3(32'h39ff7b5f),
	.w4(32'h3953d3ef),
	.w5(32'h3981e66f),
	.w6(32'h39de46db),
	.w7(32'h39f2aa71),
	.w8(32'hb7f80210),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafea5c1),
	.w1(32'hb9b9f473),
	.w2(32'hba9e531f),
	.w3(32'hbb144a68),
	.w4(32'hba415281),
	.w5(32'hbae62d76),
	.w6(32'hbad3f105),
	.w7(32'hba73936e),
	.w8(32'hbaf02cb4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79687f),
	.w1(32'h3912639a),
	.w2(32'h3a2689bb),
	.w3(32'hb8172624),
	.w4(32'h3918e411),
	.w5(32'h3a3256e9),
	.w6(32'h39c1eea4),
	.w7(32'h39814cb9),
	.w8(32'h3a7e41d0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b9e05),
	.w1(32'h3a4e9e17),
	.w2(32'h3a7093da),
	.w3(32'h3a1932a9),
	.w4(32'h3a80ad7f),
	.w5(32'h3a8d15df),
	.w6(32'h39bc967c),
	.w7(32'h3a434a82),
	.w8(32'h3a340864),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906732f),
	.w1(32'h3adbbcf6),
	.w2(32'h3b694e8f),
	.w3(32'h3a8780eb),
	.w4(32'h3b445a6f),
	.w5(32'h3b88c2a8),
	.w6(32'h3b359462),
	.w7(32'h3b6c2dc8),
	.w8(32'h3ba87eab),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb239ec6),
	.w1(32'hbae7dc1f),
	.w2(32'hbb511cc7),
	.w3(32'hbb45e662),
	.w4(32'hbb3d970a),
	.w5(32'hbb6861bb),
	.w6(32'hbb6269ed),
	.w7(32'hbadea10e),
	.w8(32'hbb383a96),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39398cb3),
	.w1(32'h3a8a2769),
	.w2(32'h3a112dbe),
	.w3(32'hb81a527a),
	.w4(32'h3a744543),
	.w5(32'h3a1644bf),
	.w6(32'hb9992cd3),
	.w7(32'h3a373b7a),
	.w8(32'h3a718744),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a425343),
	.w1(32'h3a5b3648),
	.w2(32'h3a53e7e0),
	.w3(32'h3a3c96af),
	.w4(32'h3a4dbb2b),
	.w5(32'h3a54871c),
	.w6(32'h39fa4692),
	.w7(32'h3a312cd1),
	.w8(32'h3a634138),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983d169),
	.w1(32'h39951cad),
	.w2(32'h3ab1f38a),
	.w3(32'hb9f60f98),
	.w4(32'h3a510bb2),
	.w5(32'h3b17a4e7),
	.w6(32'hba0ad2a6),
	.w7(32'h3a8eb5bc),
	.w8(32'h3b1caccd),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9429f0e),
	.w1(32'h39a59b69),
	.w2(32'h3a034d79),
	.w3(32'hb93201ba),
	.w4(32'h3a04c00a),
	.w5(32'h3a81324c),
	.w6(32'hb8ba57af),
	.w7(32'h39f0a57f),
	.w8(32'h3a403fcf),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a87b9b),
	.w1(32'hb7aadcc7),
	.w2(32'hb8cb2305),
	.w3(32'h39c03c56),
	.w4(32'hb766703f),
	.w5(32'h389b3131),
	.w6(32'h3908faa7),
	.w7(32'h38b44e18),
	.w8(32'h3922cc0d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4fbe8),
	.w1(32'hb8cff1bb),
	.w2(32'hb9df8341),
	.w3(32'hb90f248d),
	.w4(32'h3966c38c),
	.w5(32'h392e392d),
	.w6(32'h38a0d749),
	.w7(32'h384858c2),
	.w8(32'h38f0cbd3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00f5b8),
	.w1(32'hbad2894a),
	.w2(32'hbb281beb),
	.w3(32'hbb16859e),
	.w4(32'hbb04871d),
	.w5(32'hbb19b296),
	.w6(32'hbb454fa9),
	.w7(32'hbaedf0e9),
	.w8(32'hbb00ae13),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2b2d0),
	.w1(32'hbade6fad),
	.w2(32'hbb18a559),
	.w3(32'hbafc6efe),
	.w4(32'hbac696b2),
	.w5(32'hbb1b8950),
	.w6(32'hbb2a4d0a),
	.w7(32'hbac7d0ee),
	.w8(32'hbb06c0b1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c250bd),
	.w1(32'h3a206812),
	.w2(32'h3a84cae4),
	.w3(32'hb957321f),
	.w4(32'h3a699b94),
	.w5(32'h3ac210e5),
	.w6(32'h3a3ca4d9),
	.w7(32'h3a6d96ba),
	.w8(32'h3ad4fa83),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be4bb8),
	.w1(32'hb80c5fd3),
	.w2(32'h3947d88f),
	.w3(32'h3a0cdf33),
	.w4(32'h39be66f6),
	.w5(32'h38e9b4aa),
	.w6(32'h3800a4ac),
	.w7(32'h395300ec),
	.w8(32'h38a4f91f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb722bc7b),
	.w1(32'h3a3d0b13),
	.w2(32'h3a277877),
	.w3(32'h38b41d0f),
	.w4(32'h3a65b364),
	.w5(32'h3a6e0017),
	.w6(32'h3a441a9d),
	.w7(32'h3a5a8d51),
	.w8(32'h3a8d34b4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4767d7),
	.w1(32'hba18f430),
	.w2(32'hba894f59),
	.w3(32'hb9f9b4c9),
	.w4(32'hba8b1e90),
	.w5(32'hbaaccd2c),
	.w6(32'hba567d57),
	.w7(32'hba3e49e2),
	.w8(32'hb9be5463),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac67137),
	.w1(32'hba569b06),
	.w2(32'hbab44a20),
	.w3(32'hbadd973a),
	.w4(32'hba68db10),
	.w5(32'hba892a83),
	.w6(32'hbad11f06),
	.w7(32'hba962a15),
	.w8(32'hba620b39),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b3dbf),
	.w1(32'h3959c231),
	.w2(32'h38b5d293),
	.w3(32'h39bf80a2),
	.w4(32'h390e734e),
	.w5(32'h38e1d39a),
	.w6(32'h382066f4),
	.w7(32'h393dd6f5),
	.w8(32'h39d8d948),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397fda16),
	.w1(32'h38e6460b),
	.w2(32'h360c51f5),
	.w3(32'h39bc0b6c),
	.w4(32'h38e180aa),
	.w5(32'hb82bcec9),
	.w6(32'h3805831c),
	.w7(32'h39110b1e),
	.w8(32'h3994326c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38984275),
	.w1(32'h3934235a),
	.w2(32'h37d94b9d),
	.w3(32'h38c8a46d),
	.w4(32'h39462716),
	.w5(32'h33ff0291),
	.w6(32'h38b7852f),
	.w7(32'h393fca8f),
	.w8(32'h39b455de),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6e7c1),
	.w1(32'h384338c9),
	.w2(32'h38b47182),
	.w3(32'h390a4b4d),
	.w4(32'hb91b96b5),
	.w5(32'hb867c236),
	.w6(32'hb86eeeb3),
	.w7(32'h391ae239),
	.w8(32'h39b0fcce),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d74d3),
	.w1(32'hba873c18),
	.w2(32'hbaee8e88),
	.w3(32'hba2c4e8c),
	.w4(32'hba972a14),
	.w5(32'hbacc41e5),
	.w6(32'hba9783a0),
	.w7(32'hba996e5f),
	.w8(32'hba88a4f2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3872749e),
	.w1(32'h382723c8),
	.w2(32'hb78abe70),
	.w3(32'h3927a712),
	.w4(32'h39d4fa36),
	.w5(32'h39f03abb),
	.w6(32'h39d5cf11),
	.w7(32'h39371695),
	.w8(32'h39d6f36e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bcdcd0),
	.w1(32'h3a3618a9),
	.w2(32'h39dddcb4),
	.w3(32'h39295bdf),
	.w4(32'h3a00cbe7),
	.w5(32'h39f3525b),
	.w6(32'hb87fbb1e),
	.w7(32'h39b2ded8),
	.w8(32'h39dc60af),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3a698),
	.w1(32'h38c1985f),
	.w2(32'hb9e43d41),
	.w3(32'h38457da2),
	.w4(32'h39fb14e8),
	.w5(32'h399aa476),
	.w6(32'h3940cbc4),
	.w7(32'h39a01eb3),
	.w8(32'h3a157bbe),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5b333),
	.w1(32'hb80a6e8b),
	.w2(32'h396f21e6),
	.w3(32'h390b9a74),
	.w4(32'hb890fd47),
	.w5(32'h38b64520),
	.w6(32'h383cedc9),
	.w7(32'h3865df22),
	.w8(32'h389a86da),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54be9f),
	.w1(32'h39259e74),
	.w2(32'hb8ba67b7),
	.w3(32'h3a2bb982),
	.w4(32'hb7db2737),
	.w5(32'hb83adf5b),
	.w6(32'h394fd780),
	.w7(32'h394aa1bb),
	.w8(32'h394c4330),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e67c61),
	.w1(32'h38e0b8f4),
	.w2(32'hb83802d2),
	.w3(32'h38af7f99),
	.w4(32'h39e87dfc),
	.w5(32'h39e424c8),
	.w6(32'h39923801),
	.w7(32'h39443a45),
	.w8(32'h39bde976),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3953b8bc),
	.w1(32'hb6117b76),
	.w2(32'h38321eea),
	.w3(32'h39ef54b5),
	.w4(32'h38c0442f),
	.w5(32'h391eba97),
	.w6(32'hb7d955f5),
	.w7(32'h38ee3147),
	.w8(32'h38d55e92),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ded33),
	.w1(32'hba14f681),
	.w2(32'hba91a9e3),
	.w3(32'hba94f411),
	.w4(32'hba4bbc5a),
	.w5(32'hba8a85c0),
	.w6(32'hba878c68),
	.w7(32'hba5c2394),
	.w8(32'hbaa3077d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bac86),
	.w1(32'hba773296),
	.w2(32'hbafbea96),
	.w3(32'hbaab2cce),
	.w4(32'hba6cb03e),
	.w5(32'hbb0496fc),
	.w6(32'hbac5b7fe),
	.w7(32'hba57e174),
	.w8(32'hbaab0902),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376c2660),
	.w1(32'h36b15b00),
	.w2(32'h38ab3713),
	.w3(32'hb8945b61),
	.w4(32'h384aa12c),
	.w5(32'h38b410ab),
	.w6(32'hb83e2a08),
	.w7(32'h36c2f1da),
	.w8(32'h38676539),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94bcef8),
	.w1(32'h3751628c),
	.w2(32'hb8194d44),
	.w3(32'hb925f4dd),
	.w4(32'hb84c1076),
	.w5(32'hb8f02c75),
	.w6(32'h387e1d66),
	.w7(32'h38d8d07a),
	.w8(32'hb4a4ccca),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ed3ef),
	.w1(32'hb7d1bbac),
	.w2(32'hb8f014e1),
	.w3(32'hb88f0197),
	.w4(32'h379be521),
	.w5(32'hb8d470e0),
	.w6(32'h38945b50),
	.w7(32'h38da3d3d),
	.w8(32'h366e69bb),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803926),
	.w1(32'hba5d610b),
	.w2(32'hba480662),
	.w3(32'hba93d3d6),
	.w4(32'hba5dcda5),
	.w5(32'hba4399d1),
	.w6(32'hba960497),
	.w7(32'hba2d26d1),
	.w8(32'hba55f026),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8995744),
	.w1(32'hb97b26fd),
	.w2(32'hb8191e9c),
	.w3(32'hb9223bd0),
	.w4(32'hb923ebf1),
	.w5(32'h39715def),
	.w6(32'h3a2b90bd),
	.w7(32'h39ca0d71),
	.w8(32'h396a51d2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba791e07),
	.w1(32'h3997b155),
	.w2(32'h39c505f6),
	.w3(32'hba3d600f),
	.w4(32'h39ab7890),
	.w5(32'hb936988c),
	.w6(32'hba6295f2),
	.w7(32'hb8a52d9c),
	.w8(32'hb9c1ab3c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8532b9),
	.w1(32'hba34302b),
	.w2(32'hba7d4f74),
	.w3(32'hba6d2a91),
	.w4(32'hba18b56c),
	.w5(32'hba28cc3f),
	.w6(32'hba5cf709),
	.w7(32'hb916d233),
	.w8(32'hb9c63161),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba720242),
	.w1(32'hb98ff3ce),
	.w2(32'hb91f9eb4),
	.w3(32'hba0b458f),
	.w4(32'hb96624c7),
	.w5(32'hba224e71),
	.w6(32'hb9243132),
	.w7(32'h395acaa2),
	.w8(32'h39bb8641),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f08b6),
	.w1(32'h390bd919),
	.w2(32'hb9b3bfcb),
	.w3(32'hba71520b),
	.w4(32'hb81696af),
	.w5(32'hb8c11f66),
	.w6(32'hba7302b8),
	.w7(32'hb9cb9722),
	.w8(32'h3834c1c6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0168f8),
	.w1(32'hb98f8607),
	.w2(32'hba07dba1),
	.w3(32'hba1e1ec3),
	.w4(32'hb80ed5cf),
	.w5(32'hb9057f80),
	.w6(32'hb9303979),
	.w7(32'h3995f891),
	.w8(32'h378395af),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ca472),
	.w1(32'hba58a8e7),
	.w2(32'hba8b8fc1),
	.w3(32'hbaa54ebe),
	.w4(32'hba6b9095),
	.w5(32'hba9a63a8),
	.w6(32'hbaaa8d34),
	.w7(32'hba83c377),
	.w8(32'hba90e36f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba242402),
	.w1(32'hb9d10a82),
	.w2(32'hba008e74),
	.w3(32'hba11ba6e),
	.w4(32'hb9d1b6ce),
	.w5(32'hb9f9de23),
	.w6(32'hba205e78),
	.w7(32'hb99f0780),
	.w8(32'hb9e7f474),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa664e6),
	.w1(32'hba27630a),
	.w2(32'hbaa61aa4),
	.w3(32'hba4fd9b1),
	.w4(32'hb9da95ba),
	.w5(32'hba2a0a78),
	.w6(32'hb9a9e3e0),
	.w7(32'hb907f404),
	.w8(32'hb9ed7a82),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386184af),
	.w1(32'h3a62673d),
	.w2(32'h3a2c24be),
	.w3(32'hb6c1ed76),
	.w4(32'h3a810f48),
	.w5(32'h3a9a927d),
	.w6(32'h3a1bd190),
	.w7(32'h3acabfb4),
	.w8(32'h3acb9144),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af759a),
	.w1(32'h351e2685),
	.w2(32'h36053401),
	.w3(32'h3888a822),
	.w4(32'h362d5c62),
	.w5(32'h36b7e244),
	.w6(32'hb3df308c),
	.w7(32'h36a6e3ee),
	.w8(32'h3734a5d6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61cb054),
	.w1(32'hb7cbcc96),
	.w2(32'h3768a8b5),
	.w3(32'h360c78f4),
	.w4(32'hb7f427db),
	.w5(32'h36db80f2),
	.w6(32'hb7d7421b),
	.w7(32'h3773467c),
	.w8(32'h384a6173),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80b1cea),
	.w1(32'hb9508f54),
	.w2(32'hb93a43ef),
	.w3(32'hb913a5c4),
	.w4(32'hb8805296),
	.w5(32'hb77804ff),
	.w6(32'hb9777bf9),
	.w7(32'h369f70a7),
	.w8(32'hb80b2295),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff4846),
	.w1(32'h3a68fdf0),
	.w2(32'h3a059e46),
	.w3(32'h38262b3d),
	.w4(32'h3a9be3ba),
	.w5(32'h3a9ecbea),
	.w6(32'h39f91f9f),
	.w7(32'h3ac4056d),
	.w8(32'h3af871da),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6e4c4),
	.w1(32'hbad9a586),
	.w2(32'hbb2b91f2),
	.w3(32'hbaf071a8),
	.w4(32'hbabf0471),
	.w5(32'hbb15dd2a),
	.w6(32'hbaf7f0e5),
	.w7(32'hbaab161f),
	.w8(32'hbb097f5d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370dedc8),
	.w1(32'hb7a07af1),
	.w2(32'h380146d6),
	.w3(32'h371102ca),
	.w4(32'hb6d4461a),
	.w5(32'h38483093),
	.w6(32'hb793271e),
	.w7(32'h3809f1a1),
	.w8(32'hb60a54dc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8a6dc),
	.w1(32'hba5e926d),
	.w2(32'hbad2e9d2),
	.w3(32'hbab3ba21),
	.w4(32'hba7cf3cf),
	.w5(32'hbada1a1d),
	.w6(32'hbac9bcb4),
	.w7(32'hba718eba),
	.w8(32'hbabbb11d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba983ba0),
	.w1(32'hba915ff4),
	.w2(32'hbac63971),
	.w3(32'hbacfa811),
	.w4(32'hbab9ee47),
	.w5(32'hbabfa1b2),
	.w6(32'hbaf875c9),
	.w7(32'hba8e77f1),
	.w8(32'hbaa1d230),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5efad4),
	.w1(32'h3a3bf116),
	.w2(32'h3a57c3ce),
	.w3(32'hba8cd33e),
	.w4(32'hb88924cb),
	.w5(32'hb8edbb15),
	.w6(32'hbab32d82),
	.w7(32'hb9868e7d),
	.w8(32'hb94eeac1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9aa7c),
	.w1(32'h39ba84f2),
	.w2(32'hba00cd84),
	.w3(32'hb89b97a0),
	.w4(32'h39722405),
	.w5(32'hb9ab2c53),
	.w6(32'h3868fd51),
	.w7(32'h39d9518a),
	.w8(32'hb91c59b4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f18cbc),
	.w1(32'h3a6dcbb4),
	.w2(32'h3a46b897),
	.w3(32'h3a254ce8),
	.w4(32'h3a68b6b1),
	.w5(32'h3a856ff8),
	.w6(32'h3a839cb6),
	.w7(32'h3a6b4384),
	.w8(32'h3a8ac9f8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39945c1b),
	.w1(32'h39c6cf2c),
	.w2(32'h39af4a55),
	.w3(32'h39a344d5),
	.w4(32'h394d603a),
	.w5(32'h39e14b2f),
	.w6(32'h39dd7e7b),
	.w7(32'h39cecec1),
	.w8(32'h3a0ecbaf),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98a81e),
	.w1(32'hba7de9a2),
	.w2(32'hbaa4845c),
	.w3(32'hbaba9faf),
	.w4(32'hba714630),
	.w5(32'hba8d63e9),
	.w6(32'hbab032ef),
	.w7(32'hba4d389d),
	.w8(32'hba957c38),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a138578),
	.w1(32'h3a753e4f),
	.w2(32'h3a966682),
	.w3(32'h3aa7a9ef),
	.w4(32'h3abe57ed),
	.w5(32'h3adcbe95),
	.w6(32'h3ade0f70),
	.w7(32'h3adef2e3),
	.w8(32'h3adb1dfc),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395ed765),
	.w1(32'h3953fc08),
	.w2(32'h39b1d013),
	.w3(32'h39b97976),
	.w4(32'h39b8e3d8),
	.w5(32'h3a083b16),
	.w6(32'h390e83e9),
	.w7(32'h39f231c7),
	.w8(32'h3a37443b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dc1855),
	.w1(32'h389ec647),
	.w2(32'h3934f859),
	.w3(32'h37181748),
	.w4(32'h39125646),
	.w5(32'h393ae029),
	.w6(32'hb7ff90df),
	.w7(32'h38d28978),
	.w8(32'h38026985),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37433e8e),
	.w1(32'h37db304a),
	.w2(32'h372fc117),
	.w3(32'h3826653b),
	.w4(32'h36a888e6),
	.w5(32'hb645d4ed),
	.w6(32'hb843272e),
	.w7(32'hb79e1a32),
	.w8(32'hb77852f3),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8edf301),
	.w1(32'h39772950),
	.w2(32'hb9d73371),
	.w3(32'hb8c5c727),
	.w4(32'h3947ed6e),
	.w5(32'hba00ba6e),
	.w6(32'hb91f9600),
	.w7(32'hb7e7c8dc),
	.w8(32'hb9a6ffff),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3782d672),
	.w1(32'hb88eb299),
	.w2(32'hb8a6de45),
	.w3(32'h36f7788d),
	.w4(32'hb8a9c9c1),
	.w5(32'hb8a0ca54),
	.w6(32'hb8881228),
	.w7(32'hb870c436),
	.w8(32'h38817b2e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba601f79),
	.w1(32'hba1a73aa),
	.w2(32'hba494d8e),
	.w3(32'hba7189ee),
	.w4(32'hba348259),
	.w5(32'hba89d527),
	.w6(32'hba7210d0),
	.w7(32'hba351f23),
	.w8(32'hba3b6f99),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3870aac3),
	.w1(32'hb8c8dafc),
	.w2(32'hb8479111),
	.w3(32'h3889c5fa),
	.w4(32'hb87617f0),
	.w5(32'hb81097ea),
	.w6(32'hb81a1f16),
	.w7(32'hb83170a2),
	.w8(32'hb8291e4d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f52a9),
	.w1(32'h39a697a7),
	.w2(32'h393ee65a),
	.w3(32'h3a6198f8),
	.w4(32'h399da2ec),
	.w5(32'h392eee41),
	.w6(32'h3a470aef),
	.w7(32'h39e55d99),
	.w8(32'h39696ae6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384cc7c4),
	.w1(32'h38bc7730),
	.w2(32'h39010a30),
	.w3(32'h38a16987),
	.w4(32'h38d32958),
	.w5(32'h38d2d6f6),
	.w6(32'h384599ba),
	.w7(32'h38be53ab),
	.w8(32'h388c25b7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38137d6c),
	.w1(32'hb7e8746e),
	.w2(32'hb86298c2),
	.w3(32'hb865eb10),
	.w4(32'hb87a3c89),
	.w5(32'hb804a786),
	.w6(32'h386e0315),
	.w7(32'hb7b13840),
	.w8(32'h372c0fc1),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fa893),
	.w1(32'h3931caca),
	.w2(32'h39613d00),
	.w3(32'hba2c09b9),
	.w4(32'h39d8407a),
	.w5(32'h3a20061a),
	.w6(32'hb959e9d0),
	.w7(32'h3a62dd1e),
	.w8(32'h3a7f3c02),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1aa6e),
	.w1(32'hba4aae5d),
	.w2(32'hbaa939f5),
	.w3(32'hbae2fad0),
	.w4(32'hbaaaba9d),
	.w5(32'hbadf5690),
	.w6(32'hbac1a224),
	.w7(32'hb9b140c0),
	.w8(32'hba928c68),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39befa97),
	.w1(32'h38cd5a96),
	.w2(32'h3905c847),
	.w3(32'h398ec098),
	.w4(32'h386c9db8),
	.w5(32'h392d604a),
	.w6(32'h3966796e),
	.w7(32'h391fc3f9),
	.w8(32'h39c78510),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb154cc2),
	.w1(32'hbabd817b),
	.w2(32'hbb0de6b6),
	.w3(32'hbb215e87),
	.w4(32'hbafb5706),
	.w5(32'hbafe9ea8),
	.w6(32'hbb202fca),
	.w7(32'hbacbdce3),
	.w8(32'hbaebc4cd),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d039af),
	.w1(32'hb9c7a0df),
	.w2(32'hb9f5d3ad),
	.w3(32'hba090001),
	.w4(32'hba00c040),
	.w5(32'hb9ecb6f6),
	.w6(32'hba106a41),
	.w7(32'hb9b74fcb),
	.w8(32'hb9a0101c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7bca8),
	.w1(32'hba2566cb),
	.w2(32'hba96942d),
	.w3(32'hba34e3b7),
	.w4(32'hb9e0db1f),
	.w5(32'hba84dbae),
	.w6(32'hba47a905),
	.w7(32'hb92701e6),
	.w8(32'hba0e9045),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac3502),
	.w1(32'h385e53d9),
	.w2(32'h390b1448),
	.w3(32'hb8f75bd1),
	.w4(32'h39b16cf1),
	.w5(32'h39c467c9),
	.w6(32'h39819e25),
	.w7(32'h3a2a8f55),
	.w8(32'h3a0ce73c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2f615),
	.w1(32'hb9a3081d),
	.w2(32'hba8f0f33),
	.w3(32'hbae62c3b),
	.w4(32'hba6bf94d),
	.w5(32'hbac3df75),
	.w6(32'hbafbe8a2),
	.w7(32'hba17cf97),
	.w8(32'hbaac11f7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dd1f1d),
	.w1(32'h3818dd8c),
	.w2(32'h38269198),
	.w3(32'h39397d22),
	.w4(32'h3838fdd2),
	.w5(32'h38b819cf),
	.w6(32'hb8a02a7c),
	.w7(32'h3887980f),
	.w8(32'h394e3509),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909aba2),
	.w1(32'h39355cc3),
	.w2(32'hba0d07e1),
	.w3(32'hb94d595e),
	.w4(32'hb7cc4161),
	.w5(32'hba11f902),
	.w6(32'hb94e8c43),
	.w7(32'h3950e476),
	.w8(32'hb91e2e92),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76fa543),
	.w1(32'hb85271de),
	.w2(32'hb7aefb0e),
	.w3(32'hb7429f8d),
	.w4(32'hb840f9e2),
	.w5(32'hb799b65f),
	.w6(32'hb829017f),
	.w7(32'hb80207e7),
	.w8(32'hb824e0c6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de936c),
	.w1(32'h37f6743b),
	.w2(32'h377ee1cb),
	.w3(32'h38a1fca1),
	.w4(32'h387b60c3),
	.w5(32'hb7743d06),
	.w6(32'h38a830aa),
	.w7(32'h38d806b4),
	.w8(32'hb3a34b19),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc50eb),
	.w1(32'h3920c588),
	.w2(32'hb98908cf),
	.w3(32'h3885e368),
	.w4(32'h38b0f81a),
	.w5(32'hb9441e81),
	.w6(32'h38df8c54),
	.w7(32'hb949b78c),
	.w8(32'hb8563823),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe64a2),
	.w1(32'hb9c87bab),
	.w2(32'hba213334),
	.w3(32'hb912d83f),
	.w4(32'hb98a9ade),
	.w5(32'hb9ca4191),
	.w6(32'hb953fe45),
	.w7(32'hb89ded2f),
	.w8(32'hb986d3df),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7125d34),
	.w1(32'hb85a0ca5),
	.w2(32'h38826327),
	.w3(32'hb71d0c72),
	.w4(32'hb7f5dbdc),
	.w5(32'h3895233c),
	.w6(32'hb864c0ca),
	.w7(32'h3862ec89),
	.w8(32'hb7fd666e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8623c6d),
	.w1(32'hb86227dc),
	.w2(32'hb87d7f0b),
	.w3(32'hb6fdcfe5),
	.w4(32'hb87d7200),
	.w5(32'hb895bb20),
	.w6(32'hb6be3706),
	.w7(32'hb79b3fcb),
	.w8(32'h34d63b3c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954ecbc),
	.w1(32'hb9694781),
	.w2(32'hb8dfd24f),
	.w3(32'hb9236a4a),
	.w4(32'hb91c50a2),
	.w5(32'hb8d17f4b),
	.w6(32'hb8dc25a2),
	.w7(32'h394e258b),
	.w8(32'hb88fe7cd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990c0ec),
	.w1(32'h393dcc88),
	.w2(32'h39f48732),
	.w3(32'hb88428db),
	.w4(32'h39f29352),
	.w5(32'h39dc6739),
	.w6(32'hb92a51c1),
	.w7(32'h39b6ffd9),
	.w8(32'h3a40c0ad),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370798ce),
	.w1(32'hb8bbf4cf),
	.w2(32'h39985edb),
	.w3(32'hb8bdc53d),
	.w4(32'hb7f2ee1b),
	.w5(32'h39852443),
	.w6(32'hb94f0e8c),
	.w7(32'h38e2749f),
	.w8(32'h38f84cbf),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93aa92e),
	.w1(32'hb8ad7d54),
	.w2(32'hb8fa01cf),
	.w3(32'hb8f003b0),
	.w4(32'hb919cf37),
	.w5(32'hb86a8b0a),
	.w6(32'hb8c4863c),
	.w7(32'hb8db82bd),
	.w8(32'h3887e80b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6061b),
	.w1(32'hba764c25),
	.w2(32'hbb5b0822),
	.w3(32'hbb2011ff),
	.w4(32'hbb197f64),
	.w5(32'hbb8dd594),
	.w6(32'hbb621270),
	.w7(32'hbb0e91cf),
	.w8(32'hbb852f6b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb087eec),
	.w1(32'hba9f3827),
	.w2(32'hba83aa0d),
	.w3(32'hbac34d32),
	.w4(32'hba05768c),
	.w5(32'h397521ac),
	.w6(32'hba8657df),
	.w7(32'h390fde90),
	.w8(32'h39c43782),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7db247f),
	.w1(32'h38221acb),
	.w2(32'h38cf1471),
	.w3(32'hb7932d09),
	.w4(32'h3709bec7),
	.w5(32'h38623993),
	.w6(32'hb71d5059),
	.w7(32'h37bf10d8),
	.w8(32'h38e0289d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379aa6b0),
	.w1(32'h38aa961a),
	.w2(32'hb91b335d),
	.w3(32'hb555216c),
	.w4(32'h382411db),
	.w5(32'hb925cbde),
	.w6(32'h389ca9f8),
	.w7(32'hb9033634),
	.w8(32'h38a33b75),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75d72a6),
	.w1(32'hb9331ba8),
	.w2(32'hb92b5dd7),
	.w3(32'hb83a11c5),
	.w4(32'hb978c3b1),
	.w5(32'hb966dff0),
	.w6(32'hb90e43d6),
	.w7(32'hb920fa57),
	.w8(32'hb8dc32cb),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b0a931),
	.w1(32'hb7319f19),
	.w2(32'hb740358b),
	.w3(32'h36cd152c),
	.w4(32'hb7958ea2),
	.w5(32'hb774b944),
	.w6(32'hb745e30f),
	.w7(32'hb7225d72),
	.w8(32'hb705c84e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b9575),
	.w1(32'hb79cf9ad),
	.w2(32'hb8fb6cbf),
	.w3(32'hba031598),
	.w4(32'hb9a04e62),
	.w5(32'hb9500fcc),
	.w6(32'hba0f38ac),
	.w7(32'hb9400d60),
	.w8(32'hb92f2209),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba324d37),
	.w1(32'h3a3e2d54),
	.w2(32'h3a3ec99e),
	.w3(32'hb8a6f30a),
	.w4(32'h3a3ff052),
	.w5(32'h3aad793f),
	.w6(32'hb8e53503),
	.w7(32'h3a67a8dc),
	.w8(32'h3acfe822),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb2c33),
	.w1(32'hbac6bfcf),
	.w2(32'hbb275242),
	.w3(32'hbaf3ce99),
	.w4(32'hbab0beda),
	.w5(32'hbac971f9),
	.w6(32'hbaf403cd),
	.w7(32'hba204493),
	.w8(32'hba9701ea),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7851957),
	.w1(32'hb9607952),
	.w2(32'hb99557fc),
	.w3(32'hb771d728),
	.w4(32'hb98de756),
	.w5(32'hba105a88),
	.w6(32'hb8868aeb),
	.w7(32'hb8834911),
	.w8(32'h3742a001),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad9f1c),
	.w1(32'hba524c0b),
	.w2(32'hba81ee0b),
	.w3(32'hbab01f32),
	.w4(32'hba50bc8f),
	.w5(32'hba6d1460),
	.w6(32'hbad1a7d4),
	.w7(32'hba55a4de),
	.w8(32'hba829b97),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941e800),
	.w1(32'hb9062ad9),
	.w2(32'hb8d2005c),
	.w3(32'hb98dc906),
	.w4(32'hb8e95ec7),
	.w5(32'hb8dfff38),
	.w6(32'hb9b25323),
	.w7(32'hb904e744),
	.w8(32'hb8a8e832),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ca2673),
	.w1(32'hb7077abb),
	.w2(32'h3826f170),
	.w3(32'h3782b147),
	.w4(32'hb5a18260),
	.w5(32'h38312458),
	.w6(32'hb71b3871),
	.w7(32'h37d9f860),
	.w8(32'hb69112e9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9971039),
	.w1(32'hb88dc5c4),
	.w2(32'h38cd4329),
	.w3(32'hb9853c9f),
	.w4(32'h3809c982),
	.w5(32'h39245ac2),
	.w6(32'hb9a2aa63),
	.w7(32'h373e7e08),
	.w8(32'h391b1ab4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dce9d1),
	.w1(32'hb75dbfef),
	.w2(32'h37bc70cf),
	.w3(32'h37f727f8),
	.w4(32'hb76d03df),
	.w5(32'h37ef1fba),
	.w6(32'hb6fd40f6),
	.w7(32'h37864b20),
	.w8(32'h3683eb0c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8936b9),
	.w1(32'hba415b36),
	.w2(32'hba329d16),
	.w3(32'hba0b10b5),
	.w4(32'h37a6c0d0),
	.w5(32'hba10066b),
	.w6(32'hb8a2849e),
	.w7(32'h3838fcc1),
	.w8(32'hb9a40dd2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391024a0),
	.w1(32'h3a70cd6d),
	.w2(32'h3a32109a),
	.w3(32'h3a3eedac),
	.w4(32'h3a94dc86),
	.w5(32'h3aa08c0c),
	.w6(32'h3a907e09),
	.w7(32'h3ab79c7e),
	.w8(32'h3acfce2e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64faee),
	.w1(32'hba1182f0),
	.w2(32'hba5271e2),
	.w3(32'hba23dc8c),
	.w4(32'hb9c0d5cd),
	.w5(32'hb9e129d8),
	.w6(32'hba1517db),
	.w7(32'h383b413b),
	.w8(32'hb94dc2f4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e500d2),
	.w1(32'h39024a55),
	.w2(32'h39057f9f),
	.w3(32'h38c3cce1),
	.w4(32'h38c34b2a),
	.w5(32'h3902f110),
	.w6(32'h39655eef),
	.w7(32'h38b544dc),
	.w8(32'h398fbd3c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0aa7b),
	.w1(32'hba2794a6),
	.w2(32'hba62a3bd),
	.w3(32'hbaa3e7b9),
	.w4(32'hba0b1804),
	.w5(32'hb9b18c05),
	.w6(32'hba633341),
	.w7(32'h392e1a60),
	.w8(32'h382d2241),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd51ad),
	.w1(32'hbabd9be3),
	.w2(32'hbad19a91),
	.w3(32'hbaf96953),
	.w4(32'hbae62573),
	.w5(32'hbae45a5e),
	.w6(32'hbb016ff9),
	.w7(32'hbac8b020),
	.w8(32'hbad0733d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac59204),
	.w1(32'hba891239),
	.w2(32'hbafe8da7),
	.w3(32'hba9e1950),
	.w4(32'hbab12689),
	.w5(32'hbaf70f96),
	.w6(32'hbab81a31),
	.w7(32'hba423786),
	.w8(32'hbaadaecf),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee2f9e),
	.w1(32'hb7403bf7),
	.w2(32'hb737d3db),
	.w3(32'h38e70889),
	.w4(32'h36274ca0),
	.w5(32'hb74ec63b),
	.w6(32'hb72dfc44),
	.w7(32'hb78a5431),
	.w8(32'hb7b23ee2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb814ac75),
	.w1(32'hb7ddab45),
	.w2(32'hb549328c),
	.w3(32'hb7c81850),
	.w4(32'hb7cc4e84),
	.w5(32'hb7a215cf),
	.w6(32'hb80b2ff4),
	.w7(32'hb67727c2),
	.w8(32'h374cb95b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f81302),
	.w1(32'hb79b7171),
	.w2(32'hb99c625e),
	.w3(32'hb80afc59),
	.w4(32'h38be2982),
	.w5(32'h38af9bb7),
	.w6(32'h3954d461),
	.w7(32'h3a21fdc9),
	.w8(32'h3a0997cd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9c12c),
	.w1(32'hba029cab),
	.w2(32'hb9de38c0),
	.w3(32'hbaca2bdf),
	.w4(32'hba597002),
	.w5(32'hba8bcb6e),
	.w6(32'hbab7327b),
	.w7(32'h38a7cdb0),
	.w8(32'hb905b8fa),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa31453),
	.w1(32'hba77ec94),
	.w2(32'hbaefaaba),
	.w3(32'hbaac95bf),
	.w4(32'hba4e4e5c),
	.w5(32'hbac23544),
	.w6(32'hbab89efa),
	.w7(32'hba14e74b),
	.w8(32'hbaa1a973),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984793f),
	.w1(32'hb49e1afd),
	.w2(32'h38119b54),
	.w3(32'hb9581711),
	.w4(32'hb7575c55),
	.w5(32'hb8a5f71d),
	.w6(32'hb83e6398),
	.w7(32'hb8f3c5c2),
	.w8(32'h385681c8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37093bc1),
	.w1(32'hb6e729f6),
	.w2(32'h37b501c6),
	.w3(32'h386011aa),
	.w4(32'hb7713425),
	.w5(32'h382aaa52),
	.w6(32'hb7755e51),
	.w7(32'h381220ff),
	.w8(32'h37bf3d70),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37261a14),
	.w1(32'h371949c9),
	.w2(32'h37ec8fc9),
	.w3(32'h37b3d24c),
	.w4(32'h37bf00cc),
	.w5(32'h37f327e9),
	.w6(32'h38201cc2),
	.w7(32'h388d1c0a),
	.w8(32'h3885e5ac),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399435a7),
	.w1(32'h3a0696c0),
	.w2(32'h39b416f1),
	.w3(32'hb774a7cb),
	.w4(32'h39e540bf),
	.w5(32'h3a009801),
	.w6(32'hb9bf676d),
	.w7(32'h39955dad),
	.w8(32'h38fe6007),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e2e40d),
	.w1(32'h39d8519f),
	.w2(32'hb95a57a6),
	.w3(32'hb9077d9c),
	.w4(32'h396a173a),
	.w5(32'hba8645ae),
	.w6(32'hba3b3948),
	.w7(32'hb9b14c8c),
	.w8(32'hbab1e759),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38316f5a),
	.w1(32'h39a55b1d),
	.w2(32'h39e17b94),
	.w3(32'hb91925f9),
	.w4(32'h39b81068),
	.w5(32'h39e436b5),
	.w6(32'hb97ecc58),
	.w7(32'h3903dffc),
	.w8(32'hb7f2dacf),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91228be),
	.w1(32'h392593bc),
	.w2(32'h39001dea),
	.w3(32'h3872cc25),
	.w4(32'h39aeb2f6),
	.w5(32'h39bd2491),
	.w6(32'h398f49a3),
	.w7(32'h39fdca4b),
	.w8(32'h3a188b29),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6103ef),
	.w1(32'hb9d90ef7),
	.w2(32'hba347d1c),
	.w3(32'hba273d44),
	.w4(32'hb98ed075),
	.w5(32'hb94fe54b),
	.w6(32'hb9d864fc),
	.w7(32'h39f011a3),
	.w8(32'h39a2c5e6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d657b6),
	.w1(32'h35ecc097),
	.w2(32'h36568424),
	.w3(32'h38d38b79),
	.w4(32'hb6581ae5),
	.w5(32'h367db64f),
	.w6(32'h36c66130),
	.w7(32'h351d3c11),
	.w8(32'h36c1c5f7),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371601b4),
	.w1(32'hb7ddc068),
	.w2(32'h381f063a),
	.w3(32'h376ceead),
	.w4(32'hb7e43c01),
	.w5(32'h371d9753),
	.w6(32'hb8264a10),
	.w7(32'h3541dbe6),
	.w8(32'hb836aa88),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb846ef01),
	.w1(32'hb923e314),
	.w2(32'h382dc7cd),
	.w3(32'hb8231594),
	.w4(32'hb8e30a58),
	.w5(32'h388ec2c9),
	.w6(32'hb8f5b57a),
	.w7(32'h380e02ee),
	.w8(32'h38a31375),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388995e3),
	.w1(32'h37b53ade),
	.w2(32'hb8e6884f),
	.w3(32'h387f0ba8),
	.w4(32'h36ee387c),
	.w5(32'hb8ce54b7),
	.w6(32'h37f01f4b),
	.w7(32'hb8b108f4),
	.w8(32'h381c39b5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84d767f),
	.w1(32'hb88bbc34),
	.w2(32'hb6438fd1),
	.w3(32'hb816c117),
	.w4(32'hb8311503),
	.w5(32'hb805302e),
	.w6(32'hb8d9e7c6),
	.w7(32'hb86ee6b3),
	.w8(32'h380ca861),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e7369),
	.w1(32'hb89a1373),
	.w2(32'hb9f67cb9),
	.w3(32'hba67ca8c),
	.w4(32'hb93b82b2),
	.w5(32'hba38ba40),
	.w6(32'hba4cee99),
	.w7(32'hb942be4a),
	.w8(32'hba3b862c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2dd9aa),
	.w1(32'hba053d6d),
	.w2(32'hba08cfd5),
	.w3(32'hba423cd1),
	.w4(32'hba0e4a83),
	.w5(32'hb9fdb02e),
	.w6(32'hba37af8f),
	.w7(32'hb8beca2c),
	.w8(32'hb9b4c43e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8933039),
	.w1(32'hb8435c69),
	.w2(32'h3919c150),
	.w3(32'h36761f75),
	.w4(32'hb8281e0e),
	.w5(32'h38cd232b),
	.w6(32'hb8ecb70b),
	.w7(32'h38253a52),
	.w8(32'hb8398375),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11a024),
	.w1(32'h39bb0621),
	.w2(32'h3a11179e),
	.w3(32'hba5ffb38),
	.w4(32'h37046121),
	.w5(32'h38e839fc),
	.w6(32'hba77d464),
	.w7(32'hb975d17a),
	.w8(32'hb94be976),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6211f),
	.w1(32'h395775ce),
	.w2(32'hb8e0f946),
	.w3(32'hba022b62),
	.w4(32'hb8dd59d7),
	.w5(32'hb99b62ab),
	.w6(32'hba129e0d),
	.w7(32'hb7ac3b3a),
	.w8(32'hb8ee569a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369d7b0e),
	.w1(32'h3909de93),
	.w2(32'h394b3c52),
	.w3(32'h377b9c93),
	.w4(32'h3931d83f),
	.w5(32'h3954e0e6),
	.w6(32'h381a3c5a),
	.w7(32'h39743e90),
	.w8(32'h39341a06),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a9347),
	.w1(32'hb9a0d3f1),
	.w2(32'hb9c19c66),
	.w3(32'hba253d49),
	.w4(32'hb9d24d09),
	.w5(32'hba04c80e),
	.w6(32'hba3a2855),
	.w7(32'hba0b8b23),
	.w8(32'hba0de53c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d46f91),
	.w1(32'h36d84f84),
	.w2(32'hb6dd0a27),
	.w3(32'h381168e6),
	.w4(32'h37287cf5),
	.w5(32'hb70e896b),
	.w6(32'h379aadd1),
	.w7(32'h354085fe),
	.w8(32'hb7afe1ab),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8b271),
	.w1(32'h38a5c6ae),
	.w2(32'h3920508c),
	.w3(32'h38828aca),
	.w4(32'h38d56488),
	.w5(32'h39161ec2),
	.w6(32'h38580045),
	.w7(32'h38ecf943),
	.w8(32'h390859fd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f5f61b),
	.w1(32'hb8231e33),
	.w2(32'h3625d862),
	.w3(32'h38196c8b),
	.w4(32'hb7fe9b42),
	.w5(32'h3625abaf),
	.w6(32'hb6a59082),
	.w7(32'h380053b7),
	.w8(32'h3570a845),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb552d828),
	.w1(32'hb73e836e),
	.w2(32'hb853ff59),
	.w3(32'hb5dab8d9),
	.w4(32'hb6d481c1),
	.w5(32'hb823bb3e),
	.w6(32'hb6fffa50),
	.w7(32'hb818224f),
	.w8(32'h37b3b838),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f29289),
	.w1(32'h3a64f096),
	.w2(32'h3ace867e),
	.w3(32'h3a21c557),
	.w4(32'h3a6ed9b9),
	.w5(32'h3acc1c50),
	.w6(32'h3a5b29b6),
	.w7(32'h3a669798),
	.w8(32'h3abe0377),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb5979),
	.w1(32'hba3aac9a),
	.w2(32'hbadd2170),
	.w3(32'hbb02a332),
	.w4(32'hba9b3a5d),
	.w5(32'hbb031ef2),
	.w6(32'hbaf473c2),
	.w7(32'hba6ae38d),
	.w8(32'hba99c970),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa11a48),
	.w1(32'hba410da9),
	.w2(32'hbac51a54),
	.w3(32'hbac2f480),
	.w4(32'hba8ae86b),
	.w5(32'hbac8c44c),
	.w6(32'hbace7143),
	.w7(32'hba774e9c),
	.w8(32'hba8e991c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87c3f2),
	.w1(32'hba1fccec),
	.w2(32'hba941498),
	.w3(32'hba9735a3),
	.w4(32'hba606363),
	.w5(32'hbac6b5e4),
	.w6(32'hbac56d75),
	.w7(32'hba71e4fe),
	.w8(32'hbaacc87e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932a31f),
	.w1(32'hb888c0f2),
	.w2(32'hb923ca2c),
	.w3(32'hb93b3263),
	.w4(32'hb9088531),
	.w5(32'hb900bba1),
	.w6(32'hb92f748c),
	.w7(32'hb8d692f1),
	.w8(32'hb804e9bf),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38288b91),
	.w1(32'hb8503fb8),
	.w2(32'h37bc60be),
	.w3(32'h382895ea),
	.w4(32'hb83d06f0),
	.w5(32'h37f492fd),
	.w6(32'hb8250d32),
	.w7(32'h37e9d23e),
	.w8(32'h37379768),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74addaa),
	.w1(32'hb7db3d4b),
	.w2(32'h378ea1d5),
	.w3(32'hb74d1538),
	.w4(32'hb7a8e870),
	.w5(32'h37b20af3),
	.w6(32'hb7a924c1),
	.w7(32'h37076b28),
	.w8(32'hb735769d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374f8ec6),
	.w1(32'hb77c019b),
	.w2(32'h37abd74a),
	.w3(32'h370d3463),
	.w4(32'h3703a6a1),
	.w5(32'h384aad3b),
	.w6(32'hb6fbb2bf),
	.w7(32'h380a5389),
	.w8(32'h3738650a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387c7727),
	.w1(32'h3a1c0b84),
	.w2(32'h38da87c7),
	.w3(32'h391a7c73),
	.w4(32'h3a2e8256),
	.w5(32'h399deb37),
	.w6(32'h38b0f899),
	.w7(32'h3a18e2bb),
	.w8(32'h39e6521a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d0c5e),
	.w1(32'hb907aaed),
	.w2(32'h37ae101a),
	.w3(32'hb902a0e3),
	.w4(32'hb9276a49),
	.w5(32'h3741e019),
	.w6(32'hb91169fa),
	.w7(32'hb8b02160),
	.w8(32'hb867a5c5),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399be297),
	.w1(32'h393668f6),
	.w2(32'h39c78657),
	.w3(32'h39ba10ee),
	.w4(32'h396412f2),
	.w5(32'h39cff8ae),
	.w6(32'h39d07ec3),
	.w7(32'h39cfada4),
	.w8(32'h39f20002),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d511c0),
	.w1(32'hb8c2f2ad),
	.w2(32'hb83cb8ef),
	.w3(32'hb90b5d36),
	.w4(32'hb8f439b9),
	.w5(32'hb801ff2d),
	.w6(32'hb81a84f7),
	.w7(32'hb79fc2ce),
	.w8(32'h38572801),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cb3ca7),
	.w1(32'hb82bb40e),
	.w2(32'hb7518f7e),
	.w3(32'hb7d464db),
	.w4(32'hb80ed764),
	.w5(32'hb73ec87b),
	.w6(32'hb7c2b1ac),
	.w7(32'hb71d8708),
	.w8(32'hb7bd530b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a0f54),
	.w1(32'h399161d5),
	.w2(32'h389719ad),
	.w3(32'h38670620),
	.w4(32'h39407a20),
	.w5(32'hb837a174),
	.w6(32'hb8ff9921),
	.w7(32'h3884ee42),
	.w8(32'hb83a7eec),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b89560),
	.w1(32'hb8baade4),
	.w2(32'h375fe8bc),
	.w3(32'hb88f7d95),
	.w4(32'hb891e315),
	.w5(32'h380baac1),
	.w6(32'hb88eaf34),
	.w7(32'h373a6427),
	.w8(32'hb6712f76),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c541a),
	.w1(32'hb951d6e2),
	.w2(32'hba12ef1d),
	.w3(32'hba70035f),
	.w4(32'hb9eb0cc4),
	.w5(32'hba2c92c6),
	.w6(32'hb9abe1ed),
	.w7(32'h38d604ab),
	.w8(32'h3867142f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3695c7a3),
	.w1(32'h39f42d95),
	.w2(32'h3a1fe04a),
	.w3(32'h37b27923),
	.w4(32'h3a09b14a),
	.w5(32'h3a192e50),
	.w6(32'h39beb12c),
	.w7(32'h3a0e0d6b),
	.w8(32'h3a2fc88a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72c87f),
	.w1(32'hba8f4eaa),
	.w2(32'hbb73540d),
	.w3(32'hba4cf4c3),
	.w4(32'hbb187fe1),
	.w5(32'hbb5f0518),
	.w6(32'hb9cd621b),
	.w7(32'hb9b43452),
	.w8(32'hba9a45f5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule