module layer_10_featuremap_122(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c4c555),
	.w1(32'hb77a4eb7),
	.w2(32'hb76db62f),
	.w3(32'hb769ebad),
	.w4(32'hb77fa04b),
	.w5(32'hb53bef9d),
	.w6(32'hb7361822),
	.w7(32'hb71b011b),
	.w8(32'h3668a75e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac69356),
	.w1(32'hbac7091a),
	.w2(32'hba83dd76),
	.w3(32'hba0cc099),
	.w4(32'hba793566),
	.w5(32'hba435bee),
	.w6(32'hb9b192c5),
	.w7(32'hb9bf2fc7),
	.w8(32'h39e24eea),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb628e622),
	.w1(32'hb5e6d1a0),
	.w2(32'hb5ad445e),
	.w3(32'h360ee473),
	.w4(32'h362ee17a),
	.w5(32'h3626687c),
	.w6(32'h36515460),
	.w7(32'h36706676),
	.w8(32'h36568c92),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903b191),
	.w1(32'h39d2196f),
	.w2(32'h3a07de6d),
	.w3(32'hb9bba533),
	.w4(32'h370ed5d2),
	.w5(32'hb8489265),
	.w6(32'hba034844),
	.w7(32'hb87e11f2),
	.w8(32'hba49cc10),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77bfae1),
	.w1(32'hb687a225),
	.w2(32'h372c32fe),
	.w3(32'hb6ec717d),
	.w4(32'h36f8caed),
	.w5(32'h37e5d8e9),
	.w6(32'hb6499154),
	.w7(32'h374f4639),
	.w8(32'h36ea5f3f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b00d02),
	.w1(32'h35574745),
	.w2(32'hb6781540),
	.w3(32'h3659871d),
	.w4(32'h35b5c8d9),
	.w5(32'hb60c29a1),
	.w6(32'h36be9dd2),
	.w7(32'h36b00fa8),
	.w8(32'h368841c0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17c6df),
	.w1(32'h38e7f870),
	.w2(32'hbb73a3f9),
	.w3(32'h39db2610),
	.w4(32'h399da2d4),
	.w5(32'hbb40687f),
	.w6(32'h3a3dba86),
	.w7(32'hbb18ba1b),
	.w8(32'hbb5c7c23),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86df71),
	.w1(32'h39c83198),
	.w2(32'hbaea189f),
	.w3(32'hbbe287cf),
	.w4(32'hbb19bc27),
	.w5(32'h3b0b51c2),
	.w6(32'hbc0ea4e4),
	.w7(32'hbbbcfbbc),
	.w8(32'hba9cc06b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ffb61),
	.w1(32'hb897a6e2),
	.w2(32'h3888136c),
	.w3(32'hb938df3e),
	.w4(32'hb91a046a),
	.w5(32'h37db8d34),
	.w6(32'hb9b8133e),
	.w7(32'hb9a139f0),
	.w8(32'hb92d828e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb760f045),
	.w1(32'h3a6c4128),
	.w2(32'h3a99359b),
	.w3(32'hbab7eff3),
	.w4(32'h3a738206),
	.w5(32'h3a07a7c0),
	.w6(32'hbb558f51),
	.w7(32'hbb036e77),
	.w8(32'hba09fe97),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h358e8708),
	.w1(32'h37c21c44),
	.w2(32'hb73bfdf8),
	.w3(32'hb697ea8a),
	.w4(32'h38180946),
	.w5(32'hb8336364),
	.w6(32'hb85e498d),
	.w7(32'h3690867b),
	.w8(32'hb6093edb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b592dc9),
	.w1(32'h3aca8d52),
	.w2(32'hbb3104b0),
	.w3(32'h3addfff2),
	.w4(32'h3b5d3cdc),
	.w5(32'hbaf042e4),
	.w6(32'h3aa82ac5),
	.w7(32'h3a215957),
	.w8(32'hbb333ead),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab61fbe),
	.w1(32'h3b1b304e),
	.w2(32'h3b56b43b),
	.w3(32'hbb1cb04d),
	.w4(32'h3a421743),
	.w5(32'h3a97960c),
	.w6(32'hbb352a4a),
	.w7(32'hbb3aa3e5),
	.w8(32'hb9c09873),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba899f04),
	.w1(32'hba62992a),
	.w2(32'hba91cc0e),
	.w3(32'hba3cf44b),
	.w4(32'hb7e097dc),
	.w5(32'h3ac77c2b),
	.w6(32'hba1928da),
	.w7(32'hba3769ca),
	.w8(32'h3a688b2d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a80b0f),
	.w1(32'hb9983175),
	.w2(32'h3a22d674),
	.w3(32'h3950f69c),
	.w4(32'hba90d747),
	.w5(32'hba151cdd),
	.w6(32'hb9e28f0a),
	.w7(32'h38111466),
	.w8(32'h3a29e9b2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6469ed),
	.w1(32'hbae83974),
	.w2(32'h3a9e429f),
	.w3(32'hbb2d9797),
	.w4(32'h3a09d989),
	.w5(32'h3b3840c4),
	.w6(32'hbb2f9711),
	.w7(32'hbb367248),
	.w8(32'hb9b6e748),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9d511),
	.w1(32'hb88973cd),
	.w2(32'hb8844a35),
	.w3(32'h37b2ffa0),
	.w4(32'hb5cdf0b9),
	.w5(32'h373c2380),
	.w6(32'h3885c302),
	.w7(32'h38743301),
	.w8(32'h387cd87a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f3c57),
	.w1(32'h3a9765f3),
	.w2(32'h3abaaafc),
	.w3(32'hbb1f4f13),
	.w4(32'hba4820b0),
	.w5(32'h39c14857),
	.w6(32'hbba16e85),
	.w7(32'hbc1160f4),
	.w8(32'hbba006c6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c27ad),
	.w1(32'h3a9f3b40),
	.w2(32'h3b1c72da),
	.w3(32'hbac47191),
	.w4(32'h38f5c64a),
	.w5(32'h3a15544e),
	.w6(32'hbb1981f0),
	.w7(32'hbb79dedb),
	.w8(32'hbb499ae1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376b146f),
	.w1(32'hb7ed335a),
	.w2(32'hb78f09c4),
	.w3(32'h384b9e9e),
	.w4(32'hb78e4770),
	.w5(32'hb7a5ed43),
	.w6(32'hb74b0abc),
	.w7(32'h358e0ddb),
	.w8(32'hb8fa81b9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8255d65),
	.w1(32'hb8d00719),
	.w2(32'hb801495b),
	.w3(32'h37c5b4f7),
	.w4(32'hb85fe294),
	.w5(32'h384149c6),
	.w6(32'h3744e19b),
	.w7(32'h379c0db6),
	.w8(32'h3797d67e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9927f54),
	.w1(32'hb992d2c9),
	.w2(32'hb92bbd2e),
	.w3(32'hb903c96e),
	.w4(32'hb9952201),
	.w5(32'hb9a6343a),
	.w6(32'h3984c29f),
	.w7(32'h39bef34e),
	.w8(32'h39a40aac),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adea7c4),
	.w1(32'h3b07279d),
	.w2(32'h3b21334d),
	.w3(32'hbae7f9ba),
	.w4(32'h3b0a7922),
	.w5(32'hbb3aebff),
	.w6(32'hbb15484b),
	.w7(32'hbb95e1ef),
	.w8(32'hbc1ab77f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f1e22),
	.w1(32'h3aa1f0ac),
	.w2(32'h3b031f5e),
	.w3(32'h38383ff2),
	.w4(32'h39cbcd53),
	.w5(32'hb9b77cd6),
	.w6(32'hbb279047),
	.w7(32'hbad34723),
	.w8(32'h3966f035),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e464a),
	.w1(32'h39d512b3),
	.w2(32'h3af97262),
	.w3(32'hb80cb24e),
	.w4(32'hbadafa9e),
	.w5(32'hbac74b30),
	.w6(32'h36ddd430),
	.w7(32'hbaca5afa),
	.w8(32'h39e92e37),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d71b95),
	.w1(32'h365535de),
	.w2(32'hb780018c),
	.w3(32'hb82961f7),
	.w4(32'h382affd3),
	.w5(32'h38c0982c),
	.w6(32'h38684479),
	.w7(32'h389d0b12),
	.w8(32'h376bbd2b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d9b1ab),
	.w1(32'hb80225f1),
	.w2(32'hb80ed0ae),
	.w3(32'h37b9baeb),
	.w4(32'hb6e39eda),
	.w5(32'hb7668ee3),
	.w6(32'h384df6bf),
	.w7(32'h38462a86),
	.w8(32'h37ff27b2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11644d),
	.w1(32'hbaf527bb),
	.w2(32'hbaf7078b),
	.w3(32'h3acba3bb),
	.w4(32'h3aa6e9e7),
	.w5(32'hb9b26cbe),
	.w6(32'h3b7de703),
	.w7(32'h3bad5cbc),
	.w8(32'h3bc9ce2b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38236f9f),
	.w1(32'hb9e41386),
	.w2(32'hb98053f4),
	.w3(32'h39580d04),
	.w4(32'hb9da0f16),
	.w5(32'hb9e74c24),
	.w6(32'h3a686132),
	.w7(32'h3a193ce8),
	.w8(32'h3a18ef28),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bc44b),
	.w1(32'hba2853d0),
	.w2(32'hb9b89b61),
	.w3(32'h3a76c0b5),
	.w4(32'hba000c98),
	.w5(32'hbadee6b3),
	.w6(32'h3b434bbf),
	.w7(32'h3ac43568),
	.w8(32'h3af35b67),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h348801f4),
	.w1(32'hb713a2f7),
	.w2(32'hb6990154),
	.w3(32'h371dbbd2),
	.w4(32'hb69742c8),
	.w5(32'hb5179414),
	.w6(32'h378fe702),
	.w7(32'h377449e8),
	.w8(32'h37a1854d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75689f5),
	.w1(32'hb789ba29),
	.w2(32'hb768b9f5),
	.w3(32'hb79d30b9),
	.w4(32'hb7bfee98),
	.w5(32'hb7708471),
	.w6(32'hb7c78e9e),
	.w7(32'hb714366e),
	.w8(32'hb6c7c6c4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ee7872),
	.w1(32'h39c11be9),
	.w2(32'h3a804901),
	.w3(32'hba0bcd51),
	.w4(32'h3a24e4c9),
	.w5(32'h3a6cfd13),
	.w6(32'hbaa1a879),
	.w7(32'hba5c2fed),
	.w8(32'h382f969f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e48bb),
	.w1(32'hb93f2a22),
	.w2(32'h383a295c),
	.w3(32'h3a10ddd0),
	.w4(32'h39755978),
	.w5(32'h39bab294),
	.w6(32'h3a507c2d),
	.w7(32'h3a6d3c5d),
	.w8(32'h3a8fb10a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39293bba),
	.w1(32'hb90e8547),
	.w2(32'hb92a3602),
	.w3(32'h38502e9c),
	.w4(32'h398360cc),
	.w5(32'hb96b526b),
	.w6(32'h398aefc1),
	.w7(32'h39278594),
	.w8(32'h399d1df3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8acc486),
	.w1(32'h3a328d05),
	.w2(32'hb9a4691b),
	.w3(32'hba42bea0),
	.w4(32'h38f855e5),
	.w5(32'hb9802907),
	.w6(32'hba52d471),
	.w7(32'hba5361fc),
	.w8(32'hbaf00681),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad295a4),
	.w1(32'h3ab29db5),
	.w2(32'hbaec2b37),
	.w3(32'hbba66e76),
	.w4(32'hbad32aa1),
	.w5(32'h3aa92735),
	.w6(32'hbbd03d43),
	.w7(32'h3ac21009),
	.w8(32'hbc15eccf),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8a579),
	.w1(32'hbb8cc304),
	.w2(32'hbaec564f),
	.w3(32'h3a6a6e4b),
	.w4(32'hbb37b549),
	.w5(32'hbb28d73b),
	.w6(32'h3abf7257),
	.w7(32'h3b177f47),
	.w8(32'h3b536d3c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea9e4f),
	.w1(32'hbb56ec81),
	.w2(32'hbb466ada),
	.w3(32'h3ae7b553),
	.w4(32'hbb43c4db),
	.w5(32'hbb9b54b2),
	.w6(32'h3ba663fa),
	.w7(32'h3b6cb6a5),
	.w8(32'h3b8b0d15),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aeb968),
	.w1(32'hb8af3b4e),
	.w2(32'h38bf48ad),
	.w3(32'hb9e501e3),
	.w4(32'hb972fbb6),
	.w5(32'hb883b2f5),
	.w6(32'hba0e9394),
	.w7(32'h38d75e36),
	.w8(32'h3a08f1d8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e67255),
	.w1(32'hb885950e),
	.w2(32'hb862aa35),
	.w3(32'hb8988d0c),
	.w4(32'hb82662c0),
	.w5(32'hb8328da9),
	.w6(32'hb83789c0),
	.w7(32'hb7ce4bf7),
	.w8(32'hb8476724),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fafe4e),
	.w1(32'hb89839ee),
	.w2(32'hb8231582),
	.w3(32'h38a0da07),
	.w4(32'h38137583),
	.w5(32'h37e76c72),
	.w6(32'h38e78a29),
	.w7(32'h38dae53d),
	.w8(32'h38d74ded),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391fa3a2),
	.w1(32'hba7991e1),
	.w2(32'hb9e6f00b),
	.w3(32'h3938f0de),
	.w4(32'hba553ea3),
	.w5(32'hb8b5f53e),
	.w6(32'h3a2abb9d),
	.w7(32'hb97b43f4),
	.w8(32'h39871f24),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b0201),
	.w1(32'h3a902ec0),
	.w2(32'h3af39b0a),
	.w3(32'hbab7e010),
	.w4(32'h3abbbecf),
	.w5(32'hba02c4fe),
	.w6(32'hbb2ebe8c),
	.w7(32'hbb28bc53),
	.w8(32'hba5b14b8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ac372),
	.w1(32'h3a8ecd62),
	.w2(32'h3b072f01),
	.w3(32'h3a4f7474),
	.w4(32'h38808a3b),
	.w5(32'h39f027a4),
	.w6(32'h39f3a7d8),
	.w7(32'h3982a094),
	.w8(32'h3a9d0b7b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922521c),
	.w1(32'h3b48c4be),
	.w2(32'h3b792a78),
	.w3(32'h3a0edde9),
	.w4(32'h3a82e5ea),
	.w5(32'h3b012be2),
	.w6(32'hbaca6f23),
	.w7(32'hba46aed8),
	.w8(32'h39cfdbc0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f3cb3a),
	.w1(32'h39d4c5c9),
	.w2(32'h3a8f99eb),
	.w3(32'hb98eac7c),
	.w4(32'h39e7ba4c),
	.w5(32'h39d492b1),
	.w6(32'hba629545),
	.w7(32'h3980876a),
	.w8(32'h3a1d0bd6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a640fe9),
	.w1(32'h39ca5ef2),
	.w2(32'h3aeb3083),
	.w3(32'hbb97f264),
	.w4(32'hbb0cd026),
	.w5(32'hb9138449),
	.w6(32'hbc135330),
	.w7(32'hbc364132),
	.w8(32'hbc28560a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3742f413),
	.w1(32'h380cb1de),
	.w2(32'hb6ed0a3b),
	.w3(32'h38487158),
	.w4(32'h3880c30d),
	.w5(32'h37f05d1d),
	.w6(32'h38fd081d),
	.w7(32'h38c717a4),
	.w8(32'h3811d365),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e89af5),
	.w1(32'h396208e3),
	.w2(32'h38893267),
	.w3(32'h392b4705),
	.w4(32'h396bf590),
	.w5(32'h38357c0d),
	.w6(32'h3948b9c5),
	.w7(32'h391602f1),
	.w8(32'hb7fec546),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf20cd),
	.w1(32'h38bd949e),
	.w2(32'h384ac741),
	.w3(32'h3944a596),
	.w4(32'h392088a3),
	.w5(32'h38cebb2a),
	.w6(32'h394ab03d),
	.w7(32'h392a7967),
	.w8(32'h3891126e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3d5ac),
	.w1(32'h3a5474e2),
	.w2(32'h3adedde7),
	.w3(32'hba27866f),
	.w4(32'hb91b007a),
	.w5(32'h38ea3d3b),
	.w6(32'hba30c8ea),
	.w7(32'hba60fac8),
	.w8(32'hba98f3ac),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c12bfa),
	.w1(32'h3970b160),
	.w2(32'h398f7949),
	.w3(32'hb9a6da6b),
	.w4(32'h39510bd8),
	.w5(32'h3918940b),
	.w6(32'hba068d39),
	.w7(32'hb9069409),
	.w8(32'hb9c70feb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0d678),
	.w1(32'h3a45a729),
	.w2(32'h3aabd902),
	.w3(32'hba73185c),
	.w4(32'h3af29d0b),
	.w5(32'h3ae4ec77),
	.w6(32'hbb4f52a9),
	.w7(32'hbb9fbf8b),
	.w8(32'hbba1d133),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38541b04),
	.w1(32'h39c77759),
	.w2(32'hb9582203),
	.w3(32'h3a2ec889),
	.w4(32'h39499aff),
	.w5(32'hb904fecb),
	.w6(32'h3a2add5c),
	.w7(32'h3788ac6d),
	.w8(32'h39587ae6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38143def),
	.w1(32'hb82223f9),
	.w2(32'hb74ea8ae),
	.w3(32'h386b5ba3),
	.w4(32'hb8b3bed7),
	.w5(32'hb867a975),
	.w6(32'h38f69e0c),
	.w7(32'h389ef363),
	.w8(32'h386b0ff6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72686d0),
	.w1(32'hb6df5ef1),
	.w2(32'hb3474cb8),
	.w3(32'hb7a857dd),
	.w4(32'hb7a3148b),
	.w5(32'h3591231f),
	.w6(32'hb7961df7),
	.w7(32'h36a75f05),
	.w8(32'h37d3a4ca),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38973b98),
	.w1(32'hb890668c),
	.w2(32'hb9aaa213),
	.w3(32'h392ef370),
	.w4(32'hb9694144),
	.w5(32'hb9ff97a7),
	.w6(32'h39c46e4b),
	.w7(32'hb8d1090a),
	.w8(32'hb93abccc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ebdbe),
	.w1(32'hb9e39577),
	.w2(32'hb6368c56),
	.w3(32'hb985b1b6),
	.w4(32'hba17f761),
	.w5(32'hb8ec5978),
	.w6(32'h392565be),
	.w7(32'h3762dc37),
	.w8(32'h398a8837),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a5cc0),
	.w1(32'hb8b1946b),
	.w2(32'hb89c07c3),
	.w3(32'h39afa7ff),
	.w4(32'h380b3226),
	.w5(32'hb963b272),
	.w6(32'h39af20a6),
	.w7(32'hb90f365e),
	.w8(32'h38476b34),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48591d),
	.w1(32'h3a834100),
	.w2(32'h3ac6ac5f),
	.w3(32'h39f4f7a9),
	.w4(32'h3ada93f7),
	.w5(32'h3a3bbcfc),
	.w6(32'hb990a60b),
	.w7(32'hbad6e067),
	.w8(32'hba821e9c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56b435),
	.w1(32'hbadee4a5),
	.w2(32'h39d8923d),
	.w3(32'h3a790c1d),
	.w4(32'h3a3f4159),
	.w5(32'hb861344e),
	.w6(32'h3a9538f9),
	.w7(32'hba5ffd68),
	.w8(32'h3a26f85f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e88eca),
	.w1(32'hb6a8aaea),
	.w2(32'hb6e092b1),
	.w3(32'h365ae64b),
	.w4(32'h36e750b2),
	.w5(32'h369b41df),
	.w6(32'h37884fb9),
	.w7(32'h3783408a),
	.w8(32'h3795b588),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3705f0a7),
	.w1(32'h3488713c),
	.w2(32'hb66b61f4),
	.w3(32'h374824e8),
	.w4(32'h35fd8b68),
	.w5(32'hb6c14b32),
	.w6(32'h37510e07),
	.w7(32'h35e34190),
	.w8(32'h343e0f6a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb813271a),
	.w1(32'hb8348d17),
	.w2(32'hb7a26f14),
	.w3(32'hb7dc00ed),
	.w4(32'hb75608ad),
	.w5(32'hb6a3fc08),
	.w6(32'hb7ea1431),
	.w7(32'hb783fae8),
	.w8(32'h3499bf90),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79a8716),
	.w1(32'hb7d8325a),
	.w2(32'hb76712e0),
	.w3(32'hb639925f),
	.w4(32'hb69f0020),
	.w5(32'h35a91878),
	.w6(32'h373be1ce),
	.w7(32'h37a7142c),
	.w8(32'h37657737),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05aceb),
	.w1(32'hbb9aef9e),
	.w2(32'hbafe29be),
	.w3(32'hbb15290a),
	.w4(32'h3ad201ae),
	.w5(32'h3b11b309),
	.w6(32'hbae026f1),
	.w7(32'h38d955db),
	.w8(32'h3b8c747f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0afc39),
	.w1(32'h3b07b618),
	.w2(32'h3b31327d),
	.w3(32'hbab3870e),
	.w4(32'h39dedacd),
	.w5(32'h3b0e95db),
	.w6(32'hbad3b237),
	.w7(32'hba29faf2),
	.w8(32'h396afcbe),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ac872),
	.w1(32'hb9cdc2c1),
	.w2(32'h3a9436e9),
	.w3(32'h3a92937e),
	.w4(32'h3a301eba),
	.w5(32'hba02c786),
	.w6(32'h39526028),
	.w7(32'hba1d7d63),
	.w8(32'hb9311d33),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44ad42),
	.w1(32'hb91eb7a4),
	.w2(32'h39a2c955),
	.w3(32'hba2b4ead),
	.w4(32'hbafc9b0b),
	.w5(32'hbb758353),
	.w6(32'hba6f3b1b),
	.w7(32'hba1243e5),
	.w8(32'h3a61c8b7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb793864f),
	.w1(32'hb7168637),
	.w2(32'hb7e43574),
	.w3(32'h36b0035d),
	.w4(32'hb5bce00d),
	.w5(32'hb72cfbcf),
	.w6(32'h3601a1c1),
	.w7(32'hb7354e73),
	.w8(32'hb8101f7a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83dff42),
	.w1(32'hb837777d),
	.w2(32'hb8104f46),
	.w3(32'hb783ab69),
	.w4(32'hb7747637),
	.w5(32'h345ef984),
	.w6(32'h34f83cda),
	.w7(32'h372a0035),
	.w8(32'h37428d84),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb817841f),
	.w1(32'hb79db6f4),
	.w2(32'hb56ac8ee),
	.w3(32'h34ebc338),
	.w4(32'h380dc053),
	.w5(32'h379c05ea),
	.w6(32'h37c55ed3),
	.w7(32'h37b70f55),
	.w8(32'h37dc3c67),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28d15d),
	.w1(32'h3a06bccb),
	.w2(32'h3a69c7b5),
	.w3(32'h39a71cef),
	.w4(32'h3a335ff3),
	.w5(32'h3a8ebe5b),
	.w6(32'hba12d1a1),
	.w7(32'hba6adf77),
	.w8(32'h39214f96),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb758328b),
	.w1(32'hb79e6a6e),
	.w2(32'hb7f93b28),
	.w3(32'h369ea26b),
	.w4(32'hb5a19034),
	.w5(32'hb712854c),
	.w6(32'h3772bccf),
	.w7(32'h37019547),
	.w8(32'hb611929f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d84b62),
	.w1(32'hba2bf165),
	.w2(32'hbad92b4c),
	.w3(32'hbaf2c556),
	.w4(32'hb9b1be99),
	.w5(32'h3a37861e),
	.w6(32'hbae51c68),
	.w7(32'hba9c5b71),
	.w8(32'hbb876ee5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54a754),
	.w1(32'h38a93cad),
	.w2(32'hbb05df88),
	.w3(32'hbb880c5b),
	.w4(32'hba69d291),
	.w5(32'h39d0b318),
	.w6(32'hbba60921),
	.w7(32'hbb45ad68),
	.w8(32'hbba73144),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a13d16),
	.w1(32'h3a68f80f),
	.w2(32'h3afce2b2),
	.w3(32'hbb0551cc),
	.w4(32'hbadc1731),
	.w5(32'hb94585aa),
	.w6(32'hbaf693e6),
	.w7(32'hbae77f6c),
	.w8(32'hb8ccf4e8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391676e1),
	.w1(32'h3881fcb5),
	.w2(32'h39e27701),
	.w3(32'hb95df5f8),
	.w4(32'h3a577909),
	.w5(32'h3a6e70ba),
	.w6(32'hba1d58de),
	.w7(32'hba39a426),
	.w8(32'h3a0ffe4c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbcf27),
	.w1(32'hba8a9cea),
	.w2(32'hba7664bd),
	.w3(32'hba8d19d5),
	.w4(32'h38e6ddde),
	.w5(32'hb7e1a6cf),
	.w6(32'h38e12b71),
	.w7(32'h39afd78f),
	.w8(32'h3a110f3f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26ea8b),
	.w1(32'h3987fd2f),
	.w2(32'h3a4e1ac5),
	.w3(32'h3a8b037f),
	.w4(32'h3a0fc1ba),
	.w5(32'h39f47f32),
	.w6(32'h39ed17b8),
	.w7(32'h38e5ff35),
	.w8(32'h3aaf4d2c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eaa27),
	.w1(32'h3a299c71),
	.w2(32'h3a06674a),
	.w3(32'hba60b94a),
	.w4(32'h395cc10d),
	.w5(32'h3907532c),
	.w6(32'hbaeaa597),
	.w7(32'hbb13f4d3),
	.w8(32'hbb442b64),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dbd85b),
	.w1(32'hb74df2e8),
	.w2(32'hb76726b2),
	.w3(32'hb6dba5fa),
	.w4(32'hb6114435),
	.w5(32'hb66b26f0),
	.w6(32'hb6e2188b),
	.w7(32'h365f5d92),
	.w8(32'h365ca4e1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb818ce11),
	.w1(32'hb81f92ff),
	.w2(32'hb68fe2bd),
	.w3(32'hb797a770),
	.w4(32'hb78cf75f),
	.w5(32'h35073201),
	.w6(32'h360d01ca),
	.w7(32'hb723ddfd),
	.w8(32'hb6cbaa1e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb712c6da),
	.w1(32'hb6e43dc4),
	.w2(32'h36dd476e),
	.w3(32'hb6e0251a),
	.w4(32'h36b81a0d),
	.w5(32'h377c1fa5),
	.w6(32'hb4e6d4ac),
	.w7(32'h3773297b),
	.w8(32'h3728b2c0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39431218),
	.w1(32'hb981dfc0),
	.w2(32'hb986c1b3),
	.w3(32'h38b06482),
	.w4(32'hb94d79a2),
	.w5(32'hb9c909c5),
	.w6(32'h39b50a41),
	.w7(32'h3899cf4c),
	.w8(32'h391f90c0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e9733),
	.w1(32'h37a88ec6),
	.w2(32'hb8905ff8),
	.w3(32'h3a312ad1),
	.w4(32'h374c89bf),
	.w5(32'hb90d364a),
	.w6(32'h37ae74c8),
	.w7(32'h3a9cb62a),
	.w8(32'h3a96c4be),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981a921),
	.w1(32'hb96ce5e8),
	.w2(32'hb8c66008),
	.w3(32'hb9ddc822),
	.w4(32'hb9f1b276),
	.w5(32'hb9508f36),
	.w6(32'hb8591165),
	.w7(32'hb8741cd1),
	.w8(32'h38c40086),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d3804),
	.w1(32'h3ab9afca),
	.w2(32'h3ac1983d),
	.w3(32'hba4c5d6e),
	.w4(32'h39ca1b0a),
	.w5(32'h3ae3c176),
	.w6(32'hba9dc575),
	.w7(32'hba1f6bd6),
	.w8(32'hba30ef31),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac84be2),
	.w1(32'h397a59eb),
	.w2(32'hba908aa1),
	.w3(32'hbac09e38),
	.w4(32'hb9ff3e21),
	.w5(32'hb98ecb16),
	.w6(32'hbb1a7d6a),
	.w7(32'hbb9610d9),
	.w8(32'hbb9c6b40),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b012853),
	.w1(32'hba2125df),
	.w2(32'hba3f02b3),
	.w3(32'h3a90abc8),
	.w4(32'hb9eeccd1),
	.w5(32'hba7dce7e),
	.w6(32'h3b4ac3d0),
	.w7(32'h3b128389),
	.w8(32'h3ad54dec),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db8af),
	.w1(32'hba46d419),
	.w2(32'hb9b31e75),
	.w3(32'hbb305601),
	.w4(32'h3ac5996e),
	.w5(32'h39b62e17),
	.w6(32'hbb29f2e0),
	.w7(32'hb889c5f8),
	.w8(32'hbaf55117),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef0086),
	.w1(32'hba39da33),
	.w2(32'hba38b4ac),
	.w3(32'hb9e772cc),
	.w4(32'hbb156d7a),
	.w5(32'hbb47dcb4),
	.w6(32'hba08a846),
	.w7(32'hbac80b51),
	.w8(32'hbadd3d8a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb547cfe),
	.w1(32'hbae413fe),
	.w2(32'hb8ab2a00),
	.w3(32'hbb118c4f),
	.w4(32'h3a910765),
	.w5(32'h3b4946cd),
	.w6(32'hbb1a9c36),
	.w7(32'hbac7cef4),
	.w8(32'h3ac8c903),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad66d93),
	.w1(32'hbabe8771),
	.w2(32'hba53703f),
	.w3(32'hba78d2b7),
	.w4(32'hba2b64b4),
	.w5(32'hba6eb1ae),
	.w6(32'hba0b21d8),
	.w7(32'hba3d7a8a),
	.w8(32'h3a1887ce),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8a440),
	.w1(32'hba71ae6a),
	.w2(32'hba71bd4c),
	.w3(32'hb9f39f97),
	.w4(32'hb98e0097),
	.w5(32'hbab65477),
	.w6(32'h39fa61e3),
	.w7(32'h3a8845f9),
	.w8(32'h3aaaf7e6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3804f812),
	.w1(32'h38d371a6),
	.w2(32'hb88aa9ba),
	.w3(32'h392e8fc5),
	.w4(32'h399cad93),
	.w5(32'h3930e919),
	.w6(32'h398ba27c),
	.w7(32'h3985e9f9),
	.w8(32'h3909b1bb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a871cd7),
	.w1(32'h3adf4524),
	.w2(32'h3b1b8b09),
	.w3(32'hba2a1e31),
	.w4(32'h3a71dee2),
	.w5(32'h3a52cefe),
	.w6(32'hbb1ad0e1),
	.w7(32'hbb6a87b1),
	.w8(32'hbb2523b5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2425),
	.w1(32'h3a7a4d99),
	.w2(32'hb99c7e07),
	.w3(32'h3a9bce80),
	.w4(32'h3adc5ac0),
	.w5(32'hb8f0e94a),
	.w6(32'hba3044ca),
	.w7(32'h38acc468),
	.w8(32'hbabc22ea),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ba316),
	.w1(32'h3a746d3b),
	.w2(32'h3b1b5dd4),
	.w3(32'hbbe33ed2),
	.w4(32'hbb03a0d1),
	.w5(32'h3b865042),
	.w6(32'hbc0e83d4),
	.w7(32'hbb683806),
	.w8(32'hbc4c3c6e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f9ef3),
	.w1(32'hbb2fbe72),
	.w2(32'hb9392f3e),
	.w3(32'hba6cd70d),
	.w4(32'hba95109a),
	.w5(32'hb86d576a),
	.w6(32'h3ae3b04c),
	.w7(32'h3b8f5764),
	.w8(32'h3bb1140f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e0626),
	.w1(32'h3aed15ef),
	.w2(32'h3afa7132),
	.w3(32'hba35f916),
	.w4(32'hba8841d8),
	.w5(32'hbab81529),
	.w6(32'hbb54e8bd),
	.w7(32'hbb273f9e),
	.w8(32'hba661a92),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cdea1),
	.w1(32'h39808e34),
	.w2(32'hba0a7a08),
	.w3(32'hbb1a1946),
	.w4(32'h3a98b12d),
	.w5(32'h3a02f384),
	.w6(32'hbb41ccd6),
	.w7(32'hb9879363),
	.w8(32'hbb910e79),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38af8424),
	.w1(32'h39480bea),
	.w2(32'hb826fe49),
	.w3(32'h3913270c),
	.w4(32'h39c60d15),
	.w5(32'h3970266f),
	.w6(32'h3974df0e),
	.w7(32'h399a9773),
	.w8(32'h38ed61e4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb948d02),
	.w1(32'h3b35b287),
	.w2(32'h386fcdcb),
	.w3(32'hbbda896d),
	.w4(32'hbb2b5313),
	.w5(32'h3b85f984),
	.w6(32'hbc273a02),
	.w7(32'hbac040f3),
	.w8(32'hbc6f5a40),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c23c3d),
	.w1(32'hba03655c),
	.w2(32'hbb0ed4ff),
	.w3(32'hba28f602),
	.w4(32'h38f0bc14),
	.w5(32'hbb26776b),
	.w6(32'hba9927c2),
	.w7(32'h3a39618b),
	.w8(32'hbac1ef43),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d6e8e3),
	.w1(32'hb900b3d3),
	.w2(32'hb8dbe25b),
	.w3(32'hb7872792),
	.w4(32'hb8a46c56),
	.w5(32'hb8a20f37),
	.w6(32'h390191a7),
	.w7(32'h380209bf),
	.w8(32'h388720a2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2f030),
	.w1(32'hba656e43),
	.w2(32'hba14fff8),
	.w3(32'hba39ad33),
	.w4(32'hb9a4f529),
	.w5(32'hba280932),
	.w6(32'hba58cb09),
	.w7(32'hba336688),
	.w8(32'hba1dcbf8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb813ce0b),
	.w1(32'h3aa8420a),
	.w2(32'h3ab5f40c),
	.w3(32'hbae23d6d),
	.w4(32'h395a0de1),
	.w5(32'h39aa789f),
	.w6(32'hbb2e5822),
	.w7(32'hbb269552),
	.w8(32'hbaa08b28),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34afcd),
	.w1(32'h3a8514c4),
	.w2(32'h3a39e984),
	.w3(32'h391330cf),
	.w4(32'hb7446980),
	.w5(32'hba3d397b),
	.w6(32'hb8f82703),
	.w7(32'hb9715711),
	.w8(32'h39759eb5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9e49f),
	.w1(32'hbaf1d1fa),
	.w2(32'hba259b07),
	.w3(32'h3a97963d),
	.w4(32'hbb29701e),
	.w5(32'hbac9e0d2),
	.w6(32'h3adcfcd0),
	.w7(32'hba984e61),
	.w8(32'hb8f8b226),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6473c),
	.w1(32'h3a899096),
	.w2(32'h397a6516),
	.w3(32'h3a779662),
	.w4(32'h38fc9203),
	.w5(32'hb9806373),
	.w6(32'h39597173),
	.w7(32'hba26120c),
	.w8(32'hba29e3eb),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d2ee1),
	.w1(32'h38c47fbc),
	.w2(32'h3ae4ed67),
	.w3(32'hba27fd6d),
	.w4(32'h3a01d820),
	.w5(32'h3b1eabdf),
	.w6(32'hbb1e76fd),
	.w7(32'hbafc41a7),
	.w8(32'hbaadc8be),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4897e1),
	.w1(32'hbb0fe5fd),
	.w2(32'h39e92509),
	.w3(32'hbade27a9),
	.w4(32'hb70f61d4),
	.w5(32'h3b4138c3),
	.w6(32'hbaae0322),
	.w7(32'hba82d8d0),
	.w8(32'h3aedad4f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392664e8),
	.w1(32'h3a816e5b),
	.w2(32'h3a953455),
	.w3(32'h3991007d),
	.w4(32'h38b81692),
	.w5(32'hb923951d),
	.w6(32'hba6af94f),
	.w7(32'hba65cfa4),
	.w8(32'hb931c5f9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86a8697),
	.w1(32'hb881e9f4),
	.w2(32'hb794a07a),
	.w3(32'hb8309473),
	.w4(32'hb5261048),
	.w5(32'h372c37a4),
	.w6(32'hb82e4a57),
	.w7(32'hb760549e),
	.w8(32'hb19f64fa),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f619ce),
	.w1(32'hb89cb739),
	.w2(32'hb7922d89),
	.w3(32'hb85f624f),
	.w4(32'h396a624a),
	.w5(32'h399e6f76),
	.w6(32'hb85185b3),
	.w7(32'h38d5a2b2),
	.w8(32'h38827bee),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b60f8b),
	.w1(32'h385d19b3),
	.w2(32'h37f5d7b8),
	.w3(32'hb85e8e8f),
	.w4(32'hb818ea9f),
	.w5(32'hb8151c76),
	.w6(32'hb819097e),
	.w7(32'hb84bdca2),
	.w8(32'hb878263c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38510b14),
	.w1(32'h382a371c),
	.w2(32'hb78254a2),
	.w3(32'hb64a0793),
	.w4(32'h382fba5f),
	.w5(32'h375f9a41),
	.w6(32'h381843fe),
	.w7(32'h3770f514),
	.w8(32'h38702380),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938c104),
	.w1(32'h3a981c86),
	.w2(32'h3a9c3475),
	.w3(32'h3a492c5a),
	.w4(32'h39b63371),
	.w5(32'h3926e90c),
	.w6(32'hb9caaf33),
	.w7(32'hb9d0e64d),
	.w8(32'h399ad5ed),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38984d37),
	.w1(32'hb6a4a494),
	.w2(32'h38d7ea2f),
	.w3(32'h38dc10ea),
	.w4(32'h385c8efd),
	.w5(32'h38e04792),
	.w6(32'hb9518aaa),
	.w7(32'hb9565e4d),
	.w8(32'h37d30e72),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e30c08),
	.w1(32'h3a33bb12),
	.w2(32'hb8fca04d),
	.w3(32'hbaee5e4a),
	.w4(32'h39d412ea),
	.w5(32'hbaafc774),
	.w6(32'hbb258e42),
	.w7(32'hbaafa728),
	.w8(32'hbb190782),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961158e),
	.w1(32'hba41e3a7),
	.w2(32'hba1122d9),
	.w3(32'hb8ecce28),
	.w4(32'hbae31381),
	.w5(32'hbad92579),
	.w6(32'hb8950552),
	.w7(32'hba7b3d35),
	.w8(32'h38d0166b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8909163),
	.w1(32'hb8e1e569),
	.w2(32'hb89f0ff9),
	.w3(32'hb835cfed),
	.w4(32'hb88536b3),
	.w5(32'hb80d4059),
	.w6(32'hb80a531e),
	.w7(32'hb87824ac),
	.w8(32'hb777c4c6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d7e3b8),
	.w1(32'hb91389c3),
	.w2(32'hb9183499),
	.w3(32'hb915fccd),
	.w4(32'hb8d9f93c),
	.w5(32'hb897f1ba),
	.w6(32'hb896b49d),
	.w7(32'hb78ab8b3),
	.w8(32'hb885fade),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74188d5),
	.w1(32'hb74b3d00),
	.w2(32'hb72ea844),
	.w3(32'hb50b0b12),
	.w4(32'hb6930874),
	.w5(32'hb6e1c366),
	.w6(32'h35378368),
	.w7(32'h36467fc5),
	.w8(32'h36ab8140),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886c1a8),
	.w1(32'h3966bf18),
	.w2(32'h39521909),
	.w3(32'hb9e88313),
	.w4(32'hb8d72bea),
	.w5(32'h38057e7c),
	.w6(32'hba2e7f1d),
	.w7(32'hba00b58e),
	.w8(32'hb9a1da87),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bb7de),
	.w1(32'h39c0681e),
	.w2(32'hba09aff5),
	.w3(32'h3a99fdfe),
	.w4(32'h3b2c37a9),
	.w5(32'hb877832a),
	.w6(32'hbb555991),
	.w7(32'hbb98e504),
	.w8(32'hbb6f59d5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982c13e),
	.w1(32'hb8c54b3a),
	.w2(32'h3a5199c9),
	.w3(32'hba6e153d),
	.w4(32'h3ad097dc),
	.w5(32'h3a906c80),
	.w6(32'hbb21e817),
	.w7(32'hbb162a05),
	.w8(32'hb9670d25),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916638c),
	.w1(32'hb95de1af),
	.w2(32'hb937c0be),
	.w3(32'hb934f03f),
	.w4(32'h392ef678),
	.w5(32'h39644048),
	.w6(32'hb9974be1),
	.w7(32'hb8e9d8eb),
	.w8(32'hb9ba9a80),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9acc3e),
	.w1(32'hb9d9a048),
	.w2(32'hb96e28b7),
	.w3(32'hb9c8b227),
	.w4(32'hba90e1ad),
	.w5(32'hb9f5dd29),
	.w6(32'hba2a50f6),
	.w7(32'hba6abe11),
	.w8(32'hba281a22),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d437bf),
	.w1(32'h38f1af06),
	.w2(32'h38691f43),
	.w3(32'hb88b863f),
	.w4(32'hb9d1e1c2),
	.w5(32'hb9a9ad05),
	.w6(32'hb89ee511),
	.w7(32'hb981a3a8),
	.w8(32'hb9d24868),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3891362d),
	.w1(32'h388feeaf),
	.w2(32'h3a3229a2),
	.w3(32'hb8417cd0),
	.w4(32'h39eeeac1),
	.w5(32'h3a838865),
	.w6(32'hb9c9c028),
	.w7(32'hba16a0ce),
	.w8(32'hb8ca8ec9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2eaa7),
	.w1(32'hbb0e46ec),
	.w2(32'hba0adedc),
	.w3(32'h389502c0),
	.w4(32'hba108963),
	.w5(32'h3a1c0ed3),
	.w6(32'h39dd0988),
	.w7(32'hb989357e),
	.w8(32'h3b04d6c5),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3486a1),
	.w1(32'h39c0c85b),
	.w2(32'hb9f92ba8),
	.w3(32'hbaf39f89),
	.w4(32'h3ac99c49),
	.w5(32'h3a487b1e),
	.w6(32'hbb5d6751),
	.w7(32'hbb8c27b9),
	.w8(32'hbb9c7ab4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39861f83),
	.w1(32'hb7e2a562),
	.w2(32'hb796898e),
	.w3(32'hb913ee53),
	.w4(32'hba4d10b2),
	.w5(32'hb9f0f1dc),
	.w6(32'hb90b096a),
	.w7(32'h39be8b5e),
	.w8(32'h3a388404),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8902018),
	.w1(32'h36c8225a),
	.w2(32'h3aa7bda9),
	.w3(32'hba581468),
	.w4(32'h3a0b9b21),
	.w5(32'hb8c7bfbe),
	.w6(32'hbad0244e),
	.w7(32'hbace0c36),
	.w8(32'hbae3d073),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ba9e6),
	.w1(32'hb9d68a8e),
	.w2(32'hb9b4f061),
	.w3(32'hb92c9c09),
	.w4(32'h39d392c5),
	.w5(32'hb96a81c8),
	.w6(32'hbae8129a),
	.w7(32'hbb83dc7d),
	.w8(32'hbbd190c6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3db6a),
	.w1(32'h39fe41f1),
	.w2(32'h3adea304),
	.w3(32'hba3aa1bb),
	.w4(32'h38abef10),
	.w5(32'h3a9eb356),
	.w6(32'hbaae194d),
	.w7(32'hb9201207),
	.w8(32'h39c309e2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bdae9),
	.w1(32'hb9d35bca),
	.w2(32'h393e5b6d),
	.w3(32'hba483b35),
	.w4(32'h3a100f8f),
	.w5(32'h3a734927),
	.w6(32'hba75c7ce),
	.w7(32'hb9039b06),
	.w8(32'h392ea8bc),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae2afd),
	.w1(32'h39f715ab),
	.w2(32'h3a242dc8),
	.w3(32'hb8988e9f),
	.w4(32'h38155155),
	.w5(32'h39783be3),
	.w6(32'hb9acfa23),
	.w7(32'hb99d5f38),
	.w8(32'hb8eff56c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb8259),
	.w1(32'hba953665),
	.w2(32'hba11357a),
	.w3(32'h39e954c6),
	.w4(32'hba5e6de3),
	.w5(32'hba874e39),
	.w6(32'h3b34bbb9),
	.w7(32'h3a606d74),
	.w8(32'h3a9ce129),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1b3b9),
	.w1(32'h3a2448ac),
	.w2(32'h3a48f4c7),
	.w3(32'h388e5400),
	.w4(32'h391abe24),
	.w5(32'h3995bb61),
	.w6(32'hba3302d1),
	.w7(32'hba347894),
	.w8(32'hb998f04a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9053d7b),
	.w1(32'hb83886c4),
	.w2(32'h35af0c7a),
	.w3(32'hb80bff52),
	.w4(32'hb6138e6e),
	.w5(32'h3755af48),
	.w6(32'h389dd699),
	.w7(32'h38b813a6),
	.w8(32'h387e0f6b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ea3342),
	.w1(32'hb83034a7),
	.w2(32'hb789b037),
	.w3(32'hb704507b),
	.w4(32'hb843b623),
	.w5(32'hb88ac1f2),
	.w6(32'hb79af94f),
	.w7(32'h36fc36e8),
	.w8(32'hb85415f7),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5eb17c),
	.w1(32'hb9f372d0),
	.w2(32'hba2f328a),
	.w3(32'hba1cae36),
	.w4(32'hb8623488),
	.w5(32'hb9bf90d4),
	.w6(32'hba79e38e),
	.w7(32'h380d024c),
	.w8(32'h38961956),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993259c),
	.w1(32'hb9de83e1),
	.w2(32'hba8db3f9),
	.w3(32'h3a12ed4a),
	.w4(32'hb9e6eacf),
	.w5(32'hb8143862),
	.w6(32'hba371173),
	.w7(32'h3aba55d4),
	.w8(32'hb7c75c5c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b238e17),
	.w1(32'h3b699e1c),
	.w2(32'h3b852fac),
	.w3(32'hbaeb2ca3),
	.w4(32'hb9845bae),
	.w5(32'h3ac214cc),
	.w6(32'hbb2c7f03),
	.w7(32'hbb3d69c6),
	.w8(32'hb90d6ac5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a07cd5),
	.w1(32'hb7388559),
	.w2(32'hb7ad0605),
	.w3(32'hb6d5d9bc),
	.w4(32'h36e7d569),
	.w5(32'hb700e943),
	.w6(32'hb6cd01e9),
	.w7(32'hb622e206),
	.w8(32'hb60f7892),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9314dba),
	.w1(32'h391f890f),
	.w2(32'h3a72367d),
	.w3(32'hba259d78),
	.w4(32'h3a994cf0),
	.w5(32'h3a905c08),
	.w6(32'hbb1d0a87),
	.w7(32'hba8dbcb8),
	.w8(32'h3a39ab66),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c4818),
	.w1(32'h3a6e6fee),
	.w2(32'h3a8ef7da),
	.w3(32'hb9953b6d),
	.w4(32'h39db7811),
	.w5(32'h39c4fe20),
	.w6(32'hba714114),
	.w7(32'hba49809b),
	.w8(32'hb7e22137),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2dd97),
	.w1(32'hb908c0ef),
	.w2(32'h3a5675ca),
	.w3(32'hbb6bf60f),
	.w4(32'hb9aa1ca3),
	.w5(32'hb9f06311),
	.w6(32'hbb50b8ae),
	.w7(32'hbaf53afb),
	.w8(32'hbb7505dd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ad9e2),
	.w1(32'h3a598f87),
	.w2(32'hba849041),
	.w3(32'h3b25feaf),
	.w4(32'h3a13dbed),
	.w5(32'hbadebab3),
	.w6(32'h3b4155da),
	.w7(32'h3a4d9075),
	.w8(32'h3af6fb3d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a6240),
	.w1(32'hba3a57cb),
	.w2(32'hba44ed7c),
	.w3(32'h3a01cf75),
	.w4(32'hb9e6aaee),
	.w5(32'hba2c6324),
	.w6(32'h3a2b7d31),
	.w7(32'h38f37f57),
	.w8(32'hb79f433b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3846454e),
	.w1(32'h3783f6ed),
	.w2(32'hb9025308),
	.w3(32'h394c235b),
	.w4(32'h3917b86f),
	.w5(32'h39892321),
	.w6(32'h39daad5d),
	.w7(32'h39b77294),
	.w8(32'h39d36be1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952ae8a),
	.w1(32'h3aa02a51),
	.w2(32'h3abcd314),
	.w3(32'h3a91c71f),
	.w4(32'h3a84b05c),
	.w5(32'h3a1189b7),
	.w6(32'h3aa724b8),
	.w7(32'h3acbb42a),
	.w8(32'h3ae03fed),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39502dfc),
	.w1(32'hb9ef6745),
	.w2(32'h3933395f),
	.w3(32'h3a67ae9f),
	.w4(32'hb9063d80),
	.w5(32'h3a163902),
	.w6(32'h3a27b415),
	.w7(32'h3a6d4a39),
	.w8(32'h3ae4b8b2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9443e3b),
	.w1(32'hba91992c),
	.w2(32'hba3c6c0a),
	.w3(32'hb8067a1a),
	.w4(32'hba84deda),
	.w5(32'hba284e5c),
	.w6(32'h399b951b),
	.w7(32'h3a068983),
	.w8(32'h3a3a5a1c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905c72c),
	.w1(32'hb80338e2),
	.w2(32'hb8817bb9),
	.w3(32'hb8653650),
	.w4(32'h388550e9),
	.w5(32'h391d5ad5),
	.w6(32'hb9f74339),
	.w7(32'hb9dad84b),
	.w8(32'hbaad9177),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c799a2),
	.w1(32'hb8c891f8),
	.w2(32'hb92b1c3a),
	.w3(32'hb8e75c59),
	.w4(32'hb843da3a),
	.w5(32'hb90eb7f5),
	.w6(32'h382647b8),
	.w7(32'hb97a99b5),
	.w8(32'hb9bf05df),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f7a2f),
	.w1(32'h39fa5731),
	.w2(32'h394924ff),
	.w3(32'hba4cd657),
	.w4(32'h3a3e31db),
	.w5(32'h3a099955),
	.w6(32'hbaaf436a),
	.w7(32'hbaf94daa),
	.w8(32'hbb227621),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21b322),
	.w1(32'h3966bdd3),
	.w2(32'hba15ebc4),
	.w3(32'h39a3e525),
	.w4(32'h3843523b),
	.w5(32'hb98de6e9),
	.w6(32'h398f184b),
	.w7(32'h3a1840d9),
	.w8(32'h3a13c0b4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995a7d4),
	.w1(32'h3946ab3e),
	.w2(32'h39830163),
	.w3(32'h3a7ce98f),
	.w4(32'h3a2b3f22),
	.w5(32'hb94334ee),
	.w6(32'hb7cd12fb),
	.w7(32'hba7b4aa0),
	.w8(32'h39178b00),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80cd927),
	.w1(32'hb8c0889a),
	.w2(32'hb8a12c57),
	.w3(32'hb8c190c8),
	.w4(32'hb9308d93),
	.w5(32'hb91da6bb),
	.w6(32'hb889981b),
	.w7(32'hb83bb7dd),
	.w8(32'hb7f1f190),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3232a),
	.w1(32'hb9e9e629),
	.w2(32'hbb01eb98),
	.w3(32'hb789e3ee),
	.w4(32'hba43f317),
	.w5(32'hbb27c730),
	.w6(32'hb97260f5),
	.w7(32'hbb1ee815),
	.w8(32'hbb54c0cd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35234ff2),
	.w1(32'h38188ddd),
	.w2(32'h388ed4ea),
	.w3(32'h37e9ccb1),
	.w4(32'h38a13922),
	.w5(32'h38b3a876),
	.w6(32'h382a1417),
	.w7(32'h388baed9),
	.w8(32'h38883351),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bb5a69),
	.w1(32'h388080d9),
	.w2(32'hb8402f63),
	.w3(32'h3913ae08),
	.w4(32'h38da9357),
	.w5(32'hb8cb1b7f),
	.w6(32'hb8893810),
	.w7(32'hb957eade),
	.w8(32'hb98fd330),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80771e),
	.w1(32'hba4bbac2),
	.w2(32'hb99e3c83),
	.w3(32'hb918db7a),
	.w4(32'hb94ae347),
	.w5(32'h38a245e7),
	.w6(32'h3973223d),
	.w7(32'h3a2828ce),
	.w8(32'h3accf3f6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2772a5),
	.w1(32'h3b1814af),
	.w2(32'h3ad5dcd1),
	.w3(32'hbab5cd94),
	.w4(32'h3aa6251d),
	.w5(32'h3a81fc85),
	.w6(32'hbb52e854),
	.w7(32'hbaa532c3),
	.w8(32'hbb21dba7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a528f3),
	.w1(32'hb8f9e52a),
	.w2(32'hb793a33e),
	.w3(32'hb6372dbb),
	.w4(32'hba4b5c37),
	.w5(32'hba1d72d9),
	.w6(32'h39ef79c7),
	.w7(32'h379da66e),
	.w8(32'hb84ecb27),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24e191),
	.w1(32'h3a75bb5b),
	.w2(32'h3a82c617),
	.w3(32'hb9f41d00),
	.w4(32'hb986e93c),
	.w5(32'hb8ca43ef),
	.w6(32'hb9e06c53),
	.w7(32'hba1f01ff),
	.w8(32'h39e90d0b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d1c74),
	.w1(32'hb84c3ea9),
	.w2(32'hb94b4a86),
	.w3(32'h3939b032),
	.w4(32'h39762f2e),
	.w5(32'hb90dbad0),
	.w6(32'h3a7b3182),
	.w7(32'h3a8669ab),
	.w8(32'h3ac48bce),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a139a32),
	.w1(32'h3a943069),
	.w2(32'h3b1e117b),
	.w3(32'hba26f70a),
	.w4(32'h3af902e6),
	.w5(32'hba01f877),
	.w6(32'hbab8c269),
	.w7(32'hbaa6c305),
	.w8(32'hb87cfae8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ff536),
	.w1(32'hb9ce488e),
	.w2(32'h39685b81),
	.w3(32'hba8812b8),
	.w4(32'h399a1200),
	.w5(32'h3aaca62b),
	.w6(32'hba942a07),
	.w7(32'h38407f09),
	.w8(32'h39fd61b1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a871324),
	.w1(32'h3aa8c35c),
	.w2(32'h3ad9436f),
	.w3(32'hb98f6b0b),
	.w4(32'h3ace4236),
	.w5(32'h3a5f4602),
	.w6(32'hbaf5a517),
	.w7(32'hbb1e5361),
	.w8(32'hbac66f80),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a4b0e9),
	.w1(32'hb7d794f5),
	.w2(32'h383782a3),
	.w3(32'h38ba99e0),
	.w4(32'h38be3615),
	.w5(32'h3905ddb1),
	.w6(32'h3909c6bc),
	.w7(32'h391d27b1),
	.w8(32'h391d4c95),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c41918),
	.w1(32'hba15db38),
	.w2(32'h39f9c414),
	.w3(32'hba05ca86),
	.w4(32'h3a0b3f34),
	.w5(32'h3a716277),
	.w6(32'hb8487f96),
	.w7(32'h38d557c3),
	.w8(32'h39905c17),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a51f27),
	.w1(32'hb742a1cc),
	.w2(32'hb79d0f9e),
	.w3(32'hb6c8f9e6),
	.w4(32'hb765e87a),
	.w5(32'hb756d777),
	.w6(32'hb539c0c4),
	.w7(32'hb6d611b8),
	.w8(32'hb6d0d59c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc0faa),
	.w1(32'h396fe10f),
	.w2(32'h3a089017),
	.w3(32'hb93776f4),
	.w4(32'hb8aafb1f),
	.w5(32'hb97ea1f2),
	.w6(32'hba40bfa8),
	.w7(32'hba0f79c6),
	.w8(32'hb9c6f867),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373216bb),
	.w1(32'hb98a384e),
	.w2(32'hb9dfebb7),
	.w3(32'h38b98660),
	.w4(32'hba2ae92c),
	.w5(32'hba1fb050),
	.w6(32'hb9862fa7),
	.w7(32'hb963ed53),
	.w8(32'hb9b3857b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad466f5),
	.w1(32'hbaaa1401),
	.w2(32'hb7cb4b56),
	.w3(32'hbaf4871d),
	.w4(32'hb93b0460),
	.w5(32'h3a28b99a),
	.w6(32'hbb0b5fe0),
	.w7(32'hbadecfbf),
	.w8(32'hb9676650),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d299f3),
	.w1(32'hb5944668),
	.w2(32'hb5a0e05f),
	.w3(32'hb6a534ec),
	.w4(32'hb5e5c8d1),
	.w5(32'h35e6351e),
	.w6(32'hb616f20f),
	.w7(32'h35c9a5b9),
	.w8(32'hb67362e3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379416d0),
	.w1(32'h371899ed),
	.w2(32'h377516c7),
	.w3(32'h374c758a),
	.w4(32'h379d2da4),
	.w5(32'h38000f50),
	.w6(32'h383e6a06),
	.w7(32'h38172427),
	.w8(32'h37245720),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f10f4),
	.w1(32'h3a08b2aa),
	.w2(32'hb7a45b46),
	.w3(32'h3a883fa8),
	.w4(32'h39c370d3),
	.w5(32'hbaf299df),
	.w6(32'hba2f2696),
	.w7(32'hbadccbb2),
	.w8(32'hba63be0d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3950f489),
	.w1(32'hba59d1ae),
	.w2(32'hba2d0418),
	.w3(32'h39e38963),
	.w4(32'h3a48d821),
	.w5(32'hbacfb6b3),
	.w6(32'hb7b22ac8),
	.w7(32'hb9fdfd87),
	.w8(32'hbb0ba23f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad616cc),
	.w1(32'hba1113f9),
	.w2(32'hba2f8d4a),
	.w3(32'hbb622640),
	.w4(32'hba113508),
	.w5(32'h3ad7985a),
	.w6(32'hbb89bb98),
	.w7(32'hba6019a1),
	.w8(32'hbb8bcc27),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb892a153),
	.w1(32'hb989e4c9),
	.w2(32'hb94639b5),
	.w3(32'hb92c802c),
	.w4(32'hb9098f1c),
	.w5(32'hb92d24d5),
	.w6(32'hb9889db6),
	.w7(32'hb9750a71),
	.w8(32'hb8cfc2a3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c33d4),
	.w1(32'h3b6baa68),
	.w2(32'h3be7d738),
	.w3(32'h3a8e066d),
	.w4(32'h3bc62685),
	.w5(32'h3b92f417),
	.w6(32'hb9befdb5),
	.w7(32'hbae8827a),
	.w8(32'h3b88566a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b350cf),
	.w1(32'hbb26c208),
	.w2(32'hbace6bb2),
	.w3(32'h3ad779cf),
	.w4(32'h3a821199),
	.w5(32'hb9b4150c),
	.w6(32'hb914ff18),
	.w7(32'h3a8c78d3),
	.w8(32'h3bb83615),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39902d11),
	.w1(32'hb9772e9b),
	.w2(32'hba941c72),
	.w3(32'hb9268ac0),
	.w4(32'h36ac1a80),
	.w5(32'hba02e208),
	.w6(32'hba06d188),
	.w7(32'hba1aec16),
	.w8(32'hba0b4f11),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b23e9),
	.w1(32'hb6927b4f),
	.w2(32'hb79c652b),
	.w3(32'hb81f3cd0),
	.w4(32'hb80e15cc),
	.w5(32'hb5cc5953),
	.w6(32'hb7ce9b44),
	.w7(32'hb7d9aa81),
	.w8(32'hb7d0154c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e70d0),
	.w1(32'hb5bda153),
	.w2(32'hb7e2f644),
	.w3(32'h381157e2),
	.w4(32'h385af3b1),
	.w5(32'h381afdb2),
	.w6(32'h383a4d0b),
	.w7(32'h38956f39),
	.w8(32'h38034364),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d7769d),
	.w1(32'hb721b220),
	.w2(32'hb776559b),
	.w3(32'h338b73cd),
	.w4(32'h35555fe0),
	.w5(32'hb6518c1f),
	.w6(32'h35794aa1),
	.w7(32'hb5bb1022),
	.w8(32'hb528cfac),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c5604),
	.w1(32'hb9817010),
	.w2(32'hbadbbc64),
	.w3(32'hba8ebc4b),
	.w4(32'h39a458bd),
	.w5(32'hbab1819c),
	.w6(32'hbabd81eb),
	.w7(32'hbaee2cf5),
	.w8(32'hbb2812ab),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ee5b1),
	.w1(32'h3aa2e20e),
	.w2(32'h3a2821f8),
	.w3(32'hb9f9fa3a),
	.w4(32'h33481818),
	.w5(32'hba397f88),
	.w6(32'hbadb6349),
	.w7(32'hba96048d),
	.w8(32'hbadf9a07),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb1390),
	.w1(32'h3a79c034),
	.w2(32'h3af3813a),
	.w3(32'hba9da410),
	.w4(32'hba87c23d),
	.w5(32'h39b1974b),
	.w6(32'hba6c26d6),
	.w7(32'hba4a908c),
	.w8(32'h3a62432a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9229a19),
	.w1(32'h39457bf6),
	.w2(32'h39b5622f),
	.w3(32'hb929bd12),
	.w4(32'hb99e9e63),
	.w5(32'hb94ed072),
	.w6(32'hb97c85ff),
	.w7(32'hb9fc1971),
	.w8(32'hb9abd27e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb840c405),
	.w1(32'h3a9f317f),
	.w2(32'h3b21feae),
	.w3(32'hba81c3f2),
	.w4(32'h3acd3582),
	.w5(32'h3abeaea0),
	.w6(32'hbb20108a),
	.w7(32'hbadacfeb),
	.w8(32'hbab40fb6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b543c),
	.w1(32'h3a9657f2),
	.w2(32'h3964751c),
	.w3(32'h3916940f),
	.w4(32'h39973cfe),
	.w5(32'hb9a43ad8),
	.w6(32'hb9fce4ec),
	.w7(32'h39377bef),
	.w8(32'hba9de395),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78df295),
	.w1(32'hb77bcbd3),
	.w2(32'hb74e26cc),
	.w3(32'hb4536112),
	.w4(32'h3640497b),
	.w5(32'h34189626),
	.w6(32'h36d23c3b),
	.w7(32'h37383e6f),
	.w8(32'h3619604e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa967c0),
	.w1(32'hbaddcb2d),
	.w2(32'h39a6b325),
	.w3(32'hbb11fd0e),
	.w4(32'hba57c753),
	.w5(32'h3aa599d0),
	.w6(32'hbb00bd4c),
	.w7(32'hb95cd61c),
	.w8(32'hba8c5950),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82e6fdc),
	.w1(32'hb8496038),
	.w2(32'hb841a347),
	.w3(32'h36690ea9),
	.w4(32'h328b209a),
	.w5(32'hb609b0f8),
	.w6(32'h3788154a),
	.w7(32'h37927bf0),
	.w8(32'h37b99796),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a3173),
	.w1(32'h3a90c90a),
	.w2(32'h3a7da708),
	.w3(32'hb827dd80),
	.w4(32'h39dd0025),
	.w5(32'h385a3d30),
	.w6(32'hba95cae5),
	.w7(32'hbaaf59e4),
	.w8(32'hbab03e0f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cba8da),
	.w1(32'hba903059),
	.w2(32'hba75cd1f),
	.w3(32'h3a21716a),
	.w4(32'hba6254ce),
	.w5(32'hba9a38eb),
	.w6(32'h3964a092),
	.w7(32'hb72177b1),
	.w8(32'h3a3a69f5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e5721),
	.w1(32'h39286a25),
	.w2(32'h3a91a907),
	.w3(32'hb950533b),
	.w4(32'hb9a1f955),
	.w5(32'h39b6cb13),
	.w6(32'hb915c0b1),
	.w7(32'hb979c4c2),
	.w8(32'h3a07adf3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39533dc3),
	.w1(32'hb8cf19ef),
	.w2(32'hb82576c7),
	.w3(32'h398793d1),
	.w4(32'hb89a0aa1),
	.w5(32'hb8c75a2a),
	.w6(32'h39ec56a5),
	.w7(32'h39b0ba92),
	.w8(32'h394fc5e1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea79e0),
	.w1(32'hb955e5b3),
	.w2(32'h3a5a42e3),
	.w3(32'hb9d0a6c0),
	.w4(32'hb9ed9b7b),
	.w5(32'h3a31b9c0),
	.w6(32'hba193bd5),
	.w7(32'hb9cc8afd),
	.w8(32'h3a9b74df),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e1119),
	.w1(32'hb97b6089),
	.w2(32'h3a244231),
	.w3(32'hbaa7dcbc),
	.w4(32'h39b4750b),
	.w5(32'h3a76d849),
	.w6(32'hbad51155),
	.w7(32'hba995e97),
	.w8(32'h382133e0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b028a73),
	.w1(32'h3b3c04a9),
	.w2(32'h3b39b12d),
	.w3(32'hbad1e96b),
	.w4(32'h3a0e4f32),
	.w5(32'h3a1bf026),
	.w6(32'hbad8862e),
	.w7(32'hbb29725d),
	.w8(32'hba7e247f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79d01d9),
	.w1(32'hb6ea606a),
	.w2(32'hb7cd3d64),
	.w3(32'h360c95c9),
	.w4(32'h36ca27f9),
	.w5(32'hb7a87d8a),
	.w6(32'h379042ee),
	.w7(32'h37633770),
	.w8(32'hb8063f46),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d20fd2),
	.w1(32'hb7f289c5),
	.w2(32'hb8eba5e7),
	.w3(32'h379dd215),
	.w4(32'hb8604b83),
	.w5(32'hb8f78c46),
	.w6(32'h38de0480),
	.w7(32'hb85ed8c1),
	.w8(32'hb8bb2ac7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30372f),
	.w1(32'h3b139ef5),
	.w2(32'h3a699a41),
	.w3(32'h3a0dcd95),
	.w4(32'h3aa08ed7),
	.w5(32'h3aa8e6a8),
	.w6(32'hb88e3c12),
	.w7(32'hba0f2b4c),
	.w8(32'hba7fdba3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c6613),
	.w1(32'h3b06ceff),
	.w2(32'h3b37d9bb),
	.w3(32'h3a1dd2bb),
	.w4(32'h3acc06de),
	.w5(32'h3a1d1836),
	.w6(32'hbaca2787),
	.w7(32'hba5253ca),
	.w8(32'hba7a95fa),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba973461),
	.w1(32'h3ac60cbc),
	.w2(32'h3b10cdb6),
	.w3(32'h3a1087c4),
	.w4(32'hb88c14a0),
	.w5(32'hba248d3d),
	.w6(32'hbb19cc4f),
	.w7(32'hbade7d49),
	.w8(32'hb7cd5175),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394406d6),
	.w1(32'hba833fce),
	.w2(32'hbb17904c),
	.w3(32'hba0a95a4),
	.w4(32'h3a0518b1),
	.w5(32'hb98b767e),
	.w6(32'h3af2c1b7),
	.w7(32'h3ae7c47e),
	.w8(32'h3a1cccce),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8d2ac),
	.w1(32'hb9d1fea6),
	.w2(32'hb7a57ed9),
	.w3(32'hb94e537e),
	.w4(32'hb9655388),
	.w5(32'h38d120fb),
	.w6(32'hb9a692ea),
	.w7(32'hb9443e71),
	.w8(32'h393e6cd9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ac7c8),
	.w1(32'hb9b4707e),
	.w2(32'h389d338b),
	.w3(32'hb926ad81),
	.w4(32'hb92b2b72),
	.w5(32'h3a6b50db),
	.w6(32'hb9c3b4d7),
	.w7(32'h39987105),
	.w8(32'h3a286cee),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa16341),
	.w1(32'h3b0bc5f3),
	.w2(32'hbac74f33),
	.w3(32'hbae349e3),
	.w4(32'h3aee131d),
	.w5(32'hb7252a9c),
	.w6(32'hbb5df8fa),
	.w7(32'hb9a9e1f5),
	.w8(32'hbb9ec0cb),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0faf64),
	.w1(32'h3a7c09f4),
	.w2(32'h3aec5487),
	.w3(32'hbaa2a69e),
	.w4(32'h3aa96708),
	.w5(32'hb9c1fc48),
	.w6(32'hbb3a9e34),
	.w7(32'hbba7884c),
	.w8(32'hbb7bcf49),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac915b1),
	.w1(32'h39c95548),
	.w2(32'h39964795),
	.w3(32'hbb8367a5),
	.w4(32'hb9a7ce71),
	.w5(32'h3a4c6d49),
	.w6(32'hbbc56c3b),
	.w7(32'hbb6c7135),
	.w8(32'hbbda58ea),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bad5e8),
	.w1(32'hb9c008e3),
	.w2(32'hb9b873ec),
	.w3(32'hb85d5af3),
	.w4(32'hbad4fd74),
	.w5(32'hbad1e23b),
	.w6(32'h39a70829),
	.w7(32'hb87da115),
	.w8(32'hb90e7554),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39818951),
	.w1(32'hba23c7f6),
	.w2(32'hb916b1c9),
	.w3(32'h3aaac122),
	.w4(32'hb9ee0571),
	.w5(32'hb8903c0d),
	.w6(32'h3b152841),
	.w7(32'h3ae8fb8f),
	.w8(32'h3b42842e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63abe26),
	.w1(32'hb66bbc06),
	.w2(32'hb61396bd),
	.w3(32'h35da9f99),
	.w4(32'hb4a4ce25),
	.w5(32'hb4ebc459),
	.w6(32'h369e0e5a),
	.w7(32'h36cda83f),
	.w8(32'h364a44e5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782e11d),
	.w1(32'hb75580e5),
	.w2(32'hb7422816),
	.w3(32'hb691f9f8),
	.w4(32'h360dcfcd),
	.w5(32'hb4999e27),
	.w6(32'h371b3546),
	.w7(32'h3743baa5),
	.w8(32'h371ebf72),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de36da),
	.w1(32'hb9c22b9b),
	.w2(32'hba1b8b17),
	.w3(32'h3a47a8f9),
	.w4(32'h3a66d45d),
	.w5(32'hb913e05c),
	.w6(32'hb9e01b33),
	.w7(32'hba8f4b11),
	.w8(32'hba9bdd09),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7796119),
	.w1(32'hb7453bd3),
	.w2(32'hb7237853),
	.w3(32'hb6dbf7b8),
	.w4(32'h34f9d9ba),
	.w5(32'h34ef757c),
	.w6(32'hb5e01af8),
	.w7(32'h362cd3a0),
	.w8(32'h369303a7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43bd1f),
	.w1(32'hba318712),
	.w2(32'hbaec0c57),
	.w3(32'h3994f8ae),
	.w4(32'hb9d94372),
	.w5(32'hba4c5416),
	.w6(32'hb7c93715),
	.w7(32'hb96b0724),
	.w8(32'hb99b3a37),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0659ab),
	.w1(32'h38b344f0),
	.w2(32'h3b0db6b4),
	.w3(32'h38ae9f72),
	.w4(32'h3a81853e),
	.w5(32'h3a0d4f11),
	.w6(32'hbb26d0f8),
	.w7(32'hbafb5af9),
	.w8(32'hba8eebe3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a359aac),
	.w1(32'h3a489352),
	.w2(32'h3a70806d),
	.w3(32'hba1c1add),
	.w4(32'hba13ef65),
	.w5(32'hb907d177),
	.w6(32'hb9ea2081),
	.w7(32'hba19afdc),
	.w8(32'hb9a4ab9a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7940fd5),
	.w1(32'hb784e161),
	.w2(32'hb6fe46b6),
	.w3(32'hb6271f26),
	.w4(32'h366b093b),
	.w5(32'h36ee3376),
	.w6(32'h365e0b11),
	.w7(32'h36b82a86),
	.w8(32'h37010881),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4f369),
	.w1(32'hb982af41),
	.w2(32'hb7dc43d7),
	.w3(32'hbbd1d132),
	.w4(32'hbaf37720),
	.w5(32'h3ab9d922),
	.w6(32'hbbf1f2b4),
	.w7(32'hbbc8d36d),
	.w8(32'hbc064f74),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39991f7e),
	.w1(32'h398b7c9a),
	.w2(32'h3a101b26),
	.w3(32'hb9dfda56),
	.w4(32'h3a10e782),
	.w5(32'hb931ae2a),
	.w6(32'hbabf1622),
	.w7(32'hbafc9eae),
	.w8(32'hbae261aa),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909a49e),
	.w1(32'hb8edde8b),
	.w2(32'hb8f6745e),
	.w3(32'hb88af949),
	.w4(32'hb84f5b16),
	.w5(32'hb88540ec),
	.w6(32'hb825bb61),
	.w7(32'hb7495a87),
	.w8(32'hb861af40),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c0301),
	.w1(32'h39bd90a1),
	.w2(32'hb7c38a68),
	.w3(32'hba5f6ff6),
	.w4(32'h39b3d1a5),
	.w5(32'h39aa611f),
	.w6(32'hbabf1317),
	.w7(32'hbab62f0d),
	.w8(32'hbb070873),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b15f6d),
	.w1(32'h3776b516),
	.w2(32'h36dc2d40),
	.w3(32'h3829f947),
	.w4(32'h37f37428),
	.w5(32'h37bce309),
	.w6(32'h3848545d),
	.w7(32'h383a53cd),
	.w8(32'h382d3696),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81aa611),
	.w1(32'hb812bcb6),
	.w2(32'h38097977),
	.w3(32'hb8ae5296),
	.w4(32'hb88063d8),
	.w5(32'hb79f2904),
	.w6(32'hb63314aa),
	.w7(32'h383a11a5),
	.w8(32'hb7819890),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3627cb90),
	.w1(32'hb77383f8),
	.w2(32'hb6dd367e),
	.w3(32'h376c715e),
	.w4(32'h37158db9),
	.w5(32'h3766aec8),
	.w6(32'h369eb1de),
	.w7(32'hb6efc04d),
	.w8(32'hb788ba49),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d14c73),
	.w1(32'hb7bf013c),
	.w2(32'hb7f5f91c),
	.w3(32'hb73e2296),
	.w4(32'h36a3869c),
	.w5(32'hb7ccbef7),
	.w6(32'h3794a34a),
	.w7(32'h37c4936b),
	.w8(32'h363cbd0e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa60e4),
	.w1(32'hb9738239),
	.w2(32'h39309389),
	.w3(32'hb8e15d75),
	.w4(32'hb9e8df3f),
	.w5(32'hba0ddfb5),
	.w6(32'h39a3c302),
	.w7(32'h39d5c17f),
	.w8(32'hb8275218),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912fa54),
	.w1(32'hbada2fa9),
	.w2(32'hb99fef23),
	.w3(32'hb8be250e),
	.w4(32'h3add5796),
	.w5(32'h39b0bf16),
	.w6(32'hba229d5b),
	.w7(32'h3a1a9a7a),
	.w8(32'h3aa72baa),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a6ff3),
	.w1(32'h3a548964),
	.w2(32'h3a7ee0b8),
	.w3(32'hb96f88f5),
	.w4(32'h3acccb23),
	.w5(32'h3ab56637),
	.w6(32'hba6b27b7),
	.w7(32'hba8152e5),
	.w8(32'hba5b1a6e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f95356),
	.w1(32'hb91a3b61),
	.w2(32'h38807240),
	.w3(32'hba66017b),
	.w4(32'h3af8f94b),
	.w5(32'h3a42c5fe),
	.w6(32'hbab1c4ca),
	.w7(32'hba9a033b),
	.w8(32'hba2b73d5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e37df3),
	.w1(32'h3805742e),
	.w2(32'h3838e62c),
	.w3(32'h37cb54d4),
	.w4(32'h3776ed39),
	.w5(32'h37b4ab93),
	.w6(32'h384aca86),
	.w7(32'h38274236),
	.w8(32'h381b6ef8),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e2e04),
	.w1(32'h37423cc5),
	.w2(32'hb7af0f74),
	.w3(32'hb7acfe81),
	.w4(32'h39a7bc5b),
	.w5(32'h39daf52f),
	.w6(32'h369ca0dc),
	.w7(32'h38d7d545),
	.w8(32'h394e06cb),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb736cb34),
	.w1(32'hb6f2d0f8),
	.w2(32'hb71d1b7f),
	.w3(32'hb718e66d),
	.w4(32'hb6439528),
	.w5(32'hb696ef03),
	.w6(32'hb6be89bc),
	.w7(32'hb687db16),
	.w8(32'hb6d63fac),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7079f3e),
	.w1(32'hb69ddc34),
	.w2(32'hb6f63328),
	.w3(32'h3707eee2),
	.w4(32'h36002ba0),
	.w5(32'hb6e2aaf5),
	.w6(32'h37236376),
	.w7(32'h372452c8),
	.w8(32'hb642f985),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40ac43),
	.w1(32'hba5afce0),
	.w2(32'h3a7c2fc2),
	.w3(32'h3934bd4e),
	.w4(32'h3a6f7be7),
	.w5(32'h3ab427a6),
	.w6(32'hba01fc43),
	.w7(32'hba7cb117),
	.w8(32'hba03d2c1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88de6c8),
	.w1(32'hb8429af9),
	.w2(32'hb881fd72),
	.w3(32'hb83fb00e),
	.w4(32'hb7644cc9),
	.w5(32'hb83ff680),
	.w6(32'hb841ed0a),
	.w7(32'hb804989c),
	.w8(32'hb87ad548),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381af3bb),
	.w1(32'hb986d8a0),
	.w2(32'hb8be7cfc),
	.w3(32'hb84d2177),
	.w4(32'hba00a87b),
	.w5(32'hb9aa23fd),
	.w6(32'h387b05ed),
	.w7(32'hb911748b),
	.w8(32'hb923f751),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab73353),
	.w1(32'hba63f560),
	.w2(32'h3901a136),
	.w3(32'hb9d9f6ee),
	.w4(32'hb97bd5cb),
	.w5(32'h39ce6e84),
	.w6(32'hb95d8497),
	.w7(32'h39393115),
	.w8(32'h3a739fe1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7728048),
	.w1(32'hb7614de4),
	.w2(32'hb7a0e5fd),
	.w3(32'hb75cc3e5),
	.w4(32'hb47354eb),
	.w5(32'hb79cce4a),
	.w6(32'hb682aa07),
	.w7(32'hb78095b7),
	.w8(32'hb7e66895),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b8afa),
	.w1(32'h39cf16f4),
	.w2(32'h3a4564e2),
	.w3(32'hb91c2649),
	.w4(32'h399796a5),
	.w5(32'h38831193),
	.w6(32'hba3bfe62),
	.w7(32'hbabcb5f2),
	.w8(32'hba3f8fb5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa6192),
	.w1(32'hb9783fd2),
	.w2(32'hb9866eae),
	.w3(32'hb90dc11e),
	.w4(32'hb7a834b4),
	.w5(32'h384b67c2),
	.w6(32'h37b66cf3),
	.w7(32'h39124e75),
	.w8(32'h38689acb),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ad8a),
	.w1(32'hbb9a0966),
	.w2(32'hba88bf3c),
	.w3(32'hba84c6d0),
	.w4(32'h3b0a5dc2),
	.w5(32'h3b011e0e),
	.w6(32'hba8a1bfa),
	.w7(32'hbaf04fe9),
	.w8(32'h3afdc220),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7be0639),
	.w1(32'h3be2f63c),
	.w2(32'hbc1eb9c2),
	.w3(32'h37e649f0),
	.w4(32'h3a997432),
	.w5(32'hbb3ece93),
	.w6(32'h39c701f3),
	.w7(32'hbb4578e9),
	.w8(32'hbc146365),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc500206),
	.w1(32'h3adf014c),
	.w2(32'hbb985258),
	.w3(32'hbbd0371c),
	.w4(32'hbb5cb87f),
	.w5(32'hbb4c5887),
	.w6(32'h37be866c),
	.w7(32'hbaccb3a9),
	.w8(32'h3ba40b8a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule