module layer_8_featuremap_129(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77b4e0),
	.w1(32'hbb7df3e5),
	.w2(32'hbb8e8b00),
	.w3(32'hbbceb2e9),
	.w4(32'h3bcf3e00),
	.w5(32'h3b4bf9f1),
	.w6(32'hbc3ae075),
	.w7(32'hbc1e9ca5),
	.w8(32'hbbd49e14),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddeecd),
	.w1(32'h3c481389),
	.w2(32'hbaef13c2),
	.w3(32'hbb919893),
	.w4(32'h3c707a35),
	.w5(32'h3a969446),
	.w6(32'hbbb828bb),
	.w7(32'h3b564b7e),
	.w8(32'hbc32190b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb674015),
	.w1(32'h3c019be3),
	.w2(32'h3b52abe5),
	.w3(32'hba88873a),
	.w4(32'hba104f02),
	.w5(32'h3c0142ba),
	.w6(32'h3b94f25c),
	.w7(32'h380b4fbd),
	.w8(32'hba7d0f78),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17420a),
	.w1(32'h3b476516),
	.w2(32'h3c54ab23),
	.w3(32'h3bdedede),
	.w4(32'hb9f74c8f),
	.w5(32'h3c2191e3),
	.w6(32'hbafe630a),
	.w7(32'h3d0afd3d),
	.w8(32'h3d024c5b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6465ff),
	.w1(32'hbc9b66f4),
	.w2(32'hbbb916eb),
	.w3(32'hbca90f67),
	.w4(32'hbc6ca589),
	.w5(32'hbc2affb7),
	.w6(32'hbc6a264a),
	.w7(32'h396af941),
	.w8(32'h3c1618b3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6db56c),
	.w1(32'hb9dedd8f),
	.w2(32'h3c1335e0),
	.w3(32'hbc66a6f4),
	.w4(32'h3c4178a5),
	.w5(32'hbc5f738f),
	.w6(32'hbc432421),
	.w7(32'h3c5403ba),
	.w8(32'h3cece245),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae0fad),
	.w1(32'h3ba90587),
	.w2(32'hbcbc250d),
	.w3(32'hbbd7d3f2),
	.w4(32'hbc501d9e),
	.w5(32'h3b88efbf),
	.w6(32'hbc1b0e03),
	.w7(32'hbc8c8b52),
	.w8(32'h3b95066a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6873d),
	.w1(32'h3bdfdbd7),
	.w2(32'hbc7dbbf2),
	.w3(32'hbc0005bf),
	.w4(32'h3c93159c),
	.w5(32'hbbeeb7cf),
	.w6(32'hbb55b9a2),
	.w7(32'hbbcf94b5),
	.w8(32'hbc39e6d4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c3d91),
	.w1(32'hbbf9b195),
	.w2(32'hbbbf6090),
	.w3(32'hbb7bc477),
	.w4(32'hbc7b29e0),
	.w5(32'h3c22735b),
	.w6(32'hbb2d8e90),
	.w7(32'hb89d475e),
	.w8(32'h3bcf8d56),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53694d),
	.w1(32'h3b1bc5ed),
	.w2(32'h3b4c04e6),
	.w3(32'hbb16cf76),
	.w4(32'hbc35390d),
	.w5(32'hbbdc3a8e),
	.w6(32'hbc2b2348),
	.w7(32'hbc85bea4),
	.w8(32'hbb27b7c3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9945a9),
	.w1(32'hba3db1ae),
	.w2(32'hbc0365e6),
	.w3(32'hbababd2b),
	.w4(32'h3c966979),
	.w5(32'h3ca0ef41),
	.w6(32'hbc330e17),
	.w7(32'hbbba9b1e),
	.w8(32'hbcdb3038),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b938852),
	.w1(32'h3c4eb2a7),
	.w2(32'hbc229ce7),
	.w3(32'hbb1eac12),
	.w4(32'h3c7ddefe),
	.w5(32'hbbc24c39),
	.w6(32'hbbe97ed5),
	.w7(32'hbb8b63ed),
	.w8(32'hbc8036da),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87b4ef),
	.w1(32'hbbc4cdb8),
	.w2(32'h39c0e65a),
	.w3(32'h3b0e1cf2),
	.w4(32'h398640d5),
	.w5(32'h38885307),
	.w6(32'hbc2da9a4),
	.w7(32'hb7fbd679),
	.w8(32'hb99a7d45),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36835dfb),
	.w1(32'hb6faed11),
	.w2(32'hb67233b5),
	.w3(32'h36aa43c9),
	.w4(32'hb71abc88),
	.w5(32'hb74f0186),
	.w6(32'h36acb8e8),
	.w7(32'hb73c2f40),
	.w8(32'hb7150d93),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4f2b889),
	.w1(32'hb69e0246),
	.w2(32'h36883540),
	.w3(32'hb4be3aa2),
	.w4(32'hb68bcc71),
	.w5(32'h36282fbd),
	.w6(32'h357568f5),
	.w7(32'hb666a223),
	.w8(32'h365a5d58),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h353be254),
	.w1(32'hb670d120),
	.w2(32'h363b3fea),
	.w3(32'h35b09234),
	.w4(32'hb656aaca),
	.w5(32'h35ab1856),
	.w6(32'hb51ffbfa),
	.w7(32'hb6f4f32b),
	.w8(32'hb6013744),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3811f4e3),
	.w1(32'hb9f09e39),
	.w2(32'hba01b852),
	.w3(32'h3820ebfc),
	.w4(32'hba5089d5),
	.w5(32'hba0d4d8d),
	.w6(32'hb919acaa),
	.w7(32'hb7d72f00),
	.w8(32'h3944475f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1121c3),
	.w1(32'h3a1d869e),
	.w2(32'h3a4e4eca),
	.w3(32'hb9ccca18),
	.w4(32'h3a161c18),
	.w5(32'h3a66ee4b),
	.w6(32'hb8d06900),
	.w7(32'h39988609),
	.w8(32'h3a096112),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ac647),
	.w1(32'hbc099940),
	.w2(32'hbb5789da),
	.w3(32'hb9858ab2),
	.w4(32'h3b016341),
	.w5(32'h3ba902a4),
	.w6(32'h3a7d7b8e),
	.w7(32'h3b896a84),
	.w8(32'h3b92819d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8293806),
	.w1(32'h3a744abd),
	.w2(32'h38192f0e),
	.w3(32'h39d776a9),
	.w4(32'h3a44b935),
	.w5(32'h39b3aeef),
	.w6(32'h386dbc17),
	.w7(32'h38986987),
	.w8(32'hb9ad5145),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d431d),
	.w1(32'h3ae223f3),
	.w2(32'hbaec1d6f),
	.w3(32'h3b05c347),
	.w4(32'h3ab131f5),
	.w5(32'hbab86f6f),
	.w6(32'h3a7418b5),
	.w7(32'h3ad6b584),
	.w8(32'hb7acb5cf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4b40c),
	.w1(32'h3a908fbf),
	.w2(32'h3a7d9ee9),
	.w3(32'h3998d4d7),
	.w4(32'h3a2b7aa5),
	.w5(32'h3a112a37),
	.w6(32'h38612f63),
	.w7(32'hb82b94d8),
	.w8(32'h38c0ed1d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6776f),
	.w1(32'hbb8ab96e),
	.w2(32'hbb3a12bf),
	.w3(32'h3aa64e75),
	.w4(32'h39cd8afe),
	.w5(32'h3b41b826),
	.w6(32'h3adbb381),
	.w7(32'h3b68d69d),
	.w8(32'h3ba0e190),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62c419),
	.w1(32'h3aaaded5),
	.w2(32'h3a5dd701),
	.w3(32'h3a824b37),
	.w4(32'h39b63116),
	.w5(32'hb8a7f48a),
	.w6(32'h3a1052d8),
	.w7(32'h35c8fe84),
	.w8(32'hb9c2a4e1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383cf306),
	.w1(32'h38290ddf),
	.w2(32'h37b7094e),
	.w3(32'h37a595a5),
	.w4(32'hb6ea3dbd),
	.w5(32'hb7330f20),
	.w6(32'h3784b474),
	.w7(32'hb60a5b0d),
	.w8(32'h37297719),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3760eb41),
	.w1(32'hbae6ab1d),
	.w2(32'hbb3144f0),
	.w3(32'h3999d01e),
	.w4(32'h39fc72ae),
	.w5(32'h3808ffc0),
	.w6(32'hb8ed1123),
	.w7(32'h3a8c828a),
	.w8(32'h3a3c302a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3513a95a),
	.w1(32'h35f7788b),
	.w2(32'h36ec1261),
	.w3(32'hb65b2ef8),
	.w4(32'hb5f986ec),
	.w5(32'h3645b773),
	.w6(32'hb5df983c),
	.w7(32'hb6a715ba),
	.w8(32'hb5b68474),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f4cba),
	.w1(32'hbc99e487),
	.w2(32'hbcae8c7c),
	.w3(32'hbc8bad30),
	.w4(32'hb9bee960),
	.w5(32'h3baac43b),
	.w6(32'hbc8b3978),
	.w7(32'h3c2da09e),
	.w8(32'h3ca4bc39),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22e974),
	.w1(32'hbab9bc95),
	.w2(32'hbaa127e8),
	.w3(32'h38f1ce78),
	.w4(32'h38db93f9),
	.w5(32'h3975deab),
	.w6(32'h3a5ba9b7),
	.w7(32'h3a9ffd94),
	.w8(32'h3a6feb0a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb928dab2),
	.w1(32'hb6992fd1),
	.w2(32'h39724eee),
	.w3(32'hb9940e7e),
	.w4(32'hb9088f0b),
	.w5(32'h3902520e),
	.w6(32'hb9831699),
	.w7(32'hb8d026df),
	.w8(32'h3940b11b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa1cb0),
	.w1(32'hb9879fed),
	.w2(32'hb8935ef2),
	.w3(32'hb804a4ca),
	.w4(32'hb6d7d7bf),
	.w5(32'h3933b177),
	.w6(32'hb83e0baa),
	.w7(32'h388c400a),
	.w8(32'h394feb1a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a615565),
	.w1(32'h3a5c89ff),
	.w2(32'hba1d6ccb),
	.w3(32'h39f2b119),
	.w4(32'h38e9ef49),
	.w5(32'hba8b377a),
	.w6(32'hb9816aaf),
	.w7(32'hb8f663e5),
	.w8(32'hba15bedf),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376e41cc),
	.w1(32'h3644fc3e),
	.w2(32'h379b742a),
	.w3(32'h36f0617f),
	.w4(32'hb624af52),
	.w5(32'h37221357),
	.w6(32'h36f29210),
	.w7(32'h356d79b8),
	.w8(32'h35bd9b3b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36223473),
	.w1(32'h361f57e1),
	.w2(32'h37394d66),
	.w3(32'h362aa19a),
	.w4(32'h35a9e807),
	.w5(32'h37517018),
	.w6(32'h35a03f05),
	.w7(32'hb67f5bb3),
	.w8(32'h365f62d2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa6c82),
	.w1(32'h3aaa48ad),
	.w2(32'h3a382a41),
	.w3(32'h39ddd145),
	.w4(32'h37cc3da6),
	.w5(32'hb9c88476),
	.w6(32'hb9d4edac),
	.w7(32'hbab018e0),
	.w8(32'hbae120c0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa748f4),
	.w1(32'hba2d3478),
	.w2(32'hb825c1c4),
	.w3(32'hbaadeaa9),
	.w4(32'h3a0050a3),
	.w5(32'h3abc1df2),
	.w6(32'hba1d0f7a),
	.w7(32'h3a880d5f),
	.w8(32'h3a9b027e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bee845),
	.w1(32'hb6c29c02),
	.w2(32'hb63966c2),
	.w3(32'h34a199c3),
	.w4(32'hb71e568d),
	.w5(32'hb7a80aea),
	.w6(32'hb6c59ddd),
	.w7(32'hb6af056a),
	.w8(32'hb786ea62),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f706f),
	.w1(32'hb98e71f9),
	.w2(32'h3963283d),
	.w3(32'hba36987d),
	.w4(32'hba1bada9),
	.w5(32'hb84cabc2),
	.w6(32'hb9fc8d54),
	.w7(32'hba122bd7),
	.w8(32'hb8f46358),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc5d8b),
	.w1(32'h37427957),
	.w2(32'h37a7b84b),
	.w3(32'h37abb324),
	.w4(32'h3676d52f),
	.w5(32'h3731d524),
	.w6(32'h366a4493),
	.w7(32'hb71be1e8),
	.w8(32'hb520381b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df7892),
	.w1(32'hb93d629c),
	.w2(32'hb89d29af),
	.w3(32'h39862091),
	.w4(32'hb7c5a9b9),
	.w5(32'h3950b736),
	.w6(32'hb7ba3e80),
	.w7(32'hb8360cb6),
	.w8(32'h3926fb75),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb872408),
	.w1(32'hbb33fa7e),
	.w2(32'hbb818344),
	.w3(32'hbb87afb8),
	.w4(32'hbad34247),
	.w5(32'hbb11f6ee),
	.w6(32'hbb3859fa),
	.w7(32'hba35d4df),
	.w8(32'hbb0faff8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1d2b5),
	.w1(32'hba57ccef),
	.w2(32'h38a0f4e2),
	.w3(32'hb9fee20f),
	.w4(32'h3865dbd8),
	.w5(32'h3973c23c),
	.w6(32'h390b28ee),
	.w7(32'h398d6e59),
	.w8(32'h39b12af2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39344409),
	.w1(32'h393debd2),
	.w2(32'h378f51a4),
	.w3(32'h393a5c63),
	.w4(32'h391f88e0),
	.w5(32'h373b4df7),
	.w6(32'h38ebed4a),
	.w7(32'h38790562),
	.w8(32'hb74ef2d5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e279b),
	.w1(32'hba9b3d6b),
	.w2(32'hba77669f),
	.w3(32'hba4716de),
	.w4(32'hb9867eab),
	.w5(32'h3993d048),
	.w6(32'hba474962),
	.w7(32'h3a19dc77),
	.w8(32'h3a8ada57),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b890a1),
	.w1(32'hbb966f0f),
	.w2(32'hbb1af221),
	.w3(32'h3a6dc36f),
	.w4(32'h393e7a65),
	.w5(32'h3aa37cde),
	.w6(32'h39d5179b),
	.w7(32'h3b114580),
	.w8(32'h3b3920e8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aac501),
	.w1(32'hba9b73a2),
	.w2(32'h3a14070b),
	.w3(32'hb5f19000),
	.w4(32'h3a32d512),
	.w5(32'h3a932e84),
	.w6(32'h38e4684e),
	.w7(32'h39e2d704),
	.w8(32'h39c66b43),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351534fd),
	.w1(32'hb64e9fc3),
	.w2(32'h369319f8),
	.w3(32'hb6303cd4),
	.w4(32'hb6705b4d),
	.w5(32'h3601a726),
	.w6(32'hb61c06f7),
	.w7(32'hb63821bb),
	.w8(32'h3555202e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a815598),
	.w1(32'hbb3999c0),
	.w2(32'hbb0fdba1),
	.w3(32'h39ef0070),
	.w4(32'hb9061669),
	.w5(32'h3a2e27c9),
	.w6(32'h3a4a62b4),
	.w7(32'h3aee9ace),
	.w8(32'h3b051d2e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cf678),
	.w1(32'h38e090bd),
	.w2(32'hb8cd482c),
	.w3(32'hb9014702),
	.w4(32'h391f7bec),
	.w5(32'hb8e81498),
	.w6(32'hb8a7abd2),
	.w7(32'h39045015),
	.w8(32'hb879d60a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d2d3e),
	.w1(32'hbafb25cc),
	.w2(32'hbaa04340),
	.w3(32'hba2700c6),
	.w4(32'h3859beaf),
	.w5(32'h38101536),
	.w6(32'h396d5f27),
	.w7(32'h39e00978),
	.w8(32'h399fa83c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83f047),
	.w1(32'h3a9bef67),
	.w2(32'hb9e7c7e3),
	.w3(32'h3ab8be21),
	.w4(32'h3a7a3958),
	.w5(32'hba60d470),
	.w6(32'h3ad77270),
	.w7(32'h3a5455ac),
	.w8(32'hba989dde),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9088fb),
	.w1(32'hbc225499),
	.w2(32'hbbb08cd4),
	.w3(32'hbb32b204),
	.w4(32'hbb8c674e),
	.w5(32'hba12ed02),
	.w6(32'h39b944b8),
	.w7(32'h3b05f1b7),
	.w8(32'h3b4e7b3c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a20b61),
	.w1(32'hba73548d),
	.w2(32'hba3e57fb),
	.w3(32'h39dcf965),
	.w4(32'hb9e73c77),
	.w5(32'hb927a4a9),
	.w6(32'h3a0b6dd6),
	.w7(32'h3953693b),
	.w8(32'h39f20a7f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba749856),
	.w1(32'hb9b0ca5f),
	.w2(32'h39f7bf16),
	.w3(32'hba3ca7d7),
	.w4(32'h3a6ef908),
	.w5(32'h3b1f8bd0),
	.w6(32'hb8be46c7),
	.w7(32'h39fb48f7),
	.w8(32'h3a9fdf5d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74ce77f),
	.w1(32'hb77ad5e4),
	.w2(32'h360fcdf8),
	.w3(32'hb773d41f),
	.w4(32'hb74ebc40),
	.w5(32'h36d6e17b),
	.w6(32'hb702c75b),
	.w7(32'hb6af3a52),
	.w8(32'h36c6b1fb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a583d4b),
	.w1(32'hbb14ac17),
	.w2(32'hbb6cbfb5),
	.w3(32'h39d4a5ea),
	.w4(32'h3ab5bcb7),
	.w5(32'h3af37c5d),
	.w6(32'h39984f46),
	.w7(32'h3a3c9899),
	.w8(32'h3a8cd872),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ae3de),
	.w1(32'h3a34c476),
	.w2(32'h3a1e84d4),
	.w3(32'hb95135d8),
	.w4(32'hba05c598),
	.w5(32'h39ce767b),
	.w6(32'h39f9d6a4),
	.w7(32'h391d3df3),
	.w8(32'h3918bd44),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099d84),
	.w1(32'hbb4154a0),
	.w2(32'h3928807a),
	.w3(32'hbaf51bfa),
	.w4(32'hb984630c),
	.w5(32'h3ab544f0),
	.w6(32'hba995a6b),
	.w7(32'h3a880421),
	.w8(32'h3af9b19b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1090ee),
	.w1(32'hbb0359f7),
	.w2(32'hbb2d9975),
	.w3(32'h3a23804b),
	.w4(32'hba1d002a),
	.w5(32'hb99dd240),
	.w6(32'h3a0ac92d),
	.w7(32'h3a9d2a12),
	.w8(32'h3ab6d7fd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93139ef),
	.w1(32'hba528f99),
	.w2(32'hbab371ba),
	.w3(32'hb9e2c7f0),
	.w4(32'hba8e20a8),
	.w5(32'hba62cc9b),
	.w6(32'hba242953),
	.w7(32'hb9906495),
	.w8(32'h391dfe44),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372a8a93),
	.w1(32'hb59d7ef8),
	.w2(32'h3781a27b),
	.w3(32'h371a6df5),
	.w4(32'h366d8028),
	.w5(32'h37cd3ff0),
	.w6(32'h3787f09f),
	.w7(32'h3790e5a7),
	.w8(32'h37bede76),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d20cc6),
	.w1(32'hb9ab307f),
	.w2(32'hb99d8785),
	.w3(32'h3982f3ae),
	.w4(32'hb83ae179),
	.w5(32'h389df0eb),
	.w6(32'h38d1f2c7),
	.w7(32'h36bf0cde),
	.w8(32'h390564a4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac6459),
	.w1(32'hbadfb291),
	.w2(32'hbb18bd59),
	.w3(32'hba4fe5eb),
	.w4(32'h3a4d9f54),
	.w5(32'hb842b6c2),
	.w6(32'h3a349a9b),
	.w7(32'h3a74e1c7),
	.w8(32'hb981ecfc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f3f1aa),
	.w1(32'h39468b9f),
	.w2(32'h3a18d0d7),
	.w3(32'hb93bb3a3),
	.w4(32'h389b10c8),
	.w5(32'h39bbaf5a),
	.w6(32'hb9abab73),
	.w7(32'hba011910),
	.w8(32'hb8aac412),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787d1f5),
	.w1(32'hb7ff31fa),
	.w2(32'hb7d64a85),
	.w3(32'hb6d5f297),
	.w4(32'hb6b2c268),
	.w5(32'h372fd29c),
	.w6(32'hb647b524),
	.w7(32'h36dea121),
	.w8(32'hb67b4e32),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8105a),
	.w1(32'hb7990f84),
	.w2(32'h39ec445f),
	.w3(32'hb9bf3253),
	.w4(32'h39edfa52),
	.w5(32'h3a6c579c),
	.w6(32'hb92aaba8),
	.w7(32'h3a06b04f),
	.w8(32'h3a6426d2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cce05e),
	.w1(32'hb97e0042),
	.w2(32'hba0fd090),
	.w3(32'hb82a0f03),
	.w4(32'hb9854e48),
	.w5(32'hba0f445c),
	.w6(32'h387648f6),
	.w7(32'h38fa108d),
	.w8(32'hb873fbde),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eae994),
	.w1(32'hba009c6c),
	.w2(32'hba610cba),
	.w3(32'h398f5ca8),
	.w4(32'h3a8c677e),
	.w5(32'h3a3d297e),
	.w6(32'h3a2bc03f),
	.w7(32'h3a6719a9),
	.w8(32'h38bc89ac),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37866451),
	.w1(32'h3717a54d),
	.w2(32'h37111be8),
	.w3(32'h3795f824),
	.w4(32'h37812e96),
	.w5(32'h372cdde8),
	.w6(32'h37230828),
	.w7(32'h371f73e9),
	.w8(32'h371fbe65),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea9e85),
	.w1(32'hbb9c4d7a),
	.w2(32'hbbb8d113),
	.w3(32'hbb238fab),
	.w4(32'hba9e9e8a),
	.w5(32'h3ad6c8b7),
	.w6(32'hbb56ed1a),
	.w7(32'h3b053bc8),
	.w8(32'h3bbd8b73),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a7bc7a),
	.w1(32'h37058da6),
	.w2(32'h3702612e),
	.w3(32'h35a11f43),
	.w4(32'h369a8865),
	.w5(32'h367ea2bc),
	.w6(32'hb635f170),
	.w7(32'hb59df87b),
	.w8(32'h34c7eaf5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c4a5e),
	.w1(32'h3aa852e5),
	.w2(32'hb6dcb986),
	.w3(32'hb93bebe5),
	.w4(32'h378b84e7),
	.w5(32'hba41c575),
	.w6(32'hba57e6e0),
	.w7(32'hb88b5eb1),
	.w8(32'hb970c0bc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9268957),
	.w1(32'hb8b3f40d),
	.w2(32'hb8876066),
	.w3(32'hb94da53d),
	.w4(32'hb8a4ff04),
	.w5(32'hb8926be9),
	.w6(32'hb942cbde),
	.w7(32'hb8b5ad59),
	.w8(32'hb888ddfc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7889e5),
	.w1(32'h39fc5dba),
	.w2(32'h392b5620),
	.w3(32'hba52a7d1),
	.w4(32'h3a5030d5),
	.w5(32'h3a3e5977),
	.w6(32'hba07be55),
	.w7(32'h3888fb9e),
	.w8(32'h3917b737),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37690948),
	.w1(32'h3749ff30),
	.w2(32'h3753b06c),
	.w3(32'h372ac537),
	.w4(32'h362d7c11),
	.w5(32'h3710cfd3),
	.w6(32'h360842ad),
	.w7(32'hb64aa89e),
	.w8(32'h358675fa),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc581e),
	.w1(32'hba954829),
	.w2(32'hba99f96b),
	.w3(32'h3a56f28d),
	.w4(32'hba8501d7),
	.w5(32'hb9f88c4b),
	.w6(32'h3a86b478),
	.w7(32'h39d3610d),
	.w8(32'h39db4308),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb750fe77),
	.w1(32'hb52ea782),
	.w2(32'hb90f15cd),
	.w3(32'hb7803906),
	.w4(32'hbb0e4686),
	.w5(32'hba4f4d4f),
	.w6(32'hb7105953),
	.w7(32'hbb5070db),
	.w8(32'h3c79062b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0333cc),
	.w1(32'hbb0dedf3),
	.w2(32'hbbb1dd68),
	.w3(32'h3a443d2d),
	.w4(32'hbaddf949),
	.w5(32'hb9b8fb6b),
	.w6(32'h3bebcda2),
	.w7(32'h3b81fb68),
	.w8(32'h3bfb3144),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386de3d4),
	.w1(32'h3a7de4d5),
	.w2(32'hbb20db3c),
	.w3(32'h3ad482b5),
	.w4(32'hba9dbffd),
	.w5(32'h3af8c746),
	.w6(32'h3bc0929e),
	.w7(32'h398c54ab),
	.w8(32'h3b92e06f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f39bc),
	.w1(32'hb9200ac4),
	.w2(32'h3ade6974),
	.w3(32'hb9412da3),
	.w4(32'h3bcd5ec1),
	.w5(32'h3c1da1f0),
	.w6(32'h3b3a7374),
	.w7(32'hbb86f5e2),
	.w8(32'hbc205edc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13ac8e),
	.w1(32'hbb816f62),
	.w2(32'hbb4eec1f),
	.w3(32'h3ba7659a),
	.w4(32'h3acf0444),
	.w5(32'h3a552281),
	.w6(32'hbc8ffe42),
	.w7(32'hbc465f1f),
	.w8(32'hbc5c2b66),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c0e4c),
	.w1(32'h3af9b7bc),
	.w2(32'hbc48642d),
	.w3(32'h3b6c05ee),
	.w4(32'hb8b1debe),
	.w5(32'hba2e8dc7),
	.w6(32'hbbdb08c5),
	.w7(32'hb9d6b9aa),
	.w8(32'h3b21096a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc513e45),
	.w1(32'hbbaa9eae),
	.w2(32'hbc331a06),
	.w3(32'h3a3ce246),
	.w4(32'hbacc473e),
	.w5(32'hbb6e8a66),
	.w6(32'h3a5e0f7b),
	.w7(32'h3b9069db),
	.w8(32'hb9d5b734),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64d057),
	.w1(32'hbbc31755),
	.w2(32'hbc808817),
	.w3(32'hbc014798),
	.w4(32'hbc783662),
	.w5(32'hbcd8c230),
	.w6(32'hbbd899bc),
	.w7(32'h3cbb8c9a),
	.w8(32'h3d120708),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa91884),
	.w1(32'hbc904346),
	.w2(32'hbc1bae54),
	.w3(32'hbba27309),
	.w4(32'hbad95f4c),
	.w5(32'h3b8bd948),
	.w6(32'h3cf40b39),
	.w7(32'h3c88d76d),
	.w8(32'h3ca87b8e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc205fba),
	.w1(32'hbc8db8dc),
	.w2(32'hbc776e5b),
	.w3(32'h3c8b44d3),
	.w4(32'hbbe358da),
	.w5(32'h3b13c1f2),
	.w6(32'hbabd42e9),
	.w7(32'hbbfa3fe8),
	.w8(32'hbbea6b68),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90af6f),
	.w1(32'h3c08c5c9),
	.w2(32'h3b6ceecf),
	.w3(32'h3b6eb5b7),
	.w4(32'hbb056e39),
	.w5(32'hbbddeefb),
	.w6(32'hbc0335c6),
	.w7(32'hbc2ed982),
	.w8(32'h3aa0ec2c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c428afe),
	.w1(32'h3bfafb44),
	.w2(32'hbbb4aae8),
	.w3(32'hbaa505b4),
	.w4(32'h3b0fba82),
	.w5(32'h3b973548),
	.w6(32'h3a55c983),
	.w7(32'hbbcb37c9),
	.w8(32'hbbe6232c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba797cf),
	.w1(32'h3b9d2a28),
	.w2(32'h3b2a5f58),
	.w3(32'h3b55db81),
	.w4(32'h38ae2063),
	.w5(32'hbb4c107d),
	.w6(32'h3abf2adf),
	.w7(32'hbb93e59c),
	.w8(32'hbc152d1e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac84db1),
	.w1(32'hb8f49362),
	.w2(32'h3c06ceac),
	.w3(32'hbba0a428),
	.w4(32'hbbd039da),
	.w5(32'hbb881566),
	.w6(32'hbc153d49),
	.w7(32'hbc9c9b63),
	.w8(32'hbd38c921),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce92312),
	.w1(32'h3d060fd3),
	.w2(32'hbc9fbda4),
	.w3(32'hbb17a019),
	.w4(32'hbb8da657),
	.w5(32'hbba99a7b),
	.w6(32'hbca0db77),
	.w7(32'h3c0fab35),
	.w8(32'h3a58d539),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fe0c0),
	.w1(32'hbca8e859),
	.w2(32'h3c96551d),
	.w3(32'hbbf2de5f),
	.w4(32'hbc13805a),
	.w5(32'hbbab7914),
	.w6(32'h3c5413fd),
	.w7(32'hbc8b5588),
	.w8(32'hbcc16299),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd5585e),
	.w1(32'h3c9f0fe3),
	.w2(32'h3c518de0),
	.w3(32'hbc020cc6),
	.w4(32'hbc243039),
	.w5(32'h3b2676a5),
	.w6(32'hbd0a6d64),
	.w7(32'h3c1b231f),
	.w8(32'h3cd453d5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1aacc4),
	.w1(32'hbc2e8cc2),
	.w2(32'h3cbec420),
	.w3(32'h3cab8970),
	.w4(32'h3b8da191),
	.w5(32'hbbaea86a),
	.w6(32'hbc957040),
	.w7(32'hbd0239eb),
	.w8(32'hbcdc333a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2636b0),
	.w1(32'h3c34a955),
	.w2(32'h3afebeab),
	.w3(32'h3b5c4de1),
	.w4(32'h3b9afdb1),
	.w5(32'h3bc6bf18),
	.w6(32'h3bc845dc),
	.w7(32'h3b14de7b),
	.w8(32'h3bfa2241),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd9a9a),
	.w1(32'h3b06b0cf),
	.w2(32'hb983300e),
	.w3(32'h3b708c91),
	.w4(32'hbca4c70a),
	.w5(32'hbbb25e36),
	.w6(32'h3b61e7bd),
	.w7(32'h3c23572a),
	.w8(32'h3d568e1c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafa62f),
	.w1(32'hb9d43e4e),
	.w2(32'hbc32764a),
	.w3(32'hbc32c62d),
	.w4(32'h3c5443d1),
	.w5(32'h3c23dae1),
	.w6(32'h3b7cf726),
	.w7(32'h3c07c544),
	.w8(32'h3c2cf580),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6adc5),
	.w1(32'hbcbb44ec),
	.w2(32'h3aed37e8),
	.w3(32'h399b534e),
	.w4(32'h399777dd),
	.w5(32'h3c0953de),
	.w6(32'h3cc33612),
	.w7(32'h3bb93b99),
	.w8(32'hbad42e0b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399742b0),
	.w1(32'h3b7bb1ff),
	.w2(32'h3b929263),
	.w3(32'h3c057ef2),
	.w4(32'h3b2929a2),
	.w5(32'hbaa2cf63),
	.w6(32'hb8dfcabe),
	.w7(32'h3b42258d),
	.w8(32'h3c0a197c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6a4f9),
	.w1(32'h398f2cb0),
	.w2(32'hbbad2221),
	.w3(32'h39964d76),
	.w4(32'h3c509126),
	.w5(32'hba6f45d6),
	.w6(32'hb9a0ff7d),
	.w7(32'hbc6a3e7d),
	.w8(32'h3ae62cde),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe00bde),
	.w1(32'h3b93fcba),
	.w2(32'hbc16c50c),
	.w3(32'hbc473a39),
	.w4(32'hbc9d4b13),
	.w5(32'hbb5d020e),
	.w6(32'h3b91ffbf),
	.w7(32'h3c0778ab),
	.w8(32'h3cfd9f3b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0d484),
	.w1(32'hbc3d655b),
	.w2(32'h3a622c09),
	.w3(32'hbb94a91b),
	.w4(32'hbc18f890),
	.w5(32'h3afbdae5),
	.w6(32'h3bb5eb72),
	.w7(32'h3b34e754),
	.w8(32'hb91292d3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9aac8),
	.w1(32'hbc1d118a),
	.w2(32'hbb4ad936),
	.w3(32'hbabe4ad3),
	.w4(32'hbca44a2b),
	.w5(32'hbcace0b1),
	.w6(32'hbc01ac84),
	.w7(32'h3c3daf14),
	.w8(32'h3c856339),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10d866),
	.w1(32'hbc942c9c),
	.w2(32'h3c08227a),
	.w3(32'hbc5d0df8),
	.w4(32'h3ac58a86),
	.w5(32'hbb02816a),
	.w6(32'hbc1de0a3),
	.w7(32'h3ac8e539),
	.w8(32'h3b62fe87),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93c57a),
	.w1(32'h3c0ffea6),
	.w2(32'h3ba9dd04),
	.w3(32'hbb687025),
	.w4(32'hbb77b099),
	.w5(32'hbb9565d8),
	.w6(32'h3aa3d724),
	.w7(32'h3c16c0ad),
	.w8(32'hbc30b2ce),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3479ae),
	.w1(32'hbba310d5),
	.w2(32'hba616248),
	.w3(32'h3b4378ee),
	.w4(32'h3bb9bbe4),
	.w5(32'h3aa363c7),
	.w6(32'hbc98c3c5),
	.w7(32'hbcf486d7),
	.w8(32'hbd11a5eb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a694),
	.w1(32'h3ba580ac),
	.w2(32'hbc6b54c1),
	.w3(32'hbc105bc3),
	.w4(32'h3a01ab0d),
	.w5(32'h3b0fef90),
	.w6(32'hbcc7b088),
	.w7(32'h3c799ab8),
	.w8(32'h3d59ca41),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3eb9f6),
	.w1(32'hbd344f50),
	.w2(32'hba85de46),
	.w3(32'h3ab30e74),
	.w4(32'hbb157d0e),
	.w5(32'hbb41bb75),
	.w6(32'h3c255601),
	.w7(32'hbacfa468),
	.w8(32'h3c7c196a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39e4b6),
	.w1(32'hb9b09656),
	.w2(32'h3c840978),
	.w3(32'hb9a46747),
	.w4(32'hb9f9ef5b),
	.w5(32'hbc0af5e5),
	.w6(32'h3c0c0212),
	.w7(32'hbb950bb1),
	.w8(32'hbca2d0b7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cfce1),
	.w1(32'h3c3fc34b),
	.w2(32'hba582a24),
	.w3(32'h3b5a716c),
	.w4(32'h3bbc7d01),
	.w5(32'h3bc8a6a3),
	.w6(32'hbc2b9b10),
	.w7(32'hbc97680f),
	.w8(32'h3b0a5336),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef392b),
	.w1(32'h3c2064fc),
	.w2(32'hbcedd9d0),
	.w3(32'hbc1f5c58),
	.w4(32'hbb18dc62),
	.w5(32'hbbe41028),
	.w6(32'h3b89e095),
	.w7(32'hbc0dd6a7),
	.w8(32'h3ac9d5a1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ce020),
	.w1(32'h3c448808),
	.w2(32'h3b8c89d1),
	.w3(32'hba8dc859),
	.w4(32'h3c42572c),
	.w5(32'h3c94711c),
	.w6(32'h3c32b8f9),
	.w7(32'h3c5ea6d2),
	.w8(32'hbc9e229e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe936d),
	.w1(32'h3c332245),
	.w2(32'h3a162a93),
	.w3(32'h3c66f075),
	.w4(32'hbbe79700),
	.w5(32'hbc142161),
	.w6(32'hbc7da707),
	.w7(32'hbc7bd2d2),
	.w8(32'hbcdee3fb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8f339),
	.w1(32'h3a0db30d),
	.w2(32'hbc99d8ad),
	.w3(32'hbc8376a3),
	.w4(32'hbca1727b),
	.w5(32'hbc955c9f),
	.w6(32'hbc0d537c),
	.w7(32'hbc6922b6),
	.w8(32'hbc9b74a3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb71a5d),
	.w1(32'hbbd60369),
	.w2(32'h3cd88377),
	.w3(32'hbcafdc83),
	.w4(32'h3c828390),
	.w5(32'h3ca36bec),
	.w6(32'hbc6b6b60),
	.w7(32'hbd1b455b),
	.w8(32'hbd7dafae),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0bc5ce),
	.w1(32'h3ce3d08a),
	.w2(32'h3bff1dc9),
	.w3(32'h3c7ee756),
	.w4(32'hbc3ec9f5),
	.w5(32'hbbc02b15),
	.w6(32'hbcfc5314),
	.w7(32'h3bcaa696),
	.w8(32'hbba139e2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9363a8),
	.w1(32'hbc287857),
	.w2(32'h3bab7318),
	.w3(32'h3c427b8d),
	.w4(32'hb9aa2640),
	.w5(32'hbc2eef2e),
	.w6(32'hbb382193),
	.w7(32'h3a4b450d),
	.w8(32'hbc994dd0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c9b1c),
	.w1(32'h3c304f66),
	.w2(32'hbb870850),
	.w3(32'hbbd5e220),
	.w4(32'hbb257f4a),
	.w5(32'hbb6d20f6),
	.w6(32'hbbad3c3e),
	.w7(32'h3b35d18b),
	.w8(32'h3c415a16),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a765b9a),
	.w1(32'hb9cd4363),
	.w2(32'h39a79837),
	.w3(32'hba6926dc),
	.w4(32'hba783783),
	.w5(32'hb8de8342),
	.w6(32'h3bbfee07),
	.w7(32'h3bcb8702),
	.w8(32'hbc17ce90),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcceba00),
	.w1(32'hbcccd86d),
	.w2(32'hbb744ed6),
	.w3(32'hbbf0e190),
	.w4(32'hbbcdd838),
	.w5(32'hbbe18427),
	.w6(32'hbc161d70),
	.w7(32'h39f5ba6b),
	.w8(32'hbc08cd61),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd0e9d),
	.w1(32'h3bad8e4b),
	.w2(32'hba86f37f),
	.w3(32'hbae522c2),
	.w4(32'hbb6394c7),
	.w5(32'h3b230309),
	.w6(32'hbacc6c6a),
	.w7(32'hb8cf801b),
	.w8(32'h3abb610e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8068a4),
	.w1(32'h3b2febe3),
	.w2(32'h3cf3b43c),
	.w3(32'h3b827ef6),
	.w4(32'h3c7195a4),
	.w5(32'h3c051d9d),
	.w6(32'hbab3bdb7),
	.w7(32'hbceae330),
	.w8(32'hbd002c5e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82124a),
	.w1(32'h3c19eae0),
	.w2(32'hbae08027),
	.w3(32'h3c8953cc),
	.w4(32'hba88697a),
	.w5(32'hbaf86bea),
	.w6(32'hbc9f109a),
	.w7(32'h3a890d73),
	.w8(32'h3c7b3e28),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98f3eb),
	.w1(32'hbae43469),
	.w2(32'hbb4ec5a5),
	.w3(32'hba76382b),
	.w4(32'hbc3dbed0),
	.w5(32'hbc16f9a5),
	.w6(32'h3bf925ba),
	.w7(32'h3c8d3fd6),
	.w8(32'h3c481dc8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54689f),
	.w1(32'hbab8eca3),
	.w2(32'hbab5c9af),
	.w3(32'hbb99d326),
	.w4(32'h3c15ae7f),
	.w5(32'hbc357990),
	.w6(32'hbbb109dc),
	.w7(32'hbb0e4fc1),
	.w8(32'hbb8f0b6d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94cd6e),
	.w1(32'h3c82c02e),
	.w2(32'h3a9852c8),
	.w3(32'hbbd3cf52),
	.w4(32'hbbb7b408),
	.w5(32'hbbac67ca),
	.w6(32'hbc0e2d1e),
	.w7(32'hbc0d6a77),
	.w8(32'hbb862531),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b301b54),
	.w1(32'h3c0dbda3),
	.w2(32'hbb25934c),
	.w3(32'h3b5232f9),
	.w4(32'hbbf8b76b),
	.w5(32'hbb145775),
	.w6(32'h3a84fc9a),
	.w7(32'h3bdff686),
	.w8(32'hbc3de7e5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81f89c),
	.w1(32'hbc57763a),
	.w2(32'hbc078488),
	.w3(32'hbc01cc91),
	.w4(32'hbc8d3970),
	.w5(32'hbc3c8057),
	.w6(32'hbb26ecba),
	.w7(32'h3c63b35b),
	.w8(32'h3d1c79cb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule