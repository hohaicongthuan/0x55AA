module layer_6_featuremap_116(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32a908),
	.w1(32'hbc1b302a),
	.w2(32'hbc1fd81e),
	.w3(32'hbadbcae4),
	.w4(32'hbb1f36ee),
	.w5(32'hbba66e5d),
	.w6(32'hbbcb4249),
	.w7(32'hbc02bb06),
	.w8(32'hbc07ef9f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e1ab1),
	.w1(32'hbb6f3d63),
	.w2(32'hbb58f340),
	.w3(32'hbab32a57),
	.w4(32'hbb1edc05),
	.w5(32'hbba442cb),
	.w6(32'hbb97e15a),
	.w7(32'hbba4fc85),
	.w8(32'hbbc7adc3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77caf3),
	.w1(32'h3c8263a2),
	.w2(32'hbc645f2e),
	.w3(32'h3c2b1eb7),
	.w4(32'h3c541242),
	.w5(32'h3caacb05),
	.w6(32'h3cf9e5d2),
	.w7(32'h3c5b7c4b),
	.w8(32'h3a275517),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a384a),
	.w1(32'h39468e7b),
	.w2(32'h39662a42),
	.w3(32'h3b29f60c),
	.w4(32'h3b520a11),
	.w5(32'h3a995cbb),
	.w6(32'h3b91a354),
	.w7(32'h3b01af1b),
	.w8(32'h3a3ed787),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe38a),
	.w1(32'h3b09ecf7),
	.w2(32'h3b20e616),
	.w3(32'hbc05018a),
	.w4(32'hbc1c8be7),
	.w5(32'hbbb4b08f),
	.w6(32'h398baf7f),
	.w7(32'hbb4f90fa),
	.w8(32'hbc70eb9c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b636e61),
	.w1(32'hbb8fc479),
	.w2(32'hbb8f0a60),
	.w3(32'hbab61af7),
	.w4(32'hbb830c94),
	.w5(32'hbb169e96),
	.w6(32'hbbb3ec76),
	.w7(32'hbb9aac88),
	.w8(32'hbb72094f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc266cfa),
	.w1(32'hbbd48606),
	.w2(32'hbb509717),
	.w3(32'hbb3cfd40),
	.w4(32'h3ab4f81c),
	.w5(32'hba122a03),
	.w6(32'hbc1e155e),
	.w7(32'hbbcf238f),
	.w8(32'hbb6e6a3c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cea42),
	.w1(32'h3bc38177),
	.w2(32'h3baf1b6c),
	.w3(32'hbbe18858),
	.w4(32'hbb9469f7),
	.w5(32'h3ab0c9b8),
	.w6(32'h3a8a5192),
	.w7(32'h3b5c5bc4),
	.w8(32'h3c2153d0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4fb67),
	.w1(32'hbc904e3b),
	.w2(32'hbc87ec28),
	.w3(32'h3bed541e),
	.w4(32'h3ba3ccb8),
	.w5(32'h3b67b683),
	.w6(32'h3b3ae2bb),
	.w7(32'hbbe0d49b),
	.w8(32'hbc766266),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10ec23),
	.w1(32'hba10b6d8),
	.w2(32'hbab09014),
	.w3(32'hbb148798),
	.w4(32'hb9c8d9de),
	.w5(32'h39927950),
	.w6(32'hbaf93f1d),
	.w7(32'hb96870e2),
	.w8(32'hbb436baa),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7bd1c),
	.w1(32'h3b2c9331),
	.w2(32'hbc32c244),
	.w3(32'hbb6ac3ac),
	.w4(32'hbb4af6b1),
	.w5(32'hbbe30406),
	.w6(32'h3ab4106d),
	.w7(32'hb9d15418),
	.w8(32'hbbe93596),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b3d5e),
	.w1(32'hbb2cb79f),
	.w2(32'hba55f48a),
	.w3(32'hbc42ea0b),
	.w4(32'hbc094e26),
	.w5(32'hbc12e2b2),
	.w6(32'hbbce353c),
	.w7(32'hbab0f825),
	.w8(32'hbb8f0419),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fcf08),
	.w1(32'hbb446a23),
	.w2(32'h3b650155),
	.w3(32'hbb3d161c),
	.w4(32'h3b571022),
	.w5(32'hbb646ae1),
	.w6(32'hbb4e415b),
	.w7(32'h3b3dffa5),
	.w8(32'hbb2115f4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f8fa0),
	.w1(32'hbc6dc744),
	.w2(32'hbc065a9d),
	.w3(32'hbba06e02),
	.w4(32'h3b2f6d64),
	.w5(32'hbb8d810d),
	.w6(32'h3b4ac8a7),
	.w7(32'hbbbf65a6),
	.w8(32'hbadcb3c9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11f8a3),
	.w1(32'hbb92f064),
	.w2(32'hbb3e0f59),
	.w3(32'h3b4b12fd),
	.w4(32'hb89d145e),
	.w5(32'hbb8a5ad5),
	.w6(32'h3a10b9eb),
	.w7(32'hba4bc148),
	.w8(32'hbb6e2f1c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e441b),
	.w1(32'h3a983472),
	.w2(32'hba61e88d),
	.w3(32'h3ab7078d),
	.w4(32'hb95896a7),
	.w5(32'h39ad1057),
	.w6(32'hb82b05b4),
	.w7(32'hb98f2478),
	.w8(32'hbb11b069),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc557),
	.w1(32'hbbb6e2c7),
	.w2(32'hbba03dd0),
	.w3(32'h3c7b0299),
	.w4(32'hbbacb5b3),
	.w5(32'hbaf899de),
	.w6(32'h3ba5d15e),
	.w7(32'hbbd67e61),
	.w8(32'h3b6b7f1c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7755b1a),
	.w1(32'hba3d91da),
	.w2(32'hbad77d66),
	.w3(32'h3b6b3e93),
	.w4(32'h3b119fba),
	.w5(32'hb90e0c5d),
	.w6(32'hbad66572),
	.w7(32'hbb48370e),
	.w8(32'hbb6ddfdf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91fc11),
	.w1(32'h3aebb308),
	.w2(32'hbada100f),
	.w3(32'h3aea652c),
	.w4(32'hba1fcc9f),
	.w5(32'hbb0f1c40),
	.w6(32'hb958c121),
	.w7(32'hba591575),
	.w8(32'hbb6f4176),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdccca7),
	.w1(32'hbbbd4dec),
	.w2(32'hb989d99e),
	.w3(32'hbb994568),
	.w4(32'hbbd1b9bc),
	.w5(32'hbb4213de),
	.w6(32'hbbbe6bf1),
	.w7(32'hbb66a5a2),
	.w8(32'h3c2ef03f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35db34),
	.w1(32'h3b129da9),
	.w2(32'hb9ab9164),
	.w3(32'h3ad68898),
	.w4(32'h3acd736d),
	.w5(32'h38b5c2dd),
	.w6(32'h3b427129),
	.w7(32'h3a3a582e),
	.w8(32'h3aa48ca4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba260a20),
	.w1(32'hbb3a65c1),
	.w2(32'hbc1b7596),
	.w3(32'h39ded1ff),
	.w4(32'hbc0833e8),
	.w5(32'hbbdedce9),
	.w6(32'h390ce3cb),
	.w7(32'hbc0c716d),
	.w8(32'hbb86e7c5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb056cb5),
	.w1(32'h3c2b3174),
	.w2(32'h3b402823),
	.w3(32'h3b9ece15),
	.w4(32'h3ab84965),
	.w5(32'hbaafc8bb),
	.w6(32'h3bda121f),
	.w7(32'h3a20ea43),
	.w8(32'hbc0d84a8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca639c1),
	.w1(32'hbc895983),
	.w2(32'hbc78f3c6),
	.w3(32'h3a86cbcd),
	.w4(32'h3c45872e),
	.w5(32'h3c4c85ca),
	.w6(32'hbc5a0ea4),
	.w7(32'hbc8f45fc),
	.w8(32'hbb09c1d1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1cba),
	.w1(32'hbc18bb99),
	.w2(32'hbbf05f1e),
	.w3(32'h3cee382a),
	.w4(32'h3ce95740),
	.w5(32'h3ca5cd3c),
	.w6(32'h3cb0f443),
	.w7(32'h3b92b2d8),
	.w8(32'h3abf35a5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0c5b5),
	.w1(32'h3ba933f5),
	.w2(32'hb8fd7db5),
	.w3(32'h3c300fa7),
	.w4(32'h3be9cbe0),
	.w5(32'h3b1f6f19),
	.w6(32'h3b90ebe2),
	.w7(32'h3a41034e),
	.w8(32'h3afe2d29),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ad0a),
	.w1(32'hbb8bd035),
	.w2(32'hbc64f109),
	.w3(32'h3bce2a92),
	.w4(32'h3bbe607d),
	.w5(32'h3b6903ab),
	.w6(32'h3b23e754),
	.w7(32'h3b942684),
	.w8(32'hbc36dc2e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31aaee),
	.w1(32'hbad62542),
	.w2(32'h3aba01a0),
	.w3(32'h3b034c9e),
	.w4(32'h3b8f5d5a),
	.w5(32'h3b89cf47),
	.w6(32'hbb312f28),
	.w7(32'h399a51fb),
	.w8(32'h3b3aa47b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11e51e),
	.w1(32'hba01d484),
	.w2(32'hbb015a8a),
	.w3(32'h39d6a46d),
	.w4(32'hba51549d),
	.w5(32'h3a82fe8f),
	.w6(32'h3ac3fdbe),
	.w7(32'hba384d91),
	.w8(32'h3a8c6cb5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dfc0a),
	.w1(32'hbbae0191),
	.w2(32'hbc10d579),
	.w3(32'h3c806215),
	.w4(32'h3cf24b9d),
	.w5(32'h3cbc0e1f),
	.w6(32'h3c721de2),
	.w7(32'h3c23c69f),
	.w8(32'h3c0ee21b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc865522),
	.w1(32'h3c120cb4),
	.w2(32'h3c3b1bc8),
	.w3(32'h3c7487eb),
	.w4(32'h3c07824c),
	.w5(32'h3b81d728),
	.w6(32'h3a1bb765),
	.w7(32'hbc595876),
	.w8(32'hbbdb83ac),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae983a3),
	.w1(32'h3b91cc34),
	.w2(32'h3ccf5d7d),
	.w3(32'h3bae9a77),
	.w4(32'h3accb254),
	.w5(32'hbb5cd738),
	.w6(32'h3c2191de),
	.w7(32'h3c93db37),
	.w8(32'h3b8d2726),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e45f0),
	.w1(32'h3b6ba24f),
	.w2(32'hbc3b78bf),
	.w3(32'h3b0bcab9),
	.w4(32'hbb3ba8e6),
	.w5(32'hbc41d93e),
	.w6(32'hbc2089f1),
	.w7(32'hbc8947ee),
	.w8(32'hbbb736d6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9560ea),
	.w1(32'h3bc982ce),
	.w2(32'h3b2f4c92),
	.w3(32'h3b186f77),
	.w4(32'h3c58d057),
	.w5(32'h3c448b20),
	.w6(32'hba03cb10),
	.w7(32'h3c2b6fed),
	.w8(32'h3c585a44),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9959c25),
	.w1(32'hbb8ef71b),
	.w2(32'hbba30a1d),
	.w3(32'h3ada4477),
	.w4(32'h3925cafc),
	.w5(32'hb7a72c4b),
	.w6(32'h3aa2ecbc),
	.w7(32'hba1d5bf0),
	.w8(32'h38abdaad),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc9f66),
	.w1(32'h3c0a32af),
	.w2(32'h3bf1d00e),
	.w3(32'hbc011444),
	.w4(32'hbbbbd9bf),
	.w5(32'hb9b499ee),
	.w6(32'h3c0163cc),
	.w7(32'h3c4d1355),
	.w8(32'hba80e2b1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45ae1c),
	.w1(32'h38c784a6),
	.w2(32'hbb13eeb9),
	.w3(32'hbac20224),
	.w4(32'hbb4b049f),
	.w5(32'hbb880fd3),
	.w6(32'hbb22d7eb),
	.w7(32'hbb2ad2dc),
	.w8(32'hbbb38b57),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb09968),
	.w1(32'hbbb0543c),
	.w2(32'hbb2b5e07),
	.w3(32'hbb67ea33),
	.w4(32'hbb1dbf32),
	.w5(32'hbb35c4b2),
	.w6(32'hbb830ff0),
	.w7(32'hbb8d66e8),
	.w8(32'hbb6457a0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabeb2d),
	.w1(32'hbbb4d1d0),
	.w2(32'hbca66b16),
	.w3(32'h3c2b8e2c),
	.w4(32'h3c87992a),
	.w5(32'h3c08d84b),
	.w6(32'h3c8f23dd),
	.w7(32'hbae01cfc),
	.w8(32'hbc8ff643),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9881e),
	.w1(32'hbc80736e),
	.w2(32'hbc8d319a),
	.w3(32'hbc4bd4eb),
	.w4(32'hbc9e7568),
	.w5(32'hbc344585),
	.w6(32'hbc12a5e8),
	.w7(32'hbab3dd08),
	.w8(32'hbc009af2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc29f39),
	.w1(32'hba938edb),
	.w2(32'hb954eb40),
	.w3(32'h3b3da40f),
	.w4(32'h3a63080a),
	.w5(32'hbc4911de),
	.w6(32'hbbdd3fd6),
	.w7(32'hbb11af36),
	.w8(32'hbab5e4cb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a057d),
	.w1(32'hbaa18538),
	.w2(32'hbad2b46a),
	.w3(32'h3985a4a9),
	.w4(32'h3ad57321),
	.w5(32'h37ec0d6e),
	.w6(32'hba151ed6),
	.w7(32'hb815e3bc),
	.w8(32'hb9c0a7cf),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab71dc7),
	.w1(32'hbbe19799),
	.w2(32'hbc340a9e),
	.w3(32'hbaf52502),
	.w4(32'hbbd9a70f),
	.w5(32'hbba4a126),
	.w6(32'hbb8c6286),
	.w7(32'hbbd917b4),
	.w8(32'hbc111f53),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1dd92),
	.w1(32'h3b0c6178),
	.w2(32'h3b691c4e),
	.w3(32'h3c1b17e4),
	.w4(32'h3b18f856),
	.w5(32'hbb09fc1b),
	.w6(32'h3b17f5ef),
	.w7(32'hbaa740ed),
	.w8(32'hbb44092d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2172d2),
	.w1(32'hbb8d5784),
	.w2(32'hbb859698),
	.w3(32'hbb43df28),
	.w4(32'hbbb78a22),
	.w5(32'hbb143a4c),
	.w6(32'hbaa26596),
	.w7(32'hbb21456b),
	.w8(32'hba9d8c89),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8515d0a),
	.w1(32'hbc95f606),
	.w2(32'hbcdcd66c),
	.w3(32'h3cd9fc34),
	.w4(32'h3cc33dad),
	.w5(32'h3c8565fe),
	.w6(32'h3ca03046),
	.w7(32'h3b8f5500),
	.w8(32'hbc8ffdb1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ec6ed),
	.w1(32'hbb042cbf),
	.w2(32'h3a34d16e),
	.w3(32'hbb24a6d6),
	.w4(32'h3b62e2df),
	.w5(32'h3af006e9),
	.w6(32'hbb915aae),
	.w7(32'hbab35266),
	.w8(32'hbad36740),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43feb5),
	.w1(32'h3c5d40a0),
	.w2(32'h3c13ac22),
	.w3(32'h3c799532),
	.w4(32'h3c458885),
	.w5(32'h3be1248c),
	.w6(32'h3b98a45d),
	.w7(32'h3b8318eb),
	.w8(32'h3c60b275),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ba6a),
	.w1(32'hbc1193de),
	.w2(32'hbbdb98fe),
	.w3(32'hbbfd4aed),
	.w4(32'hbc10799e),
	.w5(32'hbbe43bb2),
	.w6(32'hbbc932bc),
	.w7(32'hbbe3d80d),
	.w8(32'hbb913aa2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d4abb),
	.w1(32'hb798e39e),
	.w2(32'h3b77c5de),
	.w3(32'h3b786f20),
	.w4(32'h3a9c74e8),
	.w5(32'h3be0fc5f),
	.w6(32'h3a84ee71),
	.w7(32'h3c10b631),
	.w8(32'h3c4e23a2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5a4a0),
	.w1(32'h3b8e6775),
	.w2(32'h3aec3ccd),
	.w3(32'h3bd0ed7d),
	.w4(32'h3bf88b7d),
	.w5(32'h3baabfd0),
	.w6(32'h3bc4c2a8),
	.w7(32'h3b94fc1a),
	.w8(32'h3baac621),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4686d5),
	.w1(32'h392781ff),
	.w2(32'h3ac74902),
	.w3(32'hba89082d),
	.w4(32'hbae80385),
	.w5(32'hbb2d9884),
	.w6(32'hb8956697),
	.w7(32'hb89b5c47),
	.w8(32'h3abc2f37),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb5348),
	.w1(32'hbb66cf88),
	.w2(32'hbb936ce2),
	.w3(32'hbac40f88),
	.w4(32'h38ec09a6),
	.w5(32'h3b4d82bc),
	.w6(32'hba542eb0),
	.w7(32'hbae1a20c),
	.w8(32'h3b20c26a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b577b),
	.w1(32'hbc2609c3),
	.w2(32'hbbe625af),
	.w3(32'hbb4afe41),
	.w4(32'h3b1f30b3),
	.w5(32'h3b938666),
	.w6(32'hbb5282ae),
	.w7(32'hbb09a59e),
	.w8(32'h3b3da887),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b370acc),
	.w1(32'hbacac47c),
	.w2(32'hbba83554),
	.w3(32'hb9c040f4),
	.w4(32'h3a56c8cc),
	.w5(32'hbb00e926),
	.w6(32'hb9b30139),
	.w7(32'hbb0c4aad),
	.w8(32'hbb2000a3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a720df1),
	.w1(32'h3b6b1a8b),
	.w2(32'h3bd0706a),
	.w3(32'h3ba708fb),
	.w4(32'h3afc8892),
	.w5(32'h3a7f26c1),
	.w6(32'h3ba87ea3),
	.w7(32'h3b5865ff),
	.w8(32'h3b55d84c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7104d),
	.w1(32'hba7881cd),
	.w2(32'hbb23df8d),
	.w3(32'hbafb992f),
	.w4(32'hbb799907),
	.w5(32'hbb444523),
	.w6(32'hba098cb1),
	.w7(32'hbadc6260),
	.w8(32'hbb0e8f50),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c827b),
	.w1(32'hbc3059d8),
	.w2(32'hbc153848),
	.w3(32'hbc3762bf),
	.w4(32'hbc2610a2),
	.w5(32'hbc4f05c5),
	.w6(32'hbc1fa9ec),
	.w7(32'hbc1f6cec),
	.w8(32'hbc4099db),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b39b0),
	.w1(32'hbb643b0f),
	.w2(32'hb98ada33),
	.w3(32'hba923e66),
	.w4(32'h395eecac),
	.w5(32'hb963142d),
	.w6(32'h397a793d),
	.w7(32'hba21e1ee),
	.w8(32'hbb1b3c1e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe26287),
	.w1(32'hbbdb2027),
	.w2(32'hbb89b5a8),
	.w3(32'h389f355e),
	.w4(32'hbaff91be),
	.w5(32'hbaef628b),
	.w6(32'hba8ffa57),
	.w7(32'hbb00e368),
	.w8(32'hbab563d6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0367c2),
	.w1(32'h3bd2ddea),
	.w2(32'h3c012854),
	.w3(32'h3b8399f6),
	.w4(32'h3b350d35),
	.w5(32'h3bbb103f),
	.w6(32'h3af7c777),
	.w7(32'h3b5b4c85),
	.w8(32'h3ba974fd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b265d1e),
	.w1(32'hbb3feda6),
	.w2(32'h3aa710cd),
	.w3(32'h3ada8755),
	.w4(32'h3b0e18fc),
	.w5(32'hba95922b),
	.w6(32'h3ba80db3),
	.w7(32'h3bbdb190),
	.w8(32'h3a9f1b4a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca25c28),
	.w1(32'hbb929e92),
	.w2(32'hbae980a4),
	.w3(32'h3ceaa719),
	.w4(32'h3cc7782a),
	.w5(32'h3cbe57d7),
	.w6(32'h3cbb060b),
	.w7(32'h3cec379e),
	.w8(32'h3cfc3839),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bfc63),
	.w1(32'h39b54809),
	.w2(32'h3aef4500),
	.w3(32'h3c14560d),
	.w4(32'h3c28a6c0),
	.w5(32'h3c2ad493),
	.w6(32'h3bb9b514),
	.w7(32'h3be610f0),
	.w8(32'h3be6692d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule