module layer_6_featuremap_73(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32a26d),
	.w1(32'hbc35c7e0),
	.w2(32'hbba54149),
	.w3(32'hbbbee891),
	.w4(32'hba84d865),
	.w5(32'h3adf5735),
	.w6(32'hbb9e368e),
	.w7(32'h3be8cd02),
	.w8(32'h3c739aaf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147848),
	.w1(32'h3bead7a4),
	.w2(32'h3b85da4e),
	.w3(32'hba8c643d),
	.w4(32'h3a00da9d),
	.w5(32'h3b13dcd5),
	.w6(32'h39bd04a9),
	.w7(32'hbc08e7f8),
	.w8(32'hbc84f45a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c84ff),
	.w1(32'hbbf2344b),
	.w2(32'h3bd11393),
	.w3(32'h3bc5d6b3),
	.w4(32'h3bbfd772),
	.w5(32'hbbbfdcfc),
	.w6(32'h3cddd350),
	.w7(32'h3ca1c97c),
	.w8(32'hbc8e3a22),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff1abc),
	.w1(32'h3c326450),
	.w2(32'h3c7399b2),
	.w3(32'hbb787f2f),
	.w4(32'h3a808bdd),
	.w5(32'h3c20ca3b),
	.w6(32'h385a6a8b),
	.w7(32'hbb271ade),
	.w8(32'hba17dfaf),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccd69a),
	.w1(32'h3c3f4c98),
	.w2(32'hbc251e4e),
	.w3(32'h3990a41b),
	.w4(32'hbc4bcb22),
	.w5(32'hbc2fe029),
	.w6(32'h3c657ec1),
	.w7(32'hbbbbc345),
	.w8(32'hbc1696f7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc77e01),
	.w1(32'hba3f1032),
	.w2(32'h3bb1dc8c),
	.w3(32'h3a0a98c3),
	.w4(32'h3bb5debf),
	.w5(32'h3bec961f),
	.w6(32'h3b32003e),
	.w7(32'h3c29112a),
	.w8(32'h3c79e504),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c815a78),
	.w1(32'h3bf55de1),
	.w2(32'hbc055e5c),
	.w3(32'h3b95fedc),
	.w4(32'hbc5dbdd5),
	.w5(32'hbc83452e),
	.w6(32'h3b918948),
	.w7(32'hbc67327c),
	.w8(32'hbca061b6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc343b99),
	.w1(32'h3c0bfe69),
	.w2(32'hbc4a9763),
	.w3(32'h3b93c90e),
	.w4(32'hbbbf9036),
	.w5(32'hbb238e01),
	.w6(32'h3c148f7a),
	.w7(32'h3bf51d0c),
	.w8(32'h3b258d91),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3077d4),
	.w1(32'hbbe04d63),
	.w2(32'hbc16c808),
	.w3(32'hbc0cecd2),
	.w4(32'hbc26261c),
	.w5(32'h3b391d71),
	.w6(32'h3ca7ed57),
	.w7(32'hbc29b9bf),
	.w8(32'hbcdebc3d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe446b3),
	.w1(32'hbbcc3395),
	.w2(32'hbb8ec394),
	.w3(32'hbac6a432),
	.w4(32'hba31829d),
	.w5(32'h3b91624f),
	.w6(32'h3b086ff1),
	.w7(32'h3b492007),
	.w8(32'h3c0d3912),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86ba51),
	.w1(32'hbca71942),
	.w2(32'hbc79aed1),
	.w3(32'hbc4c1d0f),
	.w4(32'hbcd559cd),
	.w5(32'hbcf8e260),
	.w6(32'hbb7f35f1),
	.w7(32'hbc76ce32),
	.w8(32'hbce21ee7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b302240),
	.w1(32'hbc1876c9),
	.w2(32'hbbb722da),
	.w3(32'h3b2dad78),
	.w4(32'h3b611fba),
	.w5(32'h3d0b0d80),
	.w6(32'hbb313933),
	.w7(32'hbaebf5d5),
	.w8(32'h3d03ea5a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c982eb0),
	.w1(32'h3acb42b2),
	.w2(32'hbc3e8722),
	.w3(32'h39ce64c7),
	.w4(32'hbc39506a),
	.w5(32'hbaffc6da),
	.w6(32'h3bb4fdb6),
	.w7(32'hbc1b6374),
	.w8(32'hbb322761),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79ba5f),
	.w1(32'hbc1bbfb1),
	.w2(32'hbb060d75),
	.w3(32'h3c1245c1),
	.w4(32'hbbeda780),
	.w5(32'hbc0aecd3),
	.w6(32'h3cda87a0),
	.w7(32'hbc470808),
	.w8(32'hbc900070),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c7aff),
	.w1(32'hbae365dd),
	.w2(32'h3b2f4e64),
	.w3(32'hba9f6172),
	.w4(32'h3b64cf20),
	.w5(32'h3c193238),
	.w6(32'hbb2cea50),
	.w7(32'h3b4e9b57),
	.w8(32'h3bdb9ce2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4300dc),
	.w1(32'hbc486982),
	.w2(32'hbba9c7b6),
	.w3(32'hbc2f8bca),
	.w4(32'hbc1747a2),
	.w5(32'hbb19d40b),
	.w6(32'hbba6f292),
	.w7(32'hbb855151),
	.w8(32'hb9af17e1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf70f87),
	.w1(32'h3af72a8f),
	.w2(32'h3c9bf2ba),
	.w3(32'h3c322fb2),
	.w4(32'h3ae852bb),
	.w5(32'h3bcc60b9),
	.w6(32'h3cf2dfb0),
	.w7(32'h3c3d6e25),
	.w8(32'hbbb207e9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53b3a5),
	.w1(32'hbbf4fb1e),
	.w2(32'hbad27223),
	.w3(32'hbbb82c36),
	.w4(32'hbb006f50),
	.w5(32'h3b4395bd),
	.w6(32'hbb57712e),
	.w7(32'h3b28a114),
	.w8(32'h3bdbd7cf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09e929),
	.w1(32'h3a1e86ac),
	.w2(32'h3b7975cb),
	.w3(32'hbb892f9a),
	.w4(32'hbb657680),
	.w5(32'hbb780d44),
	.w6(32'h3b1260b3),
	.w7(32'h3b58702a),
	.w8(32'h3b2f765d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78cd58),
	.w1(32'hbc14e355),
	.w2(32'hbb57d63b),
	.w3(32'hbba7c742),
	.w4(32'h3a85cfcb),
	.w5(32'h3c14a489),
	.w6(32'h3af45761),
	.w7(32'h3ab87c6f),
	.w8(32'h3c13c1ad),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b310967),
	.w1(32'hbb000e6d),
	.w2(32'hba89a6b2),
	.w3(32'hbbcca0e8),
	.w4(32'hbbb46b0f),
	.w5(32'hbba0ec4a),
	.w6(32'hbc04689c),
	.w7(32'hbc0c01f0),
	.w8(32'hbb9d4bc7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9aedd0),
	.w1(32'hbc78a7e8),
	.w2(32'hba1e2b43),
	.w3(32'hbc6663ad),
	.w4(32'hbcdd04d1),
	.w5(32'hbc604042),
	.w6(32'h3bda26a7),
	.w7(32'hbc014809),
	.w8(32'hbcc69975),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f58b9),
	.w1(32'h3c5f0b4d),
	.w2(32'h3cb218f6),
	.w3(32'hba8634a7),
	.w4(32'h3bf7e899),
	.w5(32'h3c3a6b50),
	.w6(32'h3c4f04b0),
	.w7(32'h3caea3a5),
	.w8(32'h3cd90a04),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc835d47),
	.w1(32'hbd2efa74),
	.w2(32'hbcba07e5),
	.w3(32'hbca57ff3),
	.w4(32'hbd407dee),
	.w5(32'hbd3e159f),
	.w6(32'hbb8798c3),
	.w7(32'hbc568413),
	.w8(32'hbd3e600e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bd23e),
	.w1(32'h3c4bfcaa),
	.w2(32'h3c8acd22),
	.w3(32'hbc09333e),
	.w4(32'h3b188353),
	.w5(32'h3cccf846),
	.w6(32'h3c77f96b),
	.w7(32'hbbccbcd4),
	.w8(32'hbb9bbbf4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccac57d),
	.w1(32'hbc96d283),
	.w2(32'hbc581d0b),
	.w3(32'hbc876c16),
	.w4(32'hbc8bbd33),
	.w5(32'hbb1848ea),
	.w6(32'h3b140d76),
	.w7(32'hbc14502c),
	.w8(32'hbc2606de),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadcb2b),
	.w1(32'hbcdcb703),
	.w2(32'hbc2336f8),
	.w3(32'hbaf0e45d),
	.w4(32'hbc95da66),
	.w5(32'hbcc6ce12),
	.w6(32'h3ad076e4),
	.w7(32'h3bf4dcf9),
	.w8(32'hbb8b887c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fc30b),
	.w1(32'hba8c91ca),
	.w2(32'hbc2c1ac0),
	.w3(32'hbc01699a),
	.w4(32'hbca4961c),
	.w5(32'hbcab99d5),
	.w6(32'h3b7d4850),
	.w7(32'hbc7337e3),
	.w8(32'hbccb2338),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc443e9b),
	.w1(32'hbb9d5ced),
	.w2(32'hbb7244db),
	.w3(32'hbb599355),
	.w4(32'hbb287a83),
	.w5(32'hbb12df47),
	.w6(32'hbbb1e8bb),
	.w7(32'hbbb4e9db),
	.w8(32'hbbc7fdf9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc084372),
	.w1(32'hbc0086d8),
	.w2(32'hbc88650d),
	.w3(32'hbcc49aaa),
	.w4(32'h3cd05550),
	.w5(32'h3c12d11f),
	.w6(32'hbce33e5b),
	.w7(32'h3c7b5f2e),
	.w8(32'h3c708ae2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffe1a5),
	.w1(32'hbb96f2b5),
	.w2(32'hbbed8afd),
	.w3(32'hbb845780),
	.w4(32'hbb220ef9),
	.w5(32'h3bca6292),
	.w6(32'h3b8c065d),
	.w7(32'h3aa80b30),
	.w8(32'h3b328dc6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b435f),
	.w1(32'hbc322c9f),
	.w2(32'hbc01f016),
	.w3(32'hbc1c365e),
	.w4(32'hbcaef192),
	.w5(32'hbc7778f8),
	.w6(32'hbcacee03),
	.w7(32'hbcae25b8),
	.w8(32'hbc5abcce),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5855b),
	.w1(32'hbbbc7420),
	.w2(32'hbbae0fe3),
	.w3(32'hbc1099ef),
	.w4(32'hbbba7a40),
	.w5(32'hbb4fd83f),
	.w6(32'hbbbe38a2),
	.w7(32'hbbb9f635),
	.w8(32'hbc2b2a18),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963ffae),
	.w1(32'hbb937f56),
	.w2(32'hbbfc31b6),
	.w3(32'hbb1e3444),
	.w4(32'hbb32b22b),
	.w5(32'h3b018efd),
	.w6(32'hbb469e9d),
	.w7(32'h3b214de9),
	.w8(32'h3bde0998),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89dd17),
	.w1(32'hbbad1d03),
	.w2(32'h3a655408),
	.w3(32'hbb8bbf5e),
	.w4(32'h3b6b5551),
	.w5(32'h3be16a71),
	.w6(32'hbbd9bda3),
	.w7(32'h3b453900),
	.w8(32'h3c093f7e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f899b),
	.w1(32'h3bb4c631),
	.w2(32'hbb157843),
	.w3(32'hbc104389),
	.w4(32'h3c01386e),
	.w5(32'h3cb4e927),
	.w6(32'h3ad35c3f),
	.w7(32'h3a90978b),
	.w8(32'h3c3ccd39),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a9c1d),
	.w1(32'hbc481589),
	.w2(32'hbc0f070f),
	.w3(32'hbc2fc63c),
	.w4(32'hbc01433b),
	.w5(32'hbb463a51),
	.w6(32'hbc0f4ace),
	.w7(32'hbb685696),
	.w8(32'h3c0d4f09),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc926c),
	.w1(32'h3b598868),
	.w2(32'hb99617b6),
	.w3(32'hbb1d2b96),
	.w4(32'hb9d4f3ec),
	.w5(32'h3b354ca4),
	.w6(32'h3b2c7eba),
	.w7(32'hbb93e32f),
	.w8(32'hbb539e05),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa7ba9),
	.w1(32'hba01f03c),
	.w2(32'hbbe2c4c5),
	.w3(32'hbbbfc1c4),
	.w4(32'hbb6d91aa),
	.w5(32'hbbd8fd8f),
	.w6(32'h3b991f15),
	.w7(32'hbc2be74f),
	.w8(32'hbbc28720),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb81705),
	.w1(32'hbcac91fe),
	.w2(32'h3c3a2c2b),
	.w3(32'hbc59b982),
	.w4(32'hbd4595c8),
	.w5(32'hbd1908be),
	.w6(32'h3cbf0642),
	.w7(32'hbcb0eb49),
	.w8(32'hbd69234f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a09ea),
	.w1(32'hbb9e451c),
	.w2(32'hbb905b88),
	.w3(32'hbadb62b9),
	.w4(32'h3a02139d),
	.w5(32'h3bfd3e06),
	.w6(32'h3b8f5143),
	.w7(32'hbc2212fc),
	.w8(32'h3bb49be3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c1b32),
	.w1(32'hb90e2a88),
	.w2(32'h3b348b4a),
	.w3(32'hbc2615b7),
	.w4(32'hbb8112ee),
	.w5(32'h39cfdc9d),
	.w6(32'hbbfd54bf),
	.w7(32'hbc17a6c9),
	.w8(32'hbba2efdd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb117ff1),
	.w1(32'hbbd4a009),
	.w2(32'h3bfc8e07),
	.w3(32'hbb86870f),
	.w4(32'h3bcbc344),
	.w5(32'h3c7b77c7),
	.w6(32'hbc0f3791),
	.w7(32'h3bfe24bc),
	.w8(32'h3cba68f0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4a4236),
	.w1(32'h3ca54731),
	.w2(32'h3c894083),
	.w3(32'h3b8ed894),
	.w4(32'h3d37c526),
	.w5(32'h3d5618f4),
	.w6(32'h3b33e459),
	.w7(32'h3c203142),
	.w8(32'h3cd34a25),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f4d96),
	.w1(32'hbc88a6a4),
	.w2(32'hbacabb68),
	.w3(32'hbb2a1b81),
	.w4(32'hbccab20c),
	.w5(32'hbc991b9a),
	.w6(32'h3c2368c6),
	.w7(32'hbbd74e65),
	.w8(32'hbcba5240),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb6b47),
	.w1(32'hb87431d0),
	.w2(32'hbc25d79a),
	.w3(32'hbb12aa23),
	.w4(32'hbc52776f),
	.w5(32'hbc8e8da2),
	.w6(32'h3bf07a0a),
	.w7(32'hbc624a1b),
	.w8(32'hbc21db15),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc216843),
	.w1(32'h3ca538f2),
	.w2(32'h3c7182f6),
	.w3(32'h3b0f8618),
	.w4(32'h39c3d680),
	.w5(32'h3c06adb7),
	.w6(32'h3c0a5cb1),
	.w7(32'h3a39a7ec),
	.w8(32'hbb4939c3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdbab63),
	.w1(32'hbbd2b1a5),
	.w2(32'hbb690585),
	.w3(32'hbbd43df1),
	.w4(32'hbb9aba18),
	.w5(32'hbbf42070),
	.w6(32'hbc033b9d),
	.w7(32'hbc006e1d),
	.w8(32'h3aa7cb0f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe849a),
	.w1(32'h3a051daf),
	.w2(32'h3b99b245),
	.w3(32'hbc0568b5),
	.w4(32'hbbb905f2),
	.w5(32'h3a258abd),
	.w6(32'hbba50178),
	.w7(32'hbb0e11fb),
	.w8(32'h3b348b44),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38c654),
	.w1(32'h3bfa60f1),
	.w2(32'hbc3626a9),
	.w3(32'hba88773e),
	.w4(32'hbbb73cb5),
	.w5(32'hbca6e509),
	.w6(32'hbb991cb2),
	.w7(32'hbbf6a68d),
	.w8(32'hbc29f8a0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc203090),
	.w1(32'hbc081cc9),
	.w2(32'hbb7ef31e),
	.w3(32'hbc813318),
	.w4(32'hbc55be27),
	.w5(32'hbc025f82),
	.w6(32'hbc185301),
	.w7(32'hbc7c751d),
	.w8(32'hbc89bc87),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc897fa9),
	.w1(32'hbc26a741),
	.w2(32'hbbdb5167),
	.w3(32'hbca9719f),
	.w4(32'hbcb654a0),
	.w5(32'hbc98f9aa),
	.w6(32'hbc009a22),
	.w7(32'hbc957338),
	.w8(32'hbc8df62c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2079e7),
	.w1(32'hbc88918a),
	.w2(32'hbb0e77ce),
	.w3(32'hbc906aa4),
	.w4(32'hbd1cb855),
	.w5(32'hbd17f016),
	.w6(32'h3c6d3eb5),
	.w7(32'hbc96c220),
	.w8(32'hbd1e8d3b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5ba2f),
	.w1(32'h3c8ba7cc),
	.w2(32'hbb3ffbda),
	.w3(32'h3b737223),
	.w4(32'hbc44d4ae),
	.w5(32'hbcbda614),
	.w6(32'h3c0bc4a1),
	.w7(32'hbb2d5671),
	.w8(32'hbc2675bb),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6426a),
	.w1(32'hbbad3823),
	.w2(32'hbb863f36),
	.w3(32'hbb286018),
	.w4(32'hbbd7150c),
	.w5(32'hbb8f87b8),
	.w6(32'h3b118cb3),
	.w7(32'h3a00dd8b),
	.w8(32'hbb8679e0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35d33f),
	.w1(32'h3ce108c4),
	.w2(32'h3d087f2f),
	.w3(32'h3a686089),
	.w4(32'hba1d7124),
	.w5(32'h3d0165d0),
	.w6(32'h3b8b9822),
	.w7(32'hbc34d6a9),
	.w8(32'h3ca4e84a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3f302),
	.w1(32'hbc9776b3),
	.w2(32'hbc4ae557),
	.w3(32'hbc875909),
	.w4(32'hbcb05dd1),
	.w5(32'hbc9fee07),
	.w6(32'hbc58fe0e),
	.w7(32'hbc91b87d),
	.w8(32'hbc851872),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7da9cf),
	.w1(32'hbc9e9d8a),
	.w2(32'hbb98d155),
	.w3(32'hbc833c88),
	.w4(32'hbbc66488),
	.w5(32'hbc43b9fd),
	.w6(32'hbcc61844),
	.w7(32'h38951255),
	.w8(32'hbc568a7f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919f87a),
	.w1(32'h3a97bf8c),
	.w2(32'hba8bb0a1),
	.w3(32'h3b66fa02),
	.w4(32'hb979c819),
	.w5(32'hba955732),
	.w6(32'h3ba03f8c),
	.w7(32'h39870a13),
	.w8(32'hbaf8484d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba374b1b),
	.w1(32'hbc92379d),
	.w2(32'h3d228464),
	.w3(32'h3c2865c0),
	.w4(32'h3c894af7),
	.w5(32'h3ccafcfa),
	.w6(32'h3ce0037e),
	.w7(32'h3c8aa91b),
	.w8(32'h3b7dafd0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41e050),
	.w1(32'hbc5237cb),
	.w2(32'hbca281b4),
	.w3(32'hbba7533d),
	.w4(32'hbc19acd8),
	.w5(32'hbbe22f1a),
	.w6(32'hba062289),
	.w7(32'hbc8347a9),
	.w8(32'h3b0ee9f7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfd59a),
	.w1(32'h3c0354e0),
	.w2(32'h3d749427),
	.w3(32'hbcc63744),
	.w4(32'h3d432c6a),
	.w5(32'hbbefd9b5),
	.w6(32'h3c5c4175),
	.w7(32'h3d8eda22),
	.w8(32'hb91baebb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d266766),
	.w1(32'hbc9307b6),
	.w2(32'hbce28e17),
	.w3(32'hbce78108),
	.w4(32'h3d12c4ca),
	.w5(32'h3ba85c81),
	.w6(32'hbd7158ae),
	.w7(32'h3be291be),
	.w8(32'h3c9635bc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c028fae),
	.w1(32'hbca452de),
	.w2(32'hbc7eba20),
	.w3(32'hbc6eb34f),
	.w4(32'hbbff6151),
	.w5(32'hbc9b3543),
	.w6(32'hbc85d852),
	.w7(32'hbb74a6c1),
	.w8(32'hbc611ed5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule