module layer_8_featuremap_142(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bebc1),
	.w1(32'h396cdd7d),
	.w2(32'h3a1faf48),
	.w3(32'h3b90f119),
	.w4(32'h3b8c2547),
	.w5(32'h3b5fc18b),
	.w6(32'h3c0d12e2),
	.w7(32'hb95a3763),
	.w8(32'hba25d859),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0613d),
	.w1(32'h3b91114e),
	.w2(32'hbb33298e),
	.w3(32'h3b96af61),
	.w4(32'hbb42b8a2),
	.w5(32'hbb7a837c),
	.w6(32'hb96b52de),
	.w7(32'hbb1a65aa),
	.w8(32'hbbb6fd44),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc201b9e),
	.w1(32'hbc0c829a),
	.w2(32'h3a4d4b29),
	.w3(32'hbbec480f),
	.w4(32'hbbbcdd61),
	.w5(32'hbc16c6b4),
	.w6(32'hbc224aa1),
	.w7(32'h3b441abe),
	.w8(32'hbbc2b6eb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb6fbb),
	.w1(32'hbba469ee),
	.w2(32'hbbaa1be5),
	.w3(32'hbc0c1b72),
	.w4(32'hbb17aea5),
	.w5(32'h3a9850db),
	.w6(32'hbbe2e35f),
	.w7(32'hbc37f273),
	.w8(32'hbb19471e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e8952),
	.w1(32'h3c6210b7),
	.w2(32'hbb6d38b5),
	.w3(32'hbb35fd52),
	.w4(32'hbba81ce1),
	.w5(32'hbb45f922),
	.w6(32'h3a9eae49),
	.w7(32'hbb13e3b7),
	.w8(32'h39c0ede9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba75765),
	.w1(32'hb9b11361),
	.w2(32'hbb72debc),
	.w3(32'hbbb612d6),
	.w4(32'hbc08f11a),
	.w5(32'h3a84eca9),
	.w6(32'hbbc44eca),
	.w7(32'hbbea0db5),
	.w8(32'hb8e5883c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e0065),
	.w1(32'hbbb54ab0),
	.w2(32'h3ab34271),
	.w3(32'hbb27516b),
	.w4(32'hbb3a3eb8),
	.w5(32'hbb5818ad),
	.w6(32'hbb718d26),
	.w7(32'hbb498145),
	.w8(32'hbb61cc9f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98fd98),
	.w1(32'hbb4aac12),
	.w2(32'h3a754200),
	.w3(32'hbbe4c3bf),
	.w4(32'hba96d621),
	.w5(32'h3a677f05),
	.w6(32'hbbcb6dea),
	.w7(32'hbad81bb6),
	.w8(32'hbb9342fc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5cb2),
	.w1(32'hbc1af5e3),
	.w2(32'hbae31a03),
	.w3(32'hb9a8b617),
	.w4(32'hbc05327f),
	.w5(32'hbbbe124c),
	.w6(32'hbb8bf33e),
	.w7(32'hbc979b6d),
	.w8(32'hbc7338e6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb975422f),
	.w1(32'hbb3dbbdd),
	.w2(32'hbbf01817),
	.w3(32'h3b9cc0c2),
	.w4(32'h3bed756c),
	.w5(32'hbac641fc),
	.w6(32'hbc03bce6),
	.w7(32'h3a9deeb8),
	.w8(32'h3b482c09),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd14c0a),
	.w1(32'hbc4ebeda),
	.w2(32'h3b9d7452),
	.w3(32'hbaddd303),
	.w4(32'hb92c9c9f),
	.w5(32'hbb4ad48b),
	.w6(32'h3b26bea8),
	.w7(32'h3b17a046),
	.w8(32'h3b1ef22a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c189d33),
	.w1(32'h3bb49c18),
	.w2(32'hbc0006b4),
	.w3(32'h3bbaf8af),
	.w4(32'hbba921aa),
	.w5(32'hbbb7cae5),
	.w6(32'h3b920edf),
	.w7(32'hbba91c18),
	.w8(32'hbc26f300),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fd4f9),
	.w1(32'hbc02d8c8),
	.w2(32'hbb870bf9),
	.w3(32'hbb7127e7),
	.w4(32'hba0bd3a6),
	.w5(32'hbabf3584),
	.w6(32'hbbbbe21e),
	.w7(32'hbc2958d6),
	.w8(32'h3bc1089e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdd48f),
	.w1(32'h39660b32),
	.w2(32'h3a03d909),
	.w3(32'h3a92bfe2),
	.w4(32'h3aa4cc31),
	.w5(32'hbb72f40a),
	.w6(32'h3bd1cfc9),
	.w7(32'hba0302dc),
	.w8(32'hbb58b782),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6cbde),
	.w1(32'hba1118e4),
	.w2(32'hbc0cebcf),
	.w3(32'hbb4c6f2c),
	.w4(32'hbba4e3c4),
	.w5(32'hbb9dc002),
	.w6(32'hbbaee07a),
	.w7(32'hbc0d6bb8),
	.w8(32'hbb95e0a7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8056d8),
	.w1(32'h3b3dd463),
	.w2(32'hbbc0d691),
	.w3(32'hb8918b57),
	.w4(32'h3c9ad061),
	.w5(32'h3b23aabc),
	.w6(32'h398c8f8f),
	.w7(32'h3a7f1564),
	.w8(32'hbad6c41e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e9577),
	.w1(32'hbc3e1ae0),
	.w2(32'hbb8aa785),
	.w3(32'hbb7ef96e),
	.w4(32'hbc152ef9),
	.w5(32'h3cd62f67),
	.w6(32'hbb3bda1e),
	.w7(32'h3ca73167),
	.w8(32'h3c2a9c2c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca69d0),
	.w1(32'hbae7e042),
	.w2(32'hbc393e8e),
	.w3(32'hbbfacffa),
	.w4(32'h3b82115b),
	.w5(32'hbc91ec41),
	.w6(32'hbca1d60d),
	.w7(32'hbc2e82ea),
	.w8(32'h3cd4a037),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd608c1),
	.w1(32'h3bc58b04),
	.w2(32'hbc58c441),
	.w3(32'h3c258ab5),
	.w4(32'hbb50c048),
	.w5(32'hbc194ebe),
	.w6(32'hbb3de7cf),
	.w7(32'hbb950608),
	.w8(32'hbcf9287c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4580b4),
	.w1(32'h3adc75c1),
	.w2(32'hbc0cb550),
	.w3(32'hbaa6a81f),
	.w4(32'h3cb06390),
	.w5(32'h3b91b6f4),
	.w6(32'hbc055358),
	.w7(32'hbaeaa4ed),
	.w8(32'hbce4d05b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c8a1a),
	.w1(32'h3b80bc15),
	.w2(32'h39145c30),
	.w3(32'hbc08e860),
	.w4(32'h3c8e75e2),
	.w5(32'h3c6a5746),
	.w6(32'hbb4afd40),
	.w7(32'h3d17c7e8),
	.w8(32'hbc545f9a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce5095b),
	.w1(32'hbc50406d),
	.w2(32'hba10d8b9),
	.w3(32'hbca93fd8),
	.w4(32'hbbd88672),
	.w5(32'hbb605a3d),
	.w6(32'hbd05d9f1),
	.w7(32'hbb015e27),
	.w8(32'hbc955f2a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca17ffc),
	.w1(32'hbc08db99),
	.w2(32'hbcad5cf3),
	.w3(32'h3bd27410),
	.w4(32'hbc4386d0),
	.w5(32'hbd0416dc),
	.w6(32'h3c86c314),
	.w7(32'hbcc3ff2a),
	.w8(32'hbd0889ef),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72caab),
	.w1(32'h3c0ac151),
	.w2(32'hbb599a69),
	.w3(32'hbbf588e3),
	.w4(32'h3c145059),
	.w5(32'hbcb42b26),
	.w6(32'h3c6b1dc9),
	.w7(32'h3a0a01b2),
	.w8(32'hbb6827cc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3c503),
	.w1(32'hbb88ca72),
	.w2(32'hbb8b5820),
	.w3(32'hbbd2d820),
	.w4(32'hbb2827cd),
	.w5(32'hbc12bf1d),
	.w6(32'h39838cc9),
	.w7(32'hbb4b3a26),
	.w8(32'hbb7d04ee),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be81604),
	.w1(32'h3ce21e09),
	.w2(32'h3936f5bb),
	.w3(32'h3c69a247),
	.w4(32'h3cc42037),
	.w5(32'h3c477840),
	.w6(32'h3ce694a8),
	.w7(32'h3d1e365a),
	.w8(32'hbc8bea92),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3f5014),
	.w1(32'h3baacc4f),
	.w2(32'hbb651595),
	.w3(32'hbb0cf669),
	.w4(32'hbc92d1ce),
	.w5(32'h3c7e5a4b),
	.w6(32'hbcaa9a5e),
	.w7(32'h3b8cfc26),
	.w8(32'h3c358f8a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb46e5d),
	.w1(32'h3afe4ed9),
	.w2(32'h3c9b957a),
	.w3(32'hbad00a70),
	.w4(32'h3c11c8fa),
	.w5(32'hbbbee8cf),
	.w6(32'hbc673e4f),
	.w7(32'h3ca7ab23),
	.w8(32'hbce21d03),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ad330),
	.w1(32'hbce53d54),
	.w2(32'hbafbc6a9),
	.w3(32'hbcc71cbb),
	.w4(32'h3c5677fd),
	.w5(32'hbc7718b4),
	.w6(32'hbcc82129),
	.w7(32'hbc89c473),
	.w8(32'hbc29d34d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03725e),
	.w1(32'hbb7ad17d),
	.w2(32'h3c70ebde),
	.w3(32'hbc3d75de),
	.w4(32'hbc35869f),
	.w5(32'h3c95edb8),
	.w6(32'hbbe52299),
	.w7(32'hbccfd54a),
	.w8(32'h3d8d54f7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e3a38),
	.w1(32'hbce966d4),
	.w2(32'h3ba8d40c),
	.w3(32'h3c765ead),
	.w4(32'h3c1b1755),
	.w5(32'h3c1e9bbb),
	.w6(32'hbc83f3be),
	.w7(32'h3b3eb910),
	.w8(32'h3addb44c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90ad5a),
	.w1(32'h3b606a7c),
	.w2(32'hbb8705ba),
	.w3(32'h3bfc4128),
	.w4(32'h3c314f11),
	.w5(32'h3be1ca49),
	.w6(32'h3b17f3eb),
	.w7(32'hbceac459),
	.w8(32'h3c7af8db),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22df57),
	.w1(32'hbc8d6b55),
	.w2(32'hbcbe92c2),
	.w3(32'hbb47a8cf),
	.w4(32'hbccaad71),
	.w5(32'h3c6d96ab),
	.w6(32'h3c966a6c),
	.w7(32'hbcab2c14),
	.w8(32'h3a9d628f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb101e1),
	.w1(32'h3ce034d1),
	.w2(32'hba187b07),
	.w3(32'h3bad80d0),
	.w4(32'hba382d60),
	.w5(32'h3c958204),
	.w6(32'h3cac10b7),
	.w7(32'h3c8636ef),
	.w8(32'h3d3e070f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd03a3f0),
	.w1(32'hbc4f7618),
	.w2(32'h3c265f5a),
	.w3(32'h3b992f13),
	.w4(32'h3c153672),
	.w5(32'h3c1df0cf),
	.w6(32'hbc86088e),
	.w7(32'h3c28e97a),
	.w8(32'hbb84c5dc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf18d9),
	.w1(32'h3c95ff10),
	.w2(32'hbbcf9421),
	.w3(32'h3c82757c),
	.w4(32'hbccc31c7),
	.w5(32'hbcb35ef6),
	.w6(32'h3c9a4a1c),
	.w7(32'hbd313530),
	.w8(32'h3c38074e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1b35ae),
	.w1(32'h3bc21065),
	.w2(32'h3bd58bcb),
	.w3(32'h3c36b9b2),
	.w4(32'h3c050ff3),
	.w5(32'h3a6c9770),
	.w6(32'h3d5ac3c0),
	.w7(32'h3a9e00d2),
	.w8(32'hbc485fdc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c95c6),
	.w1(32'hbc2f0db1),
	.w2(32'hbbb0f637),
	.w3(32'h3bef75fd),
	.w4(32'h3bb5a1a2),
	.w5(32'hbc0c6184),
	.w6(32'hbc3134b7),
	.w7(32'hbb05054a),
	.w8(32'h3c47c86d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f0417),
	.w1(32'hbc6794fb),
	.w2(32'h3b294b40),
	.w3(32'hbc945ba8),
	.w4(32'hbbc6d93e),
	.w5(32'h3c87c1fc),
	.w6(32'hbc80213e),
	.w7(32'hbb905073),
	.w8(32'h3c041a1d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b964309),
	.w1(32'h3b7d74c4),
	.w2(32'hbb91fcba),
	.w3(32'h38b0e53e),
	.w4(32'hbb008a02),
	.w5(32'h3c569285),
	.w6(32'hbbce2776),
	.w7(32'h3c0322d4),
	.w8(32'h3c61a2df),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a959e),
	.w1(32'h3c8a2372),
	.w2(32'hba885b9e),
	.w3(32'h3ca14345),
	.w4(32'h3c892485),
	.w5(32'hbc20db4a),
	.w6(32'h3ca82496),
	.w7(32'hbb9daa75),
	.w8(32'hbc4b0c7d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbaad1b),
	.w1(32'h3c6ae3a1),
	.w2(32'h3a6e75fe),
	.w3(32'hbc180ae1),
	.w4(32'hba99b82f),
	.w5(32'hbb5070d3),
	.w6(32'hbcd333b8),
	.w7(32'h3af8611c),
	.w8(32'hbc2b6dcc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b836746),
	.w1(32'h3c80cdc1),
	.w2(32'h3b34badd),
	.w3(32'h3ba78261),
	.w4(32'hbc4323f2),
	.w5(32'hbc8a2073),
	.w6(32'hbbe5f028),
	.w7(32'hbc886211),
	.w8(32'h3a1786ce),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17d9d0),
	.w1(32'h3c243d52),
	.w2(32'hbbfbc83b),
	.w3(32'h3b62bdf5),
	.w4(32'h39066aa1),
	.w5(32'hbb016f86),
	.w6(32'h3d1529d6),
	.w7(32'hbc24cc19),
	.w8(32'h3bda6e30),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c485ab8),
	.w1(32'hba8a63a5),
	.w2(32'h3c4f3c28),
	.w3(32'h3b83d9f6),
	.w4(32'hbbe2f7f3),
	.w5(32'h3ba0014f),
	.w6(32'h3c17bd36),
	.w7(32'hb9f28a1d),
	.w8(32'h3bc0413d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bac58),
	.w1(32'hbb7a8f5d),
	.w2(32'hbb5c9ee6),
	.w3(32'hbbff0e6e),
	.w4(32'hbb870a81),
	.w5(32'hbcfa0d8b),
	.w6(32'h3a4ced4d),
	.w7(32'hbd2347c2),
	.w8(32'hb9600502),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3606d2),
	.w1(32'h3c2d55c6),
	.w2(32'hbc1098e6),
	.w3(32'h3bf7cdae),
	.w4(32'h3b593f3a),
	.w5(32'h3b4ecbc4),
	.w6(32'h3d58f86a),
	.w7(32'h3bdc0fa4),
	.w8(32'hbc406e76),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb47603),
	.w1(32'h3c19ae6f),
	.w2(32'h3c18acc7),
	.w3(32'hbc5351aa),
	.w4(32'h3c5cdfcb),
	.w5(32'hbbfdf74c),
	.w6(32'h3cab3d84),
	.w7(32'hbc01842f),
	.w8(32'hbbb2aec4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39837c),
	.w1(32'h3b8d106b),
	.w2(32'hb9a47210),
	.w3(32'hbc298c33),
	.w4(32'hbcb98fba),
	.w5(32'h3bf13fba),
	.w6(32'h3cb92072),
	.w7(32'h3c63b64d),
	.w8(32'h3ceab8f4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd226045),
	.w1(32'h3cfb927d),
	.w2(32'hbcf90ff5),
	.w3(32'hbb31a455),
	.w4(32'hbd199d76),
	.w5(32'hbc671fe0),
	.w6(32'hbcc4ee3b),
	.w7(32'hbc750459),
	.w8(32'h3c44a0f8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf17ee1),
	.w1(32'hbc779f02),
	.w2(32'h3a74b4ab),
	.w3(32'hbce10755),
	.w4(32'h3c676702),
	.w5(32'hbc95048f),
	.w6(32'hbcb776f4),
	.w7(32'h3c00006e),
	.w8(32'h3bda075f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d148287),
	.w1(32'hbc0323d6),
	.w2(32'h3b93e20f),
	.w3(32'hbc8d7dca),
	.w4(32'h3d049f01),
	.w5(32'h3cca58e9),
	.w6(32'hba7f18d8),
	.w7(32'h3d306ccc),
	.w8(32'hbcad9c71),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdbf84a),
	.w1(32'hbc8cd514),
	.w2(32'h3a632b22),
	.w3(32'hbbd7fab9),
	.w4(32'h3c25701a),
	.w5(32'h3be19b88),
	.w6(32'hbce13bf5),
	.w7(32'h3b9833b1),
	.w8(32'h3cc4488f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4509d4),
	.w1(32'hbc82e99b),
	.w2(32'hbbb55f17),
	.w3(32'hbbd1cc4a),
	.w4(32'hbaee4059),
	.w5(32'hbb3a7f7b),
	.w6(32'hbc8752d3),
	.w7(32'hbc18b976),
	.w8(32'h3b990da1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c3894),
	.w1(32'h3acf04ac),
	.w2(32'h3a33aafd),
	.w3(32'h3b4b678f),
	.w4(32'hbc14a8fe),
	.w5(32'h3c8274b1),
	.w6(32'h3bb64767),
	.w7(32'h3b876132),
	.w8(32'h3cb9e05b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2aeeb),
	.w1(32'hbca2d333),
	.w2(32'hbb9f73ee),
	.w3(32'h3cd59da4),
	.w4(32'hbbbf5b03),
	.w5(32'hbc8b0d23),
	.w6(32'hb93380c1),
	.w7(32'hbb8168b6),
	.w8(32'hbc7568d3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55b1a5),
	.w1(32'h3ac0b461),
	.w2(32'hbc71db8e),
	.w3(32'hbba21ea9),
	.w4(32'hbc72d0fd),
	.w5(32'hbbfaff46),
	.w6(32'h3bd8992c),
	.w7(32'hbc499619),
	.w8(32'h3b91d454),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf744),
	.w1(32'h3b0fe9f3),
	.w2(32'h3c53bf04),
	.w3(32'hbb5aacb1),
	.w4(32'h3cf94392),
	.w5(32'hbc473577),
	.w6(32'hbba5e2c4),
	.w7(32'h3c683a96),
	.w8(32'hbc613b71),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e9342),
	.w1(32'hbcbeed45),
	.w2(32'hbb8a3ab4),
	.w3(32'hbc9ad8e5),
	.w4(32'h3a18c71c),
	.w5(32'h3a4e0def),
	.w6(32'h3b392dcd),
	.w7(32'hbc0d4ac9),
	.w8(32'h3bfc628f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5548c8),
	.w1(32'h3a120e01),
	.w2(32'h3a35a96c),
	.w3(32'h3b528da2),
	.w4(32'h3c9c2b95),
	.w5(32'hbcb1c235),
	.w6(32'h3bc4969e),
	.w7(32'h3cd66b89),
	.w8(32'hbdad5775),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced1ed5),
	.w1(32'h3ce3b969),
	.w2(32'h3c62ea79),
	.w3(32'h3b6d0756),
	.w4(32'hbb9991c1),
	.w5(32'hbd251641),
	.w6(32'h3c404973),
	.w7(32'hbcaeb3cb),
	.w8(32'h3bfa1539),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd76586),
	.w1(32'h3c851e31),
	.w2(32'h3c02d0ea),
	.w3(32'hbb904cd7),
	.w4(32'hbb25c525),
	.w5(32'hba7711cd),
	.w6(32'h3cfb71bf),
	.w7(32'h3b5ed8d0),
	.w8(32'hbaaf2511),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05edb3),
	.w1(32'h3bc8e4cf),
	.w2(32'hbc2b774e),
	.w3(32'hb950637f),
	.w4(32'hba0cebe1),
	.w5(32'h3a8564b3),
	.w6(32'h39cec017),
	.w7(32'h3b8c6995),
	.w8(32'hbc477943),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61a7ac),
	.w1(32'hbc1e2bf4),
	.w2(32'hba82d322),
	.w3(32'hbc7a400b),
	.w4(32'h3bc299b1),
	.w5(32'hbb9eb605),
	.w6(32'hbce8a68d),
	.w7(32'hbba1e642),
	.w8(32'h3abe6983),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb9692),
	.w1(32'hba1fa690),
	.w2(32'hb91eee96),
	.w3(32'hbb220808),
	.w4(32'h3c1bc166),
	.w5(32'hbb0ccca7),
	.w6(32'h3a759dc1),
	.w7(32'h3bc6bfeb),
	.w8(32'hb92f5466),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d4ba2),
	.w1(32'h3c0cd411),
	.w2(32'hbc8a1d57),
	.w3(32'h3ba5eea9),
	.w4(32'hbb0b64bd),
	.w5(32'hbc41ae95),
	.w6(32'h3c0c2794),
	.w7(32'hbb46748d),
	.w8(32'hbb6b0e45),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba574e),
	.w1(32'h3bd2e82a),
	.w2(32'hbc25a714),
	.w3(32'hbc3d1516),
	.w4(32'hbc90888d),
	.w5(32'hba531469),
	.w6(32'h3b8f0223),
	.w7(32'hbc9d875c),
	.w8(32'h3c004f5c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0be65c),
	.w1(32'hbc004685),
	.w2(32'hbd0bb78c),
	.w3(32'h3c28b8fb),
	.w4(32'hbbab3de1),
	.w5(32'h3bc734ae),
	.w6(32'hbc52041a),
	.w7(32'hbbe5c264),
	.w8(32'h3c5c144b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30a0b5),
	.w1(32'hbb8ebc73),
	.w2(32'hbc3ef6c2),
	.w3(32'h3cb3e011),
	.w4(32'h3b6ab319),
	.w5(32'h3c66c87d),
	.w6(32'h3c8b6bc3),
	.w7(32'h3c8cecb6),
	.w8(32'hbc41de0e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc102775),
	.w1(32'h3be1a297),
	.w2(32'hbc727b5f),
	.w3(32'hbb761401),
	.w4(32'hbca69379),
	.w5(32'hbb45e818),
	.w6(32'hbc5c2136),
	.w7(32'h3bcb0dc3),
	.w8(32'h3c4aaa84),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cb5d2),
	.w1(32'hbc53e581),
	.w2(32'hbd12c200),
	.w3(32'h3b229f4c),
	.w4(32'h3c1f7293),
	.w5(32'hbcf980ed),
	.w6(32'hbb8bb4cb),
	.w7(32'hbca3007a),
	.w8(32'hbbdabe56),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fc6d1),
	.w1(32'h3c84ea0d),
	.w2(32'hbc8e7a56),
	.w3(32'hbca99cdf),
	.w4(32'hbc9eb62d),
	.w5(32'h3c812246),
	.w6(32'hbbdee6f5),
	.w7(32'hbc408cf0),
	.w8(32'h3c45ff50),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf04e21),
	.w1(32'h3d2b9ac3),
	.w2(32'hbc6b9ba1),
	.w3(32'h3b84faba),
	.w4(32'h3c145471),
	.w5(32'hba6f7b7d),
	.w6(32'h3c8ca67a),
	.w7(32'hbc00f908),
	.w8(32'h3c0e8dde),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf43e7),
	.w1(32'hbc83046b),
	.w2(32'hbbf75bb8),
	.w3(32'h3c37c8e0),
	.w4(32'h3b1c8310),
	.w5(32'h3c593aa7),
	.w6(32'h3a1b216b),
	.w7(32'h3b92bfa0),
	.w8(32'h3c9f19c3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba130fb),
	.w1(32'h3bd0f5bd),
	.w2(32'hba0f8c5f),
	.w3(32'hbc9f6ca4),
	.w4(32'hbc5a50ea),
	.w5(32'h39ab0e74),
	.w6(32'hbb8a44ba),
	.w7(32'hbbabd66b),
	.w8(32'h3cef26ac),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bea63),
	.w1(32'hbcca0dc3),
	.w2(32'hbbe6839a),
	.w3(32'h3b02f04c),
	.w4(32'hbcbc64af),
	.w5(32'h3bf28c95),
	.w6(32'h3c5d66a1),
	.w7(32'h3bdb80b4),
	.w8(32'h3b2f6d2f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012c6d),
	.w1(32'h3ccff50a),
	.w2(32'h3baca780),
	.w3(32'h3c70942e),
	.w4(32'h3b0bce5d),
	.w5(32'h3b822fc9),
	.w6(32'h3cdacc33),
	.w7(32'h3c1bf565),
	.w8(32'hbb390efc),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3f53e),
	.w1(32'hbbcbbce1),
	.w2(32'hbb6721f0),
	.w3(32'h3b0e9731),
	.w4(32'hbc5faafd),
	.w5(32'hbb067a0f),
	.w6(32'hba95e55f),
	.w7(32'hbc2b9a94),
	.w8(32'hbbf40dae),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec5e76),
	.w1(32'hbb98b328),
	.w2(32'hbbb4724a),
	.w3(32'hbb677a05),
	.w4(32'hbbe9e733),
	.w5(32'hbbfc3b84),
	.w6(32'hbb207313),
	.w7(32'hbbf2daa2),
	.w8(32'hbc15a7a0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac23f),
	.w1(32'h3b6e2ee7),
	.w2(32'hbc65398b),
	.w3(32'h3aeee08b),
	.w4(32'h3b56f842),
	.w5(32'hbaa2d69b),
	.w6(32'h3b2619cb),
	.w7(32'hbafef66a),
	.w8(32'h3b4c44c2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba955bfc),
	.w1(32'h3be5c407),
	.w2(32'hbb2e7589),
	.w3(32'h3b25b906),
	.w4(32'hbd09b014),
	.w5(32'h3c3e7e8f),
	.w6(32'h3c4b4891),
	.w7(32'hbb9ffe13),
	.w8(32'h3d91fc16),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8a247),
	.w1(32'hbcc24238),
	.w2(32'hbc1df29c),
	.w3(32'hbca2c1c9),
	.w4(32'h3a7e31a4),
	.w5(32'hba02a251),
	.w6(32'hbc4d04ce),
	.w7(32'h3c71f7b5),
	.w8(32'h3c8c2242),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cf1ab),
	.w1(32'hbae4932b),
	.w2(32'hbc6ce64e),
	.w3(32'hbc81a810),
	.w4(32'hbc32fd7b),
	.w5(32'hbc9f726f),
	.w6(32'hbd0438ce),
	.w7(32'hbb902977),
	.w8(32'h3ca708ec),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd7615e),
	.w1(32'h3b64e2a6),
	.w2(32'hbbdfe048),
	.w3(32'h3bdbaa0f),
	.w4(32'hbad79978),
	.w5(32'h3c838b87),
	.w6(32'hbb7bded8),
	.w7(32'hbc267ad2),
	.w8(32'hbbfc3fe7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b853d),
	.w1(32'h3c096abd),
	.w2(32'hbc97dc59),
	.w3(32'hb9c6677d),
	.w4(32'hbbcc3236),
	.w5(32'hbbb51751),
	.w6(32'h3c13d7ad),
	.w7(32'hbb872de3),
	.w8(32'hbc38c623),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6976e),
	.w1(32'hbbfa4034),
	.w2(32'hbc2bafbc),
	.w3(32'h3b135ea2),
	.w4(32'hba17ae6e),
	.w5(32'hba646f78),
	.w6(32'h3bb1f4e1),
	.w7(32'hbb52e480),
	.w8(32'hbc7d3873),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b8546),
	.w1(32'hbbdb79dc),
	.w2(32'h3b757502),
	.w3(32'hbbc14cfc),
	.w4(32'h3c3a2924),
	.w5(32'hbc7c7e5f),
	.w6(32'h3b84c0d6),
	.w7(32'h3c639833),
	.w8(32'hbc7ae046),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4aad26),
	.w1(32'hbc244ced),
	.w2(32'h3c3824ee),
	.w3(32'hbbd78afe),
	.w4(32'h3c840f40),
	.w5(32'h3bb8802d),
	.w6(32'hba23360c),
	.w7(32'h3cafc97b),
	.w8(32'h3be05d43),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21ce3b),
	.w1(32'h3c15bb64),
	.w2(32'hbb8656a9),
	.w3(32'h3b5a48c6),
	.w4(32'hbb5b6b29),
	.w5(32'hbbee93fe),
	.w6(32'h3c999634),
	.w7(32'hbab19d27),
	.w8(32'hbb961bd8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ee3b2),
	.w1(32'h3c68454b),
	.w2(32'h3b74a4df),
	.w3(32'h3c3d486a),
	.w4(32'hba83af60),
	.w5(32'h3ca317b8),
	.w6(32'h3c258527),
	.w7(32'h3b5ada01),
	.w8(32'h3cf3e3af),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9abd36),
	.w1(32'hbc8292a5),
	.w2(32'h3bfcc5a2),
	.w3(32'hbc9c82e2),
	.w4(32'h3c12bc92),
	.w5(32'h3bd8934e),
	.w6(32'hbc72e3b7),
	.w7(32'hbb81f4bc),
	.w8(32'hbbd40d30),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6d90b),
	.w1(32'hbb0da1b0),
	.w2(32'hbb5e5b6e),
	.w3(32'h393ca058),
	.w4(32'hbb918a19),
	.w5(32'h3c98f334),
	.w6(32'hbc6f9239),
	.w7(32'hbb574fd6),
	.w8(32'h38c35d9e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13b9dd),
	.w1(32'hbb631b6b),
	.w2(32'h3c37c979),
	.w3(32'hbc8f9cd6),
	.w4(32'h3c81c736),
	.w5(32'h3ca7ce66),
	.w6(32'hbc871e77),
	.w7(32'h3c9785cd),
	.w8(32'hbc4e7a61),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffa53c),
	.w1(32'h3cbd8eff),
	.w2(32'h3bf65502),
	.w3(32'h3b4bb110),
	.w4(32'h3b00b433),
	.w5(32'hbcfdf111),
	.w6(32'hbafa3a73),
	.w7(32'h3cb59772),
	.w8(32'hbceb33ae),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7eec1d),
	.w1(32'h3a3f5c22),
	.w2(32'h3af0c852),
	.w3(32'h3c72c26e),
	.w4(32'hbb6b1a5e),
	.w5(32'h3beff101),
	.w6(32'h3b8108fe),
	.w7(32'h392d56be),
	.w8(32'h3c274f83),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c286089),
	.w1(32'h3bc24d54),
	.w2(32'h3b545aea),
	.w3(32'h3be529a1),
	.w4(32'h3b9e3556),
	.w5(32'h3ae3e8a6),
	.w6(32'h3c042952),
	.w7(32'h3c91e356),
	.w8(32'hbcd8fd41),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe72e18),
	.w1(32'h3c182d76),
	.w2(32'h3c924672),
	.w3(32'h3ac411d7),
	.w4(32'h3ae9a21d),
	.w5(32'hbc2a12bb),
	.w6(32'h3c0bfcb1),
	.w7(32'h3c82431d),
	.w8(32'hbc055d00),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc273a23),
	.w1(32'hbc064b1d),
	.w2(32'hbd1430cd),
	.w3(32'h3c3615b8),
	.w4(32'hbd173ddc),
	.w5(32'h3b4fce66),
	.w6(32'h3bac678f),
	.w7(32'hbc93457d),
	.w8(32'h3d96481b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d606718),
	.w1(32'hbd1365e7),
	.w2(32'h3c38329b),
	.w3(32'hbce66bff),
	.w4(32'h3bcb9991),
	.w5(32'hbb9e1bb2),
	.w6(32'hbc359183),
	.w7(32'h3be45dd5),
	.w8(32'hbbfdebec),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23e82c),
	.w1(32'h3be85c4d),
	.w2(32'h3ca666cd),
	.w3(32'h3c17f04b),
	.w4(32'h3cf7f86f),
	.w5(32'hbd21c89c),
	.w6(32'h3bbcbfbe),
	.w7(32'h3d199c4d),
	.w8(32'hbd988c59),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5e759d),
	.w1(32'h3d02665a),
	.w2(32'hbb9601b9),
	.w3(32'h3c985965),
	.w4(32'h3c24df49),
	.w5(32'hbc592d34),
	.w6(32'h3c7940e6),
	.w7(32'h3b864277),
	.w8(32'hbc35e941),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e97d3),
	.w1(32'h3998792e),
	.w2(32'hbc0c27f5),
	.w3(32'hbc34558a),
	.w4(32'hbc8ecb93),
	.w5(32'hbb1e8b9e),
	.w6(32'hbc8b014e),
	.w7(32'hba160c13),
	.w8(32'h3c218083),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1a19b),
	.w1(32'hbcbed8b4),
	.w2(32'h3c29ec29),
	.w3(32'hbcddf636),
	.w4(32'hbb928872),
	.w5(32'h3c5aed63),
	.w6(32'hbc8f5f4f),
	.w7(32'h3c310132),
	.w8(32'h3bbb0289),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb716ee4),
	.w1(32'hbc8ffa0d),
	.w2(32'h3be958c3),
	.w3(32'hbc8ce65b),
	.w4(32'hbb8b8d75),
	.w5(32'hbb6bd17e),
	.w6(32'hbd122803),
	.w7(32'h3bae57dc),
	.w8(32'hbc35e83f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023d34),
	.w1(32'h39c1ba83),
	.w2(32'hbc433e3b),
	.w3(32'h3c20fb59),
	.w4(32'h3bc62af4),
	.w5(32'h3b29a25e),
	.w6(32'h3c23b4b2),
	.w7(32'hbc216fb8),
	.w8(32'hbc8037f4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b8969),
	.w1(32'hbbcbcf68),
	.w2(32'h3c678e56),
	.w3(32'h3a524e38),
	.w4(32'h3cd9552c),
	.w5(32'hbcd2a740),
	.w6(32'h3b30942c),
	.w7(32'h3cb403f5),
	.w8(32'hbccd5014),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e12ad),
	.w1(32'h3cad69c4),
	.w2(32'h3c34f042),
	.w3(32'h3d13db55),
	.w4(32'hbb40d89d),
	.w5(32'hbca9e89c),
	.w6(32'h3c5e2762),
	.w7(32'h3c026642),
	.w8(32'hbc028017),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90b67f),
	.w1(32'hbc36fe7f),
	.w2(32'h3bd475af),
	.w3(32'h3cc19ed0),
	.w4(32'h3a31baa5),
	.w5(32'h3b511d4e),
	.w6(32'h3c9abf25),
	.w7(32'h3c5a2838),
	.w8(32'hba6cae85),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae90cd8),
	.w1(32'hbac55886),
	.w2(32'h3b4fba4b),
	.w3(32'hbadd484b),
	.w4(32'hbbee25ac),
	.w5(32'h3ba5f032),
	.w6(32'hbb702462),
	.w7(32'hbc6b08d3),
	.w8(32'h3a0eeccc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc028f),
	.w1(32'hbc6fb63d),
	.w2(32'h3b317db9),
	.w3(32'h3c070bfe),
	.w4(32'h3c785e81),
	.w5(32'hbce79a86),
	.w6(32'hbc06e00e),
	.w7(32'h3c7024dc),
	.w8(32'hbdb86c86),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0283ec),
	.w1(32'h3ca40023),
	.w2(32'h3bc97d20),
	.w3(32'h3c67ab2b),
	.w4(32'h3bf5afaf),
	.w5(32'h3c2eb10e),
	.w6(32'h3d019c58),
	.w7(32'h3bf8ffde),
	.w8(32'hbc984d3e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc183034),
	.w1(32'h3c57074d),
	.w2(32'hbc571078),
	.w3(32'h3add2daf),
	.w4(32'h3bbbe4b2),
	.w5(32'hbbaffa0c),
	.w6(32'h3adcf233),
	.w7(32'hbc99374b),
	.w8(32'hbc0695ef),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab28da7),
	.w1(32'h3c997a2e),
	.w2(32'hbc445fa2),
	.w3(32'h3a9c2a32),
	.w4(32'hba62f665),
	.w5(32'hbc140627),
	.w6(32'h3cc4f41f),
	.w7(32'hbaeb7de4),
	.w8(32'h3b3a21eb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb232aa),
	.w1(32'hbbf186fe),
	.w2(32'hbcbc81f6),
	.w3(32'hbc2dffdb),
	.w4(32'hbcddf1ab),
	.w5(32'hbc00a45c),
	.w6(32'hbcf86233),
	.w7(32'hbc97ebdd),
	.w8(32'h3b114814),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc82f1a),
	.w1(32'hbcf61d99),
	.w2(32'hbc8d7e4e),
	.w3(32'hbcefcb9b),
	.w4(32'hbaa8935d),
	.w5(32'h3c2079c4),
	.w6(32'hbcdf38c4),
	.w7(32'hbbd93ae9),
	.w8(32'h3cd10f80),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe4615),
	.w1(32'h3c562f50),
	.w2(32'hbc550f79),
	.w3(32'hbc9f7bb4),
	.w4(32'hbc34802e),
	.w5(32'h3c683c89),
	.w6(32'h3aa5b372),
	.w7(32'hbc8a5245),
	.w8(32'h3c3a06f4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c113525),
	.w1(32'hbbbae3bf),
	.w2(32'h3bcc4044),
	.w3(32'h3bd307dc),
	.w4(32'hbc7b239a),
	.w5(32'h3bed2c6e),
	.w6(32'h3c24cbe5),
	.w7(32'hbc5c7c84),
	.w8(32'hbbbb997d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8dce2),
	.w1(32'hbb915d0f),
	.w2(32'h3b497a89),
	.w3(32'h3a1015e9),
	.w4(32'hbb803e9b),
	.w5(32'h3b2e678d),
	.w6(32'hbc2bbf11),
	.w7(32'h3b7ccd31),
	.w8(32'hbb84c370),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dbe71),
	.w1(32'hba9c203a),
	.w2(32'h3a9b301d),
	.w3(32'hbad1df71),
	.w4(32'h3bdce312),
	.w5(32'hbc4018c4),
	.w6(32'hbaea8717),
	.w7(32'hbbebd1e4),
	.w8(32'hbd079270),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c824a82),
	.w1(32'h3c19a16a),
	.w2(32'hbc3948c8),
	.w3(32'h3c14cf9e),
	.w4(32'hbb799d41),
	.w5(32'h3c9bd8ae),
	.w6(32'h3cb89aa6),
	.w7(32'hbc599670),
	.w8(32'h3cc22926),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bc19a),
	.w1(32'hbb52ad9d),
	.w2(32'h3b0cbb06),
	.w3(32'hbbe2943b),
	.w4(32'h3bc284d2),
	.w5(32'hbba81f80),
	.w6(32'h3c2c6522),
	.w7(32'h3c0f9c7e),
	.w8(32'hba52abab),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42949f),
	.w1(32'hbb5fd55a),
	.w2(32'hbc4d7c32),
	.w3(32'hbbcf5049),
	.w4(32'h3b94e932),
	.w5(32'h3c93f01d),
	.w6(32'hbb405dfa),
	.w7(32'h3ac7e282),
	.w8(32'h3c8c3ace),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ae986),
	.w1(32'h3c6b4c72),
	.w2(32'h3bd158fa),
	.w3(32'hbb8ee273),
	.w4(32'hbafcce65),
	.w5(32'h3b44126b),
	.w6(32'h3bee8f2d),
	.w7(32'h3c21f196),
	.w8(32'hba47fce2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9989d22),
	.w1(32'hb9e7fd5f),
	.w2(32'h3b96f4d1),
	.w3(32'hbacaf8e5),
	.w4(32'h3a7f9950),
	.w5(32'h3c98be7c),
	.w6(32'hbacf4f98),
	.w7(32'hbc3610b0),
	.w8(32'h3cd2c3c4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35670a),
	.w1(32'hb9a5187c),
	.w2(32'h3c6e88da),
	.w3(32'hbc436ff4),
	.w4(32'hbb920021),
	.w5(32'hba17091f),
	.w6(32'hbbef11d5),
	.w7(32'hbac5cd7e),
	.w8(32'hbd3b4fa3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd425596),
	.w1(32'h3c5b453e),
	.w2(32'h3ab360ee),
	.w3(32'hbbdb0175),
	.w4(32'h3bf05abd),
	.w5(32'hbb8b5337),
	.w6(32'h3d0ae4cf),
	.w7(32'h3bfa09ae),
	.w8(32'hbb43b3fb),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a5319),
	.w1(32'hbbc26706),
	.w2(32'hbc2852fa),
	.w3(32'h3b28f86a),
	.w4(32'hbc03d0af),
	.w5(32'h3bd0078b),
	.w6(32'h38c01b78),
	.w7(32'hbc5d9b92),
	.w8(32'hbc3c3dc5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82e2a3),
	.w1(32'hbb1a2a74),
	.w2(32'h3bb04ae6),
	.w3(32'hbbdb480a),
	.w4(32'h3b63b64f),
	.w5(32'h3ae67f05),
	.w6(32'hbbbf8438),
	.w7(32'h3bd2e541),
	.w8(32'hbc1c1e52),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule