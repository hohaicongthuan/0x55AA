module layer_8_featuremap_135(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b8c31),
	.w1(32'hbbc0e257),
	.w2(32'hbb7f0039),
	.w3(32'hb9f8b6f6),
	.w4(32'h3ae649f1),
	.w5(32'h3c839320),
	.w6(32'h3c0ffe90),
	.w7(32'hbc8f32f5),
	.w8(32'hbbe7c180),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe68742),
	.w1(32'hbca6b3d1),
	.w2(32'h3b422185),
	.w3(32'h3c4d1325),
	.w4(32'hba4268d2),
	.w5(32'h3a6cd249),
	.w6(32'hbc8cf68f),
	.w7(32'hbba6c409),
	.w8(32'hbb9b40fd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc882d),
	.w1(32'h3a543e3e),
	.w2(32'hbc8a61df),
	.w3(32'hbbd23b44),
	.w4(32'h3a11fdaa),
	.w5(32'hbc13c185),
	.w6(32'hbc24b19e),
	.w7(32'h3c64fb08),
	.w8(32'h3ada47cc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c584348),
	.w1(32'h3b8c203d),
	.w2(32'h3b98c43f),
	.w3(32'h3bdc59ef),
	.w4(32'h3b087e93),
	.w5(32'hbb534408),
	.w6(32'hbc487ddf),
	.w7(32'hbc8d5954),
	.w8(32'hbb9fac11),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4e986),
	.w1(32'hbc63f2ce),
	.w2(32'hbab7741f),
	.w3(32'hbc067327),
	.w4(32'hbb7b7958),
	.w5(32'hbaaa096e),
	.w6(32'h3c47e940),
	.w7(32'hbbd389d0),
	.w8(32'hbcae6a3f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c2636),
	.w1(32'hbc3d25dc),
	.w2(32'h3c8546cc),
	.w3(32'hbc795e45),
	.w4(32'h3b408c9c),
	.w5(32'h3c59bcda),
	.w6(32'h3bbeed41),
	.w7(32'hbcb9c231),
	.w8(32'hbbb0b971),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf3e3f),
	.w1(32'hbc25195c),
	.w2(32'h3c137f06),
	.w3(32'hbb9d43a5),
	.w4(32'h3ba5d794),
	.w5(32'h3c1dbb1b),
	.w6(32'h3bc6c282),
	.w7(32'h3bd0a38f),
	.w8(32'hbc3da480),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d2f89),
	.w1(32'hbbc70c42),
	.w2(32'h398d00ab),
	.w3(32'hba46edb1),
	.w4(32'hbb822882),
	.w5(32'h3bf77a16),
	.w6(32'h3bf5696c),
	.w7(32'hbc077708),
	.w8(32'h3badf946),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a4163),
	.w1(32'h3a8f9e7f),
	.w2(32'h3c0a4089),
	.w3(32'hbb7cce0d),
	.w4(32'h39a3e5fa),
	.w5(32'h391cb086),
	.w6(32'hbb226005),
	.w7(32'h3b9ea4e0),
	.w8(32'h3b96afa9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac45091),
	.w1(32'h3b2e75f2),
	.w2(32'hbbfa7aee),
	.w3(32'h3ba52bae),
	.w4(32'hbc9c1566),
	.w5(32'hbca0d502),
	.w6(32'hbc849d24),
	.w7(32'h3cbe3c48),
	.w8(32'h3c21d849),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd2142),
	.w1(32'h3c905d4d),
	.w2(32'hbd3da516),
	.w3(32'h3c8cb2c1),
	.w4(32'hbc2351bf),
	.w5(32'hbcf5a2d4),
	.w6(32'hbd655c2d),
	.w7(32'hbb7b2956),
	.w8(32'hbc9a697e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c011b20),
	.w1(32'hbbd11afd),
	.w2(32'hbae377b5),
	.w3(32'hbbcda572),
	.w4(32'h3ae43598),
	.w5(32'hbae08953),
	.w6(32'hbcee0237),
	.w7(32'hbcad3c02),
	.w8(32'hbc927cd4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2c52f),
	.w1(32'hbb4f8362),
	.w2(32'h3a0bb929),
	.w3(32'hbb5a1fbe),
	.w4(32'h3b0cda11),
	.w5(32'h3b0b82b9),
	.w6(32'hba2e8fbf),
	.w7(32'hb9e7f805),
	.w8(32'h3922b995),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90523d),
	.w1(32'h3928a143),
	.w2(32'hbbdb33de),
	.w3(32'h374891d9),
	.w4(32'hbc3fceab),
	.w5(32'h3baf978b),
	.w6(32'hbb2aeb6b),
	.w7(32'hbc315d21),
	.w8(32'h3c0295e2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b108b22),
	.w1(32'h3bade9ca),
	.w2(32'hbbc438e5),
	.w3(32'h3b5a298b),
	.w4(32'hbbeb212b),
	.w5(32'hbaf43f63),
	.w6(32'h3b8cefb6),
	.w7(32'hbbd50892),
	.w8(32'hba8b771c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66f5e3),
	.w1(32'h3b6b270e),
	.w2(32'h3bb64183),
	.w3(32'h3baf0588),
	.w4(32'h3a27afe1),
	.w5(32'hbb993311),
	.w6(32'h3bf99d61),
	.w7(32'h3bbc56d6),
	.w8(32'h3a8cd9eb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb958bd),
	.w1(32'h3b5f9107),
	.w2(32'hbc0f370c),
	.w3(32'h3c6c9848),
	.w4(32'hbc7e47d5),
	.w5(32'hbbe79084),
	.w6(32'h3bf7bffc),
	.w7(32'hb9ca57c8),
	.w8(32'h3bb6243e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b148026),
	.w1(32'hbc765ff1),
	.w2(32'hbc1acbb2),
	.w3(32'hbca42612),
	.w4(32'hba32ac1f),
	.w5(32'hbb759ae5),
	.w6(32'hba18195e),
	.w7(32'h3b0beb2d),
	.w8(32'hbc08a6b9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a037b),
	.w1(32'hbb823d1e),
	.w2(32'h3b345a4d),
	.w3(32'hbcc5088a),
	.w4(32'hbba26114),
	.w5(32'hbbab614c),
	.w6(32'hbc436e8b),
	.w7(32'h3aa31f25),
	.w8(32'h3abd7123),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0bb54),
	.w1(32'hbc86be5b),
	.w2(32'hbbc1d37b),
	.w3(32'hbc519578),
	.w4(32'hbc7fad98),
	.w5(32'h3c2c785b),
	.w6(32'hbcad63dc),
	.w7(32'hbad9a6f7),
	.w8(32'hbc8bda28),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32fb7e),
	.w1(32'h3b0d4258),
	.w2(32'h3bf26a12),
	.w3(32'h3c3c37f3),
	.w4(32'h3c44c56f),
	.w5(32'hbca1b572),
	.w6(32'hbbc47ef6),
	.w7(32'h3c35b7cd),
	.w8(32'hbd7c0df3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de78cf),
	.w1(32'h3b79cc7a),
	.w2(32'hbb8e6b22),
	.w3(32'h3c891535),
	.w4(32'h3be147dc),
	.w5(32'h3aca1703),
	.w6(32'h3c8831a7),
	.w7(32'hbc856709),
	.w8(32'h3a85cfe9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca39176),
	.w1(32'h3b43c1ad),
	.w2(32'hbb1b2f3f),
	.w3(32'hbb21a595),
	.w4(32'hbc80fa89),
	.w5(32'h3b923abb),
	.w6(32'h3bc21a73),
	.w7(32'hbb24a056),
	.w8(32'h3b88173e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba86638),
	.w1(32'hbb73c6dc),
	.w2(32'hbbeb19cb),
	.w3(32'hbc122168),
	.w4(32'hbbcc3291),
	.w5(32'h3a8995cb),
	.w6(32'hb9f3d76b),
	.w7(32'hbbd52a48),
	.w8(32'hbab9c413),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaf889),
	.w1(32'hbb514969),
	.w2(32'hba9186c8),
	.w3(32'h3a3eef0f),
	.w4(32'hbb3b5835),
	.w5(32'hbbed18e0),
	.w6(32'hb967c2f3),
	.w7(32'h3846bfb5),
	.w8(32'hbbfa2b60),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe018d9),
	.w1(32'hbbd3f6e8),
	.w2(32'hba8f7201),
	.w3(32'h3b39dded),
	.w4(32'hbbf8c37f),
	.w5(32'hbb7e1c4b),
	.w6(32'h3b30b818),
	.w7(32'hbad7d03f),
	.w8(32'hbc6b2a02),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed3b2),
	.w1(32'h3c2d86c7),
	.w2(32'hbb67c605),
	.w3(32'h3c33ffc8),
	.w4(32'h3c0452ce),
	.w5(32'h3b138ad7),
	.w6(32'h3cb33417),
	.w7(32'h3be2bf1e),
	.w8(32'hbc96acac),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae5ac7),
	.w1(32'hbc909f1a),
	.w2(32'hbc746bf0),
	.w3(32'hbc78f554),
	.w4(32'hbcbf0698),
	.w5(32'hbc880bd1),
	.w6(32'hbb170f1d),
	.w7(32'hbcef2b60),
	.w8(32'hbd322d1b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49289b),
	.w1(32'h3c044500),
	.w2(32'h3bafc182),
	.w3(32'h3c5b97c9),
	.w4(32'hbc65762e),
	.w5(32'h3afabf36),
	.w6(32'hbaab654e),
	.w7(32'h3c235182),
	.w8(32'hbc28256a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71884),
	.w1(32'h3bbdb993),
	.w2(32'h3ca16f25),
	.w3(32'hbb41d0c2),
	.w4(32'h39e6c377),
	.w5(32'hbc08ed99),
	.w6(32'h3c3e7d26),
	.w7(32'h3c857a66),
	.w8(32'hbc5debc1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8e05b),
	.w1(32'h3c7d405a),
	.w2(32'hba140425),
	.w3(32'h3ba72f2b),
	.w4(32'hbb389386),
	.w5(32'h3a2e64fb),
	.w6(32'h3c64dc67),
	.w7(32'hbaae035c),
	.w8(32'h3b075222),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38789d9e),
	.w1(32'h3a12cf67),
	.w2(32'hbbb7b03f),
	.w3(32'h3a812d50),
	.w4(32'hbc23cc82),
	.w5(32'hbaa5c11f),
	.w6(32'h3b60bacb),
	.w7(32'hbb3a9f84),
	.w8(32'hbb50fe9c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7c17f),
	.w1(32'h3c07b8b6),
	.w2(32'hbb8e679d),
	.w3(32'h3c75b97b),
	.w4(32'h3c55b05a),
	.w5(32'hbc488f18),
	.w6(32'hbbd489b4),
	.w7(32'hb94f1883),
	.w8(32'hbb9207d4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b680a),
	.w1(32'h3c5b7bf1),
	.w2(32'hbbf21b68),
	.w3(32'hbc93dbf9),
	.w4(32'hbbf2763b),
	.w5(32'hbc3f6505),
	.w6(32'hbb8a7754),
	.w7(32'h3b9dfaab),
	.w8(32'hbc9aa9a5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd16f38),
	.w1(32'hba2e3160),
	.w2(32'h3c78a646),
	.w3(32'hbc9b4a7d),
	.w4(32'h3c50c32b),
	.w5(32'h3be83789),
	.w6(32'h3c5569d5),
	.w7(32'h3c2ea9a2),
	.w8(32'h3b42efe1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c230bae),
	.w1(32'h3c071987),
	.w2(32'h3c70ea6b),
	.w3(32'h3c113300),
	.w4(32'h3c75bb1d),
	.w5(32'h3c1ae954),
	.w6(32'h3c35a22e),
	.w7(32'h3cc5a663),
	.w8(32'hba98ff96),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13ce3f),
	.w1(32'hbcf500ac),
	.w2(32'h3b9ddfe6),
	.w3(32'hbcf0de15),
	.w4(32'hbb7baa90),
	.w5(32'h3aa85f31),
	.w6(32'hbd029749),
	.w7(32'hbc4eb9b7),
	.w8(32'hbc7f92bc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc131156),
	.w1(32'hbb9892b8),
	.w2(32'hbc980d20),
	.w3(32'h3ba2eb13),
	.w4(32'hbc333553),
	.w5(32'hbacc430b),
	.w6(32'hbb103e12),
	.w7(32'hbb3e887e),
	.w8(32'h3cc47881),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76fa77),
	.w1(32'hbc74b33b),
	.w2(32'h3b29f67c),
	.w3(32'hbc980f8a),
	.w4(32'h3bf057cf),
	.w5(32'hbc20fb92),
	.w6(32'hbc40587c),
	.w7(32'h3c5d2bfe),
	.w8(32'hbcf22d2f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc602725),
	.w1(32'h3c93234d),
	.w2(32'hbb6a9382),
	.w3(32'h3b3bf2da),
	.w4(32'h3ab39cfa),
	.w5(32'h3b3edae5),
	.w6(32'h3c4eebe4),
	.w7(32'hbba789aa),
	.w8(32'hbb8762a1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5841c0),
	.w1(32'h3b3ee81d),
	.w2(32'hbab6c5e7),
	.w3(32'hbc009192),
	.w4(32'hbc0f0c48),
	.w5(32'h3a8cd3ac),
	.w6(32'hbc622918),
	.w7(32'hbc8a8bce),
	.w8(32'h3c3492f0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a6408),
	.w1(32'h3b52ba90),
	.w2(32'h3c4785fc),
	.w3(32'hbc37ad56),
	.w4(32'h3c52a96b),
	.w5(32'hbc4e6a32),
	.w6(32'hbb5ea4b6),
	.w7(32'h3c4ebd4b),
	.w8(32'hbcc76892),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc764db),
	.w1(32'hb8febc34),
	.w2(32'hbc6e77b4),
	.w3(32'h3bb6439c),
	.w4(32'h3bd55c08),
	.w5(32'h3c305625),
	.w6(32'hbbc4b851),
	.w7(32'h3bb6adbd),
	.w8(32'h3c9dafea),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad10c02),
	.w1(32'hbb42143a),
	.w2(32'hbabf62ee),
	.w3(32'hbc2b154d),
	.w4(32'hbb07ae13),
	.w5(32'hbbb01b53),
	.w6(32'hbbcd7435),
	.w7(32'hbb690016),
	.w8(32'hbb7f9a18),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd63442),
	.w1(32'hbb2a4008),
	.w2(32'hbc0b1666),
	.w3(32'hbb47ce8e),
	.w4(32'hbc1df80d),
	.w5(32'hbc5da354),
	.w6(32'hbb944008),
	.w7(32'h3b44bf07),
	.w8(32'hbc4a0c2c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d9e0f),
	.w1(32'h3c3c139f),
	.w2(32'h3bbec013),
	.w3(32'hbace3d1a),
	.w4(32'hbadf42b6),
	.w5(32'h3c824fed),
	.w6(32'h3bd5e691),
	.w7(32'hbbf3c54c),
	.w8(32'h3c32ac9c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b890d77),
	.w1(32'hbc84c3e3),
	.w2(32'h3a483c7f),
	.w3(32'hbb999098),
	.w4(32'h3bacf5d2),
	.w5(32'hbc61a465),
	.w6(32'hbcbb17e9),
	.w7(32'hbb110c64),
	.w8(32'hbc0dd4ac),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b835fc2),
	.w1(32'h3bfccd06),
	.w2(32'h3b835e71),
	.w3(32'h3aa8e7d6),
	.w4(32'hbc277b0d),
	.w5(32'h3c34adca),
	.w6(32'h3a4416d6),
	.w7(32'hbb97da93),
	.w8(32'h3caeba19),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08454e),
	.w1(32'hbc7f6909),
	.w2(32'h3b3538c9),
	.w3(32'h3b342b8c),
	.w4(32'h3c1c7356),
	.w5(32'hbc2c8190),
	.w6(32'hbc2b0322),
	.w7(32'h3c6390f6),
	.w8(32'hbcbfdb94),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43cb29),
	.w1(32'hb9b24654),
	.w2(32'hbcfc1834),
	.w3(32'h3c2db6f0),
	.w4(32'hbcc11d40),
	.w5(32'hbc2badc3),
	.w6(32'h3c6000c0),
	.w7(32'hbca90e98),
	.w8(32'h3bb8d17d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d8a5c),
	.w1(32'hbbb396d0),
	.w2(32'h3c0ad964),
	.w3(32'h3a91274d),
	.w4(32'hbbc7c53d),
	.w5(32'h3c44beb9),
	.w6(32'h3b8d4903),
	.w7(32'h3c497627),
	.w8(32'h3cffd879),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69332e),
	.w1(32'hbcfa0d5a),
	.w2(32'h3b3e60e3),
	.w3(32'h3c07db48),
	.w4(32'hbba2e75e),
	.w5(32'hbcafee9b),
	.w6(32'h3b37c553),
	.w7(32'hbc1efdae),
	.w8(32'hbc4353a1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16b188),
	.w1(32'h3c980d37),
	.w2(32'hbc3b2f08),
	.w3(32'h3b67ba7b),
	.w4(32'h3b35ae6f),
	.w5(32'h3b064719),
	.w6(32'h3c819127),
	.w7(32'hbc0dfa80),
	.w8(32'h3d199836),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ef08b),
	.w1(32'h3be9c3ae),
	.w2(32'hba6ba616),
	.w3(32'hbbac5053),
	.w4(32'hbbb0e8fa),
	.w5(32'h391b675a),
	.w6(32'hbc46633f),
	.w7(32'hbbb6dfd6),
	.w8(32'h3ab7caea),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e8926),
	.w1(32'h39892d19),
	.w2(32'h3c0384dc),
	.w3(32'hb9b09c7d),
	.w4(32'h3ba786cf),
	.w5(32'hbb40f853),
	.w6(32'hbb35f6fc),
	.w7(32'hbb0e09f3),
	.w8(32'hbc646392),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49aa33),
	.w1(32'h3bb51670),
	.w2(32'hbc6aeeab),
	.w3(32'h3b766b21),
	.w4(32'hbc625795),
	.w5(32'h3c5e12d1),
	.w6(32'hbbb634a5),
	.w7(32'hbcd23e95),
	.w8(32'h3c9760fd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b5b95),
	.w1(32'hbc8df607),
	.w2(32'hbc024f9d),
	.w3(32'hbc14a475),
	.w4(32'hbbcc871e),
	.w5(32'hbba1210e),
	.w6(32'hbca2d12e),
	.w7(32'hbc04d342),
	.w8(32'hbc16c082),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa2f2f),
	.w1(32'hbb85e7d8),
	.w2(32'h3c275898),
	.w3(32'hbb9ec720),
	.w4(32'hbc672fa4),
	.w5(32'h3c135606),
	.w6(32'h3b91c7bc),
	.w7(32'hbb09e3bb),
	.w8(32'hbb74ddb9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f06ca),
	.w1(32'hbc17a567),
	.w2(32'h39d7fe2a),
	.w3(32'h3c5b4a7c),
	.w4(32'hbb7b2dc5),
	.w5(32'hbb3b084b),
	.w6(32'h3b4f6c0c),
	.w7(32'hbb822974),
	.w8(32'h398cccae),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69525b),
	.w1(32'hba57c27c),
	.w2(32'h3b238d87),
	.w3(32'hbaff08cc),
	.w4(32'h3b888615),
	.w5(32'h3ac574fd),
	.w6(32'hbb73bcdd),
	.w7(32'hbc007909),
	.w8(32'h3bf24ab4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a0431),
	.w1(32'h3bd40241),
	.w2(32'h3bd84eaf),
	.w3(32'h3c04ae25),
	.w4(32'h3b91b990),
	.w5(32'h3d09c68f),
	.w6(32'h3c549452),
	.w7(32'h3ba00610),
	.w8(32'h3d597122),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89bb06),
	.w1(32'hbb93ab4b),
	.w2(32'hb9f201b2),
	.w3(32'hbd180d95),
	.w4(32'hbb205de0),
	.w5(32'h3a589fef),
	.w6(32'hbd096a47),
	.w7(32'hb9495b39),
	.w8(32'hbba0ad7b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea1461),
	.w1(32'hbc0f5c98),
	.w2(32'hbb54ba7c),
	.w3(32'h3c2a56ad),
	.w4(32'hbae99679),
	.w5(32'h3c3aae39),
	.w6(32'h3b1281c1),
	.w7(32'hbc56ac94),
	.w8(32'h3d0aa56e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04b9b5),
	.w1(32'hb946a20b),
	.w2(32'hbaeb394b),
	.w3(32'h3c093c7c),
	.w4(32'h3b02cb8e),
	.w5(32'hbb809928),
	.w6(32'h3bae8f7b),
	.w7(32'h3be7a193),
	.w8(32'hbb8e96c2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba036f47),
	.w1(32'h3c1ccaa1),
	.w2(32'h3a8b5126),
	.w3(32'h3c31a91a),
	.w4(32'h3bb5e2e1),
	.w5(32'h39a23bc3),
	.w6(32'h3b373eb8),
	.w7(32'h3c6a3f4b),
	.w8(32'hbc334e67),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b9641),
	.w1(32'h3c247735),
	.w2(32'hbc83f1a6),
	.w3(32'h3bfdaa9a),
	.w4(32'hbc3c1d85),
	.w5(32'hbc945d8b),
	.w6(32'h3bc38db3),
	.w7(32'hbbc08dab),
	.w8(32'hbb733b18),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7134d),
	.w1(32'hbc8bdfef),
	.w2(32'hbbabed73),
	.w3(32'hbca3864d),
	.w4(32'hbbc8a321),
	.w5(32'hbc4e473b),
	.w6(32'hbb004189),
	.w7(32'hbbd29a0b),
	.w8(32'hbc723207),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96ba06),
	.w1(32'hbc3c8788),
	.w2(32'h3c0173cf),
	.w3(32'hbbfb1ce1),
	.w4(32'h3c85db68),
	.w5(32'hbc13711a),
	.w6(32'hbc09693b),
	.w7(32'hbba957f9),
	.w8(32'hbc721927),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ee8df),
	.w1(32'h3c328b6b),
	.w2(32'h3a6d1baf),
	.w3(32'hbbcaa23e),
	.w4(32'hbafa6391),
	.w5(32'hbc3f35ce),
	.w6(32'hbc104bdf),
	.w7(32'hbc1afd39),
	.w8(32'hbb484520),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97726b),
	.w1(32'hbc00ae04),
	.w2(32'hbcc7ff5e),
	.w3(32'h3c0059e6),
	.w4(32'h3a8bfa56),
	.w5(32'hbc956d9b),
	.w6(32'hb8fc61cb),
	.w7(32'h3abc77c6),
	.w8(32'h3c2bf9f9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09fb7a),
	.w1(32'hbca2ab8b),
	.w2(32'h3b2891d8),
	.w3(32'hbc4a3071),
	.w4(32'hbb1eb265),
	.w5(32'hbb5f2ec6),
	.w6(32'hbc0df6bb),
	.w7(32'h3c4c3515),
	.w8(32'h3bbefb87),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc000423),
	.w1(32'hbb9404f6),
	.w2(32'hbc061ef5),
	.w3(32'h3aea9671),
	.w4(32'h39e4bdd3),
	.w5(32'hbca34111),
	.w6(32'h3a407b3a),
	.w7(32'h3c16c202),
	.w8(32'hbcd65129),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc951483),
	.w1(32'h3c25f050),
	.w2(32'h3b7a1426),
	.w3(32'h3ba1ebfc),
	.w4(32'hbc1cb14e),
	.w5(32'hbb3b1673),
	.w6(32'h3c1f4d19),
	.w7(32'h3a94347c),
	.w8(32'hbc15751a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2856d),
	.w1(32'h3ab87b37),
	.w2(32'hbbd4342c),
	.w3(32'h3c6e3f4d),
	.w4(32'h3aa2b9a4),
	.w5(32'hbc05e89e),
	.w6(32'hb9a81d68),
	.w7(32'hbb8d04b0),
	.w8(32'h39295e7a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7606685),
	.w1(32'h3b9e52d2),
	.w2(32'hbb9c4c9a),
	.w3(32'h3bc730bf),
	.w4(32'h3bf96bf3),
	.w5(32'h3c421b7b),
	.w6(32'h3c8cdebe),
	.w7(32'hbc20ef99),
	.w8(32'h3c7d0fe7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f8e47),
	.w1(32'hbb5a3f18),
	.w2(32'hbc82c038),
	.w3(32'h3a19f047),
	.w4(32'hbbf161be),
	.w5(32'hbb8fa762),
	.w6(32'hbbf4a31f),
	.w7(32'hbc379d76),
	.w8(32'hbb377f64),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56b497),
	.w1(32'hbc2eb596),
	.w2(32'hbb862eb3),
	.w3(32'hbc86d4c9),
	.w4(32'h3b043c1d),
	.w5(32'h3ac49391),
	.w6(32'hbc33103c),
	.w7(32'hbb6d003c),
	.w8(32'hba726c73),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbb36d),
	.w1(32'hbb0550a9),
	.w2(32'hbbfdc271),
	.w3(32'h3ac2e154),
	.w4(32'h3ac3093a),
	.w5(32'hbc1d2acd),
	.w6(32'hb890b96f),
	.w7(32'hbb4905c3),
	.w8(32'hbb8f14ae),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a154eeb),
	.w1(32'hbbb447de),
	.w2(32'hbbc1fddf),
	.w3(32'hba90171c),
	.w4(32'hbadd54d7),
	.w5(32'hbb0116f6),
	.w6(32'hbb5f2f08),
	.w7(32'hbb8a2757),
	.w8(32'hb992c7b0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b330931),
	.w1(32'h3a823815),
	.w2(32'hbbe8b141),
	.w3(32'h3895d331),
	.w4(32'h3a2b797b),
	.w5(32'h3bc3ca12),
	.w6(32'h3a572590),
	.w7(32'hbbc82f42),
	.w8(32'h3a591627),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae19d),
	.w1(32'h3c00de4d),
	.w2(32'hbc2783a4),
	.w3(32'hbb680311),
	.w4(32'h3ce7e7ef),
	.w5(32'h3b8bea0a),
	.w6(32'hbc2b4d5f),
	.w7(32'h3c9153c0),
	.w8(32'hbc329692),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc41798),
	.w1(32'hbb9d0ef1),
	.w2(32'h3c7ea07f),
	.w3(32'hba5825ce),
	.w4(32'hbb8d3e1b),
	.w5(32'h3cc33fab),
	.w6(32'hbb141258),
	.w7(32'h3ba4bb0a),
	.w8(32'hbbb3ad50),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7808f7),
	.w1(32'hbc39de5b),
	.w2(32'h3c7278f8),
	.w3(32'h3b11da6e),
	.w4(32'hbb98b818),
	.w5(32'h3c65d083),
	.w6(32'hbc692254),
	.w7(32'hbac7a6c5),
	.w8(32'hbc32714b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94a08f),
	.w1(32'hbbba30a7),
	.w2(32'hbbfb42f6),
	.w3(32'hbc4bc1b9),
	.w4(32'hbc49e2a8),
	.w5(32'hbbeb0d5f),
	.w6(32'hbc13a9d9),
	.w7(32'hbcdc23f9),
	.w8(32'hbb62d9cc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1d657),
	.w1(32'hbbb5df7a),
	.w2(32'hbbd48870),
	.w3(32'hbc2ba74e),
	.w4(32'hbbb60479),
	.w5(32'hbb51d926),
	.w6(32'h3c808b03),
	.w7(32'hbcafc8f7),
	.w8(32'h3b475db6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ca03f),
	.w1(32'hbb46c61d),
	.w2(32'hbc146bf5),
	.w3(32'h3cbebf3a),
	.w4(32'hbc467e69),
	.w5(32'hbc40d0b0),
	.w6(32'hbc395e7e),
	.w7(32'hbc14f84b),
	.w8(32'hbc0f82db),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03d05f),
	.w1(32'hbb601ecc),
	.w2(32'hbadf3830),
	.w3(32'h3ca1671e),
	.w4(32'hbcb04973),
	.w5(32'hbc17baca),
	.w6(32'h3b142fd3),
	.w7(32'hbce17ca2),
	.w8(32'h3c52246d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3bb94),
	.w1(32'hbc448bff),
	.w2(32'hbbfc96ba),
	.w3(32'h3c52012b),
	.w4(32'hbc034012),
	.w5(32'hbbf4e415),
	.w6(32'h3c1cd9bd),
	.w7(32'hbc395670),
	.w8(32'hbc117add),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e554e),
	.w1(32'hbb2f07f9),
	.w2(32'hbad4e506),
	.w3(32'hbb42bb96),
	.w4(32'h3c2f4466),
	.w5(32'h3a4a3875),
	.w6(32'hbb4ef889),
	.w7(32'h3bb0ffaf),
	.w8(32'hbbc13634),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72a932),
	.w1(32'hbc8c0c7a),
	.w2(32'hbb23ef72),
	.w3(32'hbaa58c96),
	.w4(32'h3b9ac94d),
	.w5(32'hbd0651fd),
	.w6(32'hbba814da),
	.w7(32'hbcf9e479),
	.w8(32'h3c8f989d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f6458),
	.w1(32'h3b0ca708),
	.w2(32'hbc512658),
	.w3(32'h3c2a53b8),
	.w4(32'h3cd92a46),
	.w5(32'h3cf532ea),
	.w6(32'h3c922478),
	.w7(32'h3cbc2055),
	.w8(32'hbc51c839),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5ec76),
	.w1(32'h3c2c31ff),
	.w2(32'h3bdd9c81),
	.w3(32'hbc0e8552),
	.w4(32'h3b617d5c),
	.w5(32'hbbfc4c8d),
	.w6(32'h3c7f6fb0),
	.w7(32'h3b7505f1),
	.w8(32'hbcbdf53d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42e188),
	.w1(32'hbb371325),
	.w2(32'h3bac80d7),
	.w3(32'h3b53660a),
	.w4(32'hbc8439c1),
	.w5(32'hbc72f3f2),
	.w6(32'hbbd56e98),
	.w7(32'hbc2c366b),
	.w8(32'h3d0211b3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d12bf80),
	.w1(32'h3b2aaf9c),
	.w2(32'h3c2f2386),
	.w3(32'hbbe53d19),
	.w4(32'h3bf5b5f4),
	.w5(32'h3b9edfa4),
	.w6(32'h3c3a48c4),
	.w7(32'hbc55fee8),
	.w8(32'h3c5abba6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc459267),
	.w1(32'hbbce3d46),
	.w2(32'h3abb093c),
	.w3(32'hbc064525),
	.w4(32'hba64d6a1),
	.w5(32'h3a865592),
	.w6(32'hbc932cb9),
	.w7(32'h39d94694),
	.w8(32'h3b92bcca),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0520fe),
	.w1(32'h3bd43658),
	.w2(32'hbc816b9f),
	.w3(32'h3a0152e9),
	.w4(32'h3bede29d),
	.w5(32'h3c296567),
	.w6(32'h3b6a703f),
	.w7(32'hbc143e70),
	.w8(32'hbbfbb21f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8efeef),
	.w1(32'hbc7c69f5),
	.w2(32'hbbc392f0),
	.w3(32'h3beae378),
	.w4(32'hbaacdc56),
	.w5(32'h3ae0778e),
	.w6(32'hbc39169b),
	.w7(32'hbc481c3c),
	.w8(32'h3cb431e1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca10b9e),
	.w1(32'hbbae9966),
	.w2(32'hbb97dad0),
	.w3(32'hbc166876),
	.w4(32'h3c0c4b6e),
	.w5(32'h3c0f96e4),
	.w6(32'h3c1c3672),
	.w7(32'h3c1578e9),
	.w8(32'hbc39b295),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0e0320),
	.w1(32'hbc1a4244),
	.w2(32'h3c040c19),
	.w3(32'hbbef1385),
	.w4(32'hbc6b7857),
	.w5(32'hbc918ef4),
	.w6(32'h3a1b5615),
	.w7(32'hbc325761),
	.w8(32'hbb6b6ed6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05b76e),
	.w1(32'h3c4cd57c),
	.w2(32'hbab1b8cc),
	.w3(32'h3aefed9b),
	.w4(32'hbd203194),
	.w5(32'hbc0558c0),
	.w6(32'h3bfa8c66),
	.w7(32'hbd14fdef),
	.w8(32'h3ce5ac2f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf444bf),
	.w1(32'h3b700169),
	.w2(32'hbb8db775),
	.w3(32'h3c594749),
	.w4(32'hbbb0a045),
	.w5(32'hbc29adf6),
	.w6(32'h3c93710e),
	.w7(32'hbcaca85b),
	.w8(32'hbbbd1b29),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25bed5),
	.w1(32'h3baffc79),
	.w2(32'h3af1f978),
	.w3(32'h3b80f454),
	.w4(32'h3cc508c2),
	.w5(32'h3b97da1c),
	.w6(32'h3bf41e3f),
	.w7(32'h3c86bee3),
	.w8(32'hbb6097ef),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a1e10),
	.w1(32'hbc1a3155),
	.w2(32'hbb1c2fca),
	.w3(32'hbc10a9cb),
	.w4(32'h3bd2a568),
	.w5(32'h3c3f8727),
	.w6(32'hbb4a5027),
	.w7(32'h3b71f618),
	.w8(32'h3a2ae49f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91bab9),
	.w1(32'hbcbe6ea5),
	.w2(32'hbb819bba),
	.w3(32'hbaf62fbd),
	.w4(32'h3b19ef1e),
	.w5(32'h3c8cf7b7),
	.w6(32'hbc9d18ea),
	.w7(32'hbaea7f5c),
	.w8(32'h3c646ba5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b944c7b),
	.w1(32'hba813de7),
	.w2(32'hbc4b1ba6),
	.w3(32'h3b54054b),
	.w4(32'h3b463dca),
	.w5(32'hbc315218),
	.w6(32'h3b23c710),
	.w7(32'hbbe7c01e),
	.w8(32'hbd1204d0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2e0d8),
	.w1(32'hbc007d3e),
	.w2(32'hbab3cf77),
	.w3(32'hbc8d5568),
	.w4(32'hbc8b7edb),
	.w5(32'h3c587a2d),
	.w6(32'h3b9c0e79),
	.w7(32'hbbd3848f),
	.w8(32'hbc7f315e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d5587),
	.w1(32'h3bfbd5ec),
	.w2(32'h3c82a3cc),
	.w3(32'h3be3101a),
	.w4(32'h3b2436a9),
	.w5(32'h3be3a8fc),
	.w6(32'h3bccab23),
	.w7(32'hbb0823e1),
	.w8(32'h3d1487e2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00dbe0),
	.w1(32'hbc2c1af8),
	.w2(32'hbb93265c),
	.w3(32'h3b90011e),
	.w4(32'h3b66e5fc),
	.w5(32'h3ad97681),
	.w6(32'h39f94f8c),
	.w7(32'hbadb6388),
	.w8(32'h3af19dc4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b201c85),
	.w1(32'h3b2203f1),
	.w2(32'h3c3d2841),
	.w3(32'h3acaa051),
	.w4(32'h3c9cba34),
	.w5(32'h3a8f738f),
	.w6(32'h3b584198),
	.w7(32'h3cff73f0),
	.w8(32'hba304d46),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2411fc),
	.w1(32'hbc23e60f),
	.w2(32'h3c3079fb),
	.w3(32'h3c0fde39),
	.w4(32'hbc450518),
	.w5(32'h3c22a53f),
	.w6(32'h3b89708f),
	.w7(32'hbc927b6f),
	.w8(32'h3d21487c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be94892),
	.w1(32'h3b8a7c52),
	.w2(32'hbbace7a1),
	.w3(32'h3c83677f),
	.w4(32'hbcf6bc6a),
	.w5(32'hbbeec8cb),
	.w6(32'hbbc75769),
	.w7(32'hbcdd1768),
	.w8(32'h3d13e425),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb88643),
	.w1(32'h3c8c2062),
	.w2(32'hbc3e58e7),
	.w3(32'hbb4457c1),
	.w4(32'h3c6567c7),
	.w5(32'hbc1848df),
	.w6(32'h3bfe531e),
	.w7(32'hb98f0152),
	.w8(32'h3c004c30),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b255),
	.w1(32'h3a81388e),
	.w2(32'hbc0b7426),
	.w3(32'h3bf01b8c),
	.w4(32'h3c33aaf8),
	.w5(32'h3d0958b6),
	.w6(32'h3c199c2f),
	.w7(32'h3cc076b1),
	.w8(32'hbcf33a7c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceed0fd),
	.w1(32'hbbdc4b20),
	.w2(32'hbce9931a),
	.w3(32'h38cb7f77),
	.w4(32'h3d253279),
	.w5(32'h3d1c9a31),
	.w6(32'hbbc55b1b),
	.w7(32'h3cd76935),
	.w8(32'hbc4d53df),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd60eca1),
	.w1(32'hbd2a4f96),
	.w2(32'hbaccad41),
	.w3(32'hbb9d2770),
	.w4(32'h3c951266),
	.w5(32'hbcb5765d),
	.w6(32'hbca4aed1),
	.w7(32'hbbb2414d),
	.w8(32'hbc21fee6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84d040),
	.w1(32'h3a734fa8),
	.w2(32'h3c228814),
	.w3(32'hbc3eb16c),
	.w4(32'h3c0a8d0b),
	.w5(32'hbc880dc8),
	.w6(32'hbc11aea5),
	.w7(32'h3c9f4024),
	.w8(32'h39f30bcf),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46f5f9),
	.w1(32'h3b89dfae),
	.w2(32'hbb89989b),
	.w3(32'hbacc5713),
	.w4(32'h3cd8c2a1),
	.w5(32'h3bf8ff36),
	.w6(32'hbc232381),
	.w7(32'h3be78a5d),
	.w8(32'hbccd4845),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87c92f),
	.w1(32'hbb0746ec),
	.w2(32'hbb888fcc),
	.w3(32'hbc7f9a82),
	.w4(32'h3b120be4),
	.w5(32'hbadb3ffe),
	.w6(32'h3ad6a1ea),
	.w7(32'hbb4c6d1e),
	.w8(32'hbaa95f3e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ba032),
	.w1(32'hbacd2436),
	.w2(32'hbb6489ab),
	.w3(32'hb9d921e3),
	.w4(32'hbb4411d5),
	.w5(32'h3c6c29e8),
	.w6(32'h39ad11f1),
	.w7(32'hbc48076e),
	.w8(32'h3d0ca5bd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc53a25),
	.w1(32'hbc46dfaf),
	.w2(32'hbc54c649),
	.w3(32'h3bb1ea73),
	.w4(32'h3cbe5b4a),
	.w5(32'h3be1b827),
	.w6(32'hbb3273bc),
	.w7(32'h3c7a877d),
	.w8(32'hbc8e0737),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba35a5),
	.w1(32'hbc0d7ba1),
	.w2(32'hbc077163),
	.w3(32'hbaeceb90),
	.w4(32'hbc132be2),
	.w5(32'hbb68e437),
	.w6(32'h39ced2e5),
	.w7(32'hbbc34755),
	.w8(32'hba941f41),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b788fce),
	.w1(32'h3b906db0),
	.w2(32'h3caac012),
	.w3(32'h3a7b9e0a),
	.w4(32'h3bf626f5),
	.w5(32'hbc92aea9),
	.w6(32'h3c2c4435),
	.w7(32'hbb3d282d),
	.w8(32'h3b5cf8c2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18d1c7),
	.w1(32'h3acc1726),
	.w2(32'hbba2440e),
	.w3(32'hbc2a3300),
	.w4(32'h3b1a2884),
	.w5(32'hb8fc7ca0),
	.w6(32'hbc68ef00),
	.w7(32'hbb6552d7),
	.w8(32'hba592608),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8a502),
	.w1(32'h3aabe5b2),
	.w2(32'hbb9d8320),
	.w3(32'hb988bf84),
	.w4(32'hbbce08bb),
	.w5(32'hb9b143c3),
	.w6(32'h3a867a2a),
	.w7(32'hbcb9bc78),
	.w8(32'h3c3ae246),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a25ad),
	.w1(32'h3c1c06a4),
	.w2(32'hbc893a1d),
	.w3(32'h3c8a0290),
	.w4(32'h3cba300b),
	.w5(32'hbc8a33d9),
	.w6(32'h3c2c071d),
	.w7(32'h3c0b0528),
	.w8(32'hbc894a63),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc209cb),
	.w1(32'hbba8a811),
	.w2(32'hbbeabf31),
	.w3(32'hba41d0b1),
	.w4(32'h3b60af60),
	.w5(32'h3a971d24),
	.w6(32'h3cc63035),
	.w7(32'hbb829863),
	.w8(32'hbb5ac3a1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9be05),
	.w1(32'h38071c8e),
	.w2(32'hbc1d6243),
	.w3(32'h3aaa17bf),
	.w4(32'h3c0c86ff),
	.w5(32'hbc81a19b),
	.w6(32'hbaff4fb0),
	.w7(32'hbb82aae4),
	.w8(32'hbc8a949d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc909f0b),
	.w1(32'hbc1ee145),
	.w2(32'h3aad0dec),
	.w3(32'hbad7cb68),
	.w4(32'hbc1cd6f0),
	.w5(32'h3b5b486f),
	.w6(32'hbbaa046a),
	.w7(32'h3abe4845),
	.w8(32'h3b8b9140),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule