module layer_8_featuremap_226(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15f0af),
	.w1(32'hba41cf6c),
	.w2(32'h3a94be40),
	.w3(32'h3bf55e2f),
	.w4(32'h38edb8bb),
	.w5(32'hbc080d04),
	.w6(32'h3c42fb16),
	.w7(32'hba84f3ea),
	.w8(32'hbb6cd0b5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe634c),
	.w1(32'h3c0c251c),
	.w2(32'h3bbab2ab),
	.w3(32'hbb3253b3),
	.w4(32'h3c02dda6),
	.w5(32'h3bff9307),
	.w6(32'h3c12e4d4),
	.w7(32'h3bdbf9b9),
	.w8(32'h3b9d7436),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99d3d0),
	.w1(32'h3cbf5b90),
	.w2(32'h3d0424b2),
	.w3(32'h3b3ffe45),
	.w4(32'h3c4848a1),
	.w5(32'h3c9b1cf3),
	.w6(32'h3c554ff7),
	.w7(32'h3bd455f2),
	.w8(32'h3c0310d5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5eef6),
	.w1(32'hbb98f9af),
	.w2(32'hbb74354b),
	.w3(32'h3c7005ea),
	.w4(32'hbbaeb8d9),
	.w5(32'hbb95683e),
	.w6(32'h3c2c6010),
	.w7(32'h3b8ff5fa),
	.w8(32'h3bd830bf),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba921e1),
	.w1(32'hbc132595),
	.w2(32'hbc2882cc),
	.w3(32'hbc45ea94),
	.w4(32'hbbdd7197),
	.w5(32'hbbb1f890),
	.w6(32'hbbe90873),
	.w7(32'hbc01005d),
	.w8(32'hbb685fc1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd53004),
	.w1(32'hbc174eae),
	.w2(32'hbc152b9a),
	.w3(32'hbb63a0a6),
	.w4(32'hbbcbd216),
	.w5(32'h3a8292f9),
	.w6(32'hbbfe3d3a),
	.w7(32'hbc21b8ab),
	.w8(32'hbaf35adb),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb98ec7),
	.w1(32'hbc417f9b),
	.w2(32'hbc914fba),
	.w3(32'hbb957f57),
	.w4(32'hbc28f956),
	.w5(32'hbc89f1d3),
	.w6(32'hbb4c96f4),
	.w7(32'hbc20a7cb),
	.w8(32'hbbbb7ffe),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59f507),
	.w1(32'h3c65ceaa),
	.w2(32'h3c1d8b50),
	.w3(32'hbc31aa17),
	.w4(32'h3c05142a),
	.w5(32'h3b0cbcd1),
	.w6(32'h3c3204bd),
	.w7(32'h3b872bff),
	.w8(32'hbb132e35),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55619b),
	.w1(32'h3c2682ec),
	.w2(32'h3c9ace71),
	.w3(32'hbb67d3a9),
	.w4(32'h3bc2ca79),
	.w5(32'h3c7fa1b5),
	.w6(32'h3b87c2b4),
	.w7(32'h3c4737a2),
	.w8(32'h3bb5a45d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be92e11),
	.w1(32'hbb9d289b),
	.w2(32'hbbbf7876),
	.w3(32'h3bdb84d4),
	.w4(32'h3aa36228),
	.w5(32'hbc02fcbd),
	.w6(32'hbb2d457a),
	.w7(32'hbbc1fe45),
	.w8(32'hbbc4bf05),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bc245),
	.w1(32'h3ab41bab),
	.w2(32'hbc0d0970),
	.w3(32'hbbdbb597),
	.w4(32'h3b057bf0),
	.w5(32'hb82bf854),
	.w6(32'hbb893f49),
	.w7(32'h3a32e5be),
	.w8(32'h3b8eb0f0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf43226),
	.w1(32'hbc0d2b4c),
	.w2(32'hbcab56fe),
	.w3(32'hbabe44af),
	.w4(32'hbc167947),
	.w5(32'hbc50460e),
	.w6(32'hbb171b1b),
	.w7(32'hbbcf4cab),
	.w8(32'hbc25b18d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74f024),
	.w1(32'h3b8563b5),
	.w2(32'hbc80ca6f),
	.w3(32'hbc3a1f4a),
	.w4(32'hbb081251),
	.w5(32'hbc85f717),
	.w6(32'h3b9a68ee),
	.w7(32'h3a7c749c),
	.w8(32'hbb124a76),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dc9a2),
	.w1(32'h3c3586b2),
	.w2(32'h3c14890f),
	.w3(32'hbc589272),
	.w4(32'h3b7212ee),
	.w5(32'h3b284def),
	.w6(32'h3c4dfa82),
	.w7(32'h3bc8da42),
	.w8(32'hb7404974),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ebc8e),
	.w1(32'hbb6dbf40),
	.w2(32'hba029afb),
	.w3(32'h3c23e451),
	.w4(32'h3a8a904b),
	.w5(32'h39f90a54),
	.w6(32'hbb621057),
	.w7(32'hbad3aacf),
	.w8(32'hba3d165b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81e0d4),
	.w1(32'hbb400869),
	.w2(32'hbc2734b0),
	.w3(32'h3b963ca5),
	.w4(32'hbb963a5f),
	.w5(32'hbc9582fc),
	.w6(32'h3b9451fc),
	.w7(32'hbb2a965b),
	.w8(32'hbb117f6b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb5ac6),
	.w1(32'h3c4cf7c5),
	.w2(32'h3c2162c4),
	.w3(32'hbb21700e),
	.w4(32'h3c279bef),
	.w5(32'h3c2076b5),
	.w6(32'h3c69da5e),
	.w7(32'h3c1a83a1),
	.w8(32'h3b7cbbe6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccb773),
	.w1(32'h3c9a81ad),
	.w2(32'h3ce094c6),
	.w3(32'h3c44c473),
	.w4(32'h3c269fd9),
	.w5(32'h3cd13762),
	.w6(32'h3c9ef7be),
	.w7(32'h3cc1bf76),
	.w8(32'h3c2d9eae),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c158fa4),
	.w1(32'h3c05f635),
	.w2(32'hba80b4a5),
	.w3(32'h39d5c307),
	.w4(32'hbab53a06),
	.w5(32'hbbe4acbe),
	.w6(32'hbbd602cc),
	.w7(32'hbba5168f),
	.w8(32'hbc869174),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ef5c6),
	.w1(32'h3befee1f),
	.w2(32'h3c12ad46),
	.w3(32'h3b1bfffc),
	.w4(32'h3bd70511),
	.w5(32'h3b2c8e57),
	.w6(32'h3b9fcce3),
	.w7(32'h3c13da40),
	.w8(32'h3b80d3ab),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12b469),
	.w1(32'h3b0adc69),
	.w2(32'hba7a86ce),
	.w3(32'h38a9f9b8),
	.w4(32'hba6d79b0),
	.w5(32'hbbac2500),
	.w6(32'h3be3cbea),
	.w7(32'h3c018d6d),
	.w8(32'h3c10d385),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8c4ac),
	.w1(32'hbb3c4db2),
	.w2(32'h3a9a1913),
	.w3(32'hbb347d93),
	.w4(32'h3b3fdd8d),
	.w5(32'hbb826706),
	.w6(32'hbc063b51),
	.w7(32'h3a57d861),
	.w8(32'hbb989513),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c2240),
	.w1(32'h3c3b1f13),
	.w2(32'h3b4e8cfa),
	.w3(32'hbc8473dc),
	.w4(32'h3b6efb86),
	.w5(32'hbbb160b4),
	.w6(32'hba674f62),
	.w7(32'hbaf21918),
	.w8(32'hbc576e97),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49cd56),
	.w1(32'h3a2dc25b),
	.w2(32'hbc1dc0bc),
	.w3(32'hbc17bbcc),
	.w4(32'h3b7c5321),
	.w5(32'hbb371ffb),
	.w6(32'hbb496b20),
	.w7(32'hbb74f018),
	.w8(32'hbb32e25a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb166697),
	.w1(32'hbb46a6d3),
	.w2(32'hbb8902ae),
	.w3(32'hb884d3bd),
	.w4(32'hbb7eda16),
	.w5(32'hbb3bc68b),
	.w6(32'hbbc22121),
	.w7(32'hbbec224d),
	.w8(32'hbc0db21f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1519b0),
	.w1(32'h3b0dda42),
	.w2(32'hb9e36cd5),
	.w3(32'hbbdbb1ed),
	.w4(32'h3c0a2fc2),
	.w5(32'h3b84f61f),
	.w6(32'h3b3bb176),
	.w7(32'h394bd8a5),
	.w8(32'h3ab6fca5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad51b06),
	.w1(32'h3a2d07e7),
	.w2(32'hbc1ce33a),
	.w3(32'h3a0e612a),
	.w4(32'hbb7abe2f),
	.w5(32'hbc0525e0),
	.w6(32'h3b456779),
	.w7(32'hbbd01081),
	.w8(32'hbc0a1704),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce338b5),
	.w1(32'h3b0d558c),
	.w2(32'h3c6886bb),
	.w3(32'hbc025fbb),
	.w4(32'hbc40c628),
	.w5(32'h3b1e81a4),
	.w6(32'hbb9798f7),
	.w7(32'hbc7e47fd),
	.w8(32'hbc2fb3b6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32d8b6),
	.w1(32'h3ac48791),
	.w2(32'h3b712079),
	.w3(32'hbbab1dfe),
	.w4(32'h3a6cbe14),
	.w5(32'h3aa85898),
	.w6(32'hbbe263b5),
	.w7(32'h3b28d402),
	.w8(32'hb9e42f87),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ee4ae),
	.w1(32'hbbed303f),
	.w2(32'hbbbc1137),
	.w3(32'hbc21c59e),
	.w4(32'hbbbdb413),
	.w5(32'hbb95ed01),
	.w6(32'hbc05bb78),
	.w7(32'hbbe07cc4),
	.w8(32'hb9b55d5c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2eef04),
	.w1(32'hbb9c9a13),
	.w2(32'hb9d08aa4),
	.w3(32'h3b2ac3be),
	.w4(32'hbbce74a5),
	.w5(32'hbbe24933),
	.w6(32'hbad25d3d),
	.w7(32'h398a888b),
	.w8(32'h3b8bfdd2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace994e),
	.w1(32'h3be7c2c9),
	.w2(32'h3b841f18),
	.w3(32'hbbd74518),
	.w4(32'h3bc07fa8),
	.w5(32'h3c0a5176),
	.w6(32'hbbe760fd),
	.w7(32'hbba558de),
	.w8(32'hbc3ecefa),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85ee222),
	.w1(32'h3b869beb),
	.w2(32'h3c68c53c),
	.w3(32'hba7b8a08),
	.w4(32'hb9c7acc7),
	.w5(32'h3bddc55f),
	.w6(32'h3bd5b549),
	.w7(32'h3c306d4d),
	.w8(32'h3ab6d5b4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ed995),
	.w1(32'hbbc1f2a0),
	.w2(32'hbc9625be),
	.w3(32'hba394327),
	.w4(32'hbb319d1f),
	.w5(32'hbc173f15),
	.w6(32'hbc52adbc),
	.w7(32'hbbf33e23),
	.w8(32'hbaa7a5ef),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a8d35),
	.w1(32'h3c31dee0),
	.w2(32'h3c53cb1d),
	.w3(32'hbb60f006),
	.w4(32'h3adcaa79),
	.w5(32'h3c0db4bd),
	.w6(32'h3bb3e558),
	.w7(32'h3c344a36),
	.w8(32'h3ba33a33),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba840b8),
	.w1(32'hbb505fee),
	.w2(32'hbb88825a),
	.w3(32'h3bc19426),
	.w4(32'hbbf1831c),
	.w5(32'hbb5e8b31),
	.w6(32'h3b679dcf),
	.w7(32'hba3a7d5a),
	.w8(32'h3a43ea98),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f9efc),
	.w1(32'h3b3044b9),
	.w2(32'h3bdcbd00),
	.w3(32'h3b25e2f0),
	.w4(32'h39479c84),
	.w5(32'hba0bd7c5),
	.w6(32'h3b93b349),
	.w7(32'h3bf1f534),
	.w8(32'h3bcd8ba9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c191681),
	.w1(32'h3c0c63ed),
	.w2(32'h3cc15466),
	.w3(32'h38cc12b6),
	.w4(32'h3bd6d267),
	.w5(32'h3ca59f59),
	.w6(32'h39954e43),
	.w7(32'h3c7787fa),
	.w8(32'h3c36cb9e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb62811),
	.w1(32'hba84787b),
	.w2(32'hbb8ce7cc),
	.w3(32'h3ca19c59),
	.w4(32'h3b00ea4f),
	.w5(32'hbc0617e9),
	.w6(32'hbad9ceb5),
	.w7(32'h3986f3a2),
	.w8(32'hbad0f9ca),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5db9df),
	.w1(32'hbc7fe10f),
	.w2(32'hbcf7c094),
	.w3(32'hbaa5d4e9),
	.w4(32'hbc63a04c),
	.w5(32'hbc6151de),
	.w6(32'hbbff07b9),
	.w7(32'hbc651b51),
	.w8(32'hbc2b1c52),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80aa28),
	.w1(32'h3cd02504),
	.w2(32'h3cf9705b),
	.w3(32'hbbf53aa5),
	.w4(32'h3cc3f3b3),
	.w5(32'h3cd0d4e0),
	.w6(32'h3c561860),
	.w7(32'h3c9a1786),
	.w8(32'h3c4c2015),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96486a),
	.w1(32'hbc94c20b),
	.w2(32'hbc18d590),
	.w3(32'h3c3542bd),
	.w4(32'hbc9e125a),
	.w5(32'hbc576bd4),
	.w6(32'hbbe6b1e8),
	.w7(32'hbaf2396c),
	.w8(32'h3c244cbd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19aa2a),
	.w1(32'hbc356cc4),
	.w2(32'hbc47775d),
	.w3(32'h3c1db8ac),
	.w4(32'hbc1996ea),
	.w5(32'hbc62469e),
	.w6(32'hbc0a0a69),
	.w7(32'hbc1b1265),
	.w8(32'hbbae02ac),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51f269),
	.w1(32'h3b00d043),
	.w2(32'hbb15ea5b),
	.w3(32'hbbce4637),
	.w4(32'hbbb5d0a4),
	.w5(32'hbb2716ac),
	.w6(32'hbb62c26b),
	.w7(32'hbb50d44d),
	.w8(32'hbbb249f3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4777c2),
	.w1(32'hbc0a9ce5),
	.w2(32'hbc57485f),
	.w3(32'hbc4fda26),
	.w4(32'hbc53cf2a),
	.w5(32'hbc6a4805),
	.w6(32'hbc27be22),
	.w7(32'hbc6a70d0),
	.w8(32'hbc3a2cf2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f178f),
	.w1(32'h3aef8d51),
	.w2(32'hbc281d9a),
	.w3(32'hbca2b0bd),
	.w4(32'hbafc3e60),
	.w5(32'hbc63b15d),
	.w6(32'h3bd0a8d9),
	.w7(32'hbb9b938e),
	.w8(32'hbbb978bf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf217a1),
	.w1(32'hbd649096),
	.w2(32'hbdb83b29),
	.w3(32'hbc1eb3b2),
	.w4(32'hbd0b8d3a),
	.w5(32'hbd8a44d0),
	.w6(32'hbd0b1fc0),
	.w7(32'hbd7d5a4c),
	.w8(32'hbd41024b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9a51d4),
	.w1(32'h3b643d20),
	.w2(32'hbbcce1ce),
	.w3(32'hbd653eb2),
	.w4(32'h3a2d5324),
	.w5(32'hbbafe4ce),
	.w6(32'hbaec0839),
	.w7(32'hbb719b5d),
	.w8(32'hbb16f8aa),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab10c61),
	.w1(32'h3b3840ef),
	.w2(32'h3b8941ff),
	.w3(32'h3a4b43da),
	.w4(32'h3c02ad29),
	.w5(32'h3ae08eba),
	.w6(32'h3b08bd16),
	.w7(32'hbb210c90),
	.w8(32'h3ada7501),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb948dfe6),
	.w1(32'h3c4e0a5d),
	.w2(32'h3c2c12ab),
	.w3(32'hbc3909fb),
	.w4(32'h3bf511b4),
	.w5(32'h3b30c97a),
	.w6(32'h3b8f5dd4),
	.w7(32'h3b6b4ab2),
	.w8(32'hbacae061),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0870cc),
	.w1(32'hbba97483),
	.w2(32'hbc0b46cd),
	.w3(32'h3b1343a9),
	.w4(32'hbb6ec42b),
	.w5(32'hbbfab3da),
	.w6(32'hba11a51d),
	.w7(32'hbb9b7985),
	.w8(32'hb958a429),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f0ec1),
	.w1(32'h3b5ee2ba),
	.w2(32'h399777e6),
	.w3(32'h3ae351c6),
	.w4(32'h3b67cf79),
	.w5(32'hbb191c8a),
	.w6(32'h3ba9b015),
	.w7(32'hbc0b52f4),
	.w8(32'hbb96e888),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb891f37),
	.w1(32'hbc5140c3),
	.w2(32'hbc450f6b),
	.w3(32'hbbb78a1b),
	.w4(32'hbc1a4895),
	.w5(32'hbc179d11),
	.w6(32'hbc0da16c),
	.w7(32'hbc3f66d0),
	.w8(32'hbc1950f3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b8a59),
	.w1(32'hbb05e4ea),
	.w2(32'hbbaff1e2),
	.w3(32'hbbf4ba59),
	.w4(32'h3ba870ef),
	.w5(32'hbc4a1c15),
	.w6(32'h3baa0f57),
	.w7(32'hbb6bcf39),
	.w8(32'hbb647bed),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bab45),
	.w1(32'h3a83d243),
	.w2(32'h3a777d38),
	.w3(32'hbc1bb78e),
	.w4(32'h3a846ec6),
	.w5(32'hbbc12bea),
	.w6(32'h3ae0b74d),
	.w7(32'h3a927be5),
	.w8(32'h3bcedea1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28fc45),
	.w1(32'hbbda003f),
	.w2(32'hbbc5f3ec),
	.w3(32'hbbd31630),
	.w4(32'hbc09d966),
	.w5(32'hbbaea9bd),
	.w6(32'hbc25c91d),
	.w7(32'hbb50fbdf),
	.w8(32'hbc0dd61f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfec1e6),
	.w1(32'h3ba9deab),
	.w2(32'hbbdba4e6),
	.w3(32'h3b03d528),
	.w4(32'h3b9bd9a9),
	.w5(32'hbbf48d1c),
	.w6(32'h3b3e63e8),
	.w7(32'hbbb8e459),
	.w8(32'hbb9e48e4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d4ddb),
	.w1(32'hbbae1e97),
	.w2(32'hbc047f2a),
	.w3(32'hbb855c1e),
	.w4(32'hb91fcfca),
	.w5(32'hbbf0103f),
	.w6(32'hbb7da364),
	.w7(32'hbbbb49b1),
	.w8(32'hbbf1943f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc81eff),
	.w1(32'hbbf90dc1),
	.w2(32'hbc6f55e9),
	.w3(32'hbc15783d),
	.w4(32'hbb58ce19),
	.w5(32'hbbf63973),
	.w6(32'hbc02997f),
	.w7(32'hbc456cbc),
	.w8(32'hbc0d920d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24966d),
	.w1(32'h3b736d61),
	.w2(32'h3bc83568),
	.w3(32'hbb99f3fe),
	.w4(32'h3c4c39ae),
	.w5(32'h3b93346f),
	.w6(32'hb980bed6),
	.w7(32'h3b06fe0c),
	.w8(32'hba04bdac),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0edc1),
	.w1(32'hbb891aec),
	.w2(32'hbc0b3c48),
	.w3(32'hbb415ecb),
	.w4(32'h3ab3cc47),
	.w5(32'hbc028ce3),
	.w6(32'hba05e748),
	.w7(32'hbc608bd1),
	.w8(32'hbc11eca5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3685f1),
	.w1(32'hb92cf263),
	.w2(32'h3b8c1a60),
	.w3(32'hbba3c112),
	.w4(32'hbc44a889),
	.w5(32'hbc90fd7b),
	.w6(32'h3b3736ae),
	.w7(32'h3c261910),
	.w8(32'h3b888ba8),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ff141),
	.w1(32'h3cc633e1),
	.w2(32'h3d57316b),
	.w3(32'hbc695bc6),
	.w4(32'h3c401cf8),
	.w5(32'h3d1cc8ad),
	.w6(32'h3a69c52c),
	.w7(32'h3cf9fafc),
	.w8(32'h3c953177),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d26bd74),
	.w1(32'hbc0e339a),
	.w2(32'hbc535a25),
	.w3(32'h3cc98fa0),
	.w4(32'hbc2169ca),
	.w5(32'hbc5d8fcb),
	.w6(32'hbc0ed42a),
	.w7(32'hbc3ada19),
	.w8(32'hbc4398a0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78ae88),
	.w1(32'h3b83a397),
	.w2(32'h3bdfb48d),
	.w3(32'hbc65ecef),
	.w4(32'h3b6e870c),
	.w5(32'h3bc2e09e),
	.w6(32'h3adfa24e),
	.w7(32'h3b993502),
	.w8(32'h3bc8e5af),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08bb38),
	.w1(32'hbc8e26cc),
	.w2(32'hbd01bd98),
	.w3(32'h3bc2ed52),
	.w4(32'hbc5aef56),
	.w5(32'hbca4e00f),
	.w6(32'hbbc137b5),
	.w7(32'hbc666f7f),
	.w8(32'hbc792dd2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2b122),
	.w1(32'hbc234f0e),
	.w2(32'hbcad3ef2),
	.w3(32'hbc2c13e2),
	.w4(32'hbc364719),
	.w5(32'hbc8d7171),
	.w6(32'h3b5e6c3f),
	.w7(32'hbc45ca3a),
	.w8(32'hbc431382),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2440f),
	.w1(32'hbcd8c35d),
	.w2(32'hbd3cdadd),
	.w3(32'hbc670d87),
	.w4(32'hbc674e7d),
	.w5(32'hbcefc712),
	.w6(32'hbbdfbe50),
	.w7(32'hbc952c9e),
	.w8(32'hbc15de63),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce80b6f),
	.w1(32'h3b7322fd),
	.w2(32'hb9ffbc8f),
	.w3(32'hbc6022cd),
	.w4(32'h3ac01312),
	.w5(32'h3b338785),
	.w6(32'h3bbe3d13),
	.w7(32'h3bc7974f),
	.w8(32'h3b0e5d95),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60294f),
	.w1(32'h3d082788),
	.w2(32'h3d374aa2),
	.w3(32'h3a938db6),
	.w4(32'h3c9bf798),
	.w5(32'h3ce3be3a),
	.w6(32'h3b6ec86f),
	.w7(32'h3c8373e6),
	.w8(32'h3c735879),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd07379),
	.w1(32'h3b6af696),
	.w2(32'h3afa49e1),
	.w3(32'h3b97c945),
	.w4(32'h3aa03d3d),
	.w5(32'h3bb047b2),
	.w6(32'h3b285681),
	.w7(32'hba933d65),
	.w8(32'hbc2189f7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc127643),
	.w1(32'h3ad64075),
	.w2(32'hbb7658bd),
	.w3(32'h3b4a0fdc),
	.w4(32'h38b23f2e),
	.w5(32'h3bfd4840),
	.w6(32'h3bc416df),
	.w7(32'hbafcd9e0),
	.w8(32'h3b8d5445),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c4bd0),
	.w1(32'hbbb5883f),
	.w2(32'hbb6cc484),
	.w3(32'h3b8fb1dd),
	.w4(32'hbb41ffb1),
	.w5(32'hbbc6c49f),
	.w6(32'h3b0c12df),
	.w7(32'h3b9663b7),
	.w8(32'h3b1e0a89),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f314f),
	.w1(32'hbc1346b1),
	.w2(32'hbbf10236),
	.w3(32'h383857e0),
	.w4(32'hbb572a72),
	.w5(32'hbc625c6e),
	.w6(32'hbbf7505d),
	.w7(32'hbbf10584),
	.w8(32'hbc18015a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c0f43),
	.w1(32'hbb49f6b4),
	.w2(32'hbbd92a4b),
	.w3(32'hbc94682a),
	.w4(32'hba883b15),
	.w5(32'hbc477ec7),
	.w6(32'hb91c1a7f),
	.w7(32'hbb856e7e),
	.w8(32'hb915df1d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5068a7),
	.w1(32'h3ca6837f),
	.w2(32'h3d0fa998),
	.w3(32'hbc183350),
	.w4(32'h3c68c180),
	.w5(32'h3caa3144),
	.w6(32'h3c34a279),
	.w7(32'h3ccab5bb),
	.w8(32'h3c35c652),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82d0fd),
	.w1(32'hbc15647f),
	.w2(32'hbc995e77),
	.w3(32'h3c0a6750),
	.w4(32'hbbba5b8d),
	.w5(32'hbc836d61),
	.w6(32'hbb4e83f9),
	.w7(32'hbc1f81f3),
	.w8(32'hb9e57478),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f3e52),
	.w1(32'hbbedcfeb),
	.w2(32'hbbe10609),
	.w3(32'hbbd21120),
	.w4(32'hbc2cc3dd),
	.w5(32'hbc64bafc),
	.w6(32'hbb8cee03),
	.w7(32'hbae85210),
	.w8(32'h3b70e5a7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf49aa),
	.w1(32'hbb396405),
	.w2(32'hbb9ea332),
	.w3(32'hbc0a1eef),
	.w4(32'hbbf345e3),
	.w5(32'hbc044c81),
	.w6(32'h3c1a6750),
	.w7(32'hbba512fd),
	.w8(32'hbb58d0a9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3340a1),
	.w1(32'h3b1b9529),
	.w2(32'hbb959ab2),
	.w3(32'h3b08be7c),
	.w4(32'h3ae8cd60),
	.w5(32'h3a4f2bf7),
	.w6(32'h3ae3d24e),
	.w7(32'hbb01d67b),
	.w8(32'hbb23102a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2c7cb),
	.w1(32'h3c533132),
	.w2(32'h3cbd9b6a),
	.w3(32'hbc0db5e9),
	.w4(32'h3c224956),
	.w5(32'h3c973831),
	.w6(32'h3c8de604),
	.w7(32'h3c80ef9f),
	.w8(32'h3bd90c1c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c674285),
	.w1(32'hbb8ff54c),
	.w2(32'hba282ec1),
	.w3(32'h3c138d8b),
	.w4(32'h3bf0fea4),
	.w5(32'h3bcb605c),
	.w6(32'h3b53904f),
	.w7(32'hbb786797),
	.w8(32'h3b5c9e31),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad98a53),
	.w1(32'h3ccdef66),
	.w2(32'h3d0f8450),
	.w3(32'h3c21c302),
	.w4(32'h3c718bdf),
	.w5(32'h3c9e0061),
	.w6(32'h3c39c245),
	.w7(32'h3c9b047d),
	.w8(32'h3c10a2c2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fe096),
	.w1(32'hbc428695),
	.w2(32'hbb8bd7ac),
	.w3(32'h3b8857e1),
	.w4(32'h3a8e2fd8),
	.w5(32'hba52a1a1),
	.w6(32'hbb2ced7e),
	.w7(32'hbb2863aa),
	.w8(32'hbb75ae5c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e19bc),
	.w1(32'h3cacedbb),
	.w2(32'h3d0deeda),
	.w3(32'h3aceb988),
	.w4(32'h3c59b49d),
	.w5(32'h3ca0fc60),
	.w6(32'h3c49c55d),
	.w7(32'h3c124737),
	.w8(32'hbb39c21f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a5ce5),
	.w1(32'h3b665dac),
	.w2(32'hbb325671),
	.w3(32'h3c35b456),
	.w4(32'h3b171198),
	.w5(32'hbb5c4019),
	.w6(32'h3b0719f6),
	.w7(32'h3acef929),
	.w8(32'h3c35e0be),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fb176),
	.w1(32'h3a852195),
	.w2(32'h3b10546c),
	.w3(32'hbb0e6814),
	.w4(32'h3b72efdc),
	.w5(32'h3c24b1cb),
	.w6(32'hba2139c7),
	.w7(32'hbb1c76f2),
	.w8(32'hbbcf8c49),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e11731),
	.w1(32'hbb8cad21),
	.w2(32'hba6ea678),
	.w3(32'h3bcac498),
	.w4(32'h3ba7480a),
	.w5(32'h3bea2498),
	.w6(32'hbb94a681),
	.w7(32'hbb81af2c),
	.w8(32'hbb393e4e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90be3c),
	.w1(32'h3b0a2c3d),
	.w2(32'hb9f75869),
	.w3(32'h3c088739),
	.w4(32'hbaf5dab1),
	.w5(32'hba9d5b6c),
	.w6(32'h3ae3054a),
	.w7(32'hbb4bea25),
	.w8(32'hbad8f6d6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38c70c),
	.w1(32'h3c91dc53),
	.w2(32'h3ceb47e1),
	.w3(32'hbb3e7ce0),
	.w4(32'h3c0916fc),
	.w5(32'h3c83b45a),
	.w6(32'h3b79ccd1),
	.w7(32'h3c676c8a),
	.w8(32'h3c210c03),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81b54c),
	.w1(32'hbbe9b851),
	.w2(32'hbc48d80e),
	.w3(32'h3c3e52f8),
	.w4(32'hbbc2d0ad),
	.w5(32'hbbd2d595),
	.w6(32'h3a9da14b),
	.w7(32'hbb859319),
	.w8(32'h3b3c3827),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb822b3d),
	.w1(32'hbcb6d502),
	.w2(32'hbd0d3d25),
	.w3(32'h3bd327d3),
	.w4(32'hbbd3f1d1),
	.w5(32'hbca61ee4),
	.w6(32'hbc1d2f13),
	.w7(32'hbc76a678),
	.w8(32'hbb6b5aae),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65780b),
	.w1(32'h3b5a7bd4),
	.w2(32'hbb589c18),
	.w3(32'hbb4e2c7b),
	.w4(32'h3bec5b74),
	.w5(32'h3b2846d2),
	.w6(32'h3b0bf24a),
	.w7(32'h3aadfac5),
	.w8(32'hb9b18d08),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a93fc),
	.w1(32'hbc20e16a),
	.w2(32'hbcbec336),
	.w3(32'hbb287795),
	.w4(32'hbc0370df),
	.w5(32'hbc9348cb),
	.w6(32'hbbac5385),
	.w7(32'hbc898fbd),
	.w8(32'hbc8bee39),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc36161),
	.w1(32'hbbba4a6b),
	.w2(32'hbc786bd7),
	.w3(32'hbc9cc00a),
	.w4(32'h3b604405),
	.w5(32'hbc6224ce),
	.w6(32'hba52f8ca),
	.w7(32'hbbdb688e),
	.w8(32'hbb4581a6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bdcee),
	.w1(32'hbc1f60d7),
	.w2(32'hbbaeca1b),
	.w3(32'hbba2b0f4),
	.w4(32'h3b0628c2),
	.w5(32'h3b5c1619),
	.w6(32'hbc37ff06),
	.w7(32'hbbf295d0),
	.w8(32'h3adf073e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86cc00),
	.w1(32'h3ca70ac5),
	.w2(32'h3ca0ddfa),
	.w3(32'h3c1424b3),
	.w4(32'h3b2af9d9),
	.w5(32'h3bf0aa87),
	.w6(32'hba638fec),
	.w7(32'h3c5131a5),
	.w8(32'h3c5e11ac),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25f513),
	.w1(32'h3bd53f11),
	.w2(32'h3c89c1b8),
	.w3(32'h3c1a2a52),
	.w4(32'h3bec34bd),
	.w5(32'h3c634a37),
	.w6(32'h3c11157d),
	.w7(32'h3c7c47c2),
	.w8(32'h3b7070de),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22611c),
	.w1(32'hbb3a437e),
	.w2(32'hbc1a1bee),
	.w3(32'h3c1d3850),
	.w4(32'hba8a847d),
	.w5(32'hbc1a12d7),
	.w6(32'h3b520ec7),
	.w7(32'hbad986f0),
	.w8(32'hbc149403),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44a332),
	.w1(32'hbaf4919b),
	.w2(32'hbc6a2f3d),
	.w3(32'hbbc1684d),
	.w4(32'h3a9bdf78),
	.w5(32'hbc12c618),
	.w6(32'hba86ed4e),
	.w7(32'hbc0b98d3),
	.w8(32'hbb7abab0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb7bc3),
	.w1(32'h3aea52fe),
	.w2(32'h3b901797),
	.w3(32'hbc53e91e),
	.w4(32'h3bb9dfca),
	.w5(32'h3b900fc3),
	.w6(32'h3c11a51b),
	.w7(32'h3b7885a1),
	.w8(32'h3be2ae9f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeffc8),
	.w1(32'h3bab2651),
	.w2(32'h3c767a90),
	.w3(32'hbbbcc063),
	.w4(32'h3bdb8272),
	.w5(32'h3bf3876d),
	.w6(32'hbb0c205d),
	.w7(32'h3c16e73a),
	.w8(32'h3b6df517),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e811b),
	.w1(32'hbbce455b),
	.w2(32'hbc783187),
	.w3(32'hba4a3c35),
	.w4(32'hbc18a4a5),
	.w5(32'hbc557aff),
	.w6(32'h39b47e31),
	.w7(32'hbb5e1b22),
	.w8(32'h3b642b86),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d4a8c),
	.w1(32'h3b242b6b),
	.w2(32'h39d436b7),
	.w3(32'hbb2c4b4f),
	.w4(32'h3bd5e1e8),
	.w5(32'h3c30307b),
	.w6(32'h3a943cc8),
	.w7(32'h3b161167),
	.w8(32'hbb92d424),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07e500),
	.w1(32'hbb0e4427),
	.w2(32'hbbee2f3b),
	.w3(32'h3a47b5d3),
	.w4(32'h3b9ad99f),
	.w5(32'hbac7a588),
	.w6(32'h3b87aa28),
	.w7(32'hbb979292),
	.w8(32'hbaa99643),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8987cf),
	.w1(32'hb820fc49),
	.w2(32'hbc188b9b),
	.w3(32'h3adbe75b),
	.w4(32'hba2c2662),
	.w5(32'hbb40fc3a),
	.w6(32'hbb0d0db3),
	.w7(32'hbc1368d8),
	.w8(32'hbadf317d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1450b),
	.w1(32'h3982e348),
	.w2(32'hb9708af8),
	.w3(32'hb9c1deee),
	.w4(32'h3b8a9f38),
	.w5(32'h3ba51a18),
	.w6(32'h3adea9dd),
	.w7(32'hbb7558ff),
	.w8(32'hbbc32787),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00768e),
	.w1(32'h3a60ecc4),
	.w2(32'h3addec5a),
	.w3(32'hbbc49e1c),
	.w4(32'hbbb395cf),
	.w5(32'hbb3a48d3),
	.w6(32'h3b8f6b23),
	.w7(32'hba87df93),
	.w8(32'hbbb7aaa0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3804a4),
	.w1(32'hbbd75169),
	.w2(32'hbc8b5d18),
	.w3(32'hbba4f4f6),
	.w4(32'h3b4bfbec),
	.w5(32'h39034758),
	.w6(32'h3ae737ea),
	.w7(32'hbae9c875),
	.w8(32'h3c3ec053),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9615f),
	.w1(32'hbad8d2ff),
	.w2(32'h398be11b),
	.w3(32'h3c8c941a),
	.w4(32'hbaeb3aaa),
	.w5(32'h3afaf88f),
	.w6(32'hbb0e0308),
	.w7(32'h397d7cf3),
	.w8(32'h3b37efc6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4509d),
	.w1(32'hbc3af852),
	.w2(32'hbc89c428),
	.w3(32'h3bb3db00),
	.w4(32'hbc057725),
	.w5(32'hbbd12802),
	.w6(32'h3ac26aa1),
	.w7(32'h3b26ab89),
	.w8(32'hba62a145),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc305883),
	.w1(32'hbbb6725b),
	.w2(32'hbc34f18f),
	.w3(32'hbb3577d6),
	.w4(32'hbc1ed218),
	.w5(32'hbc320677),
	.w6(32'hbb4a8be0),
	.w7(32'hbb9bb0db),
	.w8(32'hbb796289),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c21c3),
	.w1(32'h3ca53c57),
	.w2(32'h3cd1f022),
	.w3(32'hbc6a8725),
	.w4(32'h3c9d692b),
	.w5(32'h3cc6ae01),
	.w6(32'h3c9d6504),
	.w7(32'h3d03494e),
	.w8(32'h3c7b9a72),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88480a),
	.w1(32'hbbe47c92),
	.w2(32'h3a9cbdba),
	.w3(32'h3c6d535d),
	.w4(32'hbaeb6311),
	.w5(32'hbb1ddf53),
	.w6(32'h3bbe30dd),
	.w7(32'h3c0fce10),
	.w8(32'h3bacb52e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8e03b),
	.w1(32'hba9011db),
	.w2(32'hbb58d16a),
	.w3(32'hbba94635),
	.w4(32'hbbb7fa16),
	.w5(32'hbbb3bc77),
	.w6(32'hbb2c1f5e),
	.w7(32'hbbc43a16),
	.w8(32'hbb4eb504),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e3f4b),
	.w1(32'hbb1c8753),
	.w2(32'h3b0d897d),
	.w3(32'hbb263db0),
	.w4(32'hbaf4c744),
	.w5(32'h3ae5ea5d),
	.w6(32'hbb8064df),
	.w7(32'hba8fa015),
	.w8(32'hba90c123),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbd5b0),
	.w1(32'h3c865116),
	.w2(32'h3c8eace9),
	.w3(32'h3ab61cdc),
	.w4(32'h3bf98fa0),
	.w5(32'h3b896bb1),
	.w6(32'h3bcf4f7d),
	.w7(32'h3c10c5a4),
	.w8(32'h3b79769a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43aa1d),
	.w1(32'h3c87dda3),
	.w2(32'h3cb0495f),
	.w3(32'hbb726ab1),
	.w4(32'h3c27f8bc),
	.w5(32'h3c8dfecb),
	.w6(32'h3bd3b7db),
	.w7(32'h3c80d383),
	.w8(32'h3c07fc19),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9347d0),
	.w1(32'hbbbe962d),
	.w2(32'hbb9b1400),
	.w3(32'h3c3cc912),
	.w4(32'hbc113ed9),
	.w5(32'hbc32846f),
	.w6(32'hbb4e79e3),
	.w7(32'hbac8ea45),
	.w8(32'hbbc2bd5b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc24fd2),
	.w1(32'hbc4996e7),
	.w2(32'hbc3f490f),
	.w3(32'h3b1c690c),
	.w4(32'hbc483585),
	.w5(32'hbc2facc0),
	.w6(32'hbc3d2601),
	.w7(32'hbbdd796a),
	.w8(32'hbba1eb46),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc093ac3),
	.w1(32'hbbba2c6a),
	.w2(32'hbbbe7344),
	.w3(32'hbb697ef9),
	.w4(32'hbab80ac5),
	.w5(32'hbad5ef4d),
	.w6(32'hbbcacb95),
	.w7(32'hbbafe5bd),
	.w8(32'h3bb0456a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b008b08),
	.w1(32'hbb79d7c7),
	.w2(32'hbc4a77ee),
	.w3(32'h3ba3da69),
	.w4(32'hbbb060e9),
	.w5(32'hbc0a9f63),
	.w6(32'hb94f345b),
	.w7(32'hbc2c0d62),
	.w8(32'hbc749beb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46ff7c),
	.w1(32'h3a84ea58),
	.w2(32'hbc0d5397),
	.w3(32'hbbd6a3f5),
	.w4(32'h3a603805),
	.w5(32'hbb4c3229),
	.w6(32'h3b4d36fa),
	.w7(32'hbb851439),
	.w8(32'hbb57f545),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe81ae1),
	.w1(32'h3c7651f3),
	.w2(32'h3caaf83d),
	.w3(32'hbbbd21bb),
	.w4(32'h3c006a5b),
	.w5(32'h3ca89e78),
	.w6(32'h3bdda94f),
	.w7(32'h3ca562a9),
	.w8(32'h3b6dba96),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c325fd2),
	.w1(32'hba0ed0c0),
	.w2(32'h3a9b3c34),
	.w3(32'h3c28d50f),
	.w4(32'h3c0df6c9),
	.w5(32'hba19034e),
	.w6(32'hbabde7da),
	.w7(32'h3b839943),
	.w8(32'hba8d72db),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74a612),
	.w1(32'hbb00acfd),
	.w2(32'hbb9ceba8),
	.w3(32'hbc0753c3),
	.w4(32'h3b35f76b),
	.w5(32'hbaa45c4f),
	.w6(32'h3ae05d06),
	.w7(32'hbb5d4881),
	.w8(32'hbb887f43),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb270f8d),
	.w1(32'hba6dba1b),
	.w2(32'hbadfb71d),
	.w3(32'hbbb971d5),
	.w4(32'hbab9c266),
	.w5(32'hbb107301),
	.w6(32'hb9fdb3bf),
	.w7(32'hbaacabf8),
	.w8(32'hba8efc68),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabff213),
	.w1(32'hba72efd3),
	.w2(32'h3c02ae82),
	.w3(32'hbba26a1f),
	.w4(32'hbc068e10),
	.w5(32'h3ba8d622),
	.w6(32'hbbda1830),
	.w7(32'h3a9103ec),
	.w8(32'hbc36489c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule