module layer_10_featuremap_36(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23ab79),
	.w1(32'h3bbf2c11),
	.w2(32'h3bd74c11),
	.w3(32'hba8d327e),
	.w4(32'h3b1184d7),
	.w5(32'h3bf2740c),
	.w6(32'h3b00b36a),
	.w7(32'h3bcfdd1b),
	.w8(32'h3c674b20),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4993d),
	.w1(32'h3b8e079f),
	.w2(32'h3b05e60b),
	.w3(32'h3c95a62b),
	.w4(32'h3b448406),
	.w5(32'h3a0b707b),
	.w6(32'h3c86dd8f),
	.w7(32'h3c277ffa),
	.w8(32'h3ae1d6b0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4baddb),
	.w1(32'hbc479879),
	.w2(32'hbb1b34e6),
	.w3(32'hbcc7f6df),
	.w4(32'hbd0dd1c4),
	.w5(32'h3bfeb684),
	.w6(32'hbcb1d4e8),
	.w7(32'hbcda5e49),
	.w8(32'h3bfa71a6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52a0f),
	.w1(32'hbb018d61),
	.w2(32'hbc32d15e),
	.w3(32'h3c19d914),
	.w4(32'h3a654c33),
	.w5(32'hbaef5aca),
	.w6(32'h3c5673b2),
	.w7(32'h3bea2b7e),
	.w8(32'h3baff7cd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1920f7),
	.w1(32'h3bc12e3c),
	.w2(32'hbca479d6),
	.w3(32'h3ad590db),
	.w4(32'h3c17ef30),
	.w5(32'hbcdc42a3),
	.w6(32'hba483954),
	.w7(32'hbba71593),
	.w8(32'hbc402100),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7565d2),
	.w1(32'h3ba49c47),
	.w2(32'hbb1975a9),
	.w3(32'hbc19fa82),
	.w4(32'hbb3ce835),
	.w5(32'hba8a3ae4),
	.w6(32'hbc351134),
	.w7(32'hbc523fba),
	.w8(32'hba07d267),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ec015),
	.w1(32'h3acf4fb0),
	.w2(32'hba685916),
	.w3(32'h3bca22cb),
	.w4(32'h3bbc82a2),
	.w5(32'hb9c555e6),
	.w6(32'h3b9c7152),
	.w7(32'hb98595e3),
	.w8(32'h3a749886),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a072ad4),
	.w1(32'h3bc324c7),
	.w2(32'hbb2b256a),
	.w3(32'hbabc198a),
	.w4(32'h3c0d406f),
	.w5(32'h3a5e3cb6),
	.w6(32'h3ac634fb),
	.w7(32'h3c2559bd),
	.w8(32'h3bfe5147),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d10da),
	.w1(32'h3c5b533b),
	.w2(32'hbbfe7fe2),
	.w3(32'h3a09c24f),
	.w4(32'h3b9e0d35),
	.w5(32'h3b9777fa),
	.w6(32'h3a6d9372),
	.w7(32'hba95792b),
	.w8(32'hbbff2830),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a34412),
	.w1(32'hbc283874),
	.w2(32'hbb0a2d42),
	.w3(32'hb9b83ba6),
	.w4(32'hbc76d8ce),
	.w5(32'h3b67f150),
	.w6(32'hbc5e484c),
	.w7(32'hbc88195c),
	.w8(32'h3a966434),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a872496),
	.w1(32'hbb39a002),
	.w2(32'h3b9582b2),
	.w3(32'h3b4b58be),
	.w4(32'hbbc2ea39),
	.w5(32'h3be0b128),
	.w6(32'h3aa34cfe),
	.w7(32'hbbc9470b),
	.w8(32'h3c0a2f69),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab02d53),
	.w1(32'h3b3b19ea),
	.w2(32'h3ada72cc),
	.w3(32'h3c41b81f),
	.w4(32'h3bb06b7a),
	.w5(32'h3b281503),
	.w6(32'h3c493481),
	.w7(32'h3af3c2b5),
	.w8(32'h38668742),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b849520),
	.w1(32'h3ade0cdf),
	.w2(32'h3a9d38db),
	.w3(32'h3b85320e),
	.w4(32'h3bbd1f5f),
	.w5(32'h3bf040d0),
	.w6(32'h3af272c3),
	.w7(32'h3b7e49f5),
	.w8(32'h3a245fd0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bdbf0),
	.w1(32'hbab5a0a8),
	.w2(32'hbc3ab154),
	.w3(32'h3be1548b),
	.w4(32'hbbb1c135),
	.w5(32'hbbf9e81f),
	.w6(32'h3aae5088),
	.w7(32'h3bb270f4),
	.w8(32'hba92e5c1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04085f),
	.w1(32'h3b83a69d),
	.w2(32'hb93793c9),
	.w3(32'hbc7812c4),
	.w4(32'hbc16952b),
	.w5(32'hb89b5e2d),
	.w6(32'hbc054fbc),
	.w7(32'hbc1a0bfc),
	.w8(32'hbb202fdd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5370a),
	.w1(32'h3bee7aa1),
	.w2(32'h3ba131e1),
	.w3(32'h3c4708d8),
	.w4(32'h3c2cc48f),
	.w5(32'h3bd4bacd),
	.w6(32'h3b65d2e7),
	.w7(32'h3bf245c9),
	.w8(32'h3b91e426),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc57d2),
	.w1(32'h39efb9d8),
	.w2(32'hbb80b17a),
	.w3(32'h3b51392a),
	.w4(32'hbbb448b7),
	.w5(32'h3ae871a6),
	.w6(32'h3a72314a),
	.w7(32'hbbb2c560),
	.w8(32'hbc191469),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0379dd),
	.w1(32'h3bc8c331),
	.w2(32'hbb912d59),
	.w3(32'h3bcab5f4),
	.w4(32'h3c4030d1),
	.w5(32'h3b33d384),
	.w6(32'hbbe56ef9),
	.w7(32'hbba74513),
	.w8(32'h3a6b1a00),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52cbf4),
	.w1(32'hbae0aca8),
	.w2(32'hbcdbdd64),
	.w3(32'h3b6d4ba7),
	.w4(32'hbb1413cd),
	.w5(32'hbc541228),
	.w6(32'h3b9b23f0),
	.w7(32'hbab58b37),
	.w8(32'hbb8fd9e1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d4cc0),
	.w1(32'hbc925b7e),
	.w2(32'hbc0413be),
	.w3(32'hbc187952),
	.w4(32'hbc024958),
	.w5(32'hbbfa9080),
	.w6(32'h3a12df88),
	.w7(32'h3b7c0d59),
	.w8(32'h3ab1e250),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb028a3f),
	.w1(32'h3bab4615),
	.w2(32'h3c00a24b),
	.w3(32'h3bb28d63),
	.w4(32'h3c3622e8),
	.w5(32'h3c16abd3),
	.w6(32'h3c1284ee),
	.w7(32'h3b90d713),
	.w8(32'h3c3e9b4b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43b0f5),
	.w1(32'h3a268618),
	.w2(32'hbc1f2893),
	.w3(32'h3cc2e819),
	.w4(32'h3ca6dc0c),
	.w5(32'hbc973037),
	.w6(32'h3cc8113e),
	.w7(32'h3cb7c08c),
	.w8(32'hbb952685),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90be23a),
	.w1(32'h3a9849cf),
	.w2(32'hba5d55da),
	.w3(32'h3a5a9b14),
	.w4(32'h3bb3e732),
	.w5(32'h3b37147a),
	.w6(32'h3b5626cc),
	.w7(32'h3b479a5f),
	.w8(32'h3af1e1e2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a2c0d),
	.w1(32'hb9c37f0f),
	.w2(32'h39ef6d35),
	.w3(32'h3bb9b498),
	.w4(32'h3b495684),
	.w5(32'h3a98755c),
	.w6(32'h3b5d0387),
	.w7(32'h39b4cf33),
	.w8(32'h3beba973),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ed84f),
	.w1(32'h3b8da81a),
	.w2(32'hba47473d),
	.w3(32'h3bbd4933),
	.w4(32'h3b65fdf4),
	.w5(32'hbb989c7f),
	.w6(32'h3b53b424),
	.w7(32'h3b580dca),
	.w8(32'h3c114231),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a393d),
	.w1(32'hbc0c38a0),
	.w2(32'hbad0a318),
	.w3(32'hbb871bae),
	.w4(32'hbb856dfc),
	.w5(32'h3b3685a3),
	.w6(32'h3bcd01b3),
	.w7(32'h3a0c10a7),
	.w8(32'h3bea9acf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4193a1),
	.w1(32'h3b8c5e59),
	.w2(32'h3c347e6e),
	.w3(32'h3bcaaed0),
	.w4(32'h3c1aa748),
	.w5(32'h3c0478c1),
	.w6(32'h3b6f620d),
	.w7(32'h3b9d9f69),
	.w8(32'h3bbfa8f0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde8926),
	.w1(32'hbbe0d1ee),
	.w2(32'h3bdccddc),
	.w3(32'hbce82c81),
	.w4(32'hbc97c931),
	.w5(32'h3bef5172),
	.w6(32'hbc90d1c7),
	.w7(32'hbc542d5c),
	.w8(32'h3b60ac7c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa79da),
	.w1(32'h3a3ec5cf),
	.w2(32'h39f40403),
	.w3(32'h3c96facb),
	.w4(32'hbb936466),
	.w5(32'hba5fa132),
	.w6(32'h3c3ca007),
	.w7(32'hbb858434),
	.w8(32'hbbcdcdc0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4f3cc),
	.w1(32'hbb3a2bf4),
	.w2(32'h3cb4bf27),
	.w3(32'h39a8c993),
	.w4(32'hbaf7b87c),
	.w5(32'h3b91eca1),
	.w6(32'h39200eb2),
	.w7(32'h3aafc157),
	.w8(32'h3c8dd8a2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b052916),
	.w1(32'h3babb9c4),
	.w2(32'hbb677852),
	.w3(32'hbcf37485),
	.w4(32'hbcbad1dc),
	.w5(32'hbb89c018),
	.w6(32'hbc878f9d),
	.w7(32'hbc3adb14),
	.w8(32'hbaaf7e7e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71c13a),
	.w1(32'h3ade018d),
	.w2(32'hbb8ff9b0),
	.w3(32'hbb035677),
	.w4(32'hb99a88a7),
	.w5(32'h3a3e9b8e),
	.w6(32'h38880d03),
	.w7(32'h3a93440d),
	.w8(32'hbb91ba03),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0db476),
	.w1(32'hbbe025a4),
	.w2(32'hbc8b8eb3),
	.w3(32'h3a6b0ca4),
	.w4(32'hbb82cc0d),
	.w5(32'hbd1484c9),
	.w6(32'h3b95b9be),
	.w7(32'h3bba94b5),
	.w8(32'hbbf6d841),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fba8e),
	.w1(32'h3c71c3f0),
	.w2(32'hbb348dc0),
	.w3(32'hbc70420b),
	.w4(32'h3ca1e061),
	.w5(32'h3974c0e8),
	.w6(32'h3b5a2927),
	.w7(32'h3cd52bb9),
	.w8(32'hbbe4d6ab),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4b924),
	.w1(32'h3bc1531b),
	.w2(32'hbc853ff6),
	.w3(32'hbb8b183e),
	.w4(32'h3c0f4adb),
	.w5(32'hbb29cff4),
	.w6(32'h38ab8232),
	.w7(32'h3b57c20f),
	.w8(32'hbbed9832),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddb7f8),
	.w1(32'h3c09fc6c),
	.w2(32'h3c176508),
	.w3(32'h3d1ab133),
	.w4(32'h3d09e7f4),
	.w5(32'h3be3e600),
	.w6(32'h3ce01382),
	.w7(32'h3ccb30a3),
	.w8(32'h3c0145d4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2641bc),
	.w1(32'hbba3e04a),
	.w2(32'hbce8ecd5),
	.w3(32'h3b59b458),
	.w4(32'h3ab42fad),
	.w5(32'hbd124f57),
	.w6(32'h3ab578ee),
	.w7(32'h3a2a2d2d),
	.w8(32'hbc368fc1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffb747),
	.w1(32'h3cdabecd),
	.w2(32'h3a90e51d),
	.w3(32'h3c022ed7),
	.w4(32'h3d34baa2),
	.w5(32'h3bcccbfb),
	.w6(32'h3c91c9bc),
	.w7(32'h3d3f6906),
	.w8(32'h38924c91),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf2cca),
	.w1(32'hbabc1ac9),
	.w2(32'hb8c342c8),
	.w3(32'h3badc45e),
	.w4(32'h3a87c698),
	.w5(32'hba9a2e23),
	.w6(32'h3baccbcf),
	.w7(32'h3afc5a44),
	.w8(32'hbbd516f0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918b9a7),
	.w1(32'h3b547f7c),
	.w2(32'h3b3b6cb1),
	.w3(32'hbbe5af74),
	.w4(32'h3bdb12e5),
	.w5(32'h3ad19114),
	.w6(32'hbbccf5b2),
	.w7(32'h3b078430),
	.w8(32'h3b0afe6a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eb4b2),
	.w1(32'h3b107f2f),
	.w2(32'hba7f9fa0),
	.w3(32'h3bfe51f3),
	.w4(32'h3bbc312e),
	.w5(32'hbba05ffb),
	.w6(32'h3b8ee116),
	.w7(32'h3b3f9cb8),
	.w8(32'hbae6cd91),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa602ee),
	.w1(32'h3bc74e54),
	.w2(32'hbaf7c48b),
	.w3(32'hb90a0465),
	.w4(32'h3bd92224),
	.w5(32'h3aeda6ff),
	.w6(32'h3ba34f55),
	.w7(32'h3bdd4d3f),
	.w8(32'hbb98e2f7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae642b),
	.w1(32'h3b21404b),
	.w2(32'h3cf419d9),
	.w3(32'h3ab0b523),
	.w4(32'hba9c3332),
	.w5(32'h3d2dd555),
	.w6(32'h3b8d34ed),
	.w7(32'hbae3a2d7),
	.w8(32'h3cbf7ccb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb939d8f),
	.w1(32'hbd27f5e2),
	.w2(32'h3b544bf5),
	.w3(32'hbcad17dd),
	.w4(32'hbd82ee60),
	.w5(32'hbb087f10),
	.w6(32'hbcd52156),
	.w7(32'hbd64c07c),
	.w8(32'h3af8038d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60bfb5),
	.w1(32'h3b85f2c4),
	.w2(32'h3bc06c6c),
	.w3(32'hbb225b4e),
	.w4(32'h3b1845a8),
	.w5(32'h3a4a6c26),
	.w6(32'h3b32fcd5),
	.w7(32'h3b3fb797),
	.w8(32'hba3bf365),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a7e5d),
	.w1(32'hbb1253a9),
	.w2(32'hbab9acc3),
	.w3(32'hbb42ac00),
	.w4(32'h3a571151),
	.w5(32'h39a1cd1b),
	.w6(32'hba993961),
	.w7(32'h3aa089ba),
	.w8(32'hbb4eaaa9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6773c1),
	.w1(32'h3a99ee27),
	.w2(32'h3b29a185),
	.w3(32'hbaafecfd),
	.w4(32'h39c9d19c),
	.w5(32'h3b913e5e),
	.w6(32'hbb1dfa06),
	.w7(32'hbafec19d),
	.w8(32'h3a684517),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9738220),
	.w1(32'h3b80be5f),
	.w2(32'hbc9bc044),
	.w3(32'h3992c844),
	.w4(32'h3b6a5901),
	.w5(32'h3bd04372),
	.w6(32'h3ab7cf7a),
	.w7(32'h3b83ca27),
	.w8(32'hbc53fc84),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffd5f6),
	.w1(32'h398fc69e),
	.w2(32'hbb7505f2),
	.w3(32'h3d52059c),
	.w4(32'h3d28dfdb),
	.w5(32'hbb97ba88),
	.w6(32'h3d01a72c),
	.w7(32'h3cc125a2),
	.w8(32'hbc019d76),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ccad0),
	.w1(32'hbbcc870d),
	.w2(32'hbae15358),
	.w3(32'hbb72a886),
	.w4(32'hbabbea3e),
	.w5(32'hbb42d7c4),
	.w6(32'hbb53c40f),
	.w7(32'h385dfbd1),
	.w8(32'hbaf7307f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad705ef),
	.w1(32'hbbc2bce0),
	.w2(32'hb9c5ac58),
	.w3(32'hbb86bd94),
	.w4(32'h3b3ab024),
	.w5(32'h3afede99),
	.w6(32'hbbbb8dbc),
	.w7(32'h3aed97e4),
	.w8(32'h3aaa0fe1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28e801),
	.w1(32'hb920baae),
	.w2(32'hbb6330f7),
	.w3(32'h3906311a),
	.w4(32'h3ad3af4f),
	.w5(32'hbbf350b8),
	.w6(32'hbaaa03a3),
	.w7(32'h3b443d48),
	.w8(32'h3aa38c70),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c4463),
	.w1(32'hbb2aeea4),
	.w2(32'hbbc85aa3),
	.w3(32'hbae94d8e),
	.w4(32'hbb97b919),
	.w5(32'hb9fe855f),
	.w6(32'hbc14f912),
	.w7(32'hbb977567),
	.w8(32'hbbecd316),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5d247),
	.w1(32'h3b8bfb29),
	.w2(32'hbc098aa1),
	.w3(32'h3b751d41),
	.w4(32'h3ba62508),
	.w5(32'hbc32630d),
	.w6(32'hbbdf9cd9),
	.w7(32'hbb4bae89),
	.w8(32'hbb71c654),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cb4f2),
	.w1(32'hbba01498),
	.w2(32'hbbed43a5),
	.w3(32'hbc116f61),
	.w4(32'hbbae7fac),
	.w5(32'h3b0d07d7),
	.w6(32'hbbce3594),
	.w7(32'hbaa92c1c),
	.w8(32'hbb855e00),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2693a),
	.w1(32'hbbb0870b),
	.w2(32'h3b606a57),
	.w3(32'h3b84f1f8),
	.w4(32'hb9cc795c),
	.w5(32'hbb6f16f3),
	.w6(32'hbb5fa301),
	.w7(32'h3ac81d29),
	.w8(32'hbba10234),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd967aa),
	.w1(32'hbbe3cad5),
	.w2(32'h3b0bf547),
	.w3(32'h3b88a665),
	.w4(32'hbb4619fc),
	.w5(32'h3b925058),
	.w6(32'h3ab3516a),
	.w7(32'hbbcd356a),
	.w8(32'h3b85abf7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b571071),
	.w1(32'hbaad66ea),
	.w2(32'h3b4f5d59),
	.w3(32'hbb43faf8),
	.w4(32'h399eb018),
	.w5(32'h3bebdca5),
	.w6(32'hbb0314d0),
	.w7(32'h3925f7e0),
	.w8(32'hbb6a9df5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba533eb),
	.w1(32'h3bb4f79f),
	.w2(32'h3a474cd8),
	.w3(32'hbbb36121),
	.w4(32'hbb0bb9b6),
	.w5(32'h3b5da08b),
	.w6(32'hbc88024d),
	.w7(32'hbc7b32e0),
	.w8(32'h3b6b63cf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b761a),
	.w1(32'hbb709eba),
	.w2(32'h3a88c013),
	.w3(32'h3ab64a11),
	.w4(32'h3a250c53),
	.w5(32'h3b1fbd29),
	.w6(32'h3bb14b29),
	.w7(32'h3bc33e61),
	.w8(32'h3aaee782),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5085),
	.w1(32'h39fbfe58),
	.w2(32'h3b044ba8),
	.w3(32'hbc099e5c),
	.w4(32'hbb6f2650),
	.w5(32'h3bdc2874),
	.w6(32'hbb986c80),
	.w7(32'hbb853d30),
	.w8(32'hbada5d49),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed048a),
	.w1(32'hbadf7a86),
	.w2(32'hbba88495),
	.w3(32'hba2e328d),
	.w4(32'hbb7747d1),
	.w5(32'hbbb5a621),
	.w6(32'h3b8ade7e),
	.w7(32'h3b81cf6a),
	.w8(32'hbb32cf61),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedd6d4),
	.w1(32'hbb3f79fc),
	.w2(32'h3925bf28),
	.w3(32'hbba60f58),
	.w4(32'hbb79ccf0),
	.w5(32'h3ae1b796),
	.w6(32'hba41dc8f),
	.w7(32'hbba08d5a),
	.w8(32'h3bc1a048),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4ed9b),
	.w1(32'h3bd09600),
	.w2(32'hbae27129),
	.w3(32'h3bfce314),
	.w4(32'h3be16358),
	.w5(32'h3a019252),
	.w6(32'h3badaea4),
	.w7(32'h3b332d8d),
	.w8(32'hbb454397),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f5059),
	.w1(32'hbb88fea2),
	.w2(32'h3b8ba509),
	.w3(32'hbbb5d575),
	.w4(32'hbab1a5a6),
	.w5(32'h3ba30060),
	.w6(32'hb9326453),
	.w7(32'hbb2e3b5c),
	.w8(32'h3c0f541f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7ba34),
	.w1(32'hbb5e6222),
	.w2(32'h3d4ca596),
	.w3(32'h3b7f76c0),
	.w4(32'hb8c8c210),
	.w5(32'h3d1a0b86),
	.w6(32'h3bfd4daa),
	.w7(32'h3bd65bb6),
	.w8(32'h3d0a0331),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dbecb),
	.w1(32'hbd39bf94),
	.w2(32'h388a44cd),
	.w3(32'hbd9896af),
	.w4(32'hbdd5e7ef),
	.w5(32'h3ac449ce),
	.w6(32'hbd653e9d),
	.w7(32'hbd9948d8),
	.w8(32'h3af78b77),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ac5fa),
	.w1(32'hbb51d8c3),
	.w2(32'hbb688b12),
	.w3(32'h3aa5fb99),
	.w4(32'h384646eb),
	.w5(32'hbba6911c),
	.w6(32'hbb572c8d),
	.w7(32'hb9991771),
	.w8(32'hbb2b642d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb841e0f),
	.w1(32'h3a701ebc),
	.w2(32'h3bfb8454),
	.w3(32'h3ace1adf),
	.w4(32'hbb24a735),
	.w5(32'h3ba53033),
	.w6(32'h39a6bba1),
	.w7(32'h3afaca9b),
	.w8(32'h3b81b757),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1360b),
	.w1(32'h3bc26361),
	.w2(32'h3c6fb1a5),
	.w3(32'hba783640),
	.w4(32'hba749e19),
	.w5(32'h3ca49698),
	.w6(32'hba2f839b),
	.w7(32'hb80d0ce5),
	.w8(32'h3c939135),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c3a2e),
	.w1(32'h3c1730cd),
	.w2(32'h3a7b96df),
	.w3(32'h3c92470c),
	.w4(32'h3c0aa261),
	.w5(32'h3b4d7f19),
	.w6(32'h3ca153c3),
	.w7(32'h3c17c817),
	.w8(32'h3b218c0b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399450b9),
	.w1(32'h3b74bd53),
	.w2(32'hbac5b6ca),
	.w3(32'h3a83c1df),
	.w4(32'h3a198b6b),
	.w5(32'hbaf1e22e),
	.w6(32'hbb255971),
	.w7(32'hb984406a),
	.w8(32'h3b35eb20),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af6d1),
	.w1(32'h3a8e28e2),
	.w2(32'h3bd20351),
	.w3(32'hbb858fe4),
	.w4(32'hbac7d59d),
	.w5(32'hbb9c8ef3),
	.w6(32'hbb080f5c),
	.w7(32'hbb51d732),
	.w8(32'hb980c1b5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30db50),
	.w1(32'h3b8a060c),
	.w2(32'hbc16f213),
	.w3(32'hbbbdb9fb),
	.w4(32'hbaa7dd21),
	.w5(32'h3bbd8a0f),
	.w6(32'hba8945f7),
	.w7(32'hb93bae8f),
	.w8(32'hbc12f0d2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4adf2d),
	.w1(32'hbc9f0348),
	.w2(32'hbbb4e61e),
	.w3(32'h3c637461),
	.w4(32'hbbdb4a32),
	.w5(32'hbbcc254d),
	.w6(32'hb900fc86),
	.w7(32'hbc82ee59),
	.w8(32'hbba9ab90),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dcf7b),
	.w1(32'h3ad123cd),
	.w2(32'h3ad80cc0),
	.w3(32'h3a7cc15e),
	.w4(32'h3bbcf0b3),
	.w5(32'hbbaf1ed3),
	.w6(32'hbae6d917),
	.w7(32'h3b89b95d),
	.w8(32'hbba5beb6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8cde6),
	.w1(32'hbabd8fb1),
	.w2(32'h3a6e0f6b),
	.w3(32'hbb996d73),
	.w4(32'hbb62df5f),
	.w5(32'h3951a6bc),
	.w6(32'hbbe77757),
	.w7(32'hbb80e724),
	.w8(32'h3a8abf50),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b6420),
	.w1(32'h3b90bd56),
	.w2(32'hbb5177f1),
	.w3(32'hba1f0269),
	.w4(32'h3b4d8c36),
	.w5(32'hbb1870e9),
	.w6(32'h3b4648e3),
	.w7(32'hbb3757a0),
	.w8(32'h3b1f30c9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17c2f5),
	.w1(32'hba07d78d),
	.w2(32'h3c7a84b6),
	.w3(32'hbb9f998c),
	.w4(32'hb920caf7),
	.w5(32'h3c3eaa15),
	.w6(32'hbae90fcd),
	.w7(32'hbb1de696),
	.w8(32'h3c0c8a38),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb156da3),
	.w1(32'hbc0db09f),
	.w2(32'h3bc3a8c7),
	.w3(32'hbcfb71fe),
	.w4(32'hbcd64ac1),
	.w5(32'h3babfd10),
	.w6(32'hbca08d12),
	.w7(32'hbc9e3173),
	.w8(32'h3ba537c3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6f36c),
	.w1(32'h3984544e),
	.w2(32'h3d59fe4c),
	.w3(32'h3bf09bf3),
	.w4(32'hbb6309d3),
	.w5(32'h3d177161),
	.w6(32'h3b797961),
	.w7(32'h3b0cc0e5),
	.w8(32'h3d142222),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca96cd4),
	.w1(32'hbd2fcc6e),
	.w2(32'h3b93bab1),
	.w3(32'hbdc489b9),
	.w4(32'hbdef112a),
	.w5(32'h38dfac40),
	.w6(32'hbda1035b),
	.w7(32'hbdb9fc4a),
	.w8(32'h3b67c3a6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2232c),
	.w1(32'h39cf1d34),
	.w2(32'hbafb929a),
	.w3(32'h3a230550),
	.w4(32'h3b0c6482),
	.w5(32'hbb09f10a),
	.w6(32'h3a136368),
	.w7(32'h3ad8dd76),
	.w8(32'h3b179f57),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdedb2d),
	.w1(32'h398418dc),
	.w2(32'hbb439717),
	.w3(32'hbc214e1d),
	.w4(32'hbb871ef8),
	.w5(32'hbab61056),
	.w6(32'hbc075a7e),
	.w7(32'hbaea17bf),
	.w8(32'h3b35aa10),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861f782),
	.w1(32'hba84387c),
	.w2(32'hbb248b28),
	.w3(32'hbb5621d9),
	.w4(32'hba29495b),
	.w5(32'hbba586f3),
	.w6(32'hbb24e7d6),
	.w7(32'hbbad0c6a),
	.w8(32'hbad5070f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c039f7d),
	.w1(32'h3b44b0f6),
	.w2(32'h3c2c2c3c),
	.w3(32'h3c03ba4c),
	.w4(32'hb8fb4e36),
	.w5(32'h3c083c88),
	.w6(32'h3b83c4c1),
	.w7(32'h3be687aa),
	.w8(32'h3c1b75c2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c0ca5),
	.w1(32'h3bb2a2c9),
	.w2(32'h3c825947),
	.w3(32'h3ab6057c),
	.w4(32'h3bcd5c23),
	.w5(32'h3c5597db),
	.w6(32'h3abb00a6),
	.w7(32'h3be3955f),
	.w8(32'h3c1ec27a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06bcbc),
	.w1(32'hbc3a674d),
	.w2(32'hba496234),
	.w3(32'hbc639b14),
	.w4(32'hbcdda9ea),
	.w5(32'hba5942e8),
	.w6(32'hbc44f786),
	.w7(32'hbca3f87c),
	.w8(32'hbae4b16f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9573ac7),
	.w1(32'hbab4cb00),
	.w2(32'hbba706e6),
	.w3(32'hbad16331),
	.w4(32'hbb4400f2),
	.w5(32'hbbda6572),
	.w6(32'hbb0ae09e),
	.w7(32'hbb2dfe56),
	.w8(32'hba2b94cb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24d939),
	.w1(32'h3ac186a9),
	.w2(32'hbadc0e95),
	.w3(32'hbb36791e),
	.w4(32'hbb15fdf3),
	.w5(32'h3b04b6af),
	.w6(32'h3a9314b1),
	.w7(32'hbb1e38ec),
	.w8(32'h3be3161d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9717f7),
	.w1(32'hbc0ebee6),
	.w2(32'hbc3b32fb),
	.w3(32'h3ad8ac23),
	.w4(32'hbb38aee3),
	.w5(32'hba49c7d5),
	.w6(32'h3be404b3),
	.w7(32'h3c01ef81),
	.w8(32'hbb8bd289),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66355f),
	.w1(32'hbbb7743b),
	.w2(32'h3b29e1c7),
	.w3(32'h3b95db53),
	.w4(32'hba7dbdf3),
	.w5(32'h388af48c),
	.w6(32'h39055836),
	.w7(32'hbc01c78f),
	.w8(32'hba76f191),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b6614),
	.w1(32'h3baf2220),
	.w2(32'h3d40b3f4),
	.w3(32'h3a0b9ffe),
	.w4(32'h3b8c45a7),
	.w5(32'h3d3d6814),
	.w6(32'h3b5e9360),
	.w7(32'h3bd4b401),
	.w8(32'h3d087ba1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74827b),
	.w1(32'hbcda8a88),
	.w2(32'hbb8fa69e),
	.w3(32'hbd211f7b),
	.w4(32'hbd8e5082),
	.w5(32'hba4d208a),
	.w6(32'hbd0df51d),
	.w7(32'hbd68ff13),
	.w8(32'hbb20a984),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b602668),
	.w1(32'hbb42a26a),
	.w2(32'hbae28ee5),
	.w3(32'h3b7f763d),
	.w4(32'hbb467ee5),
	.w5(32'hbb88fc2b),
	.w6(32'hbb56eba8),
	.w7(32'h3a48c59a),
	.w8(32'hbbee88bb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a82da),
	.w1(32'hbc0353ed),
	.w2(32'hbbf31f64),
	.w3(32'hbbab6bea),
	.w4(32'h3b303a6e),
	.w5(32'hbbcee9ee),
	.w6(32'hbb833618),
	.w7(32'hba61afc1),
	.w8(32'hbc2e6562),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d02a),
	.w1(32'hbb0c6b55),
	.w2(32'h3a9f5ff1),
	.w3(32'hba2f3d1f),
	.w4(32'h3b552a88),
	.w5(32'hb92c7530),
	.w6(32'hbc0caf9e),
	.w7(32'h3aa77f3c),
	.w8(32'hbb4cdc2d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10914f),
	.w1(32'hba968633),
	.w2(32'hba880cd9),
	.w3(32'hbaf495d2),
	.w4(32'hbb0608a5),
	.w5(32'h3b9b5fa2),
	.w6(32'hbc19e528),
	.w7(32'hbb6342b8),
	.w8(32'h3b35bc69),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba757d3b),
	.w1(32'hb78b5081),
	.w2(32'h3bf2ada3),
	.w3(32'hbb14c39e),
	.w4(32'h3aedd398),
	.w5(32'h3be4e7e9),
	.w6(32'hbaebf74b),
	.w7(32'hba9b5454),
	.w8(32'h39ce6cf5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24b2c4),
	.w1(32'h3b9910b0),
	.w2(32'hba6ac993),
	.w3(32'hbbfaa8f4),
	.w4(32'hbb60a0e8),
	.w5(32'hbae05ff6),
	.w6(32'hbc412d43),
	.w7(32'hbb0caa7e),
	.w8(32'h3b6ae9f1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65afd6),
	.w1(32'hbb1e1d96),
	.w2(32'hbb472447),
	.w3(32'hbb2da2a4),
	.w4(32'h3a69ee8f),
	.w5(32'hba29ca25),
	.w6(32'hbaf82251),
	.w7(32'hbac8a248),
	.w8(32'hbbd31cd6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90504f),
	.w1(32'hbb47cbfe),
	.w2(32'hbb4a8332),
	.w3(32'h3b502a25),
	.w4(32'h3b710f57),
	.w5(32'hbb808297),
	.w6(32'hbace6c7c),
	.w7(32'hbb67ffe7),
	.w8(32'hba2139cc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205148),
	.w1(32'hba63be5b),
	.w2(32'h3a544552),
	.w3(32'h3ad03544),
	.w4(32'h3a310725),
	.w5(32'h3b471818),
	.w6(32'hbb746198),
	.w7(32'h3a7ec218),
	.w8(32'h3c0682c2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33e4bc),
	.w1(32'h3a02aa77),
	.w2(32'h399202cc),
	.w3(32'h39442135),
	.w4(32'h3b4d40a4),
	.w5(32'h383ea5c7),
	.w6(32'hbb46c3fc),
	.w7(32'h3a89860b),
	.w8(32'h3b07caa5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb721139a),
	.w1(32'h3b3fab26),
	.w2(32'hba765e98),
	.w3(32'hbb31a881),
	.w4(32'h3ac0d56a),
	.w5(32'h3b191586),
	.w6(32'h3b960287),
	.w7(32'h3b4d95d0),
	.w8(32'h3b12b5af),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b052ba6),
	.w1(32'h3bb5f2b4),
	.w2(32'h3b840e3a),
	.w3(32'h3b9470a6),
	.w4(32'h3b3eca91),
	.w5(32'h3b9e9033),
	.w6(32'h3b0c3c53),
	.w7(32'h3b0eac06),
	.w8(32'h3beb98db),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c111161),
	.w1(32'h3b825022),
	.w2(32'hbadd5557),
	.w3(32'h3c479214),
	.w4(32'h3b8c0118),
	.w5(32'hbb5be11a),
	.w6(32'h3c0a2195),
	.w7(32'h3c046128),
	.w8(32'hbba9ccfd),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb20587),
	.w1(32'hba43b015),
	.w2(32'hb941a8c3),
	.w3(32'hba4ccb1f),
	.w4(32'hbb22f65c),
	.w5(32'hbb0ec9cc),
	.w6(32'hbb4661ad),
	.w7(32'hbae0b087),
	.w8(32'h398cd36e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4156e0),
	.w1(32'h3b4aecda),
	.w2(32'hbb8828e7),
	.w3(32'h3a55b365),
	.w4(32'h3b03a007),
	.w5(32'hbb3ff168),
	.w6(32'h3a2922f0),
	.w7(32'h39f3bc70),
	.w8(32'hbb8dac09),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba670267),
	.w1(32'hbb54e52d),
	.w2(32'h3a23066e),
	.w3(32'h3b1eab12),
	.w4(32'h3aaada2b),
	.w5(32'h39521c83),
	.w6(32'hbb6bbb13),
	.w7(32'hbb3b7ae7),
	.w8(32'h3b37e978),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade6fcb),
	.w1(32'hbb727445),
	.w2(32'h3b301985),
	.w3(32'h3a58d83e),
	.w4(32'hbbaf1dd1),
	.w5(32'hb982802e),
	.w6(32'hbbe5b531),
	.w7(32'hbaa7c684),
	.w8(32'h3a2a9189),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6af1f),
	.w1(32'h3b9d825d),
	.w2(32'hbb39511a),
	.w3(32'h3b5d3599),
	.w4(32'hb9d42fca),
	.w5(32'hbb83ee6e),
	.w6(32'hba3b2600),
	.w7(32'h3aa8a360),
	.w8(32'hbb5cc008),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba52850),
	.w1(32'hbbec1b30),
	.w2(32'hb95e98d9),
	.w3(32'hbb4ef419),
	.w4(32'hbbd5457a),
	.w5(32'hbb50bfe3),
	.w6(32'hbbb06f81),
	.w7(32'hbb26c184),
	.w8(32'h3ba4a96e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99aa455),
	.w1(32'h3bc2e6fc),
	.w2(32'hbaaf54ac),
	.w3(32'hba1c25fe),
	.w4(32'h3923bcb5),
	.w5(32'hbba063e1),
	.w6(32'h3aeca05f),
	.w7(32'h3ad1b888),
	.w8(32'hbbabc70d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917716),
	.w1(32'hbbd04f3e),
	.w2(32'h3b875594),
	.w3(32'h37fdc87b),
	.w4(32'hbaf46abc),
	.w5(32'h3a06b1a5),
	.w6(32'hbaf46788),
	.w7(32'hbba66bdb),
	.w8(32'hbb4e0589),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34e5c),
	.w1(32'h3c06d30d),
	.w2(32'hba97c93d),
	.w3(32'h3ae7e01b),
	.w4(32'h3b6feb8a),
	.w5(32'h3b754bca),
	.w6(32'hbb65fd72),
	.w7(32'hbaacbf8d),
	.w8(32'h3bc672b8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c008315),
	.w1(32'h3be79deb),
	.w2(32'h3a771c1e),
	.w3(32'h3b8a7492),
	.w4(32'h3bf2eb50),
	.w5(32'hb9ecaced),
	.w6(32'h3b55fff5),
	.w7(32'h3b0d713d),
	.w8(32'hba8eeb8f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a0cb8),
	.w1(32'hb8782581),
	.w2(32'hbb6d8a9e),
	.w3(32'h3a834972),
	.w4(32'h3adb7835),
	.w5(32'hbb3e4237),
	.w6(32'hba5f7d03),
	.w7(32'hbae36555),
	.w8(32'hbb20b25b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0e69d),
	.w1(32'hba49064c),
	.w2(32'h3af91947),
	.w3(32'hbb3e624a),
	.w4(32'h3b534bd2),
	.w5(32'hb94ac203),
	.w6(32'hbb1a300e),
	.w7(32'hbb4aee68),
	.w8(32'hbae24738),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fc5bb),
	.w1(32'hba051216),
	.w2(32'hba9c54b5),
	.w3(32'h3a8526c3),
	.w4(32'h3a63af62),
	.w5(32'hbb4ec317),
	.w6(32'hbaab5385),
	.w7(32'hbb93f009),
	.w8(32'hbbd2dfd0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b2ca2),
	.w1(32'hba08d168),
	.w2(32'hbc877b2a),
	.w3(32'hba24764c),
	.w4(32'h396b309f),
	.w5(32'hbc91ec9d),
	.w6(32'hbbb28b26),
	.w7(32'hba89f8bc),
	.w8(32'hbc6d0826),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76c734),
	.w1(32'h3be64f50),
	.w2(32'hbbd5da53),
	.w3(32'h3c0a0634),
	.w4(32'h3cb74fb2),
	.w5(32'hbc469a1e),
	.w6(32'h3c21bd86),
	.w7(32'h3c959041),
	.w8(32'hbbe648a9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b7d9d),
	.w1(32'h3baff3bc),
	.w2(32'hb9bcb511),
	.w3(32'hbc165a50),
	.w4(32'h3b16cfc8),
	.w5(32'hbb0f389b),
	.w6(32'hbb90ed1a),
	.w7(32'h3b8fb415),
	.w8(32'h3adc1983),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb965a7),
	.w1(32'hbb4de3c8),
	.w2(32'h3c1773eb),
	.w3(32'hbbe2d937),
	.w4(32'hbac66a13),
	.w5(32'h3c20ec4e),
	.w6(32'hbb88bfb5),
	.w7(32'h398a7b7e),
	.w8(32'h3b8f8d3e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ff174),
	.w1(32'h3a735396),
	.w2(32'h3b08b4dc),
	.w3(32'h3c0ddd7d),
	.w4(32'h3b6839ec),
	.w5(32'h3a1945ab),
	.w6(32'h3b4a32a6),
	.w7(32'hbacca9f3),
	.w8(32'h3a9e997d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b5aab),
	.w1(32'hbb17f5b5),
	.w2(32'hbb3560ce),
	.w3(32'hbbc668df),
	.w4(32'hba24de27),
	.w5(32'hb6a5fb53),
	.w6(32'h37fa6429),
	.w7(32'h3b635757),
	.w8(32'h3b8d6d5f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3eac96),
	.w1(32'h3ab3fa05),
	.w2(32'hbb388811),
	.w3(32'h3a8be11f),
	.w4(32'hbc20d183),
	.w5(32'hbabd1dfc),
	.w6(32'h3a2407ae),
	.w7(32'hbbbd4126),
	.w8(32'hbb4d2e23),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39199e05),
	.w1(32'h39c7ef26),
	.w2(32'h3c0446dc),
	.w3(32'h3b4d43b3),
	.w4(32'h3ac5e265),
	.w5(32'h3c0d439e),
	.w6(32'h3b1f7834),
	.w7(32'h3b098d6f),
	.w8(32'hbbdfc816),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37fd4c),
	.w1(32'hbac4d02d),
	.w2(32'hbb1cc98a),
	.w3(32'h3bffcc96),
	.w4(32'h3b93c0e2),
	.w5(32'hb7042b0f),
	.w6(32'h3bc97a51),
	.w7(32'h3bc3bfdc),
	.w8(32'hbbc39864),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f44ab),
	.w1(32'hbac0a3a0),
	.w2(32'hba1391bc),
	.w3(32'h3bbcc1a1),
	.w4(32'h3b265077),
	.w5(32'h3b41b21c),
	.w6(32'hba2cb044),
	.w7(32'h3a712f8e),
	.w8(32'h3abc3ec8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c56d8),
	.w1(32'hba6d4007),
	.w2(32'h3a61a58e),
	.w3(32'hbab3d9e7),
	.w4(32'hbb04d756),
	.w5(32'hbb4486ad),
	.w6(32'h3baefa13),
	.w7(32'hba9a4a95),
	.w8(32'hbb40a837),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77b9c3),
	.w1(32'h39c1c8fe),
	.w2(32'hbbf9c047),
	.w3(32'hbad18a15),
	.w4(32'h3a9955b3),
	.w5(32'hbb636fbe),
	.w6(32'hbb818f1d),
	.w7(32'hb98f29fc),
	.w8(32'hbc02ec71),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bf7a3),
	.w1(32'h3b3ff52f),
	.w2(32'hb9f58cc1),
	.w3(32'hb97cd85f),
	.w4(32'h3b68c29f),
	.w5(32'h3a7ab8fe),
	.w6(32'hbb5db68d),
	.w7(32'hbbe5fc57),
	.w8(32'hbc0e1553),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5226),
	.w1(32'h3ac17f64),
	.w2(32'h3d2409d1),
	.w3(32'hb9d65a42),
	.w4(32'hba2ed48f),
	.w5(32'h3d591deb),
	.w6(32'hba2a4b5d),
	.w7(32'h3ae31917),
	.w8(32'h3cf0bb54),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63b71f),
	.w1(32'hbd0ece3e),
	.w2(32'hbb81c5b2),
	.w3(32'hbbe1c4b7),
	.w4(32'hbd8b5800),
	.w5(32'hbb8b1220),
	.w6(32'hbcb8cd6a),
	.w7(32'hbd880eb3),
	.w8(32'hbc17939d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5483f6),
	.w1(32'h3a1ec2c5),
	.w2(32'hbba08968),
	.w3(32'hb9a1064e),
	.w4(32'h3af4df99),
	.w5(32'hbbe7598b),
	.w6(32'hbbbb272d),
	.w7(32'hbb387c71),
	.w8(32'h3651f8e9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba902e46),
	.w1(32'hba7430a4),
	.w2(32'hbb266afc),
	.w3(32'h3b0ca53e),
	.w4(32'hba262bf5),
	.w5(32'h3a5fa3c3),
	.w6(32'h3b306043),
	.w7(32'h3b772e59),
	.w8(32'hbb9e2247),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44d0d0),
	.w1(32'hbb7a3d11),
	.w2(32'h3c886c35),
	.w3(32'h3a58e3d2),
	.w4(32'h3b23e5c5),
	.w5(32'h3b9e6024),
	.w6(32'hbafda433),
	.w7(32'hbb80d7dd),
	.w8(32'h3c54d3d9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc20d0),
	.w1(32'hbc206d42),
	.w2(32'hba849e5e),
	.w3(32'hbd20ff98),
	.w4(32'hbd27137f),
	.w5(32'hba7a0a7b),
	.w6(32'hbccc6c3a),
	.w7(32'hbce5860c),
	.w8(32'hbb4f63d7),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78d0cb),
	.w1(32'hbb84755d),
	.w2(32'h3ba6651c),
	.w3(32'hbae8a5e5),
	.w4(32'h3b57c5ef),
	.w5(32'h3c461292),
	.w6(32'hbbb601c9),
	.w7(32'hbb957766),
	.w8(32'h3be457fe),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b921c),
	.w1(32'h3c8fee13),
	.w2(32'h39d8445e),
	.w3(32'h3d01bb17),
	.w4(32'h3d167919),
	.w5(32'hbad4445b),
	.w6(32'h3cd37b87),
	.w7(32'h3cf53cd1),
	.w8(32'h3a84c913),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eb031),
	.w1(32'hbb25e90b),
	.w2(32'h3b29594c),
	.w3(32'hbaac86b7),
	.w4(32'hbbe81074),
	.w5(32'hb9c9f822),
	.w6(32'hbc2d3eb7),
	.w7(32'hbbfa2974),
	.w8(32'h3a335380),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396fc098),
	.w1(32'h3b530c4b),
	.w2(32'h3b8cba83),
	.w3(32'hb8b5710a),
	.w4(32'h3c11c4fe),
	.w5(32'h3a63362e),
	.w6(32'h3c02a71e),
	.w7(32'h3b590cf6),
	.w8(32'h3b5b4a52),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49ab8f),
	.w1(32'h3a47f0be),
	.w2(32'h3ccdf245),
	.w3(32'h3b4f7de7),
	.w4(32'h39ca1b32),
	.w5(32'h3c5d0d0f),
	.w6(32'h3b2b3048),
	.w7(32'h3b068bfa),
	.w8(32'h3c82ee6e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c30d3),
	.w1(32'hbce2ceb1),
	.w2(32'hbb55c8a9),
	.w3(32'hbd66a17e),
	.w4(32'hbd8f0b63),
	.w5(32'h3a52c083),
	.w6(32'hbd321c1c),
	.w7(32'hbd5e3d07),
	.w8(32'hbaea1e95),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96ca2b),
	.w1(32'h3b7106ac),
	.w2(32'hbb070558),
	.w3(32'hb9767b06),
	.w4(32'h3ae82b8b),
	.w5(32'hbb66523b),
	.w6(32'hbb76aad6),
	.w7(32'hbb92d1f2),
	.w8(32'hbbfe1591),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3486aa),
	.w1(32'h39c3ef78),
	.w2(32'hbaaa9d6b),
	.w3(32'hbb70046e),
	.w4(32'h3aefe6cd),
	.w5(32'h3b3ce0aa),
	.w6(32'h3991fa2b),
	.w7(32'hbaaf2cec),
	.w8(32'h39be0714),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5db816),
	.w1(32'h39bb663b),
	.w2(32'h3b983935),
	.w3(32'hbb1d7fa7),
	.w4(32'h3b64623c),
	.w5(32'h3b7bf6a4),
	.w6(32'h3b86438a),
	.w7(32'h3b53772b),
	.w8(32'h3ba48e32),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70425e),
	.w1(32'h37554893),
	.w2(32'hbac2a0b9),
	.w3(32'h3aa69e0b),
	.w4(32'h3a432462),
	.w5(32'hbb9d8c6f),
	.w6(32'hba65f665),
	.w7(32'hbb3cdfa9),
	.w8(32'hbb2521e6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dfeda),
	.w1(32'hbb2b1196),
	.w2(32'h39ff7483),
	.w3(32'hbb6d5214),
	.w4(32'hbc0353ed),
	.w5(32'h3a73f0c1),
	.w6(32'hbab8a1e6),
	.w7(32'hbb3fb4b0),
	.w8(32'h3b0022b2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f2bc),
	.w1(32'h3b91081b),
	.w2(32'hbc44aeee),
	.w3(32'h3b7ff86c),
	.w4(32'h3beda776),
	.w5(32'hbc985053),
	.w6(32'h3bb8a9ca),
	.w7(32'h3b4cff6f),
	.w8(32'hbc38d70a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41b0c4),
	.w1(32'h3c9fcadf),
	.w2(32'h3ab6ee41),
	.w3(32'h3c0f6c1d),
	.w4(32'h3cd7ad67),
	.w5(32'h3996b587),
	.w6(32'h3c1304db),
	.w7(32'h3cc4213d),
	.w8(32'hbb021abf),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1472c),
	.w1(32'hba2ca11e),
	.w2(32'hbbbaf6b8),
	.w3(32'hbbae78f5),
	.w4(32'h3a09fd7f),
	.w5(32'h3a9ab377),
	.w6(32'h3a7e7a54),
	.w7(32'hbbacb138),
	.w8(32'hbabe46e4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeddb77),
	.w1(32'hbb88ca4a),
	.w2(32'hbb387027),
	.w3(32'hbb510ec5),
	.w4(32'h3a87d191),
	.w5(32'hbb36f87f),
	.w6(32'hba16e457),
	.w7(32'hbb0d8514),
	.w8(32'hbaf16870),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafedb04),
	.w1(32'hba0b00e5),
	.w2(32'hb9094e8f),
	.w3(32'hbb6563f5),
	.w4(32'h3a956b91),
	.w5(32'h3823132e),
	.w6(32'hbbfe4ab3),
	.w7(32'hbb882609),
	.w8(32'h3a11253f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa25a12),
	.w1(32'hba8e56ea),
	.w2(32'hbb81f9f4),
	.w3(32'h3b8064d4),
	.w4(32'hbb02fcbe),
	.w5(32'hbc4ee961),
	.w6(32'h3b001a99),
	.w7(32'hba388c05),
	.w8(32'hbbc209ab),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc293179),
	.w1(32'h3b46b7c9),
	.w2(32'h3bae3b06),
	.w3(32'hbc9fe0f6),
	.w4(32'h3b13d6cf),
	.w5(32'hba413e41),
	.w6(32'hbc62b482),
	.w7(32'h3bd594c2),
	.w8(32'hbb7caf2d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ce421),
	.w1(32'h3c33d902),
	.w2(32'h3b4631fc),
	.w3(32'h3b6530f0),
	.w4(32'hbad7290d),
	.w5(32'h3b93b361),
	.w6(32'h3bcf1efa),
	.w7(32'h3b2563f5),
	.w8(32'h3bdcb8b0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5dfc3),
	.w1(32'hbb398c95),
	.w2(32'hbb3ccd3e),
	.w3(32'h3aee7fb9),
	.w4(32'hbb48ca2d),
	.w5(32'h3ba93c32),
	.w6(32'h3ba1bdac),
	.w7(32'hba159da0),
	.w8(32'hba30bacf),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addbb32),
	.w1(32'h3a3fb21b),
	.w2(32'h3bc119bb),
	.w3(32'h3c139a30),
	.w4(32'h3a42d620),
	.w5(32'h3c467987),
	.w6(32'h3b03e10f),
	.w7(32'h3a22f9d3),
	.w8(32'h3c7e7b2d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3e097),
	.w1(32'hbb207d16),
	.w2(32'h3b3a3533),
	.w3(32'h3bc81a0d),
	.w4(32'hbc18b49a),
	.w5(32'hbadc2619),
	.w6(32'h3c22e89b),
	.w7(32'hbbd1e170),
	.w8(32'h3b81d82a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a1ef9),
	.w1(32'hbb65dc21),
	.w2(32'h3c35de97),
	.w3(32'hbb6e6d3c),
	.w4(32'hbbc1c2b2),
	.w5(32'h3c847ff6),
	.w6(32'hbadc2231),
	.w7(32'hbaa34867),
	.w8(32'h3b66dfe2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f543b),
	.w1(32'h3b88b3d3),
	.w2(32'h3a983bf9),
	.w3(32'h3baf30a8),
	.w4(32'hbb8edd5d),
	.w5(32'h3a003cfe),
	.w6(32'hbbed39d5),
	.w7(32'hbb2d6eec),
	.w8(32'hb9f2ed0f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945311a),
	.w1(32'hb955aadf),
	.w2(32'h3c66addc),
	.w3(32'h3a821093),
	.w4(32'hbafa1a4f),
	.w5(32'h3bfe83bf),
	.w6(32'hba3e209b),
	.w7(32'hbb35537f),
	.w8(32'h3b0598aa),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c329e),
	.w1(32'h3c408096),
	.w2(32'hbb7a8c75),
	.w3(32'h3bb42e18),
	.w4(32'h3bcd32b1),
	.w5(32'hbc0cdabe),
	.w6(32'h3bfd58b1),
	.w7(32'hbb5680c0),
	.w8(32'hbb30c51a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13d797),
	.w1(32'hbbaf5492),
	.w2(32'h3ba83ada),
	.w3(32'hbb8cf56e),
	.w4(32'hbbf7bcc2),
	.w5(32'h3c2c916a),
	.w6(32'hb983124b),
	.w7(32'hbab06b83),
	.w8(32'h3c03a425),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a6190),
	.w1(32'h3ae9005b),
	.w2(32'hbac886c2),
	.w3(32'h3c49a7a4),
	.w4(32'hbc2eb4f3),
	.w5(32'h3a425814),
	.w6(32'h3b1a2917),
	.w7(32'hbc3c09fc),
	.w8(32'hbab4d29d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb588c65),
	.w1(32'hbbc27142),
	.w2(32'hb9c6b337),
	.w3(32'hbae6936b),
	.w4(32'hbb93eb96),
	.w5(32'h3b449db5),
	.w6(32'h3b81ab6e),
	.w7(32'hbbbc3a6c),
	.w8(32'hb89614d5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f54045),
	.w1(32'hbbb6949c),
	.w2(32'h3c25805b),
	.w3(32'h3b2f6666),
	.w4(32'hbbe124f4),
	.w5(32'h3c969060),
	.w6(32'h3934b056),
	.w7(32'hbc48a7f5),
	.w8(32'h3c34a6ff),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe6090),
	.w1(32'hbbc86fb9),
	.w2(32'h3a29cf07),
	.w3(32'h3c2e987d),
	.w4(32'hbc6771c3),
	.w5(32'h3b88d52c),
	.w6(32'h3c3b6321),
	.w7(32'hbc09d720),
	.w8(32'h3b4e2de0),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90b4b8),
	.w1(32'h3b26ff85),
	.w2(32'hbbd6a7fb),
	.w3(32'h3c5e682e),
	.w4(32'h3b322bc5),
	.w5(32'hbbf6268d),
	.w6(32'h3be7a047),
	.w7(32'hbacbda24),
	.w8(32'hbc07dd5a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38faf7b8),
	.w1(32'h3acf3967),
	.w2(32'h3b4a525d),
	.w3(32'hba2051f5),
	.w4(32'hba5240d2),
	.w5(32'h3b0cf6e4),
	.w6(32'hbb314d5d),
	.w7(32'hbb0a4a69),
	.w8(32'h3b0cbc6d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdb25a),
	.w1(32'hbc02dbcc),
	.w2(32'h3b50b751),
	.w3(32'h3a6d2db2),
	.w4(32'hbc6a9866),
	.w5(32'hb93930ad),
	.w6(32'h3a4a364a),
	.w7(32'hbc06ea62),
	.w8(32'h3be7fbe4),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f6438),
	.w1(32'hba49e472),
	.w2(32'hbb475997),
	.w3(32'hbb172beb),
	.w4(32'hbba3fa58),
	.w5(32'hbb1c2f18),
	.w6(32'hbbae7e5b),
	.w7(32'hbb65c7ff),
	.w8(32'hbba4d645),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b981ba5),
	.w1(32'hbb240af0),
	.w2(32'h3b3c2814),
	.w3(32'h3ad89018),
	.w4(32'h3a54e2d5),
	.w5(32'h3babe49c),
	.w6(32'h3b224f3f),
	.w7(32'h3b8db0b7),
	.w8(32'hbb89c1a0),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb86d49),
	.w1(32'hbc4345b8),
	.w2(32'hbb54fae9),
	.w3(32'h399e803c),
	.w4(32'hbbc3b4f3),
	.w5(32'hbacfe6a1),
	.w6(32'h3a1d7300),
	.w7(32'hbbf5c096),
	.w8(32'hbbc8ea99),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba906731),
	.w1(32'hbaf8cf10),
	.w2(32'h3b486ca6),
	.w3(32'hba795cf6),
	.w4(32'hbaa532e1),
	.w5(32'h3b999cd3),
	.w6(32'hbb9854f8),
	.w7(32'hbb87ac7c),
	.w8(32'h3ba48ad9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d6ea9),
	.w1(32'h3bc78021),
	.w2(32'h3a8f4bf8),
	.w3(32'h3c2aa311),
	.w4(32'h3c4dfa59),
	.w5(32'h3bb2ad74),
	.w6(32'h3b82f852),
	.w7(32'h3bfd528b),
	.w8(32'hbb2eae5b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2579e9),
	.w1(32'h3bbc62d6),
	.w2(32'h3bca4fb6),
	.w3(32'h3c35bd21),
	.w4(32'h3b363edf),
	.w5(32'h3c54e7d0),
	.w6(32'h3b5acb12),
	.w7(32'hbb2ab400),
	.w8(32'h3c6acf9c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc422f6),
	.w1(32'h3aa5239e),
	.w2(32'hbb2b4595),
	.w3(32'h3c082d9d),
	.w4(32'hbbb17062),
	.w5(32'hbb978af1),
	.w6(32'h3bb603c7),
	.w7(32'hbc5cbe4c),
	.w8(32'hbbb7c3a6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba83596),
	.w1(32'hb9933f98),
	.w2(32'h3ba3e5a3),
	.w3(32'h3c11e0f8),
	.w4(32'h3bd1ea6c),
	.w5(32'h3c3fd572),
	.w6(32'h3b103018),
	.w7(32'hbaea25fd),
	.w8(32'h3bd15ec3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d4e61),
	.w1(32'hba73330a),
	.w2(32'h3adf2bab),
	.w3(32'h3aced2b9),
	.w4(32'hbb5854db),
	.w5(32'hbb2628b4),
	.w6(32'h3b95c20d),
	.w7(32'hba197d22),
	.w8(32'hba4dd7bd),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01d558),
	.w1(32'h3c19222f),
	.w2(32'h3c26a957),
	.w3(32'hbb3d11b5),
	.w4(32'h3b96577e),
	.w5(32'h3c811bb4),
	.w6(32'h38e1fc06),
	.w7(32'hbb6ef250),
	.w8(32'h3c023e6a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b4746),
	.w1(32'hbbf94e39),
	.w2(32'h3b6f9a55),
	.w3(32'h3bb722b9),
	.w4(32'hbb96a939),
	.w5(32'h3be41d18),
	.w6(32'h3c2f1375),
	.w7(32'hbb80255b),
	.w8(32'h39c517bd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba336cdb),
	.w1(32'hbba20c39),
	.w2(32'hbb5529f1),
	.w3(32'hbb4b24d5),
	.w4(32'hbbcce508),
	.w5(32'hb962d855),
	.w6(32'h3c00e3e4),
	.w7(32'hbc1ac069),
	.w8(32'h3b3ccfb9),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c288b),
	.w1(32'h3a518d95),
	.w2(32'h3b2fee61),
	.w3(32'h3cbb3547),
	.w4(32'h3bab3d2d),
	.w5(32'h39b7fd51),
	.w6(32'h3caa41fe),
	.w7(32'h3b0b85df),
	.w8(32'h3ac39f00),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87de4),
	.w1(32'hbc4c9e14),
	.w2(32'hbb9d2929),
	.w3(32'h3befce2d),
	.w4(32'hbc6fe8e7),
	.w5(32'hbb608040),
	.w6(32'h3b8e0767),
	.w7(32'hbc9eb273),
	.w8(32'h38a37264),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67feb4),
	.w1(32'hbb567348),
	.w2(32'hbc3b72e4),
	.w3(32'h3a987303),
	.w4(32'hbad0ec3f),
	.w5(32'hbc825650),
	.w6(32'hbaddc7a5),
	.w7(32'hbbbecd0e),
	.w8(32'hbc13eff5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca55a),
	.w1(32'h3b96360b),
	.w2(32'h3c05e09f),
	.w3(32'hbba5762c),
	.w4(32'h3bf4f60c),
	.w5(32'h3c44f052),
	.w6(32'hbb6f76e2),
	.w7(32'h3c3317d3),
	.w8(32'h3c1a2034),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82e307),
	.w1(32'hbb211b26),
	.w2(32'h3bb65d8a),
	.w3(32'h3aad2e1d),
	.w4(32'hbbcfe930),
	.w5(32'hba5d77ee),
	.w6(32'h3c16cf04),
	.w7(32'hbb03b339),
	.w8(32'h3bbf98b7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8e544),
	.w1(32'h3b86e797),
	.w2(32'hbbb1366c),
	.w3(32'h3b8a2a01),
	.w4(32'h39b540ac),
	.w5(32'hbbaf211a),
	.w6(32'h3b517ecf),
	.w7(32'h3bdeece2),
	.w8(32'hba7f047d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d91c3),
	.w1(32'hba2895e6),
	.w2(32'hbaef38a8),
	.w3(32'h3b885ff9),
	.w4(32'hbaded687),
	.w5(32'hbc2be448),
	.w6(32'h3b3af9a6),
	.w7(32'hbb2286dd),
	.w8(32'hbc3faa65),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abced93),
	.w1(32'hb96be6e8),
	.w2(32'hbae9f2ed),
	.w3(32'hba62c6e7),
	.w4(32'h3aae8837),
	.w5(32'h3af8d699),
	.w6(32'hbadf364a),
	.w7(32'h3accf574),
	.w8(32'h3b4fd5ad),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba0b8d),
	.w1(32'hbc075a1e),
	.w2(32'hbc4b6ef2),
	.w3(32'hbb913ae0),
	.w4(32'hbc1f5051),
	.w5(32'hbc8ce7dd),
	.w6(32'h39de3046),
	.w7(32'hbbd71665),
	.w8(32'hbc3b9aff),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb938436),
	.w1(32'h3a97a542),
	.w2(32'h3bbb779f),
	.w3(32'hbc01f140),
	.w4(32'hbabd78f9),
	.w5(32'h3b9940d8),
	.w6(32'hbb7f8b90),
	.w7(32'h3aaef3d2),
	.w8(32'hbb8dbc17),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed1bec),
	.w1(32'h3a86155d),
	.w2(32'h3beebe55),
	.w3(32'h3c3205bd),
	.w4(32'h3b741413),
	.w5(32'hbb27f24f),
	.w6(32'h3bc43798),
	.w7(32'h3b64cdb1),
	.w8(32'hbbc2a4af),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddfc41),
	.w1(32'h3b2c8fd3),
	.w2(32'hbbedf8ec),
	.w3(32'h3a8466ad),
	.w4(32'h3b808fe1),
	.w5(32'hbc0d3b9b),
	.w6(32'h3acd51a6),
	.w7(32'h3a9918c0),
	.w8(32'hbbf67229),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8179a),
	.w1(32'hbb8bbf59),
	.w2(32'h3bb555f5),
	.w3(32'hbc0571c3),
	.w4(32'hbbc0ece2),
	.w5(32'h3bf1c660),
	.w6(32'hbc0900f4),
	.w7(32'hbbe4e8da),
	.w8(32'h3b7c42b9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb716c81),
	.w1(32'hba0dc158),
	.w2(32'h3ac0dd8d),
	.w3(32'hbb6961eb),
	.w4(32'h390614bb),
	.w5(32'h3b378bb8),
	.w6(32'hbadeea62),
	.w7(32'hbb6b2e8f),
	.w8(32'h3b3df019),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec70d7),
	.w1(32'hbb934e6c),
	.w2(32'h3bafd874),
	.w3(32'hbbc165c4),
	.w4(32'hbbbcf279),
	.w5(32'h3b44ed9c),
	.w6(32'hba80ae1f),
	.w7(32'h3ab1d0dc),
	.w8(32'h3b86d251),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8212fc),
	.w1(32'h3b17c085),
	.w2(32'hbb170dad),
	.w3(32'h3c452a74),
	.w4(32'h39f86e1e),
	.w5(32'hbb61dcf9),
	.w6(32'h3c1cbdaf),
	.w7(32'h3b91c6b1),
	.w8(32'hbb03abf4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc215ca),
	.w1(32'hbbf7ea89),
	.w2(32'h3b910563),
	.w3(32'h3c0d2224),
	.w4(32'hbc13faea),
	.w5(32'h3bffbe84),
	.w6(32'h3bef246c),
	.w7(32'hbc708abe),
	.w8(32'h3b8d7ec4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57fdf1),
	.w1(32'hbadf8f5c),
	.w2(32'h3a85c9a4),
	.w3(32'h3be38e0f),
	.w4(32'hbb18dcf1),
	.w5(32'h3b6492ee),
	.w6(32'h3b38ca45),
	.w7(32'hbbc86883),
	.w8(32'h3b202f0a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdb5c8),
	.w1(32'hbbc3cf98),
	.w2(32'hbb8e9920),
	.w3(32'h3b908ce0),
	.w4(32'hbaa649fc),
	.w5(32'hbb495bd7),
	.w6(32'h3b18a484),
	.w7(32'hbba81d46),
	.w8(32'hbc00109d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac74ce4),
	.w1(32'hbacef487),
	.w2(32'h3b06f871),
	.w3(32'h3b551d19),
	.w4(32'h3b26fd47),
	.w5(32'h3b5f3625),
	.w6(32'h3b80c963),
	.w7(32'h3ba1a648),
	.w8(32'hbb0a8e68),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce4d40),
	.w1(32'h3b9c78e2),
	.w2(32'hba3c85d9),
	.w3(32'h3c39617b),
	.w4(32'h3be480aa),
	.w5(32'hbaa8ec66),
	.w6(32'h3c02158e),
	.w7(32'h3b4e207d),
	.w8(32'h3b036335),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a842),
	.w1(32'h3ac2d028),
	.w2(32'hb9ac021e),
	.w3(32'hba21e399),
	.w4(32'hbb969403),
	.w5(32'h38d41ddc),
	.w6(32'h3b1081c0),
	.w7(32'hbb1ea3c7),
	.w8(32'h39f92d25),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e2002),
	.w1(32'hba87df20),
	.w2(32'h3bdb8d90),
	.w3(32'h3b3e4bac),
	.w4(32'hbaf125d3),
	.w5(32'h3c264d96),
	.w6(32'hbb1e386e),
	.w7(32'hbaa2eb0e),
	.w8(32'h3ba9d43c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be77fb0),
	.w1(32'hbb39224f),
	.w2(32'hb988d9a8),
	.w3(32'h3c57fe2b),
	.w4(32'hbb8ecf56),
	.w5(32'hbb008dcf),
	.w6(32'h3c39bb01),
	.w7(32'hbbd7f502),
	.w8(32'h3accede9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50c2ce),
	.w1(32'hbaec13e9),
	.w2(32'h3c8fbb8b),
	.w3(32'h3a2df31c),
	.w4(32'hbb9bd811),
	.w5(32'h3ccf9f14),
	.w6(32'h3b6a4f3d),
	.w7(32'hbb1860fd),
	.w8(32'h3cfc366a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49ec69),
	.w1(32'hba88f74a),
	.w2(32'h3b665a32),
	.w3(32'h3c9685c5),
	.w4(32'h398bb7c8),
	.w5(32'h3baeac63),
	.w6(32'h3ca10ae2),
	.w7(32'hbb03689a),
	.w8(32'h3b97a24d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976258e),
	.w1(32'h3ad55cad),
	.w2(32'hbb6b3350),
	.w3(32'h3be4b89d),
	.w4(32'hbc0ec876),
	.w5(32'h3b42215e),
	.w6(32'h3b11c9cf),
	.w7(32'hbc1a33b9),
	.w8(32'h3b261d92),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba65529),
	.w1(32'h3b8cbb10),
	.w2(32'h3c2298d0),
	.w3(32'h3b92260d),
	.w4(32'h3a61872f),
	.w5(32'h3c256daf),
	.w6(32'h3c0569d1),
	.w7(32'h3bec1068),
	.w8(32'h3c7fc7e7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc91b62),
	.w1(32'hbb921f94),
	.w2(32'hbb420175),
	.w3(32'hba98da4f),
	.w4(32'hbc5bacdd),
	.w5(32'hbaa16d8f),
	.w6(32'h3b9b1713),
	.w7(32'hbc257310),
	.w8(32'h3a9b306a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf67176),
	.w1(32'hbc42fe4c),
	.w2(32'h3ae271ea),
	.w3(32'h3b4d53bc),
	.w4(32'hbc5b8f02),
	.w5(32'h3b714700),
	.w6(32'h3c071065),
	.w7(32'hbc122d1f),
	.w8(32'h3b98bdcc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14129e),
	.w1(32'h3a2eb4df),
	.w2(32'h3b2f175a),
	.w3(32'h3b5f094e),
	.w4(32'hbaa34f71),
	.w5(32'hbb1b280b),
	.w6(32'h3af835dc),
	.w7(32'hb937ba1d),
	.w8(32'hbb91e6d4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c5f63),
	.w1(32'h3baf710f),
	.w2(32'h3b6419ad),
	.w3(32'h3c246b80),
	.w4(32'hbb7933b5),
	.w5(32'h3c760475),
	.w6(32'h3bb91f07),
	.w7(32'h3a75d2fa),
	.w8(32'h3c11bcb4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a005b),
	.w1(32'hbc1b8d15),
	.w2(32'hbc2cb1b5),
	.w3(32'h3a4633e1),
	.w4(32'hbc3d6ff5),
	.w5(32'hbc288722),
	.w6(32'h3b0b9e48),
	.w7(32'hbc4c7119),
	.w8(32'h3aa82c28),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8a4d5),
	.w1(32'h39d50958),
	.w2(32'hbcb435b1),
	.w3(32'hbb408a50),
	.w4(32'h3afd2af1),
	.w5(32'hbcffc599),
	.w6(32'h3c0ecdee),
	.w7(32'h3bb34ea1),
	.w8(32'hbcb8f379),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde61c9),
	.w1(32'h3c16bbe1),
	.w2(32'hba58b8c0),
	.w3(32'hbc614385),
	.w4(32'h3c4b8706),
	.w5(32'h3b7bccf3),
	.w6(32'hbbc9ab3c),
	.w7(32'h3c55d7ac),
	.w8(32'h3b343e10),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31b363),
	.w1(32'hbb11403a),
	.w2(32'hbad8f4cf),
	.w3(32'hbb121a43),
	.w4(32'hbb24fc03),
	.w5(32'h3a432dd2),
	.w6(32'hbad202f1),
	.w7(32'hbb61f318),
	.w8(32'h384708f3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b533781),
	.w1(32'h3b3c577c),
	.w2(32'hbb31cafb),
	.w3(32'h3bca67ac),
	.w4(32'h3b9ea3ea),
	.w5(32'hbb77bd90),
	.w6(32'h3ba414be),
	.w7(32'h3b5dc0b0),
	.w8(32'hbbe8b7a0),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10f2dc),
	.w1(32'h3a207a69),
	.w2(32'hba7538ad),
	.w3(32'h3b5ea4cc),
	.w4(32'h3b1e37da),
	.w5(32'h3c810c44),
	.w6(32'h3ae633dd),
	.w7(32'hbb8797e4),
	.w8(32'hbb2c8386),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba440cbc),
	.w1(32'hb9c2c184),
	.w2(32'h3c614062),
	.w3(32'h3bacaa72),
	.w4(32'h3a74c4f2),
	.w5(32'h3c4afbe4),
	.w6(32'h3b3ca761),
	.w7(32'h3b512abe),
	.w8(32'h3c5ee8de),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27530e),
	.w1(32'h3a588ae5),
	.w2(32'h3b5fc735),
	.w3(32'h3c2362fa),
	.w4(32'h3afb972d),
	.w5(32'h3b85d011),
	.w6(32'h3c20f10e),
	.w7(32'hbb4c5200),
	.w8(32'h3b12d318),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36d023),
	.w1(32'h3c245ab8),
	.w2(32'hbaafa44b),
	.w3(32'h3ba5ba02),
	.w4(32'h3bb4fb20),
	.w5(32'h3a9d6d3c),
	.w6(32'h3c41d79b),
	.w7(32'h3b5ef82e),
	.w8(32'h3ab5b162),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896fcc9),
	.w1(32'h3ae04c9b),
	.w2(32'hba724ecd),
	.w3(32'h3b8fd151),
	.w4(32'hbbc02a37),
	.w5(32'hbbcf8883),
	.w6(32'h3bc238ec),
	.w7(32'hbc022c14),
	.w8(32'hbc2f025d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b852118),
	.w1(32'h3b8d9d8e),
	.w2(32'hbac2509d),
	.w3(32'h3c02e346),
	.w4(32'h3aeb0757),
	.w5(32'h3aba499f),
	.w6(32'h3bbccfd7),
	.w7(32'h3b598ef4),
	.w8(32'h3adf8f53),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54cb1),
	.w1(32'hb993e198),
	.w2(32'h3b3c6de0),
	.w3(32'h3be5e3c6),
	.w4(32'h3bae3245),
	.w5(32'h3ab13461),
	.w6(32'h3b7eaf1d),
	.w7(32'h3b85f259),
	.w8(32'hbb8f795b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5186b),
	.w1(32'h3b8359b3),
	.w2(32'hba9106ab),
	.w3(32'h3c07f277),
	.w4(32'hba9fb9d4),
	.w5(32'h3ac6b8d6),
	.w6(32'h3b649f78),
	.w7(32'h3a1f2926),
	.w8(32'h3b486710),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dfbdb),
	.w1(32'hbbc95175),
	.w2(32'h3b056f33),
	.w3(32'h3b43a791),
	.w4(32'hbc0978b2),
	.w5(32'h3c4f077f),
	.w6(32'h3b8f7804),
	.w7(32'hbbb31e68),
	.w8(32'h3c0583a7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b6d3a),
	.w1(32'hba7d9210),
	.w2(32'h3af3d506),
	.w3(32'h3bf21aaf),
	.w4(32'hbbb5c0fa),
	.w5(32'h3989b79e),
	.w6(32'h3c093010),
	.w7(32'hbc05a3dc),
	.w8(32'hba9ca1a9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b643b36),
	.w1(32'h3ade6be1),
	.w2(32'h3b147af6),
	.w3(32'h3a10f213),
	.w4(32'h3bae2cff),
	.w5(32'h3bb6db21),
	.w6(32'hbb9fbfc7),
	.w7(32'h3a822bc6),
	.w8(32'h3b92f290),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8902a0),
	.w1(32'hbaa598c1),
	.w2(32'h3c12912d),
	.w3(32'hba8671a4),
	.w4(32'hbb1d2c0b),
	.w5(32'h3c4756dd),
	.w6(32'h3adf86af),
	.w7(32'hbb9883ea),
	.w8(32'h3c399acb),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac5260),
	.w1(32'hbc07ca09),
	.w2(32'h3bda1cff),
	.w3(32'hbb1be643),
	.w4(32'hbc584a84),
	.w5(32'h3c456b17),
	.w6(32'h3a8b2d3a),
	.w7(32'hbc408eef),
	.w8(32'h3ac0d6c3),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ab146),
	.w1(32'h3b17bbbd),
	.w2(32'h3b58c6f0),
	.w3(32'h3c5e8e82),
	.w4(32'hbafb9036),
	.w5(32'h3bea5f4e),
	.w6(32'h3c114c63),
	.w7(32'h3a1f83d4),
	.w8(32'h3be8a9f3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a3e55),
	.w1(32'h3b5b0dbf),
	.w2(32'h3b977a97),
	.w3(32'h3c511dc8),
	.w4(32'h3a9a5d68),
	.w5(32'h3b9bc842),
	.w6(32'h3c600660),
	.w7(32'h3b901285),
	.w8(32'h3b498006),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e4fd9),
	.w1(32'h3b7d79f4),
	.w2(32'h3a4404f5),
	.w3(32'h3c234405),
	.w4(32'h3b9aa4c2),
	.w5(32'h3a6ab919),
	.w6(32'h3b15212a),
	.w7(32'hbb001aee),
	.w8(32'h3ad832f9),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb7738),
	.w1(32'h3b577b0a),
	.w2(32'h3b242a12),
	.w3(32'h3c2a2ba6),
	.w4(32'h3be8bf1d),
	.w5(32'h3a8352ce),
	.w6(32'h3bff2ce4),
	.w7(32'hb9ea54c4),
	.w8(32'hbb5739a5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac17a02),
	.w1(32'hbb00d6df),
	.w2(32'h3c0e25e2),
	.w3(32'hbb88b5de),
	.w4(32'hbb99acff),
	.w5(32'h3ca28e91),
	.w6(32'hbb2bf6a1),
	.w7(32'hbc0139e0),
	.w8(32'h3c64e57d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66f68e),
	.w1(32'hb9537978),
	.w2(32'h3ba6f0b7),
	.w3(32'h3c25933f),
	.w4(32'hbbb63ab9),
	.w5(32'h3bc62677),
	.w6(32'hbae2b608),
	.w7(32'hbb84c792),
	.w8(32'hbab45387),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3371c8),
	.w1(32'h3a36efd2),
	.w2(32'h3b19fffa),
	.w3(32'h3bbd358e),
	.w4(32'hbb3098fa),
	.w5(32'hba87abf0),
	.w6(32'h3a353c55),
	.w7(32'hbb44696f),
	.w8(32'hbc0ab8ce),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dca9b),
	.w1(32'hbbbe58af),
	.w2(32'h3b4c3a5e),
	.w3(32'h3b1e1d78),
	.w4(32'hb9fa0670),
	.w5(32'hb909fe10),
	.w6(32'hbb0179b0),
	.w7(32'hbb59ef37),
	.w8(32'hbbd6cf05),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3f7d5),
	.w1(32'hbaaf9ed4),
	.w2(32'hbacee4ff),
	.w3(32'hba975222),
	.w4(32'hbbbc637d),
	.w5(32'hb9f38bf4),
	.w6(32'hbb98043a),
	.w7(32'hbb26b449),
	.w8(32'hbb80a7d1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0930b1),
	.w1(32'hbb563d1c),
	.w2(32'h3baac626),
	.w3(32'h3b1c47d4),
	.w4(32'hbb807621),
	.w5(32'h3b741fca),
	.w6(32'h3bc22849),
	.w7(32'h3b7822ff),
	.w8(32'hbadc4e03),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fe62a),
	.w1(32'hbb07766f),
	.w2(32'h3bd194e6),
	.w3(32'h3af68879),
	.w4(32'hbbec1d74),
	.w5(32'h3ba9e78f),
	.w6(32'hbb16b2ee),
	.w7(32'hbbf7e528),
	.w8(32'h3b8ef5fd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6da86a),
	.w1(32'h3a692ce0),
	.w2(32'hbb0d1aa1),
	.w3(32'h3c899140),
	.w4(32'h3ba37a68),
	.w5(32'hba2b78c4),
	.w6(32'h3c0c1023),
	.w7(32'h3a9ed672),
	.w8(32'hbbb977e5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbafc1b),
	.w1(32'hbb41688b),
	.w2(32'hbb7dceb9),
	.w3(32'h3b4360c0),
	.w4(32'hb9f3e104),
	.w5(32'h3a917e0a),
	.w6(32'h3b3b8f73),
	.w7(32'hba090b2b),
	.w8(32'hb9c8c37a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b12da),
	.w1(32'hbb16f283),
	.w2(32'h3a798d1e),
	.w3(32'h3b682ad3),
	.w4(32'h3b237985),
	.w5(32'h3b5858d4),
	.w6(32'h3b4b2bb7),
	.w7(32'hb96362f5),
	.w8(32'h3a9ed091),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a32d60),
	.w1(32'hba412858),
	.w2(32'h3b31cdf9),
	.w3(32'h3a207d4b),
	.w4(32'hbac0901c),
	.w5(32'h3b7df8b9),
	.w6(32'hba182317),
	.w7(32'hbaf4cea6),
	.w8(32'h3b48ace9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed6d5a),
	.w1(32'hbae20aac),
	.w2(32'hbbd90ba2),
	.w3(32'h3b451080),
	.w4(32'hbacaee6c),
	.w5(32'hbb1469d7),
	.w6(32'h3b62b127),
	.w7(32'hb95ecd31),
	.w8(32'hbbabc14b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc291c9c),
	.w1(32'hbbd4edfc),
	.w2(32'h3b658f5c),
	.w3(32'h3b52b6a8),
	.w4(32'hbbbbac7d),
	.w5(32'h3b8945f3),
	.w6(32'h3ad60595),
	.w7(32'hbbca9cab),
	.w8(32'h3b21eaee),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65cd50),
	.w1(32'hbb829332),
	.w2(32'h3b29848b),
	.w3(32'hbb9a883a),
	.w4(32'hbbf3d738),
	.w5(32'h3ae18d6f),
	.w6(32'hbb3c4969),
	.w7(32'hbbb245ca),
	.w8(32'h3bb91eba),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb0941),
	.w1(32'h38c664d9),
	.w2(32'h3b82892d),
	.w3(32'h3be43816),
	.w4(32'hbada54d2),
	.w5(32'h3aaa1749),
	.w6(32'hbb62bdb8),
	.w7(32'hbbceda4a),
	.w8(32'h3a875c41),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6795e2),
	.w1(32'hba3a1348),
	.w2(32'hbb647bbc),
	.w3(32'h3c4c53ce),
	.w4(32'h3a588701),
	.w5(32'h3bcb22c9),
	.w6(32'h3bf6d41f),
	.w7(32'h3b6bf1fb),
	.w8(32'h3c2541c4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc978a),
	.w1(32'hbbae5b04),
	.w2(32'h3c4b5ddb),
	.w3(32'h3bf3b46b),
	.w4(32'hbbb6ccc6),
	.w5(32'h3ca7c3f2),
	.w6(32'h3b8d1c2e),
	.w7(32'hbbe1c71d),
	.w8(32'h3c066da4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule