module layer_8_featuremap_102(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8851f3),
	.w1(32'hbbf6cec2),
	.w2(32'h3d1028f1),
	.w3(32'hbc0e0999),
	.w4(32'h3cf1e6cd),
	.w5(32'h3d6c9297),
	.w6(32'hbc1c97cb),
	.w7(32'h3d7198d6),
	.w8(32'h3d39475d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a38a5),
	.w1(32'hbc4a01fa),
	.w2(32'hbcb434df),
	.w3(32'h3b1bf7ff),
	.w4(32'hbc2491f5),
	.w5(32'hbc407f9f),
	.w6(32'hbcc2c38e),
	.w7(32'hbc713a1d),
	.w8(32'hbc84a132),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3b93a),
	.w1(32'h3d19a80b),
	.w2(32'h3bbf1fd4),
	.w3(32'h3c553ae0),
	.w4(32'hbb83542b),
	.w5(32'hbbc2b584),
	.w6(32'h3d0caf75),
	.w7(32'hbb62bbb4),
	.w8(32'hbc794b13),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99e6dd),
	.w1(32'h3b3c31f0),
	.w2(32'h3cc93aa9),
	.w3(32'hbc9cc55f),
	.w4(32'hbbbe3cad),
	.w5(32'h3a85e70f),
	.w6(32'h3c2398f3),
	.w7(32'h3cb18a54),
	.w8(32'h3c3fec8c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35d1e1),
	.w1(32'hbc3b3efb),
	.w2(32'h3cc69ac0),
	.w3(32'h3c08c068),
	.w4(32'h3b9c5a6d),
	.w5(32'hbb60307e),
	.w6(32'h3c2645c6),
	.w7(32'h3b550f15),
	.w8(32'hbb7389ab),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80d78c),
	.w1(32'hbca112bc),
	.w2(32'hbcd1cd81),
	.w3(32'hbc6deb31),
	.w4(32'hbc9783a6),
	.w5(32'hbd798cbd),
	.w6(32'hbd0918f8),
	.w7(32'hbcff6430),
	.w8(32'hbd168f5d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccebf9b),
	.w1(32'h3ceb4dbb),
	.w2(32'h3c991a1a),
	.w3(32'h3c5a880d),
	.w4(32'hbbe6db37),
	.w5(32'hbc2c4a4d),
	.w6(32'h3cf8d75b),
	.w7(32'h3b1f8c64),
	.w8(32'h3c0186d3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbee8ac),
	.w1(32'h3c9b8cb1),
	.w2(32'hbb4c6040),
	.w3(32'hbce4eaff),
	.w4(32'h3c4dc518),
	.w5(32'h3c3fd708),
	.w6(32'h3c1bd507),
	.w7(32'h3cda3c41),
	.w8(32'hbc2f91d9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e64a0),
	.w1(32'hbb94d229),
	.w2(32'h3cbd4055),
	.w3(32'h3b0b6108),
	.w4(32'h3c50af4b),
	.w5(32'h3a9aa4fb),
	.w6(32'hbc0a8986),
	.w7(32'h3d0b89b5),
	.w8(32'h3ba31f63),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1df786),
	.w1(32'hbc5e3c35),
	.w2(32'h3c4651e4),
	.w3(32'hbd06e112),
	.w4(32'h3c823bb0),
	.w5(32'h3cad95d9),
	.w6(32'hbcfe517d),
	.w7(32'h3c0ef9e2),
	.w8(32'h3ca5d9da),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a5f1b),
	.w1(32'h3c0d7aa2),
	.w2(32'h3d1093a3),
	.w3(32'h3acffc62),
	.w4(32'h3cb56055),
	.w5(32'h3d20b37c),
	.w6(32'h3caecd0c),
	.w7(32'h3d0aa911),
	.w8(32'h3d50510d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96bd84),
	.w1(32'hbd08989d),
	.w2(32'h3a7648b3),
	.w3(32'hbcd88b53),
	.w4(32'h3b3c0441),
	.w5(32'h3bde6747),
	.w6(32'hbcbe4ca8),
	.w7(32'h3c7a0f41),
	.w8(32'h3c58a433),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba65713),
	.w1(32'h3b1b5090),
	.w2(32'hbba4dda7),
	.w3(32'hba718917),
	.w4(32'h3ba7ef19),
	.w5(32'hba0ba26e),
	.w6(32'h3979b45c),
	.w7(32'hbb497dd0),
	.w8(32'hbc1ee8c6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b219811),
	.w1(32'h3b4dd927),
	.w2(32'hba9a660c),
	.w3(32'h3a8fd20e),
	.w4(32'h3a7ab71d),
	.w5(32'hbb22315c),
	.w6(32'h3bb2855b),
	.w7(32'hbc100a5e),
	.w8(32'hbbd252fc),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae19f60),
	.w1(32'hba79b118),
	.w2(32'h3b11a235),
	.w3(32'hba0a6b34),
	.w4(32'h3be55ab7),
	.w5(32'hba727c65),
	.w6(32'hb966007c),
	.w7(32'hbab4d5fa),
	.w8(32'hbba86ac4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cdfde),
	.w1(32'hbb164382),
	.w2(32'h3c11941b),
	.w3(32'hba7df14d),
	.w4(32'hbc2ca3f6),
	.w5(32'h3c320372),
	.w6(32'hbb7cc1ff),
	.w7(32'h3c71d0c3),
	.w8(32'h3ca3b1c7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d0578),
	.w1(32'h3cb36461),
	.w2(32'h3c75d632),
	.w3(32'hbb0b6451),
	.w4(32'hbc8c91f3),
	.w5(32'hb97862c9),
	.w6(32'hbd00c299),
	.w7(32'hbb89fd3a),
	.w8(32'hba12bcfc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd108036),
	.w1(32'hbcb54420),
	.w2(32'hbc2305ab),
	.w3(32'h39e805d5),
	.w4(32'h3c48066e),
	.w5(32'hbc0335a5),
	.w6(32'h3bd93775),
	.w7(32'hbc08c515),
	.w8(32'hbbb45947),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd36c3d6),
	.w1(32'hbcdc5ab4),
	.w2(32'h3d328bdf),
	.w3(32'hbd586e74),
	.w4(32'hbc221507),
	.w5(32'h3d8b4492),
	.w6(32'h3ce00dee),
	.w7(32'h3d907222),
	.w8(32'h3d9397d4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee1664),
	.w1(32'hbc9c937e),
	.w2(32'h3b89135e),
	.w3(32'hbc11da68),
	.w4(32'h3c1cf29d),
	.w5(32'h3c310a0f),
	.w6(32'hbb8b6709),
	.w7(32'hbab66bf8),
	.w8(32'hbcfb8af5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba38d7e),
	.w1(32'hbb6d2cdc),
	.w2(32'hbac9b69f),
	.w3(32'hbb2169a6),
	.w4(32'h3b1be93a),
	.w5(32'hbd0e3949),
	.w6(32'h3b16b1cb),
	.w7(32'hbc92e5af),
	.w8(32'h3be09768),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fc39e),
	.w1(32'h3caa74a8),
	.w2(32'h3c45a7ed),
	.w3(32'hba0e3c4d),
	.w4(32'hbc59ba46),
	.w5(32'hba3ecb8a),
	.w6(32'hbcb258d6),
	.w7(32'hbca56d2e),
	.w8(32'hbc49263e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3a09f0),
	.w1(32'hbd736144),
	.w2(32'h3d257192),
	.w3(32'hbc89a19e),
	.w4(32'h3c99cd3b),
	.w5(32'h3d8fdfb7),
	.w6(32'h3b8858f7),
	.w7(32'h3d2e8ac2),
	.w8(32'h3dc71018),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ffb0c),
	.w1(32'h3c05f8c2),
	.w2(32'h3c112663),
	.w3(32'hbb156535),
	.w4(32'h3c8c8fec),
	.w5(32'h3c0ab685),
	.w6(32'hbc8be7c4),
	.w7(32'hbaa2b1de),
	.w8(32'hbaaf2563),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c129db0),
	.w1(32'h3bda5c6e),
	.w2(32'hbac3c903),
	.w3(32'h3a75a3ee),
	.w4(32'hbc072c26),
	.w5(32'hbc3b416a),
	.w6(32'h3bd5952c),
	.w7(32'hbb961857),
	.w8(32'hbab7eaa8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc955049),
	.w1(32'hbc2a872f),
	.w2(32'h3d0d3a21),
	.w3(32'hbc548135),
	.w4(32'hbd00983e),
	.w5(32'h3c27aa06),
	.w6(32'h3b054b72),
	.w7(32'hba331dab),
	.w8(32'h3d567c24),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fe12d),
	.w1(32'hbd62bb5b),
	.w2(32'hbbcb4126),
	.w3(32'h3d474110),
	.w4(32'hb9124784),
	.w5(32'h3c1bffd0),
	.w6(32'h3ba03c78),
	.w7(32'h3bddef04),
	.w8(32'hbc7a6886),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdcddfbd),
	.w1(32'h3d2f2992),
	.w2(32'hbbc4304a),
	.w3(32'hbd9a88ec),
	.w4(32'hbd0e8045),
	.w5(32'hbd3b1c01),
	.w6(32'hbd6ed9de),
	.w7(32'hbd2564fa),
	.w8(32'h3d844968),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09d758),
	.w1(32'hbc1b7d40),
	.w2(32'h3cd4913c),
	.w3(32'hbb0f7de3),
	.w4(32'hbb3a0f0e),
	.w5(32'h3d06e241),
	.w6(32'h3c409b3a),
	.w7(32'h3cf04521),
	.w8(32'h3d1d38f2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1fb54),
	.w1(32'hbd0f23cd),
	.w2(32'h3b3c3ba3),
	.w3(32'h3ae1cb13),
	.w4(32'hbb4a84f3),
	.w5(32'hbbc14a44),
	.w6(32'h3d090091),
	.w7(32'hbc34489d),
	.w8(32'h3ce9c094),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fd465),
	.w1(32'h3ca56520),
	.w2(32'h3c16f181),
	.w3(32'h3bbdc19f),
	.w4(32'h3c053dee),
	.w5(32'h3b9f3f92),
	.w6(32'hbc79dff7),
	.w7(32'h3b4363e0),
	.w8(32'h3b211c79),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcd58d),
	.w1(32'hba0ee32f),
	.w2(32'hbcd5a1d4),
	.w3(32'h3be1758c),
	.w4(32'h3b65622c),
	.w5(32'hbb7ee529),
	.w6(32'hb8164043),
	.w7(32'hbc5ece73),
	.w8(32'hbcdbcbf7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2415f2),
	.w1(32'hbc2f5471),
	.w2(32'h3c452cf8),
	.w3(32'hbc673c83),
	.w4(32'hbb2c87e3),
	.w5(32'hbc7dbd59),
	.w6(32'hbc32792e),
	.w7(32'hbc8ca21d),
	.w8(32'h3ca41409),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164bb4),
	.w1(32'hbcc298bb),
	.w2(32'hbbcfc607),
	.w3(32'h3c9e0c03),
	.w4(32'h3c3ad791),
	.w5(32'hbc1a0f4f),
	.w6(32'h3c8fac0e),
	.w7(32'hbb864318),
	.w8(32'hbc98f7d9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57e86b),
	.w1(32'h3cf8fe7f),
	.w2(32'h3b0ffe53),
	.w3(32'hbbb1f453),
	.w4(32'h3b4f78df),
	.w5(32'hbbc2a8f2),
	.w6(32'h3c05e30f),
	.w7(32'hbc6bfcde),
	.w8(32'hbc15060f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbae546),
	.w1(32'hbc521b5b),
	.w2(32'h3ca89b51),
	.w3(32'hbbffa78b),
	.w4(32'hbb45c5c8),
	.w5(32'h3c2a6de1),
	.w6(32'hbc5bc59c),
	.w7(32'hbbc29586),
	.w8(32'h3c289829),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ef5e2),
	.w1(32'hbca920f7),
	.w2(32'h3c9bbf8a),
	.w3(32'h3c5504b0),
	.w4(32'hbbb161ad),
	.w5(32'h3bfa2bfb),
	.w6(32'h3bc122ca),
	.w7(32'hbc3e8aef),
	.w8(32'hbb7ffb53),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5c41c),
	.w1(32'hbd323840),
	.w2(32'hbc4cc0ef),
	.w3(32'h3a7389fa),
	.w4(32'hbb920731),
	.w5(32'hbc72aedb),
	.w6(32'hbc11e748),
	.w7(32'h3b8295f5),
	.w8(32'hbc919c1f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fdddc),
	.w1(32'h3b18a27c),
	.w2(32'h3c453170),
	.w3(32'hbbedb327),
	.w4(32'hbca86a79),
	.w5(32'hbc20e6b9),
	.w6(32'h3a21a9f3),
	.w7(32'hbbac5837),
	.w8(32'hbc930f6f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5163b3),
	.w1(32'hbd574195),
	.w2(32'hb9891235),
	.w3(32'h3cbc5468),
	.w4(32'hbbcbf389),
	.w5(32'h3b8498f9),
	.w6(32'hbc07e692),
	.w7(32'h3bd42086),
	.w8(32'h3c70101e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd32f623),
	.w1(32'hbc888900),
	.w2(32'hbc6d48c3),
	.w3(32'hbd0e4587),
	.w4(32'h3a63ab51),
	.w5(32'h3c482e2b),
	.w6(32'h381915c5),
	.w7(32'h3cea4154),
	.w8(32'hbd143dd3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7ccd1),
	.w1(32'hbab167e9),
	.w2(32'hbcaf6051),
	.w3(32'hbd09b778),
	.w4(32'h3a1d9837),
	.w5(32'h3b39f4af),
	.w6(32'hbc25c8c5),
	.w7(32'hb83c0711),
	.w8(32'hbbf0da76),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32e02e),
	.w1(32'h3d204c4d),
	.w2(32'h3c5eca97),
	.w3(32'hbcf91b76),
	.w4(32'hbc866608),
	.w5(32'hbc4f76cb),
	.w6(32'hbc17e5a9),
	.w7(32'hbb90c32a),
	.w8(32'h3c9db33a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd8208),
	.w1(32'hbc8969b8),
	.w2(32'h3c000952),
	.w3(32'h3c4216a0),
	.w4(32'hba83e613),
	.w5(32'h3c35b245),
	.w6(32'hbb1641a3),
	.w7(32'h3c137fd2),
	.w8(32'h3c95394a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c6ec2),
	.w1(32'hbbce3b87),
	.w2(32'h3c86cc09),
	.w3(32'hbb2b5b5f),
	.w4(32'hbcfc82ae),
	.w5(32'h3d10f1d0),
	.w6(32'h3c90ab6a),
	.w7(32'h3cf9755a),
	.w8(32'h3d1b2347),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6324e3),
	.w1(32'hbd36edd0),
	.w2(32'h3cdf37d2),
	.w3(32'hbc59f2e7),
	.w4(32'hbc06bf66),
	.w5(32'h3c37eaaa),
	.w6(32'hbc438ccd),
	.w7(32'h3bfe6daf),
	.w8(32'h3cd774da),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56734c),
	.w1(32'hbbd9cdd6),
	.w2(32'h3ca30b10),
	.w3(32'h3c3b1c5d),
	.w4(32'hbcabbc2e),
	.w5(32'h3bceae1c),
	.w6(32'hbb5412f5),
	.w7(32'h3983a51a),
	.w8(32'h3c6e5be0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9c35d),
	.w1(32'hbd83056f),
	.w2(32'h3d285c2e),
	.w3(32'h3c13ffea),
	.w4(32'hbd1e8166),
	.w5(32'h3d20ea7f),
	.w6(32'h3b4ff7b1),
	.w7(32'h3c8f0eb9),
	.w8(32'h3d517314),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03f92c),
	.w1(32'hbd5d4846),
	.w2(32'hbd12d78c),
	.w3(32'h3c917e90),
	.w4(32'h3c2175d9),
	.w5(32'h3af21934),
	.w6(32'h3c8ebcfa),
	.w7(32'h3b628e11),
	.w8(32'hbcc473f7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d6a4),
	.w1(32'h3c6b0937),
	.w2(32'hbc729fc5),
	.w3(32'hbd03f846),
	.w4(32'hbca1c63f),
	.w5(32'h3c430de3),
	.w6(32'hbc17c59a),
	.w7(32'h3b5e8d16),
	.w8(32'hbc65607f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60ac04),
	.w1(32'hbd06f28f),
	.w2(32'hbd68c29a),
	.w3(32'hbd1e4c88),
	.w4(32'h3c2cf5df),
	.w5(32'hbd20b1b2),
	.w6(32'hbbe17ab0),
	.w7(32'hbc5d9c24),
	.w8(32'hbc9c20f2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0df1d1),
	.w1(32'h3cd49c53),
	.w2(32'h3cb6e43d),
	.w3(32'hbd9fb395),
	.w4(32'hbd0a6eaf),
	.w5(32'h3c8ff4ed),
	.w6(32'hbca91de5),
	.w7(32'h3c4bea6d),
	.w8(32'h3d6d6070),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06dedf),
	.w1(32'hbbe6f858),
	.w2(32'hbc61fd29),
	.w3(32'h3bf48fb1),
	.w4(32'h3ca41e1a),
	.w5(32'h3b8f853c),
	.w6(32'hbc4c6f8d),
	.w7(32'h3b85e5cb),
	.w8(32'hba1bc546),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce002e0),
	.w1(32'hbc98d7b3),
	.w2(32'h3842a435),
	.w3(32'hbcb260be),
	.w4(32'h3c3e5fe5),
	.w5(32'h3d1706be),
	.w6(32'h3d262210),
	.w7(32'h3c8ab2db),
	.w8(32'h3c9e1c0f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6620c6),
	.w1(32'h3b0004ae),
	.w2(32'h3bd601c1),
	.w3(32'h3aa5ad53),
	.w4(32'hbc9ab7e7),
	.w5(32'h3ba645b9),
	.w6(32'h3bd82bcb),
	.w7(32'h3c80df3e),
	.w8(32'h3c341cae),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee2d2a),
	.w1(32'hbd883daa),
	.w2(32'h3a9534f1),
	.w3(32'h3c33766f),
	.w4(32'h3b435fba),
	.w5(32'h3c98cab7),
	.w6(32'hbc72883e),
	.w7(32'h3d18ffac),
	.w8(32'h3cfc99c5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b3c01),
	.w1(32'hbc209c1f),
	.w2(32'hbb24766e),
	.w3(32'hbb3bfc1f),
	.w4(32'h3b98ec8b),
	.w5(32'h3c0c138f),
	.w6(32'h3c0f8de6),
	.w7(32'h3b950066),
	.w8(32'hbb39db7a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d36f3),
	.w1(32'hbbc7146d),
	.w2(32'h3c5bccb8),
	.w3(32'hbcf2db76),
	.w4(32'hbc4cd7a5),
	.w5(32'h3c772c43),
	.w6(32'hbc829d4b),
	.w7(32'h3b735ff8),
	.w8(32'h3cd52296),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce38216),
	.w1(32'h3bc2fa8c),
	.w2(32'h3bd945a0),
	.w3(32'hbbcc0b95),
	.w4(32'hbb988144),
	.w5(32'h3c6cf435),
	.w6(32'hbafa7cbd),
	.w7(32'h3ab3475b),
	.w8(32'h3ccd6318),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b348551),
	.w1(32'h3b4f53b9),
	.w2(32'h3b6e21fb),
	.w3(32'hb9f09e50),
	.w4(32'hbb8ecb25),
	.w5(32'hbc3cce31),
	.w6(32'h3b75fd3b),
	.w7(32'hbc6eeffb),
	.w8(32'h3d004d75),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64fbf9),
	.w1(32'hbc15ee70),
	.w2(32'hbd002f5b),
	.w3(32'h3b84200f),
	.w4(32'h3cc589d2),
	.w5(32'h3a748674),
	.w6(32'hbbd9e431),
	.w7(32'h3bd1d88c),
	.w8(32'hbc55512f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca514ca),
	.w1(32'h3ce27d0d),
	.w2(32'h3a9b9f64),
	.w3(32'hbd10bee8),
	.w4(32'hbc00c3be),
	.w5(32'hba855001),
	.w6(32'h3c5752ab),
	.w7(32'h3b9f5858),
	.w8(32'h3c177c7e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd35c41),
	.w1(32'hbcb6ad66),
	.w2(32'h3b739a78),
	.w3(32'hbc81dbff),
	.w4(32'h3c035a7a),
	.w5(32'h3cd1b876),
	.w6(32'h3b819130),
	.w7(32'h3d15a150),
	.w8(32'h3ba2393b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a5990),
	.w1(32'hbb58902d),
	.w2(32'hbac2eb52),
	.w3(32'h3c02b740),
	.w4(32'h3c05ff4e),
	.w5(32'h392712fd),
	.w6(32'h3b5761a0),
	.w7(32'hbb414bc2),
	.w8(32'hbb9b6427),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8642ec),
	.w1(32'h3ae5ede6),
	.w2(32'h3cab8db4),
	.w3(32'h3c4bec97),
	.w4(32'h3bb2c4f3),
	.w5(32'hbabda8ce),
	.w6(32'h396ae8c1),
	.w7(32'h3cb15bd3),
	.w8(32'h3c7ae659),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55f8d0),
	.w1(32'hbbf28f37),
	.w2(32'h3bfe889a),
	.w3(32'h3c59c8e5),
	.w4(32'h3c2630bb),
	.w5(32'hbb3ddfe0),
	.w6(32'hbbe1a2cd),
	.w7(32'h3b8c33df),
	.w8(32'h3c309758),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d2d1c),
	.w1(32'h3c802e21),
	.w2(32'hbc89de62),
	.w3(32'hba79eff8),
	.w4(32'hbca78eb7),
	.w5(32'hbce80b29),
	.w6(32'h3bb4890c),
	.w7(32'h3b85dae4),
	.w8(32'hbcb29225),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c5a1ef),
	.w1(32'hbd3773b0),
	.w2(32'hbd33ffaf),
	.w3(32'h3c5b1dbf),
	.w4(32'h3b67a8b1),
	.w5(32'hbc85e846),
	.w6(32'h3c361785),
	.w7(32'h3c9a1464),
	.w8(32'hbc3fa597),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf75c28),
	.w1(32'h3d40c5d7),
	.w2(32'hbb84faae),
	.w3(32'hbcc75e6e),
	.w4(32'hbbfd1667),
	.w5(32'h3b2c9317),
	.w6(32'hbb98d199),
	.w7(32'hbc3f68ed),
	.w8(32'hbcbd5b91),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23bfb5),
	.w1(32'hbc815408),
	.w2(32'hbc7c7a10),
	.w3(32'hbc22eff9),
	.w4(32'h3aa53cd6),
	.w5(32'h3c529737),
	.w6(32'hbd05008b),
	.w7(32'h3b54d102),
	.w8(32'h3d512f74),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cef1176),
	.w1(32'h3d655dc9),
	.w2(32'hbc94f957),
	.w3(32'hbd28f7bd),
	.w4(32'h3be8f796),
	.w5(32'h3cacdfdd),
	.w6(32'h3c77c397),
	.w7(32'h3d100647),
	.w8(32'h3bb14a43),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c111b82),
	.w1(32'h3d222ea2),
	.w2(32'hbbab84f8),
	.w3(32'hbcddc250),
	.w4(32'h3ba28413),
	.w5(32'h3ca60a19),
	.w6(32'h3ad17119),
	.w7(32'h3ca05152),
	.w8(32'hbabfcf08),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399782b5),
	.w1(32'h3d10a3d4),
	.w2(32'hbca139e5),
	.w3(32'h3c5325a8),
	.w4(32'h3bae9cd4),
	.w5(32'hbba43582),
	.w6(32'h3bb51038),
	.w7(32'hb7b00f64),
	.w8(32'hbca33f7e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24bb4f),
	.w1(32'h3b89e252),
	.w2(32'hbd2d5705),
	.w3(32'hbc8a1a49),
	.w4(32'h3d32915b),
	.w5(32'hbae4d603),
	.w6(32'h3c26111f),
	.w7(32'h3be21935),
	.w8(32'hbbefe7ed),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ef097),
	.w1(32'h3d8a20de),
	.w2(32'h3cf01f6c),
	.w3(32'hbd43d4a5),
	.w4(32'hbc4922e9),
	.w5(32'h3c85a6de),
	.w6(32'h3b523f1d),
	.w7(32'hbcab732e),
	.w8(32'h3c19f95f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3d56c),
	.w1(32'hbd3aff75),
	.w2(32'hbcb2182c),
	.w3(32'h3c15bb1e),
	.w4(32'h3c5548c3),
	.w5(32'hbc9ccd10),
	.w6(32'h3cacc900),
	.w7(32'h3bacc3ff),
	.w8(32'hbbb61e38),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e1ba9),
	.w1(32'hbc68fabe),
	.w2(32'h3b4b2c85),
	.w3(32'h3b004db5),
	.w4(32'h3a24850a),
	.w5(32'h3bb3c9f5),
	.w6(32'h3b7e3522),
	.w7(32'h3bd20c4c),
	.w8(32'hbb93b06f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb50a65),
	.w1(32'hbb691e52),
	.w2(32'h3c040c4e),
	.w3(32'hbc03f6b4),
	.w4(32'hbb33747b),
	.w5(32'h3c09eada),
	.w6(32'hbab9a772),
	.w7(32'h3c80581e),
	.w8(32'h3c917c94),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc871107),
	.w1(32'hbb7665cb),
	.w2(32'h3c3c0032),
	.w3(32'hbc3d87d1),
	.w4(32'hbaf19f21),
	.w5(32'h3cab78bd),
	.w6(32'hbc48abe7),
	.w7(32'h3bf2a69b),
	.w8(32'h3c821130),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b341704),
	.w1(32'h3b46573c),
	.w2(32'h3b5d36a0),
	.w3(32'h3b4b3568),
	.w4(32'h3be87648),
	.w5(32'hb98ff9d3),
	.w6(32'h3a7dcb94),
	.w7(32'h3ccf4891),
	.w8(32'hbb8b584f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b083112),
	.w1(32'h3c25b4b1),
	.w2(32'hbc8de1c0),
	.w3(32'h3bccf781),
	.w4(32'h3b1fadea),
	.w5(32'hbcabd2ee),
	.w6(32'h3c2aa77b),
	.w7(32'h3cd7bae0),
	.w8(32'h3ceb67e7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08e00c),
	.w1(32'hbc88cac4),
	.w2(32'hbbb2146c),
	.w3(32'hbcad53a5),
	.w4(32'hbb8a36ed),
	.w5(32'h3a931357),
	.w6(32'hbd1c339d),
	.w7(32'hbcd72708),
	.w8(32'hbafcad6a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea2b4b),
	.w1(32'hbbf9baeb),
	.w2(32'hbc6bbd66),
	.w3(32'h3badda22),
	.w4(32'hbc00c96c),
	.w5(32'hbad7763e),
	.w6(32'h3b66d320),
	.w7(32'h3bea1c1c),
	.w8(32'h3c40e9a3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0cf22),
	.w1(32'hbcc2db68),
	.w2(32'hbd3b70d0),
	.w3(32'hbd642c2f),
	.w4(32'hbb98fc48),
	.w5(32'hbcd4a970),
	.w6(32'hbccf4cdd),
	.w7(32'h3cc53039),
	.w8(32'hbd5ef447),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd33edcb),
	.w1(32'hbc530bee),
	.w2(32'h3c9b6bfd),
	.w3(32'hbc4e4498),
	.w4(32'h3bc45b7a),
	.w5(32'h3ce63558),
	.w6(32'h3ad83e1d),
	.w7(32'h3d34638f),
	.w8(32'h3d5918c2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbafb2d),
	.w1(32'hbc652691),
	.w2(32'hba3cce81),
	.w3(32'hbc393e48),
	.w4(32'hbb7cfcc0),
	.w5(32'h3a7fb8c9),
	.w6(32'hbd00622b),
	.w7(32'hbcd21bf4),
	.w8(32'h3d2a19d3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7aa5c),
	.w1(32'hbc734027),
	.w2(32'h3b970a74),
	.w3(32'hbbf92641),
	.w4(32'hbc063821),
	.w5(32'hbbee32d1),
	.w6(32'hbc6037fe),
	.w7(32'h3ac21f85),
	.w8(32'hbc813f21),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc1ab9),
	.w1(32'hba235080),
	.w2(32'h3bb09163),
	.w3(32'h3c414fec),
	.w4(32'hbbdcba23),
	.w5(32'hbc1c3944),
	.w6(32'h3c694edf),
	.w7(32'hba118dc4),
	.w8(32'h3a761d09),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8884),
	.w1(32'hb859317d),
	.w2(32'hbb8a2ff4),
	.w3(32'hbb0e1bb9),
	.w4(32'h3ab5b766),
	.w5(32'hba279eb0),
	.w6(32'h3b92db9c),
	.w7(32'hbaefa1ce),
	.w8(32'h3bfcdf33),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e9a3d),
	.w1(32'hbbd85ac4),
	.w2(32'hbc1ab943),
	.w3(32'h3b70085b),
	.w4(32'hbc0912a8),
	.w5(32'hbc20e1f4),
	.w6(32'hba57f4cc),
	.w7(32'h3c709b8b),
	.w8(32'h3d1e34a8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf60cf3),
	.w1(32'hbba186ae),
	.w2(32'h3bdf4829),
	.w3(32'h3bf7dc57),
	.w4(32'hbaa44c15),
	.w5(32'h3bc865f3),
	.w6(32'h3bcc12b8),
	.w7(32'h3ae0e02c),
	.w8(32'hbc321e9f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26b955),
	.w1(32'hbb9d3994),
	.w2(32'h3c1be19b),
	.w3(32'h3c323a8f),
	.w4(32'h3bcc15c7),
	.w5(32'hbd19c012),
	.w6(32'h3be5c7d1),
	.w7(32'h3bd539ea),
	.w8(32'hbcd89ece),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92668b),
	.w1(32'h3ca0eb29),
	.w2(32'h3b81336c),
	.w3(32'h3cafa778),
	.w4(32'hbc5119b1),
	.w5(32'h3a43ce5c),
	.w6(32'hb88cba6c),
	.w7(32'hbcaa42b7),
	.w8(32'h3be948e3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad7125),
	.w1(32'hbb5b4aa3),
	.w2(32'hbc4a0983),
	.w3(32'h3b93ab4e),
	.w4(32'hbc1529e6),
	.w5(32'h3ca53313),
	.w6(32'hbc4c43e1),
	.w7(32'hbb814c60),
	.w8(32'h3d3c1a20),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c605342),
	.w1(32'hbc763db2),
	.w2(32'h3aa1e908),
	.w3(32'h3a7d9416),
	.w4(32'h3be9acf9),
	.w5(32'h3a83aaf9),
	.w6(32'hbc5d4eaf),
	.w7(32'h3ba66277),
	.w8(32'hbb148242),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb830e43),
	.w1(32'hbc41ea43),
	.w2(32'h3ad50ade),
	.w3(32'hbbe5ccfa),
	.w4(32'hbbcab2cf),
	.w5(32'hbc5b99ad),
	.w6(32'hbbe5c529),
	.w7(32'h3c607545),
	.w8(32'hbbfd5a75),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9571f3),
	.w1(32'hbc3f1607),
	.w2(32'h3cadb8bd),
	.w3(32'h3b6a030f),
	.w4(32'h3c530d7c),
	.w5(32'h3cd46c95),
	.w6(32'hbbcf1fec),
	.w7(32'h3c046904),
	.w8(32'hbc7dbc4c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf022ae),
	.w1(32'hbc695eec),
	.w2(32'hbc148faf),
	.w3(32'hbc8733ca),
	.w4(32'hbb4c2483),
	.w5(32'h3be20403),
	.w6(32'hbbe1f127),
	.w7(32'hbab32615),
	.w8(32'h3d919dc4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3ec21c),
	.w1(32'hbc59f318),
	.w2(32'h37f2ca66),
	.w3(32'hbc9bcc2b),
	.w4(32'h3bfbb0e4),
	.w5(32'h3a6e35e7),
	.w6(32'hbc80f924),
	.w7(32'h3b76e4c3),
	.w8(32'hbb2b4a5a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b6c51),
	.w1(32'h3c63f7dc),
	.w2(32'hbc815343),
	.w3(32'h3be21a4c),
	.w4(32'hbc185e46),
	.w5(32'h3ce6b030),
	.w6(32'h3bbf64bc),
	.w7(32'hbd3380ca),
	.w8(32'h3cb21e4a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f1a7c),
	.w1(32'h3cccda7e),
	.w2(32'hbc372303),
	.w3(32'h3b4df84e),
	.w4(32'hb8f5bc4b),
	.w5(32'h3b982fae),
	.w6(32'h3cbfa662),
	.w7(32'hbb6ed65e),
	.w8(32'hbc35aaf7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35efea),
	.w1(32'h3b998058),
	.w2(32'h3bd0ac73),
	.w3(32'h3c0e5d3c),
	.w4(32'hbca9d22a),
	.w5(32'h3c633935),
	.w6(32'h3ab7cf01),
	.w7(32'hba6ce884),
	.w8(32'h3cc22e07),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa19ff8),
	.w1(32'hbc1061cb),
	.w2(32'hbc94754d),
	.w3(32'hbcacd833),
	.w4(32'hbbf9ce31),
	.w5(32'hbb02e2a8),
	.w6(32'hbbdff638),
	.w7(32'hbbed2e2b),
	.w8(32'h3d3cb5ca),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d2ee7),
	.w1(32'h3bd875fc),
	.w2(32'h3b7510f5),
	.w3(32'h3c878a56),
	.w4(32'h3c5a97d2),
	.w5(32'hbc29436b),
	.w6(32'hbc7d5787),
	.w7(32'hbadd49d6),
	.w8(32'hbc2804b9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2bad7),
	.w1(32'hb95e8e48),
	.w2(32'h3b9ae632),
	.w3(32'hbbb9180d),
	.w4(32'h3c6a1c8c),
	.w5(32'h39a0b099),
	.w6(32'hbae3f942),
	.w7(32'h3cc55b87),
	.w8(32'hbcd86eea),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb391209),
	.w1(32'hbb9f8429),
	.w2(32'h3cc4a2c4),
	.w3(32'hbc0935d9),
	.w4(32'hbbf06d1d),
	.w5(32'h3cf1ad66),
	.w6(32'hbc5be453),
	.w7(32'hbbb5fd5d),
	.w8(32'h3c205ce0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca14cd9),
	.w1(32'h3bd54606),
	.w2(32'h3bd1708d),
	.w3(32'h3ab075cc),
	.w4(32'h3bc34d0a),
	.w5(32'h3cc79112),
	.w6(32'h3c64b88b),
	.w7(32'hbbcb36ff),
	.w8(32'h3ccdaabe),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c640e),
	.w1(32'hbb5c058a),
	.w2(32'h3ae7fec2),
	.w3(32'hbaeb0de7),
	.w4(32'hba41b0a4),
	.w5(32'h3bdf9f27),
	.w6(32'h39d05f43),
	.w7(32'h3a76c661),
	.w8(32'hbc009be4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77655d),
	.w1(32'h3b28d549),
	.w2(32'hbadb7bdf),
	.w3(32'h3a201e59),
	.w4(32'hbb62e80c),
	.w5(32'hbabb54a8),
	.w6(32'h3ac52a5f),
	.w7(32'h39ab8e4e),
	.w8(32'h3c9fc0a1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fa9e3),
	.w1(32'hbc6f176b),
	.w2(32'h3bd50264),
	.w3(32'hbc5ebaad),
	.w4(32'hbc5f96c1),
	.w5(32'h3cdc373c),
	.w6(32'hbc49d315),
	.w7(32'h3c3c3151),
	.w8(32'hbc7f9612),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd051f91),
	.w1(32'h3c7c3478),
	.w2(32'h3c085308),
	.w3(32'h3c7a49eb),
	.w4(32'h3b2ae041),
	.w5(32'hbc8c6d42),
	.w6(32'h3d0df2e5),
	.w7(32'hbc1436cf),
	.w8(32'hbc63a32d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca724ad),
	.w1(32'h3c3c3eff),
	.w2(32'hbd3907ff),
	.w3(32'h3bb52854),
	.w4(32'hbc9211e5),
	.w5(32'h3abc3748),
	.w6(32'hbc97a200),
	.w7(32'hbcc3759d),
	.w8(32'h3d375d5c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d0353),
	.w1(32'h3ce198ac),
	.w2(32'h3ca4448b),
	.w3(32'hbba2729d),
	.w4(32'hba5e66be),
	.w5(32'h3c322671),
	.w6(32'h3c3bc1da),
	.w7(32'h3be80254),
	.w8(32'hbd2b76b3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc494fb),
	.w1(32'h3c07cd7c),
	.w2(32'hbcb74858),
	.w3(32'hbabac4bf),
	.w4(32'hbcc1a873),
	.w5(32'hbc9e0f54),
	.w6(32'h3cc9734e),
	.w7(32'hbc321dc3),
	.w8(32'hbc4e7e23),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3d96c),
	.w1(32'hbcfa1008),
	.w2(32'hbb9e066b),
	.w3(32'hbcecb90f),
	.w4(32'hbc9858b6),
	.w5(32'hb97fba74),
	.w6(32'hbc4c12e5),
	.w7(32'hbacfc398),
	.w8(32'hbcea4b6b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc15a35),
	.w1(32'h3bea073c),
	.w2(32'h3b842b67),
	.w3(32'h3c93c0e6),
	.w4(32'h3cb2b457),
	.w5(32'hbad77866),
	.w6(32'h3c52707f),
	.w7(32'h3d112018),
	.w8(32'h3c464968),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1bbba),
	.w1(32'hbb85e600),
	.w2(32'h3bd41753),
	.w3(32'hbb163641),
	.w4(32'h3cb4a1e9),
	.w5(32'hbc0deab7),
	.w6(32'hbcb64d40),
	.w7(32'h3ca1eb60),
	.w8(32'hbcc85426),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19f761),
	.w1(32'hbc987b4c),
	.w2(32'hbadd037d),
	.w3(32'hbbb81e45),
	.w4(32'hbb92db91),
	.w5(32'h3baa83ff),
	.w6(32'hbc66aa9b),
	.w7(32'h3bc4ed1c),
	.w8(32'h3be8ece0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fb23c),
	.w1(32'hbb14e307),
	.w2(32'h3ad1c6ce),
	.w3(32'hbb5ce64c),
	.w4(32'h3b270b4a),
	.w5(32'h3bc4e6fe),
	.w6(32'hbadbcfa7),
	.w7(32'h3b9356d3),
	.w8(32'hbc07688c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c288383),
	.w1(32'hbbf89266),
	.w2(32'h3bfe367b),
	.w3(32'hbcaaad57),
	.w4(32'hbc12522d),
	.w5(32'h3c8c2c4b),
	.w6(32'hbbbecc68),
	.w7(32'h3be63443),
	.w8(32'hbc3003c8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6da9f),
	.w1(32'h3b7131da),
	.w2(32'hbc072043),
	.w3(32'hbc72d9a3),
	.w4(32'h3b3b43e3),
	.w5(32'h3cb28a83),
	.w6(32'h3ac4680c),
	.w7(32'hbbcc22f9),
	.w8(32'h3beb77f5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb713999),
	.w1(32'hba377c9f),
	.w2(32'hbca6a161),
	.w3(32'h3c1d9320),
	.w4(32'hbd0f5074),
	.w5(32'hbc2da8dc),
	.w6(32'h3c4643d8),
	.w7(32'hbc9f30f7),
	.w8(32'hb9b8b756),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc317ab),
	.w1(32'h3b81cfb2),
	.w2(32'hba9c82c8),
	.w3(32'h3ccd24ac),
	.w4(32'hbb197eda),
	.w5(32'h3b806907),
	.w6(32'h3c1adee2),
	.w7(32'hba8f5dea),
	.w8(32'hbbc98bf7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3892b9d1),
	.w1(32'h3b777278),
	.w2(32'h3c9a8637),
	.w3(32'hb9eca4e8),
	.w4(32'h3b89d342),
	.w5(32'hbbe5ca7a),
	.w6(32'h3b000ee0),
	.w7(32'h3c9c0f7d),
	.w8(32'hbd723359),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf45f06),
	.w1(32'h3bf68c52),
	.w2(32'hbd1c921e),
	.w3(32'h3bc76923),
	.w4(32'hbc0137ac),
	.w5(32'h3d3e8a34),
	.w6(32'h3c99f946),
	.w7(32'hbcdad0da),
	.w8(32'h3d8957ea),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4aabb),
	.w1(32'hbca09cb0),
	.w2(32'hbcc1ed55),
	.w3(32'hbc26784f),
	.w4(32'hbc84e023),
	.w5(32'hbb1ed2e9),
	.w6(32'h3b73d0af),
	.w7(32'hbc2e7e63),
	.w8(32'h3c9d5ec3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66cb00),
	.w1(32'hbb018ed5),
	.w2(32'h3c881293),
	.w3(32'h3b91579a),
	.w4(32'hbc13de0b),
	.w5(32'h3ca78345),
	.w6(32'h3ae6cbbc),
	.w7(32'hbc07551a),
	.w8(32'h3c8d3d62),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5c9c4),
	.w1(32'hbcab8c12),
	.w2(32'h3a1b256e),
	.w3(32'hbc4c6fa5),
	.w4(32'hbcd78aa3),
	.w5(32'h3b971999),
	.w6(32'hbce50e29),
	.w7(32'hbb8f8b0a),
	.w8(32'h3c061eb0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule