module layer_10_featuremap_28(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4a164),
	.w1(32'hbc6cbe37),
	.w2(32'h3b3dc748),
	.w3(32'h3be38a3e),
	.w4(32'hbb10864a),
	.w5(32'hbbafb987),
	.w6(32'h3baab67e),
	.w7(32'h3b4d297b),
	.w8(32'hba7650dc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee4490),
	.w1(32'h3c1e4f97),
	.w2(32'hbb96f899),
	.w3(32'hbc45121b),
	.w4(32'h3ab94cff),
	.w5(32'hba410beb),
	.w6(32'hbb71ffba),
	.w7(32'hbc071f46),
	.w8(32'hbab11e45),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f4993),
	.w1(32'hbabcc9c7),
	.w2(32'h3c643f62),
	.w3(32'h3c620299),
	.w4(32'h3aa1c2fe),
	.w5(32'h3a02267d),
	.w6(32'h3bd7d46b),
	.w7(32'hbb597a03),
	.w8(32'hbc7843df),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45283c),
	.w1(32'h3b47fd98),
	.w2(32'hba85de52),
	.w3(32'h3c41ad35),
	.w4(32'h3b5e1a36),
	.w5(32'h3a054128),
	.w6(32'hbc9c8269),
	.w7(32'hbcae5003),
	.w8(32'h3a53d3dc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd13f9),
	.w1(32'hbad5f2c8),
	.w2(32'hbba13154),
	.w3(32'hba46a36d),
	.w4(32'h3bd541e8),
	.w5(32'h3b4bfaf0),
	.w6(32'h3b3b1424),
	.w7(32'h3a1a6f25),
	.w8(32'h3b54d948),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59c03f),
	.w1(32'h39e1d138),
	.w2(32'hbab43a47),
	.w3(32'hbb5d73bc),
	.w4(32'h3b91bdda),
	.w5(32'hba6d9d48),
	.w6(32'h3ab8e13f),
	.w7(32'h3c499cb0),
	.w8(32'hbba0ee9e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ab84b),
	.w1(32'hbbf9e849),
	.w2(32'hbb4c8ffa),
	.w3(32'h3ae3f509),
	.w4(32'hbb8a0a34),
	.w5(32'h3baa2ade),
	.w6(32'h3a0e3e4e),
	.w7(32'hbac4a2f8),
	.w8(32'h3c3786e2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78d12e),
	.w1(32'hbba653c6),
	.w2(32'h3b01be52),
	.w3(32'hbb18de13),
	.w4(32'hbb3ef95b),
	.w5(32'h3b3dabb3),
	.w6(32'hbac8a6cb),
	.w7(32'h3a604052),
	.w8(32'hba5a4a6f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55f052),
	.w1(32'hbb44dd06),
	.w2(32'h3a9d8eee),
	.w3(32'hbac10817),
	.w4(32'hbabb408d),
	.w5(32'hbb2be022),
	.w6(32'h3b92eba5),
	.w7(32'h3a880b3e),
	.w8(32'h3b52e244),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a042b84),
	.w1(32'h3ab6acb7),
	.w2(32'h3a185068),
	.w3(32'h3a003395),
	.w4(32'h3c280825),
	.w5(32'hbabe3a68),
	.w6(32'h3a393836),
	.w7(32'h3bb3c859),
	.w8(32'h3b3ee5a2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00fca3),
	.w1(32'hba032889),
	.w2(32'h3c88b113),
	.w3(32'hbb63d525),
	.w4(32'hba4e8a07),
	.w5(32'h3c612e86),
	.w6(32'h3a039c09),
	.w7(32'h39b3b405),
	.w8(32'hbc10dd2e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9358f),
	.w1(32'h3bb1c643),
	.w2(32'h3bc336f2),
	.w3(32'h3c2ef74e),
	.w4(32'h3b0acbce),
	.w5(32'h3bb596e0),
	.w6(32'hbba88e15),
	.w7(32'hbc2d3929),
	.w8(32'h3c148de2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7691d),
	.w1(32'h3c2dd737),
	.w2(32'h3bdf206a),
	.w3(32'h3be44093),
	.w4(32'h3c173aff),
	.w5(32'hba4a1372),
	.w6(32'h3bc9c1ef),
	.w7(32'h3b8286a0),
	.w8(32'hbad8d5be),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff949f),
	.w1(32'hbb7bf62f),
	.w2(32'hbc0ddee0),
	.w3(32'h3aee7b36),
	.w4(32'h3b0aa524),
	.w5(32'h3b766ae5),
	.w6(32'h3a2c8f62),
	.w7(32'h3b6026dc),
	.w8(32'h3bea1fd6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91e54f),
	.w1(32'hbc7a675c),
	.w2(32'hbb41303f),
	.w3(32'hbaaef860),
	.w4(32'h3ba8d01a),
	.w5(32'hbb897cef),
	.w6(32'hbabd5062),
	.w7(32'hbc0ea87b),
	.w8(32'h3b3df0ea),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cf8e5),
	.w1(32'h3a92db26),
	.w2(32'hbab08a35),
	.w3(32'hba975cd7),
	.w4(32'hba507599),
	.w5(32'hbbd24545),
	.w6(32'h3b6a101d),
	.w7(32'h3aab4852),
	.w8(32'hbb2d78fe),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b3f32),
	.w1(32'h3ac25b3b),
	.w2(32'hb9b21654),
	.w3(32'hba512942),
	.w4(32'h381cf904),
	.w5(32'hbb71dff3),
	.w6(32'h3b04dffa),
	.w7(32'h3a9bbb61),
	.w8(32'hbb172fae),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a397386),
	.w1(32'h3b75a02f),
	.w2(32'h3ba357da),
	.w3(32'hbb6489ee),
	.w4(32'h3b3a0358),
	.w5(32'h391af55a),
	.w6(32'hbb6a4995),
	.w7(32'h3ba53d2e),
	.w8(32'hb9be5624),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc7d6e),
	.w1(32'h3c072597),
	.w2(32'h3c34c453),
	.w3(32'h3b746489),
	.w4(32'h3b91269f),
	.w5(32'hbac4b328),
	.w6(32'hbad8c70c),
	.w7(32'hbbb2df65),
	.w8(32'hb92741cc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95156a),
	.w1(32'hbc0f4457),
	.w2(32'hba8558dc),
	.w3(32'h3b1f1925),
	.w4(32'h3af199d2),
	.w5(32'h3a7934e0),
	.w6(32'hbbbfe312),
	.w7(32'hbb732064),
	.w8(32'hba998eb9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc3ab7),
	.w1(32'h3b1e0872),
	.w2(32'hbb02950d),
	.w3(32'h3bbdaf34),
	.w4(32'h3b909953),
	.w5(32'hbc447588),
	.w6(32'h3b6b18fc),
	.w7(32'h3bdbadea),
	.w8(32'hbbf5434e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d13e6),
	.w1(32'h3c76abe5),
	.w2(32'h3b20f307),
	.w3(32'hb93dc5a0),
	.w4(32'h3c940c97),
	.w5(32'h3b5a8321),
	.w6(32'hbc80169b),
	.w7(32'hbb7903b1),
	.w8(32'h3bc186b7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd173e3),
	.w1(32'hb9c0b856),
	.w2(32'h3aa4ecf1),
	.w3(32'h3c2b0ce3),
	.w4(32'h3bd0d56e),
	.w5(32'h3b8b57a4),
	.w6(32'hbb0b41a0),
	.w7(32'hbb322759),
	.w8(32'h3b96ba76),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e95c8),
	.w1(32'hb8c67578),
	.w2(32'h3b5e5280),
	.w3(32'h36ea0d54),
	.w4(32'h3a6ac7d6),
	.w5(32'hbb3fda33),
	.w6(32'hbb1b0e31),
	.w7(32'hbade350e),
	.w8(32'hbab7d300),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dfe9f),
	.w1(32'hbc003724),
	.w2(32'hbb0d05c1),
	.w3(32'hbba104ee),
	.w4(32'hbc899f31),
	.w5(32'hbc46a742),
	.w6(32'h3aa30cd1),
	.w7(32'hbc462acc),
	.w8(32'hbc941e0d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22f79a),
	.w1(32'h3c5e4055),
	.w2(32'hbb5a09e2),
	.w3(32'hbc1d1e33),
	.w4(32'h391defb2),
	.w5(32'hbbac04ab),
	.w6(32'hbc20ac62),
	.w7(32'hbbf0c9f1),
	.w8(32'hbb27cd07),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9403a9),
	.w1(32'h390ec8bd),
	.w2(32'hba2bb113),
	.w3(32'hbb6c1da6),
	.w4(32'hbaea3317),
	.w5(32'hb8ffdb8b),
	.w6(32'h3b24ff17),
	.w7(32'h3bbd0c98),
	.w8(32'hba6f9dd2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e22f8),
	.w1(32'h3bd352dd),
	.w2(32'h3b809cf8),
	.w3(32'h3b4e5c25),
	.w4(32'h3ba78959),
	.w5(32'h3ad76679),
	.w6(32'h3c34a1a1),
	.w7(32'h3c78aa35),
	.w8(32'h3c123f5a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c268ad0),
	.w1(32'hbac27220),
	.w2(32'hbb707986),
	.w3(32'h3c078165),
	.w4(32'h3970dc2c),
	.w5(32'h3be881a2),
	.w6(32'h3bb9b518),
	.w7(32'h3a1583aa),
	.w8(32'hbc01f6e0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f6926),
	.w1(32'hbc23063c),
	.w2(32'hbb8b8f8f),
	.w3(32'h3a7b08d9),
	.w4(32'hbb4b1c31),
	.w5(32'hbbce756b),
	.w6(32'hbaba15c1),
	.w7(32'h3bc64f16),
	.w8(32'hbb4291d9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75a2a9),
	.w1(32'h3bb50646),
	.w2(32'hba74fe71),
	.w3(32'h3b487f2f),
	.w4(32'h3be07ed6),
	.w5(32'h3b6632d1),
	.w6(32'hbb123aa6),
	.w7(32'h3a84ac8f),
	.w8(32'h39cffd31),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b61cf),
	.w1(32'hbc0be62d),
	.w2(32'hbba86d53),
	.w3(32'h3b62f9b0),
	.w4(32'hbb843ecd),
	.w5(32'h3be6f17e),
	.w6(32'h3c0d3c13),
	.w7(32'h3ba5d96f),
	.w8(32'h3cacc6fd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d02c5),
	.w1(32'hbbcd5efc),
	.w2(32'h3ab3de27),
	.w3(32'hbab459fc),
	.w4(32'hbbcdc4a7),
	.w5(32'hba799f58),
	.w6(32'h3ccef100),
	.w7(32'h3c6b1e0a),
	.w8(32'h39140be9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e71de),
	.w1(32'hbbb21a12),
	.w2(32'hbc373844),
	.w3(32'hbbd20ef0),
	.w4(32'hbbab57d5),
	.w5(32'hbc1ad111),
	.w6(32'hbbc9b0e2),
	.w7(32'hbb9d0a7d),
	.w8(32'hbc8798bf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c077d56),
	.w1(32'h3bb337f2),
	.w2(32'h3aaeae39),
	.w3(32'hbc1f7b7c),
	.w4(32'hbb98d1d6),
	.w5(32'h3a67c224),
	.w6(32'hbc1f0b4f),
	.w7(32'h3ad6c389),
	.w8(32'h3bc6b777),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0def7f),
	.w1(32'hbb18a0ec),
	.w2(32'h3c20579f),
	.w3(32'h3a1f8891),
	.w4(32'hbada0519),
	.w5(32'h3c36516c),
	.w6(32'h3b772bf2),
	.w7(32'h3a8ad2fe),
	.w8(32'h3c34a9c5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b08b5),
	.w1(32'hbc75f97e),
	.w2(32'h3c602433),
	.w3(32'hbc92a459),
	.w4(32'hbcd6f81b),
	.w5(32'hbc1ebc53),
	.w6(32'hbbd096b3),
	.w7(32'hbc4e23eb),
	.w8(32'hbb3d9a96),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c6f33),
	.w1(32'hbbc0ed54),
	.w2(32'hbc36ab44),
	.w3(32'hbb30e86d),
	.w4(32'hbab2e3bd),
	.w5(32'h3b2c4329),
	.w6(32'hb92cde9a),
	.w7(32'h3b7356af),
	.w8(32'h3c5b8c43),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30b312),
	.w1(32'hbbc58da2),
	.w2(32'hbb0c2313),
	.w3(32'h3b9e7f03),
	.w4(32'h3b8e7ecc),
	.w5(32'hbbd82af7),
	.w6(32'h3c62acc3),
	.w7(32'h3c999240),
	.w8(32'h3be4ca9e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c500391),
	.w1(32'h3cbeac3b),
	.w2(32'hbb5309f0),
	.w3(32'hbbbcc098),
	.w4(32'h3c4d9eb7),
	.w5(32'hbb9c27b1),
	.w6(32'hbc6e9589),
	.w7(32'hb930c015),
	.w8(32'hbbbd1116),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04fc49),
	.w1(32'hbb645537),
	.w2(32'h3a34cbe8),
	.w3(32'hbc148f87),
	.w4(32'hbb96f726),
	.w5(32'hbbdd9bb8),
	.w6(32'hbc1178f1),
	.w7(32'hbb799b4a),
	.w8(32'hbb5f5e7d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b467165),
	.w1(32'h3bdd1d8a),
	.w2(32'hbb71bfe2),
	.w3(32'hbb213619),
	.w4(32'h3be4bc60),
	.w5(32'hbbceb45a),
	.w6(32'hbb2746fe),
	.w7(32'h3c043c25),
	.w8(32'h3b8b6881),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc354e42),
	.w1(32'hbc80b333),
	.w2(32'h3afea06c),
	.w3(32'hbbac73da),
	.w4(32'hbc24e578),
	.w5(32'h3bb758be),
	.w6(32'h3b212660),
	.w7(32'h39227dbb),
	.w8(32'h3bf6d377),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7c450),
	.w1(32'h3b9ac138),
	.w2(32'h3b2d7dca),
	.w3(32'h3c04f82d),
	.w4(32'h3bedaad1),
	.w5(32'h3bec2fcd),
	.w6(32'h3c074ae8),
	.w7(32'h3c0496cf),
	.w8(32'hbb71576c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23f77e),
	.w1(32'h3bb84c9b),
	.w2(32'hbbcef13f),
	.w3(32'h3b6fffd1),
	.w4(32'h3c3f1fb6),
	.w5(32'h3842e4c1),
	.w6(32'hbc240ba5),
	.w7(32'h3b5bc156),
	.w8(32'hbc221d9c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd5401),
	.w1(32'h3ac0af83),
	.w2(32'h3bb2ead9),
	.w3(32'hbbcf4285),
	.w4(32'h3a7dc7ad),
	.w5(32'h3c0267ad),
	.w6(32'hbb9f5084),
	.w7(32'hbbaf6ba2),
	.w8(32'h3b1db131),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8dd7f),
	.w1(32'hbc18b37d),
	.w2(32'h39add0e4),
	.w3(32'h3b88b696),
	.w4(32'hbbeff16e),
	.w5(32'h3ae1963c),
	.w6(32'h3b93614c),
	.w7(32'hbac5bd0c),
	.w8(32'hbbafc9f6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b752dda),
	.w1(32'h3c3d4bf2),
	.w2(32'h3c5d6b18),
	.w3(32'h3b888451),
	.w4(32'h3b909e8f),
	.w5(32'h3c7eac8c),
	.w6(32'hbbe47dac),
	.w7(32'h38e05d3f),
	.w8(32'h3c34a350),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0a0f8),
	.w1(32'hba03f79e),
	.w2(32'h3b74ce22),
	.w3(32'h3aaf2b67),
	.w4(32'h3ab203d9),
	.w5(32'hbba8df50),
	.w6(32'h3b45c6df),
	.w7(32'h3b92504e),
	.w8(32'hbc2ff34c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c4aae),
	.w1(32'h3ca7831a),
	.w2(32'hbb7d1d64),
	.w3(32'hbbab77ad),
	.w4(32'h3b80788e),
	.w5(32'hbbb781f7),
	.w6(32'hbc525e16),
	.w7(32'hbb29218b),
	.w8(32'hbb7112b3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaceb8b),
	.w1(32'hbbf39bde),
	.w2(32'hbc65f323),
	.w3(32'hbb9f6db1),
	.w4(32'h3b8e4734),
	.w5(32'hbc0fc108),
	.w6(32'h3b529ede),
	.w7(32'h3adbe0da),
	.w8(32'hbbefde5b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab74437),
	.w1(32'h3c1cd4fe),
	.w2(32'hbb57de21),
	.w3(32'hbba5ce0a),
	.w4(32'h3bb6d23e),
	.w5(32'hbba85c90),
	.w6(32'hbbdb1969),
	.w7(32'hbbf99f46),
	.w8(32'h3c110843),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7bf25),
	.w1(32'hbb3b0534),
	.w2(32'hbb4a8121),
	.w3(32'h3c2e2e65),
	.w4(32'hbb124855),
	.w5(32'h3b6da94f),
	.w6(32'h3c54a62a),
	.w7(32'hbac0a023),
	.w8(32'h3a8a1baf),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ec639),
	.w1(32'hbafb8726),
	.w2(32'h3cde471e),
	.w3(32'h3c3e6c06),
	.w4(32'h3c1a44c9),
	.w5(32'h3c17292f),
	.w6(32'h3c2d4063),
	.w7(32'h3c96b58a),
	.w8(32'hbbde7215),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf62565),
	.w1(32'h3ca7944c),
	.w2(32'hbb02e97b),
	.w3(32'h3c8e45c9),
	.w4(32'h3cef8076),
	.w5(32'hbbe17354),
	.w6(32'hbc2d5107),
	.w7(32'h3bf1be41),
	.w8(32'hbbf572d7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b280f04),
	.w1(32'h3b7f5f3a),
	.w2(32'h3c46e98a),
	.w3(32'hbb9417e8),
	.w4(32'hba02781f),
	.w5(32'h3ca9362e),
	.w6(32'hbbb30ff7),
	.w7(32'hbb3c9c72),
	.w8(32'h3c8646e9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8317af),
	.w1(32'hbbdd7875),
	.w2(32'hba56b5e7),
	.w3(32'h3bd543e6),
	.w4(32'hbb8f52c0),
	.w5(32'hbac8654a),
	.w6(32'h3c0bde19),
	.w7(32'h3c03f503),
	.w8(32'hbbaa28c3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81852a),
	.w1(32'h3afafbdd),
	.w2(32'hbae2a5a8),
	.w3(32'hbbb28211),
	.w4(32'hbb388675),
	.w5(32'hbab55e97),
	.w6(32'hbc026163),
	.w7(32'hba3c640a),
	.w8(32'h393fce43),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc58018),
	.w1(32'h3afae013),
	.w2(32'h3b25525d),
	.w3(32'hbba299f9),
	.w4(32'h3ab37e47),
	.w5(32'h3ac5d5e6),
	.w6(32'hbb7daa83),
	.w7(32'h3b7cd221),
	.w8(32'h3ba46dfe),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b181757),
	.w1(32'h3c030794),
	.w2(32'h3b91a860),
	.w3(32'hbb27b2ed),
	.w4(32'hba6957cd),
	.w5(32'h3a2a7777),
	.w6(32'h3b7cc48a),
	.w7(32'h3bbf9cb6),
	.w8(32'hbc24f66b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fade5),
	.w1(32'h3c852706),
	.w2(32'hbb6f58ba),
	.w3(32'h3c2abb71),
	.w4(32'h3c1ec6da),
	.w5(32'h3b115061),
	.w6(32'hbb105416),
	.w7(32'hbc063276),
	.w8(32'h3b8ea98c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39874400),
	.w1(32'hba13b796),
	.w2(32'hbc037ad0),
	.w3(32'h3b43e6e3),
	.w4(32'hba2d7755),
	.w5(32'hbc3e0376),
	.w6(32'h3c0e9d2e),
	.w7(32'h3c35cc08),
	.w8(32'hbbe3d970),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2a09d),
	.w1(32'hbafe1e94),
	.w2(32'hbb2086a8),
	.w3(32'hbc6ca558),
	.w4(32'hbbaf55e8),
	.w5(32'hbbcb6f90),
	.w6(32'hbc792266),
	.w7(32'hbbcc91c7),
	.w8(32'hbbd8a7fe),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2ce35),
	.w1(32'h3a97743f),
	.w2(32'h3b16e8f3),
	.w3(32'h3b7b0407),
	.w4(32'h3b51fcf9),
	.w5(32'h3bfd1134),
	.w6(32'h3b0d1a0a),
	.w7(32'h3b776a93),
	.w8(32'h3a90dc4f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b20a6),
	.w1(32'h3b1b5f04),
	.w2(32'h3a3871c5),
	.w3(32'h39353777),
	.w4(32'h3a683995),
	.w5(32'h3aedc293),
	.w6(32'h3acfb36a),
	.w7(32'h3b649380),
	.w8(32'hb9f24735),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0ab94),
	.w1(32'h3bc29159),
	.w2(32'h3b81399e),
	.w3(32'h3bc1b8a2),
	.w4(32'h3bcaa243),
	.w5(32'h3c076f1c),
	.w6(32'h3b3e37d6),
	.w7(32'h3b898ed1),
	.w8(32'h3c0770a1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8d041),
	.w1(32'h3bf30abb),
	.w2(32'h3c0611a8),
	.w3(32'h3a03398a),
	.w4(32'h3b312f48),
	.w5(32'hbac090b0),
	.w6(32'h3c752482),
	.w7(32'h3c5a5f5e),
	.w8(32'h3c1eb544),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0693c3),
	.w1(32'hbafa7818),
	.w2(32'h3b851fed),
	.w3(32'hbb5cf16d),
	.w4(32'h3bf09603),
	.w5(32'h3c708a38),
	.w6(32'h3aaf5727),
	.w7(32'h3baa853a),
	.w8(32'hbade2d5e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb3298),
	.w1(32'h398d03a9),
	.w2(32'h3b5b94c3),
	.w3(32'h3b5f40af),
	.w4(32'hba79f4d5),
	.w5(32'hb816153e),
	.w6(32'h3b0ade38),
	.w7(32'h3acf7bcf),
	.w8(32'hbae87cc9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70a3c4),
	.w1(32'h3a9c6890),
	.w2(32'hbbfee57e),
	.w3(32'h3c589f23),
	.w4(32'h3b7dd2e7),
	.w5(32'hbc183735),
	.w6(32'h3c1337ab),
	.w7(32'h3b3dc657),
	.w8(32'hbc1680dc),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af549bc),
	.w1(32'h3bd911a9),
	.w2(32'h3b9a8144),
	.w3(32'hbb6ed49b),
	.w4(32'h3ae85a01),
	.w5(32'h3bda4cfe),
	.w6(32'hbad009be),
	.w7(32'hbb63c019),
	.w8(32'hbaa6c2c8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cf6eb),
	.w1(32'h394fd38f),
	.w2(32'hba884c6a),
	.w3(32'h3c130a7d),
	.w4(32'h3bba39b1),
	.w5(32'h3b364f08),
	.w6(32'h3a3a1e74),
	.w7(32'h3b762d41),
	.w8(32'hbb95fdb9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ce438),
	.w1(32'hbc33b447),
	.w2(32'h39f52dd8),
	.w3(32'hbbfae960),
	.w4(32'hbb6247f1),
	.w5(32'hbc8187a3),
	.w6(32'hbb249681),
	.w7(32'hbbadbbab),
	.w8(32'hbc402952),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4ec44),
	.w1(32'h3b52604f),
	.w2(32'h3b39ed41),
	.w3(32'hbc073bc0),
	.w4(32'hbb8b9454),
	.w5(32'h3b25ab5f),
	.w6(32'hbc40803d),
	.w7(32'hbc2999ab),
	.w8(32'h3ac3a639),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3dd33),
	.w1(32'hb9e78a96),
	.w2(32'hbba7cd8d),
	.w3(32'hbb7f0be9),
	.w4(32'hba52f071),
	.w5(32'hbbd7401f),
	.w6(32'hbb93f0c6),
	.w7(32'hba988ed5),
	.w8(32'hbb5799c4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b8678),
	.w1(32'hbb928c17),
	.w2(32'h3bad2c12),
	.w3(32'hbc5b1337),
	.w4(32'hbc37353f),
	.w5(32'h3ba7ab77),
	.w6(32'hbbfb4744),
	.w7(32'hbbc92fa9),
	.w8(32'h3bcfed98),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0017b7),
	.w1(32'h3c0afd53),
	.w2(32'h3bdee450),
	.w3(32'h3bc15608),
	.w4(32'h3a9cfc7b),
	.w5(32'h3ba2aeaf),
	.w6(32'hb8d5fdc2),
	.w7(32'hbb0b8cac),
	.w8(32'hbb2e660e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7c95),
	.w1(32'hbc029d4f),
	.w2(32'h3c81dc26),
	.w3(32'h3af79aee),
	.w4(32'h3a33fd66),
	.w5(32'h3be1a308),
	.w6(32'h3a86eef7),
	.w7(32'hba2165d4),
	.w8(32'hbb085862),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf3505),
	.w1(32'h3c1acaa5),
	.w2(32'hba790adb),
	.w3(32'h3cdbf5f7),
	.w4(32'h3ca521e0),
	.w5(32'h39b3c8f2),
	.w6(32'h3c35099f),
	.w7(32'h3c9f6cb8),
	.w8(32'h3939018d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb98c68),
	.w1(32'h3b356755),
	.w2(32'h3bd3d782),
	.w3(32'h3b9196c3),
	.w4(32'hbae4beef),
	.w5(32'hb9bc8abe),
	.w6(32'h3c2b7197),
	.w7(32'h3b40055a),
	.w8(32'h3b89de0d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6194c),
	.w1(32'h3b353bee),
	.w2(32'hbb150ade),
	.w3(32'h39a089b4),
	.w4(32'hba0c3e63),
	.w5(32'hbb820984),
	.w6(32'hba0473a5),
	.w7(32'h3b407653),
	.w8(32'hbb93c52e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5858f),
	.w1(32'h3b8a8436),
	.w2(32'h3c540075),
	.w3(32'h3b5f0641),
	.w4(32'h3bf33231),
	.w5(32'h3c0b35fd),
	.w6(32'hbaebdd16),
	.w7(32'h3a940111),
	.w8(32'hb8ffa763),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8c6a6),
	.w1(32'h3bde060a),
	.w2(32'hb936f34a),
	.w3(32'hbc1586fa),
	.w4(32'h3a7ab850),
	.w5(32'h3c2691ef),
	.w6(32'hbc600a3d),
	.w7(32'hbb8d653f),
	.w8(32'h3bfeb043),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3faccd),
	.w1(32'h3ad4de91),
	.w2(32'hbb4994e3),
	.w3(32'h3c48af2e),
	.w4(32'hbbf92571),
	.w5(32'hbbb364fd),
	.w6(32'h3c04ac88),
	.w7(32'hbb3d1e5d),
	.w8(32'hbbdf36b6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc514212),
	.w1(32'hbc950fb5),
	.w2(32'h3bad45fb),
	.w3(32'hbc54984a),
	.w4(32'hbc815a38),
	.w5(32'hbb171810),
	.w6(32'hbb2bb25e),
	.w7(32'hbbae9fbd),
	.w8(32'hbb2f6be6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7526c5),
	.w1(32'hbbf611b4),
	.w2(32'h391096f8),
	.w3(32'hbb788ac8),
	.w4(32'hbb3ec97a),
	.w5(32'hb9ce326d),
	.w6(32'hb9d5b6f5),
	.w7(32'h3a4244c7),
	.w8(32'hbb869ec7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1de9a),
	.w1(32'hbac30744),
	.w2(32'hbaca2310),
	.w3(32'h3b653337),
	.w4(32'hb8b0f3d3),
	.w5(32'hbb27f627),
	.w6(32'hb99a730a),
	.w7(32'h3b400efa),
	.w8(32'hbb3c0221),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0ccfe),
	.w1(32'h3aa889c8),
	.w2(32'hba6f236c),
	.w3(32'h3b168548),
	.w4(32'h3b7d385f),
	.w5(32'h3b5d39a4),
	.w6(32'h3b3aa14e),
	.w7(32'h3b9e5bd2),
	.w8(32'h3c103eb8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4089bc),
	.w1(32'hbc1eb802),
	.w2(32'hbb92d60c),
	.w3(32'h3be2ed60),
	.w4(32'hbb9cfbe8),
	.w5(32'h3a8d6286),
	.w6(32'h3b419bf9),
	.w7(32'hbb882052),
	.w8(32'hbbef4f9b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf08789),
	.w1(32'h3a653d0e),
	.w2(32'h3bbd7b4f),
	.w3(32'h3b9a629d),
	.w4(32'h3c0b37cb),
	.w5(32'h3c2c2717),
	.w6(32'hbbd07123),
	.w7(32'h3a96166c),
	.w8(32'h3bd236b1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66c655),
	.w1(32'h3aa6e3db),
	.w2(32'h3b5b47bd),
	.w3(32'h3bc5c398),
	.w4(32'h3be1dd42),
	.w5(32'h3bc7eee5),
	.w6(32'h3be9bd3a),
	.w7(32'h3bf2db96),
	.w8(32'h3bfdd51f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa12a55),
	.w1(32'h3b03dc9c),
	.w2(32'hbbad8ead),
	.w3(32'hbb561ac2),
	.w4(32'hbb46ea13),
	.w5(32'hbc1c672a),
	.w6(32'h3ace5981),
	.w7(32'hba87876c),
	.w8(32'hba8ff964),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4d2c2),
	.w1(32'hbc028d95),
	.w2(32'hbbe85725),
	.w3(32'hbbb9f91e),
	.w4(32'hbba542d5),
	.w5(32'hbb361e50),
	.w6(32'h39a4eb01),
	.w7(32'hbae00b66),
	.w8(32'hbb90d14e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cd2d4),
	.w1(32'h3a3a712c),
	.w2(32'h39fa8faf),
	.w3(32'hbba3055e),
	.w4(32'h3abdb0c3),
	.w5(32'h3b00589e),
	.w6(32'hbc0a9d9e),
	.w7(32'hbb620bfd),
	.w8(32'h3c0bc319),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803c89),
	.w1(32'hbc463f20),
	.w2(32'hbbe89eb1),
	.w3(32'h3a7de179),
	.w4(32'hbb9bada2),
	.w5(32'hbc32f4b1),
	.w6(32'h3c1a6532),
	.w7(32'h3b2f7b1f),
	.w8(32'h3b105cfe),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc758bd1),
	.w1(32'hbbd55126),
	.w2(32'hbbaf12c6),
	.w3(32'hbc4c8691),
	.w4(32'hbc16e2bd),
	.w5(32'hbc377bbe),
	.w6(32'h3c498f58),
	.w7(32'h3c4e9eb6),
	.w8(32'hbb8b6fc9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1013c),
	.w1(32'h3bcff15c),
	.w2(32'hbb9ff491),
	.w3(32'hbb5bfa61),
	.w4(32'h3b90684a),
	.w5(32'h39b98f08),
	.w6(32'hbc11f47d),
	.w7(32'h3a360b8a),
	.w8(32'hba841df3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffca69),
	.w1(32'hbc1f4742),
	.w2(32'h3b22b402),
	.w3(32'h3b45e404),
	.w4(32'hbc19251e),
	.w5(32'h3b0a0bc6),
	.w6(32'h3bb9bb59),
	.w7(32'hbbbc823f),
	.w8(32'hbc0569dd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be92e3b),
	.w1(32'h3be680a7),
	.w2(32'h3bfe819f),
	.w3(32'hbc550c00),
	.w4(32'hbc0cb9a0),
	.w5(32'h3a094e73),
	.w6(32'hbc01276a),
	.w7(32'h3ae0fc93),
	.w8(32'h3c46e808),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe89167),
	.w1(32'hbbcf22fa),
	.w2(32'hbabe24b2),
	.w3(32'hbb35dd78),
	.w4(32'hbc115f78),
	.w5(32'hbbc6ea5c),
	.w6(32'hbb797784),
	.w7(32'hbc16393a),
	.w8(32'hbc6a67ec),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc860668),
	.w1(32'hbca9d5ac),
	.w2(32'hbb57e73d),
	.w3(32'hbc010646),
	.w4(32'hbc3c6b1f),
	.w5(32'hbb7bee7b),
	.w6(32'hbbc79d53),
	.w7(32'hbb5eb89c),
	.w8(32'hbbf3b2e2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cbf44),
	.w1(32'hbc1a14d0),
	.w2(32'hbb67d971),
	.w3(32'hbc30afc2),
	.w4(32'hbc897366),
	.w5(32'hbc21717e),
	.w6(32'hbbd35963),
	.w7(32'hbc62973e),
	.w8(32'hbc256a84),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5b801),
	.w1(32'h3be1f2f9),
	.w2(32'h3c34b90a),
	.w3(32'hbbd92c55),
	.w4(32'hbb04ac7f),
	.w5(32'hbba088e6),
	.w6(32'hbbbfbd27),
	.w7(32'hb7ce36c2),
	.w8(32'h3b4c538b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a071ee8),
	.w1(32'h3be424df),
	.w2(32'h3a77cf2d),
	.w3(32'h3bbaae54),
	.w4(32'h3c1782da),
	.w5(32'h3b868e72),
	.w6(32'h3bd90106),
	.w7(32'h3c27e02e),
	.w8(32'hbb9e1f99),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab27d34),
	.w1(32'hbbba4d39),
	.w2(32'h3c30ceaa),
	.w3(32'h3b3fc3d1),
	.w4(32'hbb88bd83),
	.w5(32'hbc693aaf),
	.w6(32'h3a8c57ff),
	.w7(32'hbc479a9d),
	.w8(32'hbcbe9c60),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c909904),
	.w1(32'h3c1bc9bf),
	.w2(32'h3b6b79f5),
	.w3(32'h3c28cd13),
	.w4(32'h3c2812cb),
	.w5(32'h3b94c425),
	.w6(32'hbadd0e10),
	.w7(32'h3baf3872),
	.w8(32'h3b68c866),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36e1a6),
	.w1(32'hb9d21c46),
	.w2(32'h3abf8af3),
	.w3(32'h3c21a4e5),
	.w4(32'h3b495a2a),
	.w5(32'h3c069654),
	.w6(32'h3b80fa16),
	.w7(32'h3b61dbf5),
	.w8(32'h3c7715db),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8c88e),
	.w1(32'hbb85308b),
	.w2(32'hbc1937c9),
	.w3(32'hbb8151ca),
	.w4(32'hbc00079b),
	.w5(32'h3b8b1f48),
	.w6(32'h3b7e7fa1),
	.w7(32'h3a158814),
	.w8(32'h3bec7480),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7971a2),
	.w1(32'h3b8fb5ee),
	.w2(32'h3b6fc434),
	.w3(32'hbbbe1c64),
	.w4(32'h3b1cd5cc),
	.w5(32'h3b5dca2f),
	.w6(32'hb9152365),
	.w7(32'h3baae628),
	.w8(32'hbba87570),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea334),
	.w1(32'hbab95a50),
	.w2(32'hbbbb53d5),
	.w3(32'h3c03928f),
	.w4(32'h3bd18f32),
	.w5(32'hbc303e58),
	.w6(32'hbad7141e),
	.w7(32'h3b79fc54),
	.w8(32'hbb8aa511),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc032a19),
	.w1(32'hbbe888be),
	.w2(32'hb9dfae08),
	.w3(32'hbbe9e9fd),
	.w4(32'hbc1601c3),
	.w5(32'hbabbe137),
	.w6(32'hbc103284),
	.w7(32'hb961af45),
	.w8(32'hbba1b1c4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78ef1f),
	.w1(32'h3b1fdb8d),
	.w2(32'h3b28a6b6),
	.w3(32'h3935718d),
	.w4(32'h3b141d71),
	.w5(32'hbbfa81a9),
	.w6(32'hbbe1367e),
	.w7(32'h3b7b4949),
	.w8(32'hbb83e32f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3aade8),
	.w1(32'hba9d3466),
	.w2(32'hbb9e0ef0),
	.w3(32'hbbfa5c5d),
	.w4(32'hba459d2b),
	.w5(32'h3c3a9a58),
	.w6(32'hbc5d4a14),
	.w7(32'hbc2743ab),
	.w8(32'h3bc96b3b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16d4e0),
	.w1(32'hbb8f2b3f),
	.w2(32'h3b2389bc),
	.w3(32'h3bd857f0),
	.w4(32'hbc0305b7),
	.w5(32'hbbcb321e),
	.w6(32'h3ca1c5b3),
	.w7(32'hbad702f8),
	.w8(32'h3af45171),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12c7bd),
	.w1(32'h3b5868ff),
	.w2(32'h3a29f75d),
	.w3(32'hbc20c669),
	.w4(32'hbc51df63),
	.w5(32'h3b2c46b6),
	.w6(32'hbb948ded),
	.w7(32'hbb7b5558),
	.w8(32'h3b80379a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba699ac3),
	.w1(32'h3bc179e8),
	.w2(32'hb82aa4c7),
	.w3(32'hba8ad741),
	.w4(32'h3a2d330b),
	.w5(32'h3ad7e4cd),
	.w6(32'h3b893af9),
	.w7(32'h3b73d864),
	.w8(32'hbb13ff7a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1474f4),
	.w1(32'hbb188d1e),
	.w2(32'h3b1a73ec),
	.w3(32'h3af30dc5),
	.w4(32'h3b933b30),
	.w5(32'hbb75e31f),
	.w6(32'hbb0f0ee3),
	.w7(32'h38136420),
	.w8(32'h3b2bf2fc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace458c),
	.w1(32'h3b756576),
	.w2(32'hbb949951),
	.w3(32'hbb907112),
	.w4(32'hbb6cd7c0),
	.w5(32'hba1da59f),
	.w6(32'h3b1f09f2),
	.w7(32'h3b478afd),
	.w8(32'hbbbec194),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc193b72),
	.w1(32'hbbaf365b),
	.w2(32'h3a9d174d),
	.w3(32'hbb90e6da),
	.w4(32'h3ab84979),
	.w5(32'h3bf71954),
	.w6(32'h3bf80833),
	.w7(32'h3aa32146),
	.w8(32'h39adef6e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1fe47),
	.w1(32'hbc16f25c),
	.w2(32'hbbc42c81),
	.w3(32'hbb4fd88c),
	.w4(32'hbbc115ef),
	.w5(32'hbc22bae2),
	.w6(32'hb9986111),
	.w7(32'hbbb16b4d),
	.w8(32'hbc79c89c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98f0d5),
	.w1(32'h3b8a3619),
	.w2(32'h3b1ad8c8),
	.w3(32'hbc5749ae),
	.w4(32'hbc0d1e60),
	.w5(32'h3aa061e9),
	.w6(32'hbc3dbfc1),
	.w7(32'hbc87a03c),
	.w8(32'h3a3a42fb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eda28),
	.w1(32'h3bc82793),
	.w2(32'h3b327744),
	.w3(32'h3b5fd1df),
	.w4(32'h3b8d408c),
	.w5(32'h3b3a370e),
	.w6(32'hba02b771),
	.w7(32'h3abec4e8),
	.w8(32'h3b0fc6b8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae21403),
	.w1(32'hbbfe8ae3),
	.w2(32'h3b96ba5e),
	.w3(32'hbb074322),
	.w4(32'hbb5a8309),
	.w5(32'hbb545035),
	.w6(32'h3ad2e18d),
	.w7(32'h3a89a82b),
	.w8(32'hbcb7b908),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb470b2),
	.w1(32'h3c6b5c1d),
	.w2(32'h3ae9dd6c),
	.w3(32'h3cc09f54),
	.w4(32'h3caf6fb8),
	.w5(32'hbb7f956b),
	.w6(32'h392852f8),
	.w7(32'h3bae9ae0),
	.w8(32'hbbba1808),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c8bbd),
	.w1(32'h3bc6a931),
	.w2(32'h3bbbccba),
	.w3(32'h3b649fc2),
	.w4(32'h3b1c51f9),
	.w5(32'hbb0b7518),
	.w6(32'hbb22b1c3),
	.w7(32'hba1d2301),
	.w8(32'hbc645544),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56b5e1),
	.w1(32'h3c8005d0),
	.w2(32'h3b81d1cb),
	.w3(32'h3bc0f152),
	.w4(32'h3c4f7252),
	.w5(32'hbb61dfa9),
	.w6(32'hbbc07045),
	.w7(32'h3aa55e3c),
	.w8(32'hbb0c9761),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb331356),
	.w1(32'hbbda932a),
	.w2(32'hbab5be36),
	.w3(32'h3b273491),
	.w4(32'hbb090e67),
	.w5(32'hb982fba2),
	.w6(32'hbb0ad5e0),
	.w7(32'h3a82b6e8),
	.w8(32'h3acbb393),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc352201),
	.w1(32'hbc39f135),
	.w2(32'h3a8c9af9),
	.w3(32'hba7d0bbf),
	.w4(32'hbb0b9186),
	.w5(32'h3d1a7e3c),
	.w6(32'h3b9f0849),
	.w7(32'hba93728c),
	.w8(32'h3cc873f7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31ec04),
	.w1(32'hbc1a1dff),
	.w2(32'hba13b69d),
	.w3(32'h3ac6492f),
	.w4(32'hbb808727),
	.w5(32'h3b961994),
	.w6(32'h3c5ec799),
	.w7(32'hb8ae73c1),
	.w8(32'h3bfacac3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ba062),
	.w1(32'h3c1cd3b3),
	.w2(32'h3b4746b2),
	.w3(32'hbbca3335),
	.w4(32'hbbc18551),
	.w5(32'hbbf30680),
	.w6(32'h3b0cf7d6),
	.w7(32'hbae983aa),
	.w8(32'hbc7664c1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c2956),
	.w1(32'h3b4617b9),
	.w2(32'hb9845ac5),
	.w3(32'hbc47d5e0),
	.w4(32'h3b5600e4),
	.w5(32'hbc121309),
	.w6(32'hbcc4972a),
	.w7(32'hbc73aacc),
	.w8(32'hbc45be83),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb805a70),
	.w1(32'hbb8f2542),
	.w2(32'hbb7bd0d0),
	.w3(32'hbc075b37),
	.w4(32'hbc5f65bb),
	.w5(32'h3a3775c6),
	.w6(32'hbc44303d),
	.w7(32'hbbe7c8e6),
	.w8(32'h3bdbb803),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae52412),
	.w1(32'hbb862839),
	.w2(32'h3b04e499),
	.w3(32'hbb682747),
	.w4(32'h3c2c631b),
	.w5(32'h3ab6f558),
	.w6(32'h3b289083),
	.w7(32'h3bea36b4),
	.w8(32'h3ae59f9e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80aa91),
	.w1(32'h3bc0a293),
	.w2(32'h3895f85d),
	.w3(32'hba80ab36),
	.w4(32'h3baea658),
	.w5(32'hbba2a161),
	.w6(32'hbbcbaa27),
	.w7(32'h3b1144a9),
	.w8(32'hbb4eaad9),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b034c4a),
	.w1(32'h3bef3324),
	.w2(32'h3b3293b5),
	.w3(32'h389d37a5),
	.w4(32'h3bc70afc),
	.w5(32'hbb278e90),
	.w6(32'h3a39c99e),
	.w7(32'h3ba2e1f2),
	.w8(32'h3c09f152),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc068910),
	.w1(32'hbb8d9b95),
	.w2(32'h3b000c9a),
	.w3(32'hbc3869e9),
	.w4(32'hbc3833ec),
	.w5(32'h3c1f0bb6),
	.w6(32'h3b29f0a0),
	.w7(32'hba103e23),
	.w8(32'hba80909d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd916c5),
	.w1(32'hbc0466a3),
	.w2(32'h3b942eac),
	.w3(32'h3c8f9f16),
	.w4(32'h3b811a97),
	.w5(32'h3c029e0d),
	.w6(32'h3c0d5141),
	.w7(32'h3bf720c3),
	.w8(32'h3bd01c3d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af523fa),
	.w1(32'h3ba1cbf2),
	.w2(32'h3ac56a74),
	.w3(32'hba512556),
	.w4(32'hbb9cc5a6),
	.w5(32'h3ae0e250),
	.w6(32'hbb361c00),
	.w7(32'hbb8c1732),
	.w8(32'h3a69c05c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff4fc3),
	.w1(32'hbb9cae7d),
	.w2(32'hbac18a8c),
	.w3(32'hbb3c6eed),
	.w4(32'hbb9f90e8),
	.w5(32'hbc567e19),
	.w6(32'hbbacc522),
	.w7(32'hbbde91c7),
	.w8(32'hbc7f8a50),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43f527),
	.w1(32'hbb813de3),
	.w2(32'hbace5aae),
	.w3(32'hbc3b9eda),
	.w4(32'hbc3aafca),
	.w5(32'hbb357245),
	.w6(32'hbc2f64b3),
	.w7(32'hbc081701),
	.w8(32'hbbb92ee0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba249188),
	.w1(32'hb993b2ac),
	.w2(32'h3bc2b0cc),
	.w3(32'hbb4a99b2),
	.w4(32'hbb3ef365),
	.w5(32'h3b13d35a),
	.w6(32'hbbdc18ed),
	.w7(32'hbbce0b82),
	.w8(32'h3a8f4b0b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36dbb1),
	.w1(32'h3b8aab58),
	.w2(32'h3b88606c),
	.w3(32'h385ffc08),
	.w4(32'h3c18f13c),
	.w5(32'hbc0220a2),
	.w6(32'h3b9f1f46),
	.w7(32'h3c20c9e2),
	.w8(32'hbc04396c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf794),
	.w1(32'hbb3baf4b),
	.w2(32'hbb37b9cb),
	.w3(32'h3b2cd006),
	.w4(32'h3c3762d8),
	.w5(32'hb9eb617a),
	.w6(32'hbc1351b6),
	.w7(32'h3b4f7b50),
	.w8(32'h3be6728b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbfd05),
	.w1(32'h3bb0f315),
	.w2(32'hbb9eb9f9),
	.w3(32'hbc353842),
	.w4(32'hbbbecdfe),
	.w5(32'hbb6789ab),
	.w6(32'hba885494),
	.w7(32'hbaed2720),
	.w8(32'hbb94788f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b5ff8),
	.w1(32'h3b0638b0),
	.w2(32'hbb01dce4),
	.w3(32'h39d406c6),
	.w4(32'h3b3924d7),
	.w5(32'hbaec4383),
	.w6(32'hbb43cc0c),
	.w7(32'hb8ede11b),
	.w8(32'hbb253d9f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90081c),
	.w1(32'h3c0f6d02),
	.w2(32'h3ade61ab),
	.w3(32'h3bdf675e),
	.w4(32'h3c052099),
	.w5(32'h3bb10e69),
	.w6(32'h3c00ac27),
	.w7(32'h3bf137aa),
	.w8(32'hbb02773e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84cb36),
	.w1(32'hba8e7c8f),
	.w2(32'h3bea71bf),
	.w3(32'h3940341d),
	.w4(32'hbb83b510),
	.w5(32'h3b0c5993),
	.w6(32'hba2da19a),
	.w7(32'hbba316a8),
	.w8(32'hbb87c77e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04b010),
	.w1(32'hba721a2d),
	.w2(32'h3b4e7ce5),
	.w3(32'h3cab20f8),
	.w4(32'h3c414e9c),
	.w5(32'h3b63b076),
	.w6(32'h3bb5173b),
	.w7(32'h3c430a57),
	.w8(32'h3b078f89),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e3ca9),
	.w1(32'h3b063543),
	.w2(32'hbc71ada2),
	.w3(32'h3b679305),
	.w4(32'h3b952363),
	.w5(32'hbab40fde),
	.w6(32'h3b7f31bb),
	.w7(32'h3b580dee),
	.w8(32'hbb6403d0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc673048),
	.w1(32'hbc08c665),
	.w2(32'hbbd1f694),
	.w3(32'hbb6d9533),
	.w4(32'hbbec3721),
	.w5(32'h3b3491c3),
	.w6(32'hbb08c965),
	.w7(32'hbbe19527),
	.w8(32'h3b672a25),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc058810),
	.w1(32'hbb0f5fa7),
	.w2(32'h3add920d),
	.w3(32'hbc2a1270),
	.w4(32'hbc54d471),
	.w5(32'hb9f66190),
	.w6(32'h3adc5512),
	.w7(32'hbbda525b),
	.w8(32'hbb38b9b9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b862c09),
	.w1(32'h3be69836),
	.w2(32'h3c2069dc),
	.w3(32'hbab77f8a),
	.w4(32'h3b22ee3b),
	.w5(32'h3c1fa6ba),
	.w6(32'hbb2c41d6),
	.w7(32'hbaa416ac),
	.w8(32'h3bf0516b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b879b5e),
	.w1(32'h3bf4fb9e),
	.w2(32'h3baccdcd),
	.w3(32'h3c5bb26d),
	.w4(32'h3b83ea97),
	.w5(32'h3be25e46),
	.w6(32'h3c25442e),
	.w7(32'h3c18305a),
	.w8(32'h3c8bad46),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b899ae3),
	.w1(32'hbc97b7ac),
	.w2(32'hbb4fd179),
	.w3(32'h3c9a323f),
	.w4(32'hbaaad903),
	.w5(32'h3b672973),
	.w6(32'h3c68f830),
	.w7(32'h3c0ea3b0),
	.w8(32'hbb88112a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89e5d7),
	.w1(32'h3bb35242),
	.w2(32'h39d6e302),
	.w3(32'hbaef6a6b),
	.w4(32'h3b8fafd1),
	.w5(32'h3aadf848),
	.w6(32'h3a124b8d),
	.w7(32'hba070eb8),
	.w8(32'h3a092ef7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf00cd),
	.w1(32'h392cacac),
	.w2(32'hbab0703f),
	.w3(32'hba5ba9e1),
	.w4(32'h39d39d98),
	.w5(32'h3acebe6d),
	.w6(32'hbae116e5),
	.w7(32'hba13c84c),
	.w8(32'h3adbcdc8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fc426),
	.w1(32'h3a269196),
	.w2(32'hbbe44c33),
	.w3(32'hbc4e9484),
	.w4(32'h3c45d331),
	.w5(32'h3a37d90a),
	.w6(32'hbc585023),
	.w7(32'h3c6188c0),
	.w8(32'h3ca48dc4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ab05d),
	.w1(32'h3d480674),
	.w2(32'hbb8ae411),
	.w3(32'hbcd1d94d),
	.w4(32'h3d9547fd),
	.w5(32'hbac1b709),
	.w6(32'h3b3d1ad4),
	.w7(32'h3cab3f1f),
	.w8(32'hbb333359),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18c9cf),
	.w1(32'h3b1e218d),
	.w2(32'hbb1b87b5),
	.w3(32'h3b813451),
	.w4(32'h3b584374),
	.w5(32'hbc089ef1),
	.w6(32'h39fa4c2d),
	.w7(32'hbae64180),
	.w8(32'h3add47c2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3192e2),
	.w1(32'h3c9406bf),
	.w2(32'h3b93df5d),
	.w3(32'hbc59369e),
	.w4(32'h3c543b87),
	.w5(32'hbba91b38),
	.w6(32'hbc682611),
	.w7(32'h3c400f38),
	.w8(32'hb9a18b51),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c22c),
	.w1(32'h3a138ebf),
	.w2(32'hba5ea60f),
	.w3(32'hbc0bf251),
	.w4(32'hbb582cde),
	.w5(32'h3b0a0f2e),
	.w6(32'hbc5f2c42),
	.w7(32'hbc082d3b),
	.w8(32'h3ab25d0e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a4461),
	.w1(32'h3a486c68),
	.w2(32'h3bf6c6f8),
	.w3(32'hb958c1fd),
	.w4(32'h3b253927),
	.w5(32'h3bb26df0),
	.w6(32'hbbaf19b6),
	.w7(32'h3ad84b55),
	.w8(32'h3b23e124),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c45c0),
	.w1(32'hbc580699),
	.w2(32'hbb5d92f7),
	.w3(32'h3a463adf),
	.w4(32'hbc4e2d86),
	.w5(32'hbbae9bf1),
	.w6(32'hbb7ec489),
	.w7(32'hbcaefd0b),
	.w8(32'hba85b48d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b8dd1),
	.w1(32'h3a3e4ef1),
	.w2(32'hbaf487be),
	.w3(32'hba8af3a7),
	.w4(32'h3b488ba5),
	.w5(32'hbcbdc35b),
	.w6(32'hbb0b14f2),
	.w7(32'h3b909487),
	.w8(32'hbc0814be),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e19dd),
	.w1(32'hbc1ff245),
	.w2(32'h3b1e04b3),
	.w3(32'h3cd464f0),
	.w4(32'hbb5afbc7),
	.w5(32'h3c45afbd),
	.w6(32'h3c63b52b),
	.w7(32'hbc1403af),
	.w8(32'h3c27183f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae20393),
	.w1(32'h3bd2bef0),
	.w2(32'h3a93b9f2),
	.w3(32'h3bd48906),
	.w4(32'h3c18469d),
	.w5(32'h3c11edf2),
	.w6(32'h3a73b754),
	.w7(32'h3b8d4682),
	.w8(32'h3c8d75eb),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78b0d3),
	.w1(32'h3c7919c7),
	.w2(32'h3ad0f048),
	.w3(32'hbcacaeb6),
	.w4(32'hbbb8baa4),
	.w5(32'h3940db82),
	.w6(32'hbb73c170),
	.w7(32'hbc430550),
	.w8(32'h39a3d53d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf17b43),
	.w1(32'hbba80e14),
	.w2(32'h391bd2fb),
	.w3(32'h3cac8f7d),
	.w4(32'hbc07ad66),
	.w5(32'h3a9fc732),
	.w6(32'h3c98d491),
	.w7(32'hbc040ee1),
	.w8(32'hbafdb60e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc428e30),
	.w1(32'hbbbaaea0),
	.w2(32'h3c19ab2e),
	.w3(32'hbb9dd1e0),
	.w4(32'h3b9797dc),
	.w5(32'h3c368d87),
	.w6(32'hbc0bc7a5),
	.w7(32'h3af0965f),
	.w8(32'h3b06279d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b801d36),
	.w1(32'hbc2ae12f),
	.w2(32'hbb37c38e),
	.w3(32'h3b670723),
	.w4(32'hbd1a4578),
	.w5(32'hbc38b98f),
	.w6(32'h3b949d48),
	.w7(32'hbd186468),
	.w8(32'hb94663c9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc761373),
	.w1(32'h3bf7d95f),
	.w2(32'hbb831d89),
	.w3(32'hbbda5720),
	.w4(32'h3c81d007),
	.w5(32'hbc0c5bc9),
	.w6(32'h3b65eda4),
	.w7(32'h3c0b89b2),
	.w8(32'hbae728bd),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0d59b),
	.w1(32'hba0f094b),
	.w2(32'h3c74c4b6),
	.w3(32'hbc2013f6),
	.w4(32'h3b3562f1),
	.w5(32'h3d0bde07),
	.w6(32'hbb5e2365),
	.w7(32'h3b41c501),
	.w8(32'h3ce403ad),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf16f64),
	.w1(32'h3cd52aba),
	.w2(32'h3c4d7b1a),
	.w3(32'hbcd677ce),
	.w4(32'h3d618bf1),
	.w5(32'h383d42c6),
	.w6(32'hbc634c1f),
	.w7(32'h3c954a59),
	.w8(32'h3c303ab6),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36a2fd),
	.w1(32'h3c8f8f06),
	.w2(32'h3c072563),
	.w3(32'hbcdc296a),
	.w4(32'h3d176e85),
	.w5(32'h3b8b83bc),
	.w6(32'hbcf1076b),
	.w7(32'h3ce48a59),
	.w8(32'hbbb05411),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e1aea),
	.w1(32'hbb684e9f),
	.w2(32'h3ae03cd1),
	.w3(32'h3c2d1e9f),
	.w4(32'hbb595dad),
	.w5(32'h3bda2788),
	.w6(32'h3bbc52a3),
	.w7(32'hbb6ba79b),
	.w8(32'h3b04a7d5),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc375bb9),
	.w1(32'hbc89286e),
	.w2(32'h3ab3c114),
	.w3(32'hbc9f5fac),
	.w4(32'hbcb3d2fb),
	.w5(32'h3b2d0acd),
	.w6(32'hbcb401e3),
	.w7(32'hbcd1b4bb),
	.w8(32'h3b8171d1),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab00e55),
	.w1(32'h39b301d5),
	.w2(32'hbb526d55),
	.w3(32'hbaa26be7),
	.w4(32'hbb8a7de5),
	.w5(32'hbc057d0f),
	.w6(32'h3b75424c),
	.w7(32'h3a2277e6),
	.w8(32'h3c1cf16e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a016ae6),
	.w1(32'h3c855599),
	.w2(32'h3bb13b7e),
	.w3(32'h3b286d18),
	.w4(32'h3c9c02f0),
	.w5(32'hbc875aa2),
	.w6(32'hbb73682d),
	.w7(32'h3c46f3c1),
	.w8(32'h3a2cf9e8),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb23c62),
	.w1(32'hbc0f5dde),
	.w2(32'hba9e9ff1),
	.w3(32'hbbe5cfe1),
	.w4(32'h3ad9fdc5),
	.w5(32'hbc2c343a),
	.w6(32'hbc34d50f),
	.w7(32'hbc2f4492),
	.w8(32'h3b689865),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b091d46),
	.w1(32'hbc90e5e1),
	.w2(32'hb9d7d212),
	.w3(32'hb839c289),
	.w4(32'hbbd97a23),
	.w5(32'hbbf45d66),
	.w6(32'h3ac120ae),
	.w7(32'h3a536de9),
	.w8(32'hbbf655b2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c721b1e),
	.w1(32'hbb8b6be5),
	.w2(32'h3a07e335),
	.w3(32'hbbd0411d),
	.w4(32'h398b892c),
	.w5(32'h3b70a10a),
	.w6(32'hbc9bf070),
	.w7(32'hbb9a3fe0),
	.w8(32'h3bc2ae96),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ed827),
	.w1(32'hbbad3474),
	.w2(32'hbc240e76),
	.w3(32'h3b35e897),
	.w4(32'hbc04edc6),
	.w5(32'hbb5883d0),
	.w6(32'hbac0e899),
	.w7(32'hbc1d8cec),
	.w8(32'h3c27e0e1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13349e),
	.w1(32'h3d0ada2e),
	.w2(32'h3c45aa26),
	.w3(32'hbc84e18d),
	.w4(32'h3d142f97),
	.w5(32'h3ba6113e),
	.w6(32'hbb5ee847),
	.w7(32'h3b19b657),
	.w8(32'hbb050192),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d3ddb),
	.w1(32'hb952ebf1),
	.w2(32'hba2c20ce),
	.w3(32'hbc937f59),
	.w4(32'h3a29a9b4),
	.w5(32'h3b2be4ce),
	.w6(32'hbc6223ad),
	.w7(32'h3b945db9),
	.w8(32'h3bfb24a8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39241040),
	.w1(32'hba50a027),
	.w2(32'h3b21e75e),
	.w3(32'h39903dbe),
	.w4(32'hbc80e56b),
	.w5(32'hbb3d9a18),
	.w6(32'hbb045cea),
	.w7(32'hbc248c7d),
	.w8(32'hbaeae5fa),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58abd6),
	.w1(32'hbb9ae903),
	.w2(32'h392140ff),
	.w3(32'h3c44e4e9),
	.w4(32'hbc005dfa),
	.w5(32'hbc0f19af),
	.w6(32'h3c2129a4),
	.w7(32'hbb1e7031),
	.w8(32'hbc48ed17),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac94ff),
	.w1(32'h3c566743),
	.w2(32'h3b3a20b2),
	.w3(32'hbba8cc8c),
	.w4(32'h3c610bb0),
	.w5(32'h3aa99e68),
	.w6(32'hbbee2a6e),
	.w7(32'h3c6ae607),
	.w8(32'h3b893683),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ea163),
	.w1(32'h3b61feb2),
	.w2(32'h3bf7f350),
	.w3(32'h3c703326),
	.w4(32'h3b9ce7e1),
	.w5(32'h3bad7060),
	.w6(32'h3ba1c315),
	.w7(32'h3ae5acf5),
	.w8(32'h3b5babc8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a638825),
	.w1(32'hb9f732e7),
	.w2(32'h3b2238be),
	.w3(32'hbc07b351),
	.w4(32'h3c10d47b),
	.w5(32'hbbb943d1),
	.w6(32'hbb825a83),
	.w7(32'h3c9ef2f1),
	.w8(32'hb9bed378),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8100b),
	.w1(32'hba840a2e),
	.w2(32'h3b660375),
	.w3(32'h3be00795),
	.w4(32'h3b53d290),
	.w5(32'hba52b6d3),
	.w6(32'h3c044683),
	.w7(32'hbabe5a0c),
	.w8(32'h3bca72fa),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62330b),
	.w1(32'hbba89f8d),
	.w2(32'hbb8db6eb),
	.w3(32'h36b43ae2),
	.w4(32'h3b81c144),
	.w5(32'h3b9f3a9c),
	.w6(32'h3abe21ea),
	.w7(32'h3b10c944),
	.w8(32'h3aa131e5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccc235),
	.w1(32'hbb9cf0c0),
	.w2(32'h3a0db889),
	.w3(32'h3b682a99),
	.w4(32'h3b587ba6),
	.w5(32'hbc73d6e3),
	.w6(32'hbb5c7ae9),
	.w7(32'hbc08a2e0),
	.w8(32'hbb9e41c7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b69a8),
	.w1(32'h3bdc6536),
	.w2(32'h3bb76a31),
	.w3(32'hbc276104),
	.w4(32'h3c604de0),
	.w5(32'h3bc1797a),
	.w6(32'hbca22592),
	.w7(32'h3c634bca),
	.w8(32'h3b77df87),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba199edf),
	.w1(32'hb82e834b),
	.w2(32'h3bb41f7b),
	.w3(32'hba59d65f),
	.w4(32'hbac45ef4),
	.w5(32'h3b8055d0),
	.w6(32'hbb76d0bd),
	.w7(32'hbac5c0ba),
	.w8(32'h3c13c665),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ad3f5),
	.w1(32'hbaff3f84),
	.w2(32'h3a9ab684),
	.w3(32'hbc1afbea),
	.w4(32'h3b04ed4f),
	.w5(32'h3bb958f0),
	.w6(32'hbc1fcf11),
	.w7(32'hbb8fa8ec),
	.w8(32'h3b6bc15e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b4bf2),
	.w1(32'hbc0c686f),
	.w2(32'hbb812f1e),
	.w3(32'h3aebdc98),
	.w4(32'hbb8b6010),
	.w5(32'hbc0e3f36),
	.w6(32'hbb6ed20b),
	.w7(32'hbc1ca1ff),
	.w8(32'hbb2c620e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e9bdc),
	.w1(32'hbc292826),
	.w2(32'h3b4575df),
	.w3(32'hbc5311bd),
	.w4(32'hbacc53fc),
	.w5(32'h3b62356c),
	.w6(32'hbca0d61f),
	.w7(32'hbb0a0a97),
	.w8(32'h3bdba187),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76d770),
	.w1(32'h3bc569d5),
	.w2(32'h3bee0f7f),
	.w3(32'h3c075cf4),
	.w4(32'h3ba44b30),
	.w5(32'h3c87163d),
	.w6(32'h3c05b4e6),
	.w7(32'h3bbc98e8),
	.w8(32'h3c6de6e7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac71204),
	.w1(32'h3c13ca77),
	.w2(32'hbb8b92bb),
	.w3(32'h3b7d59ec),
	.w4(32'h3bcc38af),
	.w5(32'h3aa403f9),
	.w6(32'hbb2e10d9),
	.w7(32'h3af2a7c9),
	.w8(32'hbb472518),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8d274),
	.w1(32'hbb9f8b13),
	.w2(32'hbbb0e64d),
	.w3(32'hbbdd2e52),
	.w4(32'h39ab510f),
	.w5(32'hbbb952ab),
	.w6(32'hbc1ee7f3),
	.w7(32'hbaa74948),
	.w8(32'hba22e456),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e694c),
	.w1(32'hbc2fcd47),
	.w2(32'h3c16f94d),
	.w3(32'h3ab3c1ae),
	.w4(32'hba2e0e98),
	.w5(32'h3bc03057),
	.w6(32'hbb09f961),
	.w7(32'hbbd98b0f),
	.w8(32'h3bf1c520),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17c666),
	.w1(32'h3cd17caa),
	.w2(32'hbaa14af6),
	.w3(32'hbc62c057),
	.w4(32'h3c78fe0b),
	.w5(32'hba832f7b),
	.w6(32'hbbed8d5e),
	.w7(32'h3cbf1ebb),
	.w8(32'h3aeb24f1),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9522d3),
	.w1(32'h3be01992),
	.w2(32'hbc04beb8),
	.w3(32'h3bab314c),
	.w4(32'h3b3237e4),
	.w5(32'hbb8601d4),
	.w6(32'h3bd1fa37),
	.w7(32'h3b49a584),
	.w8(32'hbb93db8b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41df3e),
	.w1(32'hbc8e4b66),
	.w2(32'hbc2243ce),
	.w3(32'hbc0e75ca),
	.w4(32'hbc4a9093),
	.w5(32'hbb4b86a6),
	.w6(32'hbc61c6a2),
	.w7(32'hbb08b752),
	.w8(32'hbb858129),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae43f35),
	.w1(32'h3c04c3fa),
	.w2(32'hba417b21),
	.w3(32'hbc1e6f7d),
	.w4(32'h3c0a13b3),
	.w5(32'hbc32b63c),
	.w6(32'hbcd909f5),
	.w7(32'h3aa5dd78),
	.w8(32'hbbc50f4a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbacde8),
	.w1(32'h3c05d954),
	.w2(32'h39d82eb1),
	.w3(32'hba236200),
	.w4(32'h3cc29c9f),
	.w5(32'h3c13f6a0),
	.w6(32'hbc34cb0f),
	.w7(32'h3c1ebad2),
	.w8(32'hbb177a66),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafff2b),
	.w1(32'hbacd7b3b),
	.w2(32'hbbc24c73),
	.w3(32'hbb752004),
	.w4(32'hbc265690),
	.w5(32'hbbb81403),
	.w6(32'h3ba34a66),
	.w7(32'hbcab1645),
	.w8(32'hbbfcd1bb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7cf13),
	.w1(32'h3a928be7),
	.w2(32'hbacae611),
	.w3(32'h39ed92fa),
	.w4(32'h3b09e66a),
	.w5(32'h3b1d141a),
	.w6(32'hbb4c8b39),
	.w7(32'h399f0296),
	.w8(32'hbc00ba1b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ec848),
	.w1(32'h3b0241fd),
	.w2(32'h3b996286),
	.w3(32'h3a9f6c1f),
	.w4(32'hbae87dba),
	.w5(32'h3a14fa48),
	.w6(32'hbbb053b4),
	.w7(32'hbbab07af),
	.w8(32'h3a9fdd98),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba548545),
	.w1(32'h3b0e4a60),
	.w2(32'hbb169385),
	.w3(32'hbb031436),
	.w4(32'h3b9e6c82),
	.w5(32'hbbfd6eaf),
	.w6(32'hbbb0d923),
	.w7(32'h3a2281fd),
	.w8(32'hbbec4981),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb7ad05),
	.w1(32'h3c90d21d),
	.w2(32'h3bbd202d),
	.w3(32'h3d3acd98),
	.w4(32'h3d0ce469),
	.w5(32'h3b937993),
	.w6(32'h3cef9641),
	.w7(32'h3d0ea7ec),
	.w8(32'h3aaacaca),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24d4a2),
	.w1(32'hbc99a806),
	.w2(32'h3b8278c0),
	.w3(32'hbb36a981),
	.w4(32'hbc857eab),
	.w5(32'h3baf7fe9),
	.w6(32'hbc037fcc),
	.w7(32'hbc555748),
	.w8(32'hbbcb4abd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e0336),
	.w1(32'hb9b6198f),
	.w2(32'h3bf9ed0a),
	.w3(32'h3b1d2588),
	.w4(32'h3b9cf056),
	.w5(32'h3a8e2afd),
	.w6(32'h3b8308df),
	.w7(32'hba5421f9),
	.w8(32'hbac443db),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad38397),
	.w1(32'hbc95120d),
	.w2(32'hbb3ada1b),
	.w3(32'h3c58f1ad),
	.w4(32'hbc2a8ac5),
	.w5(32'hbbd271f9),
	.w6(32'h3bf79f15),
	.w7(32'hbc321986),
	.w8(32'hbc40d8c4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f30ea),
	.w1(32'h3bac890c),
	.w2(32'h3b388ebb),
	.w3(32'hbc028415),
	.w4(32'hbb6dd2fe),
	.w5(32'hbbc4e43f),
	.w6(32'h3ae005de),
	.w7(32'h3c476f10),
	.w8(32'h3c1e6bb5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2565e4),
	.w1(32'h380023dc),
	.w2(32'hbb59a53e),
	.w3(32'h3abfbba3),
	.w4(32'h3934109e),
	.w5(32'hba8d7068),
	.w6(32'hbac66acc),
	.w7(32'h3b04883a),
	.w8(32'hbb16e922),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf577f),
	.w1(32'hbbd19183),
	.w2(32'h3c66527e),
	.w3(32'hba8f6759),
	.w4(32'h3b4f71f6),
	.w5(32'h3c109934),
	.w6(32'hbca8e53b),
	.w7(32'h3ade43a9),
	.w8(32'h3b757b8a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8cc1),
	.w1(32'hbc30fd90),
	.w2(32'h3c57ac3c),
	.w3(32'h3b8173bd),
	.w4(32'hbcec71f7),
	.w5(32'h3c49f561),
	.w6(32'h3a04523b),
	.w7(32'hbc8b7dc4),
	.w8(32'h3c6f7346),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e0f76),
	.w1(32'h3c86371c),
	.w2(32'h3b261b22),
	.w3(32'h3b58912f),
	.w4(32'h3c031e40),
	.w5(32'hbb3c6ea1),
	.w6(32'hbb28d1eb),
	.w7(32'h3acda12b),
	.w8(32'hbb5fa277),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76d276),
	.w1(32'hbb349c26),
	.w2(32'hbb0f01df),
	.w3(32'hbb3e714c),
	.w4(32'hbba1a40f),
	.w5(32'hb9d2e0a1),
	.w6(32'hbb9f8fa9),
	.w7(32'hbb5efab1),
	.w8(32'h3a123d80),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21fd1c),
	.w1(32'hbba34286),
	.w2(32'hbb61d60b),
	.w3(32'hbaa84d1b),
	.w4(32'h3803b7c5),
	.w5(32'hbbb6181b),
	.w6(32'h3b4255bc),
	.w7(32'h3ba246c6),
	.w8(32'hbac0957f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8077db),
	.w1(32'hba98b475),
	.w2(32'hbb29f417),
	.w3(32'h3b2ca4ef),
	.w4(32'hba63e4bc),
	.w5(32'hbc37a5dc),
	.w6(32'h3b85f9b0),
	.w7(32'h3b904be9),
	.w8(32'hbb3f3743),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86ca0d),
	.w1(32'h3aceed50),
	.w2(32'h3c3de3a4),
	.w3(32'hbb7bfcf3),
	.w4(32'h3a2f23bd),
	.w5(32'hba18c896),
	.w6(32'hbc68a8a2),
	.w7(32'h3b5fd7be),
	.w8(32'hbbb80568),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c351a60),
	.w1(32'h3cd3430d),
	.w2(32'hbb74edb8),
	.w3(32'h3c045cd9),
	.w4(32'h3d9bdb8c),
	.w5(32'hbaa9e971),
	.w6(32'hbce1f8a8),
	.w7(32'h3d7971bd),
	.w8(32'hbb85d450),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc345e68),
	.w1(32'hbab7deda),
	.w2(32'hb9a90e7b),
	.w3(32'hbc1f9718),
	.w4(32'h39aede1e),
	.w5(32'h3c1aea54),
	.w6(32'hbc47de6d),
	.w7(32'h3bfeb357),
	.w8(32'h3a8a6c1c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc172095),
	.w1(32'hbbb06085),
	.w2(32'h3b905c22),
	.w3(32'h3bb5e23d),
	.w4(32'h3bd7f8b1),
	.w5(32'h3b2136b0),
	.w6(32'h3bcd7496),
	.w7(32'h3b92f429),
	.w8(32'h3bc7eb19),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa3deb),
	.w1(32'hbb6ebd96),
	.w2(32'hba01dd64),
	.w3(32'hbc183eab),
	.w4(32'h3b67e427),
	.w5(32'h3b92421f),
	.w6(32'hbc55b64d),
	.w7(32'h3bddbef3),
	.w8(32'h3a8c19d9),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1165cf),
	.w1(32'h3b7159c6),
	.w2(32'hbc1cee48),
	.w3(32'h3bdd9eea),
	.w4(32'h3c51d500),
	.w5(32'hbbf0d24b),
	.w6(32'hbb3793f6),
	.w7(32'h3b21f680),
	.w8(32'hba507fdb),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55e2d9),
	.w1(32'h3c8ab94c),
	.w2(32'hbb4d88dc),
	.w3(32'hbc9cb2f8),
	.w4(32'h3ce8348f),
	.w5(32'hbc33b69b),
	.w6(32'hbc4a2bf8),
	.w7(32'h3c3ed77f),
	.w8(32'hbc02e80a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9528d3),
	.w1(32'h3c573e61),
	.w2(32'h3b29fd84),
	.w3(32'hbc9d2ce5),
	.w4(32'h3cd7bdad),
	.w5(32'h3baf8bc7),
	.w6(32'hbca54fc4),
	.w7(32'h3cb1e694),
	.w8(32'h3bfa80ba),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc188daa),
	.w1(32'h3b899c37),
	.w2(32'h3b0643e2),
	.w3(32'hbc0458fa),
	.w4(32'hbb25cf46),
	.w5(32'h3ac509c3),
	.w6(32'h3a9dafbd),
	.w7(32'hbb11613c),
	.w8(32'hb9ac60ff),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb461557),
	.w1(32'hbadcc008),
	.w2(32'h3b41c2d3),
	.w3(32'hb9ea4f3e),
	.w4(32'hba21f026),
	.w5(32'hbb95cdc1),
	.w6(32'hbab70fd8),
	.w7(32'h3b993e22),
	.w8(32'hbbcfeb91),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24533d),
	.w1(32'hbc12d1ef),
	.w2(32'hb9b0b981),
	.w3(32'h3c0b65f6),
	.w4(32'hbb08ec95),
	.w5(32'h3aeed5db),
	.w6(32'h3b8c21b6),
	.w7(32'h3b97feae),
	.w8(32'h3b60f98b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8fef3),
	.w1(32'h3c13c52d),
	.w2(32'h3aca150b),
	.w3(32'h3a51307f),
	.w4(32'h3bb85d30),
	.w5(32'h3b50ea9c),
	.w6(32'h3b521ace),
	.w7(32'h3be14f29),
	.w8(32'h3b1154dc),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad20b85),
	.w1(32'h3b4fa699),
	.w2(32'hbc3459f4),
	.w3(32'hbb5e98c8),
	.w4(32'h3b0eaf72),
	.w5(32'hbbbfae07),
	.w6(32'hbae2ec0b),
	.w7(32'h3b631d2f),
	.w8(32'hb9dd231d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d569f4),
	.w1(32'hbb60de89),
	.w2(32'hbbc13d31),
	.w3(32'h3a93dd3f),
	.w4(32'hbc072646),
	.w5(32'h3b1c944b),
	.w6(32'h3ac01e0e),
	.w7(32'hbb8efefc),
	.w8(32'hbb23218d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc903f),
	.w1(32'h3c077910),
	.w2(32'h3b350cd1),
	.w3(32'hbb2a584e),
	.w4(32'h3a1c8d49),
	.w5(32'hbb66f57a),
	.w6(32'h397b328f),
	.w7(32'hbc464272),
	.w8(32'h3c12b23f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf77ff3),
	.w1(32'h3ca21f2f),
	.w2(32'h3b531915),
	.w3(32'hbc17e9cb),
	.w4(32'h3c9b72f0),
	.w5(32'hb9c1aaad),
	.w6(32'h3a936226),
	.w7(32'h3c04f938),
	.w8(32'hbba1708a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88f78b),
	.w1(32'h3c0bbddf),
	.w2(32'hb8d23c95),
	.w3(32'hbb797dc7),
	.w4(32'h3bc21fe9),
	.w5(32'hba233880),
	.w6(32'h3bae2372),
	.w7(32'h3c74a445),
	.w8(32'hbb29d717),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c864165),
	.w1(32'h3c257cc4),
	.w2(32'h3b90e530),
	.w3(32'h3c8b7f0c),
	.w4(32'h3c57802b),
	.w5(32'h3b94207f),
	.w6(32'h3c0b078b),
	.w7(32'h3c6443b6),
	.w8(32'h3c0ab169),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07cfb8),
	.w1(32'hbbef8a58),
	.w2(32'h3882080f),
	.w3(32'hbb9a6752),
	.w4(32'hbc895864),
	.w5(32'hba9bba40),
	.w6(32'hbbabd147),
	.w7(32'hbcdcb366),
	.w8(32'hba8f4e67),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b9661),
	.w1(32'h3bb17bf3),
	.w2(32'h3c3d54e1),
	.w3(32'hbb220430),
	.w4(32'h3b9230f5),
	.w5(32'h3c7ce63a),
	.w6(32'h3c21b4b1),
	.w7(32'h3b3cec42),
	.w8(32'h3c69fde7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d29f6),
	.w1(32'h3ba7d87c),
	.w2(32'hbad8af6d),
	.w3(32'hbc6aa44b),
	.w4(32'hba183546),
	.w5(32'hba7d873d),
	.w6(32'hbc3a7b20),
	.w7(32'h3a99c858),
	.w8(32'h3b60541c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6576a),
	.w1(32'h3b32b5d4),
	.w2(32'h3b46f5cf),
	.w3(32'h3bb16ac3),
	.w4(32'h3c0c680d),
	.w5(32'h3b9d5b71),
	.w6(32'h3aba160f),
	.w7(32'h3b21eaee),
	.w8(32'h3b905845),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749d58),
	.w1(32'hbbbbe0c2),
	.w2(32'h3b131275),
	.w3(32'h3bcd4cc8),
	.w4(32'hbb44a3ac),
	.w5(32'h3b48d7ca),
	.w6(32'h3c15c27d),
	.w7(32'h3c023271),
	.w8(32'h3b790e74),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf4f8e),
	.w1(32'hbb675e40),
	.w2(32'hbb19bbaa),
	.w3(32'h3b727035),
	.w4(32'h3b180925),
	.w5(32'hbb8c3b04),
	.w6(32'h3b900e37),
	.w7(32'h3b19eff7),
	.w8(32'h3babdc51),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47318e),
	.w1(32'h3bd6f72f),
	.w2(32'hbc40b0bb),
	.w3(32'hbc9407f0),
	.w4(32'h3ca0df1d),
	.w5(32'hbc73e686),
	.w6(32'hbc6f7500),
	.w7(32'h3c4076df),
	.w8(32'hbbd1a569),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbae511),
	.w1(32'h3caa20b8),
	.w2(32'hbbd23aff),
	.w3(32'hbc6cc4e8),
	.w4(32'h3cea23ba),
	.w5(32'hbac05900),
	.w6(32'hbcb6f96d),
	.w7(32'h3cdbf5aa),
	.w8(32'hbb7a02f3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6096be),
	.w1(32'hbb1cce25),
	.w2(32'hba8ee1cd),
	.w3(32'hbc00b2d3),
	.w4(32'h3bc0e3c9),
	.w5(32'hba4229ef),
	.w6(32'hbb830fb5),
	.w7(32'h3c917759),
	.w8(32'hbb0a3dec),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5313ee),
	.w1(32'hbaa5f75e),
	.w2(32'hbab92ffa),
	.w3(32'hb8a2e946),
	.w4(32'hbbd38c5d),
	.w5(32'hba5f1015),
	.w6(32'h3ad15e2e),
	.w7(32'hbbb874d5),
	.w8(32'hbb66b139),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81dc95),
	.w1(32'hbb99b439),
	.w2(32'hba4a7b70),
	.w3(32'hb9d141c5),
	.w4(32'hbaf9983a),
	.w5(32'h3c065e1e),
	.w6(32'hbb37a2b6),
	.w7(32'hbbc63043),
	.w8(32'h3a448dab),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6eacfb),
	.w1(32'hbbd74363),
	.w2(32'h3b17b7a8),
	.w3(32'hbcd0cf53),
	.w4(32'hbc7b0a08),
	.w5(32'h3bd97408),
	.w6(32'hbc91f8f6),
	.w7(32'hbc1f3dcf),
	.w8(32'h3bd1dff7),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf46a5),
	.w1(32'hbb23832e),
	.w2(32'h3bd7cdc9),
	.w3(32'hbb1b58ee),
	.w4(32'hb9cda928),
	.w5(32'hbbaab146),
	.w6(32'hb94ef724),
	.w7(32'h3aad12b5),
	.w8(32'hbb686e5c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f7440),
	.w1(32'hbc13f045),
	.w2(32'hbb5ee1bb),
	.w3(32'h3ba8b506),
	.w4(32'hbc1abad1),
	.w5(32'hbc66d491),
	.w6(32'hbc0d865f),
	.w7(32'hbc162d5a),
	.w8(32'hb9b04b91),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8f544),
	.w1(32'hba84028b),
	.w2(32'h3ac1b3ba),
	.w3(32'h3be42e91),
	.w4(32'h3c766e97),
	.w5(32'hbb774a21),
	.w6(32'hbbc2362f),
	.w7(32'hbb822409),
	.w8(32'hbb9a9364),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a5e42),
	.w1(32'hbc682ccb),
	.w2(32'h3b504aac),
	.w3(32'hbb8dd551),
	.w4(32'hbc308bad),
	.w5(32'hbb500c65),
	.w6(32'hbc298e55),
	.w7(32'hbc368cf3),
	.w8(32'hbc4bfe09),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule