module layer_8_featuremap_49(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba886e7a),
	.w1(32'hb9c6fdd9),
	.w2(32'hb9db6e82),
	.w3(32'hbb038f3f),
	.w4(32'hbaa22a6c),
	.w5(32'hba40f533),
	.w6(32'hbacd1dfd),
	.w7(32'hba40580f),
	.w8(32'h39932ed8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40bf9e),
	.w1(32'hbadbe459),
	.w2(32'hbb21e269),
	.w3(32'hbaf0a3f3),
	.w4(32'hba54a397),
	.w5(32'hbb25a809),
	.w6(32'hba9a3b68),
	.w7(32'hb9947b8e),
	.w8(32'hba942e5f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba197699),
	.w1(32'hba373043),
	.w2(32'h39242766),
	.w3(32'hb9c0fe7c),
	.w4(32'hba89e588),
	.w5(32'hba8dab78),
	.w6(32'hba3be261),
	.w7(32'hb9b193b1),
	.w8(32'hbaf0f74d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f7c7e),
	.w1(32'hb9f86d79),
	.w2(32'h3b42fcfc),
	.w3(32'hb921ab5e),
	.w4(32'hba8ad9e5),
	.w5(32'h3a317cab),
	.w6(32'hbac6bd86),
	.w7(32'hb96261b8),
	.w8(32'h388f6b3d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57c1bd),
	.w1(32'hbb3d0536),
	.w2(32'hbb0e2fc3),
	.w3(32'hbaa9df25),
	.w4(32'hba57a743),
	.w5(32'hba4b0822),
	.w6(32'h39eadd4a),
	.w7(32'h3a81f472),
	.w8(32'hba0fc649),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada8225),
	.w1(32'h3b38b3ff),
	.w2(32'h3b373f3a),
	.w3(32'h3a3eb210),
	.w4(32'h3a99e254),
	.w5(32'h3ad19635),
	.w6(32'hba03d7a3),
	.w7(32'hb82076b7),
	.w8(32'hb99471de),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9642cdd),
	.w1(32'hb8b89dad),
	.w2(32'hb9a05336),
	.w3(32'h399a36d9),
	.w4(32'h39e0e3e5),
	.w5(32'h3a0f60de),
	.w6(32'h39aaa7dc),
	.w7(32'h393335da),
	.w8(32'hb8b81b09),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba946cfa),
	.w1(32'h3a031bb7),
	.w2(32'hbaca7d11),
	.w3(32'hbb420cda),
	.w4(32'hbb5a0080),
	.w5(32'hbba4dca3),
	.w6(32'hb96d41e6),
	.w7(32'hbae126ec),
	.w8(32'hbb1b4d06),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc965a),
	.w1(32'hbb966a1b),
	.w2(32'hbb89931d),
	.w3(32'hbb651089),
	.w4(32'hbaaa7da1),
	.w5(32'hbaaedf7a),
	.w6(32'hbaa0858a),
	.w7(32'hba0fee67),
	.w8(32'hbb55bace),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb169aa),
	.w1(32'hbb7e6f28),
	.w2(32'hba96d617),
	.w3(32'hbb5c896d),
	.w4(32'hbb14caf8),
	.w5(32'hbaae430a),
	.w6(32'hbb72b48e),
	.w7(32'hbac20e6b),
	.w8(32'h3a4e06db),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f72a6),
	.w1(32'hb91922db),
	.w2(32'hba29e478),
	.w3(32'h3ac09798),
	.w4(32'h3a5d6cdc),
	.w5(32'hba23bbff),
	.w6(32'h3ac8b52a),
	.w7(32'h3ac39a72),
	.w8(32'hb9937b34),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9bb7e),
	.w1(32'hb9f862f3),
	.w2(32'hba826f0e),
	.w3(32'hba23d1d2),
	.w4(32'hb9068966),
	.w5(32'hb9b2e702),
	.w6(32'hba3ccf2e),
	.w7(32'hba3d4473),
	.w8(32'hba08e9a5),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac75c57),
	.w1(32'hba9587c5),
	.w2(32'hb95e12e5),
	.w3(32'hbab8f94d),
	.w4(32'hba99fb72),
	.w5(32'hba1f6d16),
	.w6(32'hba9f9d08),
	.w7(32'hbb114112),
	.w8(32'hbb06b967),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1dc05),
	.w1(32'h3aa8ff69),
	.w2(32'h3ad98eec),
	.w3(32'h3ab133f4),
	.w4(32'h3aea4a05),
	.w5(32'h3b4b6274),
	.w6(32'h376b9dc9),
	.w7(32'h3a84c1f1),
	.w8(32'h3af98dcc),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922856b),
	.w1(32'hb6ca7e8c),
	.w2(32'h394a20af),
	.w3(32'h3a1b08ed),
	.w4(32'h39d1b2dd),
	.w5(32'h3a26d83d),
	.w6(32'h398719c3),
	.w7(32'h3980b6b7),
	.w8(32'hba14f9af),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955fa07),
	.w1(32'h3a3a954d),
	.w2(32'h39856610),
	.w3(32'h39bf81b1),
	.w4(32'h39babd76),
	.w5(32'hb84ab684),
	.w6(32'h39dce37a),
	.w7(32'h3a5eb7df),
	.w8(32'hbb31ea3a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00cb98),
	.w1(32'hbb3213a9),
	.w2(32'h3b7ba2a2),
	.w3(32'hbb5b7cd5),
	.w4(32'hbb129af4),
	.w5(32'h3b232a19),
	.w6(32'hbb83a385),
	.w7(32'hbb16e830),
	.w8(32'h38261483),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac65a7d),
	.w1(32'hba36db3f),
	.w2(32'h3972ea41),
	.w3(32'hba475028),
	.w4(32'hbae50893),
	.w5(32'hb96b140f),
	.w6(32'h3a7c86bc),
	.w7(32'h38b345b6),
	.w8(32'h3a7d632c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a6e5),
	.w1(32'hbb81f1d0),
	.w2(32'hbb8fcbb1),
	.w3(32'hbb7e8047),
	.w4(32'hbb8dccf7),
	.w5(32'hbb9f4b31),
	.w6(32'h3a523550),
	.w7(32'hba1d6144),
	.w8(32'hbbad27da),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb375558),
	.w1(32'hbb06a3de),
	.w2(32'h3a6a94c4),
	.w3(32'hb99e32ec),
	.w4(32'hbbd6dfa8),
	.w5(32'hbb5ebb74),
	.w6(32'h3bd1a8a4),
	.w7(32'h3c0eb07a),
	.w8(32'h3c053361),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0f2ed),
	.w1(32'h391bdd13),
	.w2(32'hba887cc8),
	.w3(32'h3a95660a),
	.w4(32'h3a882304),
	.w5(32'h3a75b236),
	.w6(32'hba6d6baa),
	.w7(32'hbb453e9c),
	.w8(32'hb99cafbf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18a143),
	.w1(32'hbbb4bb5b),
	.w2(32'hbb60a8b6),
	.w3(32'hbbf00a82),
	.w4(32'hbbfa2c2b),
	.w5(32'hbb98916a),
	.w6(32'hbba63435),
	.w7(32'hbbabf309),
	.w8(32'h3a16a5fd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf4f1d),
	.w1(32'hbb346b2d),
	.w2(32'hbba03b45),
	.w3(32'h3b8ff74c),
	.w4(32'hb9bb7f92),
	.w5(32'hbb2c9b79),
	.w6(32'h3c16ce2f),
	.w7(32'h3bcded86),
	.w8(32'h3b99bc88),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2828b9),
	.w1(32'hbad3af57),
	.w2(32'hbb05fbcd),
	.w3(32'hbb04d536),
	.w4(32'hbb0407b8),
	.w5(32'hbb20e991),
	.w6(32'hb89d1ce3),
	.w7(32'hba1777d2),
	.w8(32'hbb033e8b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73f53e),
	.w1(32'h3bd4a5a2),
	.w2(32'h3b02bba8),
	.w3(32'hb9332ab0),
	.w4(32'h3b812cd4),
	.w5(32'h3a044963),
	.w6(32'h393f1ff5),
	.w7(32'hb8c89862),
	.w8(32'h3a80d72c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb308cf2),
	.w1(32'hbb039a09),
	.w2(32'hbbc8cc3c),
	.w3(32'h39da6319),
	.w4(32'hba35a0fa),
	.w5(32'hbb875797),
	.w6(32'h3a655756),
	.w7(32'h391cb155),
	.w8(32'h39c4ac5e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39688cab),
	.w1(32'h37aa4718),
	.w2(32'hbb07affb),
	.w3(32'h3ab390ce),
	.w4(32'h3aaaa7f8),
	.w5(32'hba862b9d),
	.w6(32'h3a0bc9b8),
	.w7(32'hbab6c2a4),
	.w8(32'h3a787d6f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb561547),
	.w1(32'hbace7edf),
	.w2(32'hbbfc1c08),
	.w3(32'hbb69fa06),
	.w4(32'hb9b5a365),
	.w5(32'hbc0b1a40),
	.w6(32'hbab449c2),
	.w7(32'hbafde4dc),
	.w8(32'hbb8d39bd),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75fb48),
	.w1(32'h3b704f79),
	.w2(32'hbb97e89e),
	.w3(32'hbb8abf50),
	.w4(32'h3a947095),
	.w5(32'hbb244a65),
	.w6(32'h3a002664),
	.w7(32'hb9e1c232),
	.w8(32'hba0f7354),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9530335),
	.w1(32'hb92c6cbb),
	.w2(32'hb9112e8d),
	.w3(32'h3a37694b),
	.w4(32'h39fdd94a),
	.w5(32'h3a30bd44),
	.w6(32'h3a621c47),
	.w7(32'h3a7cfd8d),
	.w8(32'h39ef88d4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57c397),
	.w1(32'hbba447c6),
	.w2(32'h3b3dc429),
	.w3(32'hbb7a4bc2),
	.w4(32'hbbc15b9a),
	.w5(32'hbb46d355),
	.w6(32'hbbccdb62),
	.w7(32'hbbc1fea2),
	.w8(32'hbb18466d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3cd53),
	.w1(32'hba966b0e),
	.w2(32'hbb6c7256),
	.w3(32'hbb1529f4),
	.w4(32'hb9c899a5),
	.w5(32'hbb20460c),
	.w6(32'hba1ae9ec),
	.w7(32'hbb0f7cff),
	.w8(32'hbac194a9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e5d00),
	.w1(32'hba1c262a),
	.w2(32'h3b66b247),
	.w3(32'hb85deff6),
	.w4(32'hba89592d),
	.w5(32'h3a97c7b6),
	.w6(32'hbb05e408),
	.w7(32'h39e7dfd6),
	.w8(32'hba7245bf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ba16f),
	.w1(32'hbb49104f),
	.w2(32'hbacd7783),
	.w3(32'hbb0cc02c),
	.w4(32'hbbc9a0e9),
	.w5(32'hbb3d5bee),
	.w6(32'h38d30c72),
	.w7(32'hb8cf312b),
	.w8(32'h398e026b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9429f5),
	.w1(32'h396bccd1),
	.w2(32'h3a60c012),
	.w3(32'h3ad8dac0),
	.w4(32'h3aea8753),
	.w5(32'h3b3361b9),
	.w6(32'h3a721374),
	.w7(32'h3b26a91d),
	.w8(32'h3b15494d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a2196),
	.w1(32'h38dfb953),
	.w2(32'hbaf365a1),
	.w3(32'h3a16ee8e),
	.w4(32'hba928861),
	.w5(32'hbb046887),
	.w6(32'h3a98a03c),
	.w7(32'hba8bb6cd),
	.w8(32'hbb0da91e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6f33f),
	.w1(32'h3a83ef9e),
	.w2(32'h3a5cb75d),
	.w3(32'hba421673),
	.w4(32'h3a0c9c94),
	.w5(32'h397cabfc),
	.w6(32'h3a91467d),
	.w7(32'h3a89658f),
	.w8(32'h3aaf5e43),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac07065),
	.w1(32'hbabcc6a0),
	.w2(32'hbaad9881),
	.w3(32'hb816e80d),
	.w4(32'h38d187fd),
	.w5(32'h38f92de1),
	.w6(32'h3a9b7402),
	.w7(32'h3b19073b),
	.w8(32'h3b2bf030),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ce0b4),
	.w1(32'h3a0c7843),
	.w2(32'h3a158524),
	.w3(32'h3a79176f),
	.w4(32'h3a1b0662),
	.w5(32'h3a4a4a31),
	.w6(32'h3a074d9d),
	.w7(32'h39768fc0),
	.w8(32'h3a11305f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39949bc9),
	.w1(32'h3ab1b43b),
	.w2(32'h36d57cc3),
	.w3(32'h392919f9),
	.w4(32'h3a957659),
	.w5(32'hb91d0c8a),
	.w6(32'h3a84d22c),
	.w7(32'hb9b00fab),
	.w8(32'hb9a65d30),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903d23d),
	.w1(32'hb96f4507),
	.w2(32'hbaac0bfa),
	.w3(32'h3a45357c),
	.w4(32'h3a87125f),
	.w5(32'hba039ed8),
	.w6(32'h3a29bf78),
	.w7(32'h39482edc),
	.w8(32'hba3b10f3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb550007),
	.w1(32'hbb9fe18e),
	.w2(32'hbb9392a0),
	.w3(32'hbb49d417),
	.w4(32'hbb90b5e8),
	.w5(32'hbb8f0c86),
	.w6(32'hbba0bdd9),
	.w7(32'hbb88c103),
	.w8(32'h3b80570f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dcb16),
	.w1(32'hbb5730b6),
	.w2(32'hbb441880),
	.w3(32'h3bb98c67),
	.w4(32'hbb83642e),
	.w5(32'hbbb24840),
	.w6(32'hba21b75c),
	.w7(32'hba34cdfb),
	.w8(32'hbacae216),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4ca5c),
	.w1(32'hbb8e480b),
	.w2(32'hbb6a2d53),
	.w3(32'hba814b87),
	.w4(32'hbb5165ea),
	.w5(32'hbb40a09e),
	.w6(32'hbb3ee2f4),
	.w7(32'hbb23cf95),
	.w8(32'hba0da3f2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe34e41),
	.w1(32'hbc1315cf),
	.w2(32'hbc0dd0c9),
	.w3(32'hbbb9b22b),
	.w4(32'hbc1d619f),
	.w5(32'hbc1fc8c4),
	.w6(32'hbb985712),
	.w7(32'hbbab412a),
	.w8(32'hbbfd1a3a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ef3ba),
	.w1(32'hbb84bbf6),
	.w2(32'hbb99b98d),
	.w3(32'hbae186f4),
	.w4(32'hbb23a67e),
	.w5(32'hbb382722),
	.w6(32'hbb899be2),
	.w7(32'hbb9bfac6),
	.w8(32'h3ac2463c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b719619),
	.w1(32'hbb974cb1),
	.w2(32'hbb246f9d),
	.w3(32'h39822658),
	.w4(32'hbbdcf7b4),
	.w5(32'hbb491611),
	.w6(32'hba69503a),
	.w7(32'hbb879317),
	.w8(32'hbb0a2dce),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1722f3),
	.w1(32'hbb83d40c),
	.w2(32'hbad81ec4),
	.w3(32'h3ae54c27),
	.w4(32'hbb95622e),
	.w5(32'hbb7866f6),
	.w6(32'h3a4850e2),
	.w7(32'h39ab429b),
	.w8(32'hba962425),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7462),
	.w1(32'h3ac7e40d),
	.w2(32'h39755b19),
	.w3(32'hbb994752),
	.w4(32'h39ef596b),
	.w5(32'hba447405),
	.w6(32'hb9f65e8f),
	.w7(32'hbaeec8ff),
	.w8(32'hbaf8bd3b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82de78),
	.w1(32'hbbc7e18c),
	.w2(32'hbbae1572),
	.w3(32'hbb139e22),
	.w4(32'hbb827e93),
	.w5(32'hbb8f7c9b),
	.w6(32'hbb87c210),
	.w7(32'hbb51a07c),
	.w8(32'hbad5ebb4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb145bbe),
	.w1(32'hbb1a1aa6),
	.w2(32'hbb0b2733),
	.w3(32'hbad66025),
	.w4(32'hbad781b9),
	.w5(32'hba3f610c),
	.w6(32'hbb2ab802),
	.w7(32'hbade4e99),
	.w8(32'hbab3dccc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75e259),
	.w1(32'hbb826781),
	.w2(32'hbb43048d),
	.w3(32'hbbca68ea),
	.w4(32'hbc40a0ac),
	.w5(32'hbc2fdd94),
	.w6(32'hbb872730),
	.w7(32'hbb89707b),
	.w8(32'hbbbc869f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a1633),
	.w1(32'h3c60cb99),
	.w2(32'h3b45bc93),
	.w3(32'hbbae3f92),
	.w4(32'h3b8225ce),
	.w5(32'hbb8f7de9),
	.w6(32'h3c1abe9e),
	.w7(32'h3af8684d),
	.w8(32'hbb0f204f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f53b2f),
	.w1(32'h3a8fceb8),
	.w2(32'hb7b5b32f),
	.w3(32'hb9560025),
	.w4(32'h3b1e8b93),
	.w5(32'h3b14b88e),
	.w6(32'hb9f70ef6),
	.w7(32'hbb581b6b),
	.w8(32'hbba358ce),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1529e),
	.w1(32'hbb8fb2cf),
	.w2(32'hbb3b2f9a),
	.w3(32'h3a69bf30),
	.w4(32'hbb3d2f26),
	.w5(32'hbb94f5d8),
	.w6(32'hba440fc4),
	.w7(32'hbb22665e),
	.w8(32'h3b72a62b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4a738),
	.w1(32'hbb11cb6f),
	.w2(32'hbb956357),
	.w3(32'hb9e91947),
	.w4(32'hbae4cdf9),
	.w5(32'hbb821179),
	.w6(32'h3a9cbff5),
	.w7(32'hba5b9b35),
	.w8(32'hbb97f558),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966e067),
	.w1(32'h3a856803),
	.w2(32'h3b1524aa),
	.w3(32'hb9e53c1a),
	.w4(32'hb932f3e8),
	.w5(32'hb9e5e92c),
	.w6(32'hbaaea11a),
	.w7(32'h3a9a3c93),
	.w8(32'h3ad98d86),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d18b4),
	.w1(32'hbac22075),
	.w2(32'hba7f7245),
	.w3(32'hba40bd28),
	.w4(32'hbbea0838),
	.w5(32'hbc2804da),
	.w6(32'hbb422999),
	.w7(32'hbb7d5536),
	.w8(32'hbbab7960),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a478d21),
	.w1(32'h3945fd8e),
	.w2(32'hb9fcf326),
	.w3(32'hb93cf8b4),
	.w4(32'hba53d9cc),
	.w5(32'hbafd3ea5),
	.w6(32'hb9a8a131),
	.w7(32'hba8d17b2),
	.w8(32'hbafc726b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b105819),
	.w1(32'h3b753578),
	.w2(32'hbb03e882),
	.w3(32'h3a678a53),
	.w4(32'h3ae8b1a5),
	.w5(32'hba859af0),
	.w6(32'h3ae54b50),
	.w7(32'hbb8fb3b6),
	.w8(32'hbb34be1c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56f280),
	.w1(32'h3b7a2de6),
	.w2(32'h3b80054d),
	.w3(32'hbb0772fe),
	.w4(32'hba40f38d),
	.w5(32'hba6bbb3e),
	.w6(32'hbb19ec98),
	.w7(32'hbaf368ff),
	.w8(32'hbad018d2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7de75f),
	.w1(32'hbb590ddc),
	.w2(32'hbb69c840),
	.w3(32'hbabe2070),
	.w4(32'hbb621d1e),
	.w5(32'hbb771f8b),
	.w6(32'hbb0ca847),
	.w7(32'hbb474693),
	.w8(32'h3ac323be),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3970dc),
	.w1(32'hbb66777b),
	.w2(32'hbb80b7de),
	.w3(32'h3a553ca8),
	.w4(32'hbb20c3d5),
	.w5(32'hbb881bc6),
	.w6(32'hba934f41),
	.w7(32'hbb1507b0),
	.w8(32'hbbc77add),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4270c),
	.w1(32'hbaa5228e),
	.w2(32'hbbb951f8),
	.w3(32'hbb6842db),
	.w4(32'hbc0764c5),
	.w5(32'hbc160c59),
	.w6(32'hbbad6cea),
	.w7(32'hbb0aeea8),
	.w8(32'hbb1e02ec),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaaae5),
	.w1(32'hbb6b31d2),
	.w2(32'hbb1fcd63),
	.w3(32'hbaa9e6f1),
	.w4(32'hbb562911),
	.w5(32'hbb3493cd),
	.w6(32'hbb829ed2),
	.w7(32'hbb6e23a4),
	.w8(32'hbabceb14),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca94cb),
	.w1(32'hbb6ed79e),
	.w2(32'hbb51a94c),
	.w3(32'hbaa679da),
	.w4(32'hbb52b7c2),
	.w5(32'hbb801272),
	.w6(32'hbad18de0),
	.w7(32'hbb064c51),
	.w8(32'hbb1d7e46),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c513a),
	.w1(32'hbb106b42),
	.w2(32'hbb090e09),
	.w3(32'hb9ef3b0c),
	.w4(32'hbb252c8b),
	.w5(32'hbb83abdd),
	.w6(32'hba762ccd),
	.w7(32'hba937c66),
	.w8(32'hbb071066),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65e207),
	.w1(32'hba89f27b),
	.w2(32'hba48cb2c),
	.w3(32'h3ac5daa7),
	.w4(32'hbaba2581),
	.w5(32'hb9a0adab),
	.w6(32'hbb026254),
	.w7(32'hbb41e2c6),
	.w8(32'hba5b159f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad9cc3),
	.w1(32'hbaa37a5a),
	.w2(32'hbb19bff9),
	.w3(32'h3ab486f3),
	.w4(32'hba53de17),
	.w5(32'hbae85479),
	.w6(32'hbaabbd5a),
	.w7(32'hbb0913c2),
	.w8(32'h3a85c0c9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80608c),
	.w1(32'hbb51986d),
	.w2(32'hbb439426),
	.w3(32'h3b81b245),
	.w4(32'hbb85019d),
	.w5(32'hbbc5a9a3),
	.w6(32'h3a086307),
	.w7(32'h37719399),
	.w8(32'hba5b591d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed9cf5),
	.w1(32'hbb7e7539),
	.w2(32'hbb764ed4),
	.w3(32'hbb089a7e),
	.w4(32'hbb522a6f),
	.w5(32'hbb3b431b),
	.w6(32'hbb8d0bf5),
	.w7(32'hbb84c71d),
	.w8(32'hbab24276),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad40561),
	.w1(32'hbb6221a7),
	.w2(32'hbb799b5b),
	.w3(32'hba9e8d95),
	.w4(32'hbb4e6774),
	.w5(32'hbb7618ca),
	.w6(32'hbb0e2f4f),
	.w7(32'hba674ee7),
	.w8(32'hba649092),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf740db),
	.w1(32'hbba5a0a0),
	.w2(32'hbb9cc8de),
	.w3(32'hbad5cc0a),
	.w4(32'hbb73a54e),
	.w5(32'hbb6748f3),
	.w6(32'hbb89c5a9),
	.w7(32'hbb8e94a9),
	.w8(32'hba4cb02c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379a03f1),
	.w1(32'h3b27162f),
	.w2(32'h3ac2fef5),
	.w3(32'hbb2a3775),
	.w4(32'hba62b0fe),
	.w5(32'h385834c1),
	.w6(32'h3a4610db),
	.w7(32'h3abe5bce),
	.w8(32'hba8b944c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2931f2),
	.w1(32'hbb88ecc2),
	.w2(32'hbb896684),
	.w3(32'hbb0af181),
	.w4(32'hbb68cf7b),
	.w5(32'hbb6cba46),
	.w6(32'hbb6f70dc),
	.w7(32'hbb670e71),
	.w8(32'hbab24635),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ecfb7),
	.w1(32'hba9b6fc3),
	.w2(32'hbaa68076),
	.w3(32'h3a3db4b2),
	.w4(32'hba28822a),
	.w5(32'hbad5fcd7),
	.w6(32'hba25f055),
	.w7(32'h390ca3b4),
	.w8(32'hb9ba56a7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0ce59),
	.w1(32'hbb5998b6),
	.w2(32'hbb6444ef),
	.w3(32'hba9ec8a5),
	.w4(32'hbb382b19),
	.w5(32'hbb34d891),
	.w6(32'hbb4091b0),
	.w7(32'hbb4da736),
	.w8(32'h3ab8940f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abce377),
	.w1(32'hbb7da903),
	.w2(32'hbb715c6d),
	.w3(32'h3ad609ea),
	.w4(32'hbba4361d),
	.w5(32'hbbdb5f03),
	.w6(32'hbb13aa3f),
	.w7(32'hbacfb4f3),
	.w8(32'h3ab197d6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bbdcc),
	.w1(32'hb98defbf),
	.w2(32'h3a769c66),
	.w3(32'h3b955896),
	.w4(32'h3a6146aa),
	.w5(32'hba00fa18),
	.w6(32'h38e77295),
	.w7(32'h39f9d117),
	.w8(32'h3a564ad0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba775187),
	.w1(32'hbac99a4d),
	.w2(32'hbad9445f),
	.w3(32'hb9715456),
	.w4(32'hba7d33a4),
	.w5(32'hba6d09c2),
	.w6(32'hba22dace),
	.w7(32'hba5fa241),
	.w8(32'h3a8ea9ef),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c123685),
	.w1(32'h3c0f0f2f),
	.w2(32'h3b9cc8e6),
	.w3(32'hbbe3a237),
	.w4(32'hbb47e74b),
	.w5(32'hbb601d90),
	.w6(32'h3b4860d0),
	.w7(32'h3ac7a4cb),
	.w8(32'hbaa187cc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d31e3),
	.w1(32'hbb31c4ff),
	.w2(32'hbb43fc38),
	.w3(32'hbb14e5c7),
	.w4(32'hbb0c2ef9),
	.w5(32'hbadd5820),
	.w6(32'hbaa586e5),
	.w7(32'hb9d54a70),
	.w8(32'hba5be7f6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6d446),
	.w1(32'hbc08f850),
	.w2(32'hbc0725c6),
	.w3(32'hbb4b11bc),
	.w4(32'hbbe9adcd),
	.w5(32'hbbfea2ad),
	.w6(32'hbb3a229b),
	.w7(32'hbb1f4321),
	.w8(32'hbbd05891),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d956e),
	.w1(32'h3a95fdbf),
	.w2(32'hbb51eb46),
	.w3(32'hbc1960a4),
	.w4(32'hb9dff18c),
	.w5(32'hbb8cfae6),
	.w6(32'h3ae4cc25),
	.w7(32'hb9bbd1d5),
	.w8(32'h38958626),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398caab2),
	.w1(32'h3aea7259),
	.w2(32'h3a1d151f),
	.w3(32'h3b3e51e5),
	.w4(32'h3b97f6ef),
	.w5(32'h3b1a6db4),
	.w6(32'h3b9c6116),
	.w7(32'h3bc3a7de),
	.w8(32'h3b38b222),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14286c),
	.w1(32'hbaff2a75),
	.w2(32'hbb511edb),
	.w3(32'h3b83f739),
	.w4(32'hbad6da26),
	.w5(32'hbb6951ac),
	.w6(32'h3b1af526),
	.w7(32'hbb013189),
	.w8(32'hbbe9a14d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b157e),
	.w1(32'h3aed0373),
	.w2(32'h398f5e9a),
	.w3(32'hbbb941c4),
	.w4(32'h3a02778b),
	.w5(32'hb9c30b1b),
	.w6(32'hb80a6eef),
	.w7(32'hbb10baac),
	.w8(32'hbac3371f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba804a58),
	.w1(32'hbb4cf5e3),
	.w2(32'hbb38db79),
	.w3(32'hb9daf525),
	.w4(32'hbb31627c),
	.w5(32'hbb33b339),
	.w6(32'hbb64ebc5),
	.w7(32'hbb4d9da3),
	.w8(32'hbb5bbbbd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba244219),
	.w1(32'h3b22482f),
	.w2(32'hbb154d84),
	.w3(32'hbb04db9b),
	.w4(32'h3a716bf3),
	.w5(32'hbb0f138c),
	.w6(32'h39905944),
	.w7(32'hbb602a50),
	.w8(32'hbbc1f082),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44acf8),
	.w1(32'h394c6b4e),
	.w2(32'hbaf133ba),
	.w3(32'hbb9465a3),
	.w4(32'h398c240e),
	.w5(32'hbab4c6aa),
	.w6(32'h39a872bc),
	.w7(32'hbb1a320e),
	.w8(32'hbbd39456),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7374ad),
	.w1(32'h3a507dcc),
	.w2(32'hb8d87bb4),
	.w3(32'hbbc24ab9),
	.w4(32'hba86c2f5),
	.w5(32'hbabe0c6c),
	.w6(32'hbabe257f),
	.w7(32'hbb5a40c3),
	.w8(32'hbb20246f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c5ab8),
	.w1(32'h3b727564),
	.w2(32'h3a8b3746),
	.w3(32'h3ae32744),
	.w4(32'h3b7dfcd9),
	.w5(32'h3ad895b0),
	.w6(32'hb974fb5b),
	.w7(32'hbb46269a),
	.w8(32'hbbd37af1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8e556),
	.w1(32'hba8f70fe),
	.w2(32'h3b6e63b5),
	.w3(32'hbb7c1cba),
	.w4(32'hbb2b33e8),
	.w5(32'hba92e206),
	.w6(32'hbb411449),
	.w7(32'h3b6340e9),
	.w8(32'h3acdf1c4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcde5f2),
	.w1(32'hbbc128fa),
	.w2(32'hbb9534de),
	.w3(32'hbba9927a),
	.w4(32'hbbad247e),
	.w5(32'hbb8b5074),
	.w6(32'hbb50a47e),
	.w7(32'hbb2ccca2),
	.w8(32'hbb433b96),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89db7b),
	.w1(32'hbb94d5b1),
	.w2(32'hbba7f221),
	.w3(32'hbba875f8),
	.w4(32'hbbdddbad),
	.w5(32'hbc118196),
	.w6(32'h39ff28fd),
	.w7(32'h3a7b40b1),
	.w8(32'h3b847422),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be10802),
	.w1(32'h3c21525b),
	.w2(32'h3b7a44c6),
	.w3(32'h3c261fb6),
	.w4(32'h3c84e173),
	.w5(32'h3c292811),
	.w6(32'h3b97a127),
	.w7(32'hbb825afc),
	.w8(32'hbb17bcaa),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d638bd),
	.w1(32'hbbacfd13),
	.w2(32'hb80d8efd),
	.w3(32'h39d342b9),
	.w4(32'hbbc5dba9),
	.w5(32'hbb715256),
	.w6(32'h3b6b499c),
	.w7(32'h3bccd751),
	.w8(32'h3b371de8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f9481),
	.w1(32'hba3f0791),
	.w2(32'hbb2d3bcd),
	.w3(32'hbae30012),
	.w4(32'hbb630a48),
	.w5(32'hbb135579),
	.w6(32'h3b5d38b9),
	.w7(32'h3aeee6df),
	.w8(32'h3aa3fbe2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2033d1),
	.w1(32'hbaf220bd),
	.w2(32'hbaafac55),
	.w3(32'h3b21a3ee),
	.w4(32'hbb2d21d5),
	.w5(32'hbb5e0bcb),
	.w6(32'hbb079707),
	.w7(32'hbac3bc22),
	.w8(32'hbae2d488),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9115c5),
	.w1(32'hbb75a34c),
	.w2(32'hbb818b08),
	.w3(32'hba407e5a),
	.w4(32'hbb3c28a5),
	.w5(32'hbb569025),
	.w6(32'hbb80c354),
	.w7(32'hbb86acf2),
	.w8(32'hba8b7a18),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147171),
	.w1(32'h3bad57cb),
	.w2(32'h3a02192b),
	.w3(32'hba2ddb58),
	.w4(32'h3ad67032),
	.w5(32'hb9bd0df3),
	.w6(32'h3b284fad),
	.w7(32'hbb7dc0a9),
	.w8(32'hbacadfb7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3465d),
	.w1(32'hbbdf3f18),
	.w2(32'hbbb475b5),
	.w3(32'hbb5c451a),
	.w4(32'hbb8fbd3f),
	.w5(32'hbb88cd94),
	.w6(32'hbba05d63),
	.w7(32'hbb9867ae),
	.w8(32'h3b295c8a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c2c2),
	.w1(32'h3a86451c),
	.w2(32'h3b1a1c01),
	.w3(32'h3c232342),
	.w4(32'h3b745662),
	.w5(32'h3b099087),
	.w6(32'h3ab0f845),
	.w7(32'h3ae6b716),
	.w8(32'hba144d46),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41aa23),
	.w1(32'h3b071bf9),
	.w2(32'hbad3625b),
	.w3(32'hbb155180),
	.w4(32'h39889e92),
	.w5(32'hba623dff),
	.w6(32'h3a6a3a62),
	.w7(32'hb920a35b),
	.w8(32'hb9e9fa30),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97ab5f),
	.w1(32'h3a4bcaaa),
	.w2(32'h3999a6be),
	.w3(32'hbb10ab8a),
	.w4(32'h39c227fc),
	.w5(32'hb8955b99),
	.w6(32'hb970e01d),
	.w7(32'hba6c6053),
	.w8(32'hb99d42d6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a3c15),
	.w1(32'h3b3877d8),
	.w2(32'h3ad9475c),
	.w3(32'h3b9def1d),
	.w4(32'h3a4d22bb),
	.w5(32'hb888d3d4),
	.w6(32'h3bb4b5e8),
	.w7(32'h3b4e2e69),
	.w8(32'h3b226a85),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf40916),
	.w1(32'hbb39b965),
	.w2(32'hb985726e),
	.w3(32'hb9b735b4),
	.w4(32'hbb02eb87),
	.w5(32'hba018ff9),
	.w6(32'h3920bbfe),
	.w7(32'hb9afbd49),
	.w8(32'h3b0c3bb7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb088cac),
	.w1(32'hbb0afcc1),
	.w2(32'hba40a5f9),
	.w3(32'h391a7755),
	.w4(32'hbaa94a7d),
	.w5(32'hb9d8a9c7),
	.w6(32'h3a9ebbc2),
	.w7(32'h3a7fd31f),
	.w8(32'h3af66c54),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f93d4),
	.w1(32'h3910b233),
	.w2(32'h3985daa3),
	.w3(32'hba142c4c),
	.w4(32'h39d9a175),
	.w5(32'hb8196ddd),
	.w6(32'hbad59c97),
	.w7(32'hbaad46a3),
	.w8(32'hbabb2b78),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cb442),
	.w1(32'hbb45faf8),
	.w2(32'hbb033f15),
	.w3(32'hba76c640),
	.w4(32'h3a57b565),
	.w5(32'h39b9c6cd),
	.w6(32'h3a5116c1),
	.w7(32'h3b12766e),
	.w8(32'h3b19725f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba348ecb),
	.w1(32'h39692ad1),
	.w2(32'hb99282cf),
	.w3(32'h3a02ed0e),
	.w4(32'h3b62d80e),
	.w5(32'h3b9ab753),
	.w6(32'hb9c7c2f4),
	.w7(32'h3ae92c9d),
	.w8(32'h3b6c6dc4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee7aa0),
	.w1(32'h3a098598),
	.w2(32'h3aca9898),
	.w3(32'hba10750d),
	.w4(32'h3ac1e247),
	.w5(32'h3b08fbff),
	.w6(32'h394c0564),
	.w7(32'h3af6c9f2),
	.w8(32'h3b0f3eac),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390fbc4c),
	.w1(32'hbaabb5be),
	.w2(32'h395466e2),
	.w3(32'hba9cba0c),
	.w4(32'hba452f45),
	.w5(32'hbaca1f23),
	.w6(32'hba43e1e4),
	.w7(32'hba347716),
	.w8(32'hbade0c1e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b816d5),
	.w1(32'h3627bf45),
	.w2(32'hb899edf5),
	.w3(32'hb8bacc56),
	.w4(32'hb8fc9eff),
	.w5(32'hb9961d9a),
	.w6(32'hb91a1859),
	.w7(32'hb9ae17f1),
	.w8(32'hba0db47a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81dc32c),
	.w1(32'hb9422445),
	.w2(32'hb8f12c06),
	.w3(32'hb9021801),
	.w4(32'hb9c88c46),
	.w5(32'hb9875875),
	.w6(32'hb832de6b),
	.w7(32'hb8e00ee7),
	.w8(32'hb8d2de61),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e728a),
	.w1(32'h3ad87e75),
	.w2(32'h3acb1932),
	.w3(32'h3b07cddb),
	.w4(32'h3b202567),
	.w5(32'h3afeee8d),
	.w6(32'h3aefaa24),
	.w7(32'h3b10f935),
	.w8(32'h3a170481),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dd11f0),
	.w1(32'hb8a0bca2),
	.w2(32'hb98552a0),
	.w3(32'hb9febcf1),
	.w4(32'h3a5183e0),
	.w5(32'h39c4a4d1),
	.w6(32'hba030c33),
	.w7(32'hb9eff7d3),
	.w8(32'hb9f776c9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bee197),
	.w1(32'hb8fa2592),
	.w2(32'hb918357a),
	.w3(32'hba344142),
	.w4(32'hb9e4b3bb),
	.w5(32'hb988bc98),
	.w6(32'hba057119),
	.w7(32'hb9b0d0d6),
	.w8(32'hb9755dde),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38000883),
	.w1(32'h36f70522),
	.w2(32'h35c7a580),
	.w3(32'h37f9e3fe),
	.w4(32'h373ae678),
	.w5(32'hb407f55c),
	.w6(32'h37af109d),
	.w7(32'h362a0169),
	.w8(32'hb726dfae),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373146e9),
	.w1(32'hb898bb5b),
	.w2(32'hb8e3d0c7),
	.w3(32'hb7c62c8e),
	.w4(32'hb813c965),
	.w5(32'hb83476ff),
	.w6(32'hb78b9df8),
	.w7(32'hb7c59fb3),
	.w8(32'hb80a92b2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1b9f8),
	.w1(32'h39598555),
	.w2(32'hb96c9df3),
	.w3(32'h3aaf70c1),
	.w4(32'h39f43995),
	.w5(32'hb9dddd1f),
	.w6(32'h3a85a00a),
	.w7(32'h39a8d450),
	.w8(32'hba0e0a30),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c2f70),
	.w1(32'h3aa353e4),
	.w2(32'h396021e2),
	.w3(32'h3aa8b40e),
	.w4(32'h3ad1fffd),
	.w5(32'h3a6af250),
	.w6(32'h3a4cce00),
	.w7(32'h3ad99010),
	.w8(32'h3a581064),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a582f),
	.w1(32'h3a2af3a7),
	.w2(32'h3a0c9456),
	.w3(32'h376c17fe),
	.w4(32'h37f32b3d),
	.w5(32'h39cc9775),
	.w6(32'hb9122bce),
	.w7(32'hba3db376),
	.w8(32'hbab2c4db),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e8fae),
	.w1(32'h3acfed99),
	.w2(32'h3aabee87),
	.w3(32'h399b0773),
	.w4(32'h3aab7095),
	.w5(32'h39c796d3),
	.w6(32'hba5492d4),
	.w7(32'hba882f30),
	.w8(32'hbae26daa),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01253e),
	.w1(32'hba7b892d),
	.w2(32'hba1a5dc9),
	.w3(32'hba8ae3ea),
	.w4(32'hba47e0a7),
	.w5(32'hb9e0c245),
	.w6(32'hba264da6),
	.w7(32'h3994e59a),
	.w8(32'h393369c1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01f345),
	.w1(32'hba84a3de),
	.w2(32'hba0e8a15),
	.w3(32'hbb2950dc),
	.w4(32'hbae60a3a),
	.w5(32'hba932c11),
	.w6(32'hbb434604),
	.w7(32'hbb09f111),
	.w8(32'hbaf72e99),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad89938),
	.w1(32'h3ad60191),
	.w2(32'h3a910ac5),
	.w3(32'h3aca9edd),
	.w4(32'h3b0ed5c6),
	.w5(32'h3ae8ffe4),
	.w6(32'h3ac52f6a),
	.w7(32'h3afca3f3),
	.w8(32'h3af9fa30),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997d84c),
	.w1(32'h39bf2de7),
	.w2(32'h3a693065),
	.w3(32'h39d2bd47),
	.w4(32'h3963f8a0),
	.w5(32'h3a447ee6),
	.w6(32'h3946877d),
	.w7(32'hb991546e),
	.w8(32'h3a1ec0d3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule