module layer_10_featuremap_291(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c1bb3a),
	.w1(32'hb99b8c4a),
	.w2(32'hb927c877),
	.w3(32'h3a0dfc03),
	.w4(32'h39d2c0a8),
	.w5(32'hba807df9),
	.w6(32'hb88a8ca0),
	.w7(32'hb9311bf7),
	.w8(32'hbaf98579),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf98867),
	.w1(32'hbaf48a4a),
	.w2(32'hbabde94f),
	.w3(32'hbae8a06f),
	.w4(32'hbb018fe4),
	.w5(32'h3aee5f85),
	.w6(32'hbb07a448),
	.w7(32'hbb0bc373),
	.w8(32'h3a15cf53),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927628b),
	.w1(32'hba3afb3b),
	.w2(32'hbaaf1292),
	.w3(32'h3a9fe432),
	.w4(32'h3a849d0c),
	.w5(32'h3a2133e6),
	.w6(32'h39e1bb77),
	.w7(32'hba3af2c2),
	.w8(32'h39c593fd),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bb31f),
	.w1(32'hb8d4076e),
	.w2(32'h381412c2),
	.w3(32'h39e40834),
	.w4(32'h3a0b07be),
	.w5(32'h3a8bd6d7),
	.w6(32'h379a8ece),
	.w7(32'h3940398d),
	.w8(32'h3a860f17),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02b2fe),
	.w1(32'h3a5be933),
	.w2(32'hb9ee3f1f),
	.w3(32'h3ac58022),
	.w4(32'h39c10cb6),
	.w5(32'h3a9c6836),
	.w6(32'h3aceb18c),
	.w7(32'h3989d3bd),
	.w8(32'h3a5e16e4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f7155),
	.w1(32'h3a1c3d53),
	.w2(32'h39912e43),
	.w3(32'h3a9b8509),
	.w4(32'h3a3225bd),
	.w5(32'h3ae226cf),
	.w6(32'h3a2cbfec),
	.w7(32'h39417686),
	.w8(32'h3ad616ac),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaabdd0),
	.w1(32'h3ac3d692),
	.w2(32'h3a782426),
	.w3(32'h3aff9c4a),
	.w4(32'h3aa7c2d1),
	.w5(32'h3aa81d3c),
	.w6(32'h3b14882b),
	.w7(32'h3ab9021c),
	.w8(32'h3a3581cc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7307b),
	.w1(32'h39e03557),
	.w2(32'h38034bd4),
	.w3(32'h3b01dc1f),
	.w4(32'h3a9033fa),
	.w5(32'h3a94cea7),
	.w6(32'h3a93d10e),
	.w7(32'h3a59795c),
	.w8(32'h3ab14338),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5d253),
	.w1(32'h3adb3e71),
	.w2(32'h3adfebbe),
	.w3(32'h3afdc989),
	.w4(32'h3ae7e81c),
	.w5(32'h3a97a652),
	.w6(32'h3adcb15e),
	.w7(32'h3aeab7d9),
	.w8(32'h3a837a30),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a9132),
	.w1(32'hb89eb107),
	.w2(32'hba8c7e70),
	.w3(32'h3ab27e48),
	.w4(32'h39b960e1),
	.w5(32'hb9b6a772),
	.w6(32'h3a665d6c),
	.w7(32'h379631a7),
	.w8(32'h39d38f30),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5fbc7),
	.w1(32'h39f48aa9),
	.w2(32'h3a0a9f56),
	.w3(32'h3a550dbe),
	.w4(32'h39aaea79),
	.w5(32'hbb2a0f0d),
	.w6(32'h3a3dd40f),
	.w7(32'h3937d000),
	.w8(32'hba85a563),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba367b8a),
	.w1(32'h3a667ed8),
	.w2(32'h3a2b43eb),
	.w3(32'hbb1f1305),
	.w4(32'hbae952dc),
	.w5(32'h375c073a),
	.w6(32'h39b6aa56),
	.w7(32'h3a046a73),
	.w8(32'h39bbbae1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5823fe),
	.w1(32'h39a8b832),
	.w2(32'hbad64e08),
	.w3(32'hb99d6976),
	.w4(32'hbad42b9d),
	.w5(32'hb9a3b5fc),
	.w6(32'h3a116590),
	.w7(32'hb9f07bf8),
	.w8(32'h39ade548),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c9215),
	.w1(32'h399edeec),
	.w2(32'h3a104bf8),
	.w3(32'h3a854832),
	.w4(32'h39d9f85e),
	.w5(32'hbac2ec48),
	.w6(32'h3a2a0b0b),
	.w7(32'h39e42c1c),
	.w8(32'hbaae24ea),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cae77),
	.w1(32'hbaa152e8),
	.w2(32'hbac94dfd),
	.w3(32'hbaaf333d),
	.w4(32'hbacc92c7),
	.w5(32'hba70ae53),
	.w6(32'hbac5a87d),
	.w7(32'hbae51173),
	.w8(32'hba43b542),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9336ca7),
	.w1(32'hb97740cc),
	.w2(32'hbadacd2f),
	.w3(32'hb91ee04b),
	.w4(32'hbad42cf5),
	.w5(32'h398c09a2),
	.w6(32'h385aaa51),
	.w7(32'hbaf72afa),
	.w8(32'h39adb859),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990683a),
	.w1(32'h3937c544),
	.w2(32'h39bd050d),
	.w3(32'h3a74eccf),
	.w4(32'h3a156348),
	.w5(32'hba01111d),
	.w6(32'h3a639a0d),
	.w7(32'h3a23fc5d),
	.w8(32'hb9a1a7a4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba258ccc),
	.w1(32'hbaad4d06),
	.w2(32'hbb1f45b5),
	.w3(32'hba5dd2f5),
	.w4(32'hbacbbee5),
	.w5(32'hb9eb2d9f),
	.w6(32'hb9c74a94),
	.w7(32'hba8c7fb8),
	.w8(32'h3797dfba),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bdd7b),
	.w1(32'hba8a1ab0),
	.w2(32'hbb09c44f),
	.w3(32'hb9438e11),
	.w4(32'hba6c8821),
	.w5(32'h390f045f),
	.w6(32'hba05e5d1),
	.w7(32'hbabd1579),
	.w8(32'h39f57f5d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fef19),
	.w1(32'hb95a0ed1),
	.w2(32'hbaacbaa4),
	.w3(32'hba3b18cd),
	.w4(32'hbae3ba4f),
	.w5(32'h39cc4d45),
	.w6(32'hb7a8e459),
	.w7(32'hbaa0f2f7),
	.w8(32'h399ba964),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a751eb6),
	.w1(32'h3a476a23),
	.w2(32'hb9f76cc0),
	.w3(32'h39a5e417),
	.w4(32'hba3969ca),
	.w5(32'h3aaf89e1),
	.w6(32'h39e0dccc),
	.w7(32'hba4e3598),
	.w8(32'h3aaa7e09),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96d3e3),
	.w1(32'h3a80f788),
	.w2(32'h3abfd33c),
	.w3(32'h3a964575),
	.w4(32'h3ac93f49),
	.w5(32'h3ad0bed6),
	.w6(32'h3a496597),
	.w7(32'h3ab185e9),
	.w8(32'h3a915da8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25206f),
	.w1(32'h3a4cf962),
	.w2(32'h3a0a0e26),
	.w3(32'h3b1e3027),
	.w4(32'h3aaf427a),
	.w5(32'hb9c8952d),
	.w6(32'h3b022fd9),
	.w7(32'h3ab32854),
	.w8(32'h397f306b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c17cd),
	.w1(32'hbad70070),
	.w2(32'hbb04bc59),
	.w3(32'hb9a60bdb),
	.w4(32'hbaf9ee65),
	.w5(32'h3a6843df),
	.w6(32'hba1f9df6),
	.w7(32'hbaf1f52e),
	.w8(32'h3adee26e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86e265f),
	.w1(32'h38a10b43),
	.w2(32'hb9148f99),
	.w3(32'h3b073ff5),
	.w4(32'h3b2d8ba8),
	.w5(32'hba700627),
	.w6(32'h3ad78d8c),
	.w7(32'h3adc75f4),
	.w8(32'hba232c35),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63d34d),
	.w1(32'h38f20b30),
	.w2(32'hba0f812e),
	.w3(32'h3a088bbe),
	.w4(32'hb9518a6f),
	.w5(32'hbaa34d7b),
	.w6(32'h3a9ce551),
	.w7(32'h39a0cd7e),
	.w8(32'hbabfd11b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6cf40),
	.w1(32'hba62f601),
	.w2(32'hba5c101f),
	.w3(32'hba417594),
	.w4(32'hba332a18),
	.w5(32'h3a109b64),
	.w6(32'hba88afec),
	.w7(32'hba7bebd3),
	.w8(32'h393ae5a9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996524d),
	.w1(32'h39eea265),
	.w2(32'h39e7ee00),
	.w3(32'h39b1ea1e),
	.w4(32'h3a02b933),
	.w5(32'h3b1ea4b5),
	.w6(32'hb916f9b7),
	.w7(32'h3901675e),
	.w8(32'h3aed3106),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb7d29),
	.w1(32'h3b3445bb),
	.w2(32'h3b41cd2e),
	.w3(32'h3b486525),
	.w4(32'h3b4d5c40),
	.w5(32'hba65fa5c),
	.w6(32'h3b4de65d),
	.w7(32'h3b4f6ae2),
	.w8(32'hba8341fa),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bdc40),
	.w1(32'hbaab289a),
	.w2(32'hbac85f66),
	.w3(32'hba97d9d0),
	.w4(32'hbad1596c),
	.w5(32'hba387b68),
	.w6(32'hba48585c),
	.w7(32'hba8154ea),
	.w8(32'hb89b1bb4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c76a95),
	.w1(32'h3a3b8cfc),
	.w2(32'h3a85c5be),
	.w3(32'hb93ea19a),
	.w4(32'h3a125435),
	.w5(32'h39aff12b),
	.w6(32'h39d2582a),
	.w7(32'h38b2ec2a),
	.w8(32'hb8de67d8),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07daca),
	.w1(32'hb994f9fd),
	.w2(32'hb88cd131),
	.w3(32'h39d8beda),
	.w4(32'h3a21fec7),
	.w5(32'h3a11e1d3),
	.w6(32'h3a196d04),
	.w7(32'h3a029d96),
	.w8(32'h3abb58bf),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa72c9b),
	.w1(32'h3a64395d),
	.w2(32'hbaa77f15),
	.w3(32'h3ad09930),
	.w4(32'h39959b72),
	.w5(32'hba941366),
	.w6(32'h3b1a21a2),
	.w7(32'hb8a117d8),
	.w8(32'hba085d0d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e8273),
	.w1(32'hb8a33523),
	.w2(32'h38aab569),
	.w3(32'hba10dd2b),
	.w4(32'hba0e865c),
	.w5(32'hba518253),
	.w6(32'h391e977a),
	.w7(32'h38461317),
	.w8(32'hba37b948),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a8ad7),
	.w1(32'hba6171d7),
	.w2(32'hba2b19ae),
	.w3(32'hba9cc30b),
	.w4(32'hb9dd427a),
	.w5(32'h3a7f01cd),
	.w6(32'hbaa6d046),
	.w7(32'hba4b2919),
	.w8(32'h3aa87993),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d4732),
	.w1(32'h3a0cfd18),
	.w2(32'hbaa63cec),
	.w3(32'h3a902ada),
	.w4(32'hb997b777),
	.w5(32'hb9b3b5c0),
	.w6(32'h3af9048a),
	.w7(32'hb9b5c78d),
	.w8(32'h39ce22ee),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05af7c),
	.w1(32'h39a43f09),
	.w2(32'hb9d69bd9),
	.w3(32'h3a70c70d),
	.w4(32'h3aa1dd82),
	.w5(32'hba9e1076),
	.w6(32'h3b186be7),
	.w7(32'h3a9a84fa),
	.w8(32'hba730f6d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0f347),
	.w1(32'h3946cc06),
	.w2(32'h38ecee8b),
	.w3(32'hbab5afe9),
	.w4(32'hba5011f4),
	.w5(32'h3786cd16),
	.w6(32'hbab00f73),
	.w7(32'hbb032b92),
	.w8(32'hbb18487f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af944),
	.w1(32'hbadf3b5a),
	.w2(32'hb9b805a5),
	.w3(32'hbb0fb879),
	.w4(32'hba81f0c0),
	.w5(32'hb97c0c46),
	.w6(32'hbb2bde3d),
	.w7(32'hbb1e3dd0),
	.w8(32'hbab3845f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87e483),
	.w1(32'hbb09d2ef),
	.w2(32'hbb01001e),
	.w3(32'hba939011),
	.w4(32'hbac4bf81),
	.w5(32'hb972f520),
	.w6(32'hbae97c6e),
	.w7(32'hbb033b01),
	.w8(32'hb8d3b494),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e96ff4),
	.w1(32'h3acb15bd),
	.w2(32'h3b16a28d),
	.w3(32'h3a58f06c),
	.w4(32'h3aed35ec),
	.w5(32'h39966d6c),
	.w6(32'h3a6b414c),
	.w7(32'h3b17c4a6),
	.w8(32'h39fefb2d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9becf03),
	.w1(32'h39f3844d),
	.w2(32'h38e312f7),
	.w3(32'h3a84a1d1),
	.w4(32'h39f94eb0),
	.w5(32'hba905f3a),
	.w6(32'h3abc1860),
	.w7(32'h3a766bb5),
	.w8(32'hba9488d7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f5b73),
	.w1(32'hba129738),
	.w2(32'hba4f287c),
	.w3(32'hbaa72b04),
	.w4(32'hba7cc6dc),
	.w5(32'hbb0d9579),
	.w6(32'hba909de1),
	.w7(32'hba879ca6),
	.w8(32'hbb6453dc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e831b),
	.w1(32'hbb7cee48),
	.w2(32'hbb65abb1),
	.w3(32'hbb15a8c0),
	.w4(32'hbb43f612),
	.w5(32'hb9c0c984),
	.w6(32'hbb55c0b6),
	.w7(32'hbb51523d),
	.w8(32'hb97756f1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30f02c),
	.w1(32'hba752786),
	.w2(32'hba378619),
	.w3(32'h398923be),
	.w4(32'h394e43a7),
	.w5(32'hba30f34b),
	.w6(32'hba49a179),
	.w7(32'hb91210bf),
	.w8(32'hb9c08478),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa2215),
	.w1(32'hbad192e4),
	.w2(32'hbabbcab8),
	.w3(32'h39042fd7),
	.w4(32'h38578be8),
	.w5(32'hbb371707),
	.w6(32'hba22e529),
	.w7(32'hb90836fb),
	.w8(32'hbb08ca8a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170e1e),
	.w1(32'hbae1fbf1),
	.w2(32'hbaa43501),
	.w3(32'hbb007af7),
	.w4(32'hbab6a05e),
	.w5(32'h39fd6907),
	.w6(32'hbb097e89),
	.w7(32'hbaa53c03),
	.w8(32'h3a6be990),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8aba6f),
	.w1(32'h39c390f9),
	.w2(32'hb90a46e9),
	.w3(32'h3ae206df),
	.w4(32'h3aaa69b4),
	.w5(32'hbad5cbf8),
	.w6(32'h3a6c536c),
	.w7(32'h3ab0751e),
	.w8(32'hb9bdb30c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389436af),
	.w1(32'hb64795c9),
	.w2(32'hbaa71fa9),
	.w3(32'hba5b5cec),
	.w4(32'hbac7088a),
	.w5(32'h3a893ec9),
	.w6(32'hb9719400),
	.w7(32'hbab528db),
	.w8(32'h3a93f4b4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7545d1),
	.w1(32'h3a5b264d),
	.w2(32'h3a6e9eef),
	.w3(32'h3a91a7bf),
	.w4(32'h3a8e20fc),
	.w5(32'h3a03766b),
	.w6(32'h3a92ba39),
	.w7(32'h3a7cea8f),
	.w8(32'h39cf9d77),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17215b),
	.w1(32'h3867e33b),
	.w2(32'hbae62a7f),
	.w3(32'h390fc16c),
	.w4(32'hba8b657c),
	.w5(32'hb97a9120),
	.w6(32'hba2b176d),
	.w7(32'hbab89b32),
	.w8(32'h3956286b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba02bb),
	.w1(32'h3954d3ea),
	.w2(32'hba8241ad),
	.w3(32'hba0d0a46),
	.w4(32'hbae4e19a),
	.w5(32'hba55854f),
	.w6(32'h37e847b7),
	.w7(32'hba916215),
	.w8(32'h3a6f1e20),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bb834),
	.w1(32'h3b07f289),
	.w2(32'h3acf6f85),
	.w3(32'h3a03e568),
	.w4(32'h3a0d7df8),
	.w5(32'hb9ac69af),
	.w6(32'h3b17c226),
	.w7(32'h3ace6a04),
	.w8(32'h3992e3d5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f56792),
	.w1(32'hb9912e41),
	.w2(32'hbac6211d),
	.w3(32'h39f972cb),
	.w4(32'hba374d75),
	.w5(32'h3a11325c),
	.w6(32'h3ab73d7b),
	.w7(32'h3a291444),
	.w8(32'h3b426f69),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3abbff),
	.w1(32'h3b219e6c),
	.w2(32'h3a85fe32),
	.w3(32'hb7dad73e),
	.w4(32'hbadb68e5),
	.w5(32'hba3d84a4),
	.w6(32'h3b1c1718),
	.w7(32'h399eae68),
	.w8(32'hbb05121b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb430311),
	.w1(32'hbaa1aceb),
	.w2(32'hb9fb89c4),
	.w3(32'h3a47655b),
	.w4(32'h3aac7234),
	.w5(32'hba3ef7fb),
	.w6(32'h380d08fe),
	.w7(32'h39e05f4b),
	.w8(32'hba312d11),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6133f1),
	.w1(32'h379d4672),
	.w2(32'h3a9a8f60),
	.w3(32'h38b4616b),
	.w4(32'h3aab4cae),
	.w5(32'hb9f2a7e7),
	.w6(32'hb9692536),
	.w7(32'h3ab5465d),
	.w8(32'hb95c751a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afb763),
	.w1(32'hb9cdd7a5),
	.w2(32'hba64eb9e),
	.w3(32'hba42e655),
	.w4(32'hbac51b8e),
	.w5(32'h3ad27e08),
	.w6(32'h393371e1),
	.w7(32'hbaa21a7b),
	.w8(32'h3ae1bb5e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9f774),
	.w1(32'h3adae72a),
	.w2(32'h3aacbcc9),
	.w3(32'h3b07afaf),
	.w4(32'h3ae19d1f),
	.w5(32'h397564d9),
	.w6(32'h3b131e6c),
	.w7(32'h3aed04be),
	.w8(32'h395d6dc9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d5b6c),
	.w1(32'hba3fb021),
	.w2(32'h383e96eb),
	.w3(32'h3907b137),
	.w4(32'h3a5b6cf4),
	.w5(32'hba11d28b),
	.w6(32'h39ee1908),
	.w7(32'h3a76efa0),
	.w8(32'hba927cd7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba690d12),
	.w1(32'hbad3035c),
	.w2(32'hbacfb75b),
	.w3(32'hb8a6e2f7),
	.w4(32'h39d5c046),
	.w5(32'h39a4b882),
	.w6(32'hbaae7d38),
	.w7(32'hba475c09),
	.w8(32'h39c466a8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957db6e),
	.w1(32'hb970e6d9),
	.w2(32'hb991270a),
	.w3(32'h3a46bfc9),
	.w4(32'h3a27615b),
	.w5(32'hbac9937e),
	.w6(32'h3a8ede59),
	.w7(32'h3a75abbe),
	.w8(32'hba8a2ef7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b9a55),
	.w1(32'hba139237),
	.w2(32'hba4415c6),
	.w3(32'hbb1b5779),
	.w4(32'hbb039703),
	.w5(32'hba270839),
	.w6(32'hbaaa00c1),
	.w7(32'hbaac04d2),
	.w8(32'hba2a8540),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36002d),
	.w1(32'h384f9b2b),
	.w2(32'h3a847ed8),
	.w3(32'h39ab7e4d),
	.w4(32'h3aa1949e),
	.w5(32'h39676977),
	.w6(32'h398f326a),
	.w7(32'h3ab51e2d),
	.w8(32'h3a6bbb31),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba552a),
	.w1(32'h39541fab),
	.w2(32'hb9e65e02),
	.w3(32'hba7ad7ec),
	.w4(32'hbae59fdf),
	.w5(32'hb568f919),
	.w6(32'h39dfb3b8),
	.w7(32'hba476fa2),
	.w8(32'h3ad78431),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf0d74),
	.w1(32'h3b11fa84),
	.w2(32'h3b0201aa),
	.w3(32'hb99d59cc),
	.w4(32'hba2f9258),
	.w5(32'h3a4a7ab9),
	.w6(32'h3b260277),
	.w7(32'h3ae7e537),
	.w8(32'h3a23f0a1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53a215),
	.w1(32'h398c23f4),
	.w2(32'hb9b5c762),
	.w3(32'h39757a29),
	.w4(32'hb82bfafd),
	.w5(32'hbacde729),
	.w6(32'h3a29c7eb),
	.w7(32'h391506e1),
	.w8(32'hbab43f83),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ad325),
	.w1(32'hb9c18e95),
	.w2(32'hba24311b),
	.w3(32'hb9004a97),
	.w4(32'hb9801c88),
	.w5(32'h3b35d313),
	.w6(32'hba086aa2),
	.w7(32'hb9dd251e),
	.w8(32'h3b8d564f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b755b5d),
	.w1(32'h3b97ee71),
	.w2(32'h3abe027f),
	.w3(32'h3b544c0d),
	.w4(32'h3a645169),
	.w5(32'h3a0ad7b7),
	.w6(32'h3ba1a97f),
	.w7(32'h3adbc630),
	.w8(32'h395a7879),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89cd761),
	.w1(32'hba1bf3a9),
	.w2(32'hbade1d72),
	.w3(32'hba6d3186),
	.w4(32'hbad9ae84),
	.w5(32'hba0facc6),
	.w6(32'hba9ac423),
	.w7(32'hbb07bd52),
	.w8(32'hb9ed4210),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e77552),
	.w1(32'hb9c76d8c),
	.w2(32'hb9447f02),
	.w3(32'hb91bb721),
	.w4(32'hb8a3b033),
	.w5(32'hb9cf2c33),
	.w6(32'hb9f4bcb6),
	.w7(32'hb96ece42),
	.w8(32'hba0a1954),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990f724),
	.w1(32'hb98fd13e),
	.w2(32'hbab0b706),
	.w3(32'h39d82d0d),
	.w4(32'hba0502db),
	.w5(32'hba4c9a7b),
	.w6(32'h39d50a6d),
	.w7(32'hba8a09b3),
	.w8(32'h39029f59),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cdc84),
	.w1(32'hbae7e680),
	.w2(32'hbafcb07c),
	.w3(32'hba8014aa),
	.w4(32'hba7a173a),
	.w5(32'hba60ba2d),
	.w6(32'h3a185818),
	.w7(32'h388ba8ea),
	.w8(32'hba079aa3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78689b),
	.w1(32'hba85e672),
	.w2(32'hbae93e4d),
	.w3(32'hbb017637),
	.w4(32'hbb2ae557),
	.w5(32'h39d0b488),
	.w6(32'hba4b306b),
	.w7(32'hbad0c516),
	.w8(32'h39c981bd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df3bd1),
	.w1(32'hb972a3c4),
	.w2(32'hb7d0b594),
	.w3(32'hb8769423),
	.w4(32'hb907a188),
	.w5(32'hbb16861a),
	.w6(32'hb9abb341),
	.w7(32'hba0e503d),
	.w8(32'hbaddb0c0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5a2c2),
	.w1(32'hbabcc02b),
	.w2(32'hbb24e677),
	.w3(32'hbb0f4e81),
	.w4(32'hbb42d5da),
	.w5(32'hbac0a184),
	.w6(32'hba9a3df7),
	.w7(32'hbaf4f97c),
	.w8(32'hbaa4337b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907ee80),
	.w1(32'hba847e80),
	.w2(32'hb99cf639),
	.w3(32'h38ecc0db),
	.w4(32'h39069189),
	.w5(32'hba40723c),
	.w6(32'hba616752),
	.w7(32'h3927fcee),
	.w8(32'hba3f9f23),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c6cfa2),
	.w1(32'h3695dc6b),
	.w2(32'hba398347),
	.w3(32'hb920305b),
	.w4(32'hba5d00bb),
	.w5(32'hbac1262b),
	.w6(32'hb9fbb4fb),
	.w7(32'hba713cab),
	.w8(32'hba49915b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73246c),
	.w1(32'hba495d0e),
	.w2(32'hba91dea0),
	.w3(32'hba471558),
	.w4(32'hba457b60),
	.w5(32'h3a8f0cc5),
	.w6(32'hba3dcb78),
	.w7(32'hba1c796e),
	.w8(32'h3a282cc0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a516a51),
	.w1(32'h3a2a94b4),
	.w2(32'h3934b349),
	.w3(32'h3aca516c),
	.w4(32'h3a993d05),
	.w5(32'hbb3f26d4),
	.w6(32'h3a9643b1),
	.w7(32'h3a2793e8),
	.w8(32'hbb37367d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0812a6),
	.w1(32'hbaeea411),
	.w2(32'hbabc75b3),
	.w3(32'hbb081b1e),
	.w4(32'hbb040666),
	.w5(32'hba4d0550),
	.w6(32'hbb198c92),
	.w7(32'hbae851a1),
	.w8(32'hb93875e0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49da57),
	.w1(32'hba1df518),
	.w2(32'hbb1c475d),
	.w3(32'hb9fcc5ec),
	.w4(32'hbac7f291),
	.w5(32'h3b02b315),
	.w6(32'h39999e98),
	.w7(32'hba966dc4),
	.w8(32'h3aa0625e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72ac9d),
	.w1(32'h3a0550b2),
	.w2(32'h39c78eff),
	.w3(32'h3af9e538),
	.w4(32'h3ac4f21c),
	.w5(32'h39494bfd),
	.w6(32'h3aaaaf77),
	.w7(32'h39fdc467),
	.w8(32'h3881721b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb857a783),
	.w1(32'hba235e5d),
	.w2(32'hb9e47c45),
	.w3(32'hba0c8503),
	.w4(32'hb9d41f77),
	.w5(32'h3b453402),
	.w6(32'hba2b33f1),
	.w7(32'hba591c91),
	.w8(32'h3ab09d85),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dfc5d),
	.w1(32'hb901374e),
	.w2(32'hb9b2ceb8),
	.w3(32'h3b14a0d3),
	.w4(32'h3af08cd4),
	.w5(32'hb6edfcfb),
	.w6(32'h3a3a8ab2),
	.w7(32'h390e8508),
	.w8(32'hb9e28c14),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba516deb),
	.w1(32'hb9d560a7),
	.w2(32'hb759cb71),
	.w3(32'h3a036c58),
	.w4(32'h3a1106b8),
	.w5(32'hb8be8b01),
	.w6(32'h38b62bdf),
	.w7(32'h39315897),
	.w8(32'hba164c65),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c53c2),
	.w1(32'hba979015),
	.w2(32'hbb1d999e),
	.w3(32'hba4622f9),
	.w4(32'hbb06fe68),
	.w5(32'h3a04ea32),
	.w6(32'hba1a8bfe),
	.w7(32'hbb3d340e),
	.w8(32'hba6a6616),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7361f),
	.w1(32'hb9ec729c),
	.w2(32'hb9ea91fa),
	.w3(32'h3a2cff87),
	.w4(32'h39b45811),
	.w5(32'h3ac5af43),
	.w6(32'hba657424),
	.w7(32'hba91ed5e),
	.w8(32'h3a9f94b7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8393f6),
	.w1(32'h39d5861a),
	.w2(32'hb953f59f),
	.w3(32'h3ad44d09),
	.w4(32'h38e4dc08),
	.w5(32'hb9f26377),
	.w6(32'h3a7b4e46),
	.w7(32'h393dd75e),
	.w8(32'hb9fb1e00),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e322f),
	.w1(32'h392bd6bc),
	.w2(32'h387debb3),
	.w3(32'h3a60b150),
	.w4(32'h3a55215e),
	.w5(32'hb9e9b2ee),
	.w6(32'h3999c3bc),
	.w7(32'h3aaee092),
	.w8(32'h390289f6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39920359),
	.w1(32'hba8fdb5c),
	.w2(32'hba6925b8),
	.w3(32'hbb120f0e),
	.w4(32'hba730c5a),
	.w5(32'h398a0bf2),
	.w6(32'hbb07da83),
	.w7(32'hbaf42cac),
	.w8(32'h3596f2e3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986500c),
	.w1(32'hba58f9fb),
	.w2(32'hba9fe39a),
	.w3(32'hba1ab403),
	.w4(32'hba859f3a),
	.w5(32'hba74e46f),
	.w6(32'h39c92917),
	.w7(32'h3872916a),
	.w8(32'hbb14e37a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28579e),
	.w1(32'hbaff873c),
	.w2(32'hba97ea42),
	.w3(32'hb8e502fe),
	.w4(32'h39560271),
	.w5(32'hbaaf495a),
	.w6(32'hba919be0),
	.w7(32'hba9535cc),
	.w8(32'hbaccdc61),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0bd25),
	.w1(32'hbb1e43c7),
	.w2(32'hbaf3f5db),
	.w3(32'hbb179208),
	.w4(32'hbb033501),
	.w5(32'hba32478b),
	.w6(32'hbb21d634),
	.w7(32'hbb1148f1),
	.w8(32'hb984ce64),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e0f277),
	.w1(32'hba9959b6),
	.w2(32'hbada42a8),
	.w3(32'hba1b8160),
	.w4(32'hbaa48c56),
	.w5(32'hba843228),
	.w6(32'h38c0d88a),
	.w7(32'hbaa38d3e),
	.w8(32'hb9d8b3ab),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923d83a),
	.w1(32'hba67bcae),
	.w2(32'hba59510f),
	.w3(32'h3a5d9cb7),
	.w4(32'hb92b047d),
	.w5(32'hb9df7223),
	.w6(32'hb8849a0b),
	.w7(32'hba65a168),
	.w8(32'hba127516),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d75e42),
	.w1(32'hba0c809a),
	.w2(32'hb9705880),
	.w3(32'hba0b0d32),
	.w4(32'hb9d80925),
	.w5(32'hbb5b531e),
	.w6(32'hba470ce0),
	.w7(32'hb993f26c),
	.w8(32'hbb6a5cd6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb617ee3),
	.w1(32'hbb5c5218),
	.w2(32'hbad55765),
	.w3(32'hbb32679b),
	.w4(32'hbae71b92),
	.w5(32'h3a7be76f),
	.w6(32'hbb63f2b9),
	.w7(32'hbaf6c015),
	.w8(32'h3a1fb84b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1f0dd),
	.w1(32'h3b3277a6),
	.w2(32'h3b46e00e),
	.w3(32'h3b981790),
	.w4(32'h3b80d8b1),
	.w5(32'hbbb96756),
	.w6(32'h3b46301b),
	.w7(32'h3af329a7),
	.w8(32'hbb42bfb3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d79c6),
	.w1(32'hb8e423ea),
	.w2(32'hba2d8d88),
	.w3(32'hbab68338),
	.w4(32'hbb2212b5),
	.w5(32'hbbe50a7d),
	.w6(32'hba882d5b),
	.w7(32'hba8c7493),
	.w8(32'hbaf4cd4a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73eab3),
	.w1(32'h3b930c08),
	.w2(32'h3be2cd8e),
	.w3(32'hbbe4d2f2),
	.w4(32'h3a119f45),
	.w5(32'hbbc89e6e),
	.w6(32'h3b720eb5),
	.w7(32'h3bc233c8),
	.w8(32'hbb6c48ee),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d0691),
	.w1(32'hba7676f2),
	.w2(32'h3a85cdfc),
	.w3(32'hbb997f79),
	.w4(32'hbbec5fa7),
	.w5(32'h3b1fcafb),
	.w6(32'hba794a91),
	.w7(32'hbb28bd4b),
	.w8(32'h3aee7344),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e3b21),
	.w1(32'hba761a1e),
	.w2(32'h3aed1848),
	.w3(32'h3b0824fa),
	.w4(32'h3b3646f5),
	.w5(32'hbba7ff8a),
	.w6(32'h3823f127),
	.w7(32'h3b24b693),
	.w8(32'hbb26cf96),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac11872),
	.w1(32'hbb8535aa),
	.w2(32'hba205738),
	.w3(32'hbb56e3fd),
	.w4(32'hba67d0df),
	.w5(32'h3a7c5071),
	.w6(32'hbb574cb5),
	.w7(32'hb9069184),
	.w8(32'h3b9b0618),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cc2c6),
	.w1(32'h3b27125b),
	.w2(32'h3aa102c5),
	.w3(32'h3ba1862d),
	.w4(32'h3b0daeae),
	.w5(32'hbb970698),
	.w6(32'h3bfcc92d),
	.w7(32'h3bbdc8e0),
	.w8(32'hbb81e182),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb064760),
	.w1(32'hb9d6077b),
	.w2(32'h3a054bf1),
	.w3(32'hbb487d04),
	.w4(32'hbb2216dd),
	.w5(32'hba70e60a),
	.w6(32'hbb0f8637),
	.w7(32'hba49f69f),
	.w8(32'hba836648),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb946d0e),
	.w1(32'hbbbfdc04),
	.w2(32'hba141fcd),
	.w3(32'h3a7c481c),
	.w4(32'hbb233c1d),
	.w5(32'h3b21e9e3),
	.w6(32'hbb3d6473),
	.w7(32'hbb38d38a),
	.w8(32'h3bb82a63),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b713636),
	.w1(32'h3b066f52),
	.w2(32'h3a5724d2),
	.w3(32'h3b2dc61b),
	.w4(32'h3b2265eb),
	.w5(32'hba15ec2c),
	.w6(32'h3ba6f19d),
	.w7(32'h3b08c146),
	.w8(32'hba5ac6d2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b94448),
	.w1(32'h3b07045a),
	.w2(32'h3b13ec53),
	.w3(32'h3b80e6e7),
	.w4(32'h3b8d2e1f),
	.w5(32'h3bd021a1),
	.w6(32'h3aea148d),
	.w7(32'h3ae93faf),
	.w8(32'h3bda5a79),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3efab),
	.w1(32'h3c08131a),
	.w2(32'h3ba61cfe),
	.w3(32'h3c23018b),
	.w4(32'h3bce513e),
	.w5(32'hbb52f307),
	.w6(32'h3c1b145a),
	.w7(32'h3bc8fff7),
	.w8(32'hbb2e368e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402ace),
	.w1(32'h39598075),
	.w2(32'hbb0f1930),
	.w3(32'hbb3d72e9),
	.w4(32'hbb4773cc),
	.w5(32'hbae957eb),
	.w6(32'h3a163bb6),
	.w7(32'hbaff6b4f),
	.w8(32'hb9a6a0b3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba039597),
	.w1(32'hb951310f),
	.w2(32'h3b68efdb),
	.w3(32'hb9ce8b61),
	.w4(32'h37fe2253),
	.w5(32'h3ba7a798),
	.w6(32'hb92697ec),
	.w7(32'h3b389723),
	.w8(32'h3b116bb3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf90b4),
	.w1(32'hba92e584),
	.w2(32'hbb754a34),
	.w3(32'h390d8dac),
	.w4(32'hbb5bd274),
	.w5(32'hba86b398),
	.w6(32'hbb87a732),
	.w7(32'hbbb5b8de),
	.w8(32'hbb3f1b1b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace2b44),
	.w1(32'hbae0c022),
	.w2(32'hba7c1408),
	.w3(32'h3a8f3971),
	.w4(32'h39c64ffd),
	.w5(32'hbaadd38e),
	.w6(32'hba7a4bc0),
	.w7(32'hbafc7c22),
	.w8(32'hbb01d33e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ea0d6),
	.w1(32'hba073555),
	.w2(32'h3b15bef9),
	.w3(32'h3a8693f3),
	.w4(32'h3a7440f6),
	.w5(32'hbab31fc8),
	.w6(32'h3b2bf6de),
	.w7(32'h3b4c3cfa),
	.w8(32'h3982c5b3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa504c9),
	.w1(32'h3a941bf4),
	.w2(32'h3b81252f),
	.w3(32'hb934fb41),
	.w4(32'hb99b3e2f),
	.w5(32'hbb829f2a),
	.w6(32'h3b05cf9e),
	.w7(32'h3b004334),
	.w8(32'hbb5e2fcc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb147b1b),
	.w1(32'hb8e90633),
	.w2(32'h3aa77d6b),
	.w3(32'hbb5e5cc2),
	.w4(32'hba412dfe),
	.w5(32'h39cd7684),
	.w6(32'hba8dee4c),
	.w7(32'h3ac2b19e),
	.w8(32'h3aa39447),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ce337),
	.w1(32'h3b70b7f3),
	.w2(32'h3b5f59f3),
	.w3(32'h399d7ff8),
	.w4(32'hb811be5f),
	.w5(32'hb9d61bbd),
	.w6(32'hba3e83a4),
	.w7(32'h3b80cb5c),
	.w8(32'hbad0b9b4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981d6f3),
	.w1(32'h3b2b5bac),
	.w2(32'hbb34bae2),
	.w3(32'h3b7a9637),
	.w4(32'hbb40cb8d),
	.w5(32'hbb530c43),
	.w6(32'h3b065e9a),
	.w7(32'hbb53f927),
	.w8(32'hbb2d8fdd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0688a),
	.w1(32'hb9a276be),
	.w2(32'h3b68bf26),
	.w3(32'h3aa6f8f0),
	.w4(32'h3b535897),
	.w5(32'hbb02a5b6),
	.w6(32'h3a9e9d8b),
	.w7(32'h3b99aaae),
	.w8(32'hb997bf53),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a123d),
	.w1(32'hbacac4e7),
	.w2(32'h3b109e64),
	.w3(32'hb9ebe10b),
	.w4(32'h3b562742),
	.w5(32'h3b11df61),
	.w6(32'hbb0146df),
	.w7(32'h3b00f49b),
	.w8(32'h3b9bd5a1),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb18955),
	.w1(32'h3a973deb),
	.w2(32'hbb3c6e37),
	.w3(32'hbb11736a),
	.w4(32'hbb082796),
	.w5(32'h3b92fcd7),
	.w6(32'hba6d79ae),
	.w7(32'hbb24deb0),
	.w8(32'h3b308671),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24b6bb),
	.w1(32'h3997be20),
	.w2(32'hbaf88722),
	.w3(32'h3b5db85a),
	.w4(32'h3a035e0a),
	.w5(32'hba282ce1),
	.w6(32'hbad78ad8),
	.w7(32'hbbc2705d),
	.w8(32'hba2f8701),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b95bc2),
	.w1(32'hbb2151e7),
	.w2(32'hbb59c590),
	.w3(32'hbae5afbc),
	.w4(32'hba80c969),
	.w5(32'h3b7f4615),
	.w6(32'hbb1a0508),
	.w7(32'hbb354b73),
	.w8(32'h3bafea12),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f5102),
	.w1(32'h3a7f6a5d),
	.w2(32'hba75d625),
	.w3(32'h3a75d884),
	.w4(32'hba16e5bb),
	.w5(32'hbb32dc4c),
	.w6(32'h3ad7b353),
	.w7(32'hbb58fe4f),
	.w8(32'hbab8f415),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24d086),
	.w1(32'hbacc9008),
	.w2(32'hbaf6652f),
	.w3(32'hbae57d9d),
	.w4(32'h3a5003b7),
	.w5(32'h3b89500f),
	.w6(32'hbb2bdd68),
	.w7(32'hba9803b6),
	.w8(32'h3c2e3719),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eeaa8),
	.w1(32'h3a368806),
	.w2(32'hb9da50dd),
	.w3(32'h3b93579b),
	.w4(32'h3b210992),
	.w5(32'h37820cf4),
	.w6(32'h3be77bff),
	.w7(32'h3b3874b4),
	.w8(32'hb9c8f8a1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48ac43),
	.w1(32'h3a863e86),
	.w2(32'h3afc8165),
	.w3(32'hbb23f69b),
	.w4(32'hb7c41082),
	.w5(32'h3c286504),
	.w6(32'h39e9a8a0),
	.w7(32'h3b5af5a6),
	.w8(32'h3b9a9314),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2f9ec),
	.w1(32'h3b60b511),
	.w2(32'h3aa489a0),
	.w3(32'h3c096236),
	.w4(32'h3b0870ef),
	.w5(32'h3ac21b02),
	.w6(32'h3b820722),
	.w7(32'h3a75b787),
	.w8(32'h3b59e27c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ff560),
	.w1(32'hbb8723ab),
	.w2(32'hbb1def89),
	.w3(32'h3a52d134),
	.w4(32'hbafe7a25),
	.w5(32'hbb384b15),
	.w6(32'hbad2d22b),
	.w7(32'hbb312a0e),
	.w8(32'hbb365664),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22419c),
	.w1(32'h397affe6),
	.w2(32'h3ad5e5e1),
	.w3(32'h39fa00fe),
	.w4(32'hbaaee46c),
	.w5(32'hbb33684c),
	.w6(32'h3a29fce2),
	.w7(32'hbb3571e2),
	.w8(32'hbaef31ae),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1110f6),
	.w1(32'hbb311565),
	.w2(32'hbac618d7),
	.w3(32'hbb4d9dea),
	.w4(32'hbafbfc5f),
	.w5(32'hbbb360df),
	.w6(32'hbae37d6a),
	.w7(32'hbab7a9d7),
	.w8(32'h3ac22031),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ed1ca),
	.w1(32'hbaad454b),
	.w2(32'hbb896e5c),
	.w3(32'hbb867728),
	.w4(32'hbbbef5ff),
	.w5(32'hbb092bec),
	.w6(32'hbb445f7c),
	.w7(32'hbba38ca6),
	.w8(32'h3a135e45),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa54bb3),
	.w1(32'h3b22d6ab),
	.w2(32'h3b2dfff8),
	.w3(32'hb8db2841),
	.w4(32'h39deefcd),
	.w5(32'hbb43d5c6),
	.w6(32'h3aa5e673),
	.w7(32'h3ada9e06),
	.w8(32'hba1d5965),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c81cc),
	.w1(32'hbb29507c),
	.w2(32'hbb16f6bf),
	.w3(32'hbb0d1c1a),
	.w4(32'hbb3782ca),
	.w5(32'hbb8122df),
	.w6(32'h398f3057),
	.w7(32'hba99b88e),
	.w8(32'hbb7f4a21),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14acd6),
	.w1(32'hbaf5b1f2),
	.w2(32'h3936e70c),
	.w3(32'h3a8f5c01),
	.w4(32'hb9d47d48),
	.w5(32'hbadafff4),
	.w6(32'h3b46d9ea),
	.w7(32'h3b307729),
	.w8(32'hbb318c0a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc33ad),
	.w1(32'hbaa3db00),
	.w2(32'hbb6f9fc3),
	.w3(32'hbb20b927),
	.w4(32'hbb8c0acc),
	.w5(32'hb74e4e1d),
	.w6(32'hbb1f5046),
	.w7(32'hbb7c4eb9),
	.w8(32'h3b4ff0b7),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1567b9),
	.w1(32'h3b44bfb4),
	.w2(32'h3b3e9e31),
	.w3(32'h3ab78509),
	.w4(32'h3aafe747),
	.w5(32'hbb380c59),
	.w6(32'h3b3d64e6),
	.w7(32'h3b479a61),
	.w8(32'hbaaf7aa7),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad59bc0),
	.w1(32'hba90ba2c),
	.w2(32'hba060964),
	.w3(32'hbb55012e),
	.w4(32'hbb1c9452),
	.w5(32'h3ac8bf51),
	.w6(32'hbaacc74b),
	.w7(32'hbacff527),
	.w8(32'hbb0ce999),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7646a4),
	.w1(32'hbb3dda31),
	.w2(32'hb8f7aad1),
	.w3(32'h3adaf615),
	.w4(32'h3b03a0ba),
	.w5(32'h3b2ecaef),
	.w6(32'h3ae4e117),
	.w7(32'h3a8f3c1b),
	.w8(32'h3a8ec9f6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b1029),
	.w1(32'hbabcce0f),
	.w2(32'hba8f0f8a),
	.w3(32'h3be429fa),
	.w4(32'h3b4a4444),
	.w5(32'hbb8345fc),
	.w6(32'h3a5bfd0b),
	.w7(32'h3aa471ee),
	.w8(32'hbbc20754),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87cec9),
	.w1(32'hbb51b15a),
	.w2(32'hbb3ccb0d),
	.w3(32'h3a8b0ee8),
	.w4(32'hbaecfa72),
	.w5(32'hbbcf8997),
	.w6(32'hbb701c7e),
	.w7(32'hbb3c9ab4),
	.w8(32'hbbc8fbdd),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e7080),
	.w1(32'hbbe115dd),
	.w2(32'hbbb23adf),
	.w3(32'hbb94803e),
	.w4(32'hbb6941cd),
	.w5(32'h3bddfb78),
	.w6(32'hbb7d84e3),
	.w7(32'hbb9ea7a1),
	.w8(32'h3bd59290),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5261b),
	.w1(32'h3bcb62d4),
	.w2(32'hbaedf615),
	.w3(32'h3ac26d5f),
	.w4(32'hbb192633),
	.w5(32'hb9ee2a71),
	.w6(32'h3af6f42c),
	.w7(32'hbb49a655),
	.w8(32'hb9b4d673),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a0184),
	.w1(32'hba376859),
	.w2(32'hba5b2b66),
	.w3(32'h3b60536a),
	.w4(32'h3b131ed9),
	.w5(32'hbb458490),
	.w6(32'h39f98c88),
	.w7(32'h397ae391),
	.w8(32'hbb03b362),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1330c1),
	.w1(32'hb9fd3e75),
	.w2(32'hba96facf),
	.w3(32'hb8681c09),
	.w4(32'hbaeda67f),
	.w5(32'hbb108805),
	.w6(32'h37954949),
	.w7(32'hbaac1990),
	.w8(32'hbb11a071),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b638b),
	.w1(32'h3ab661b4),
	.w2(32'hb97f4a58),
	.w3(32'hb799e629),
	.w4(32'hbb34ba14),
	.w5(32'hbb9792b0),
	.w6(32'hbb0d407b),
	.w7(32'hbae00966),
	.w8(32'hbb1f1590),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a88be),
	.w1(32'hba0835fb),
	.w2(32'hbb167051),
	.w3(32'hba71506b),
	.w4(32'h3a95d7ff),
	.w5(32'h3bb02cfe),
	.w6(32'hbb3796a3),
	.w7(32'hba77ea79),
	.w8(32'h3ba6ec13),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafcee9),
	.w1(32'h3c0068ea),
	.w2(32'hbae8d97b),
	.w3(32'hb8aa1719),
	.w4(32'hbb611493),
	.w5(32'h3b02a477),
	.w6(32'h3b1156bb),
	.w7(32'hbb78659f),
	.w8(32'h3b65b27e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07efc7),
	.w1(32'h3b072d3f),
	.w2(32'h3a9e2b52),
	.w3(32'h3b36fc4b),
	.w4(32'h3b2b8198),
	.w5(32'h3b1f79d6),
	.w6(32'h3b84b6d9),
	.w7(32'h3b5bd787),
	.w8(32'h3a468ed5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0af2c8),
	.w1(32'h3a782dfd),
	.w2(32'h3a810c43),
	.w3(32'h3b17688c),
	.w4(32'h3a44d32d),
	.w5(32'h3b9081b9),
	.w6(32'h3ad69dec),
	.w7(32'h3a5daef4),
	.w8(32'h3bcbf61d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13c62f),
	.w1(32'h3af2443a),
	.w2(32'hbb64f28d),
	.w3(32'h3a134932),
	.w4(32'hbb13633d),
	.w5(32'hbb24e0da),
	.w6(32'h3a058fe8),
	.w7(32'hba867f1f),
	.w8(32'hbb40c341),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1841c5),
	.w1(32'hba800917),
	.w2(32'h395ccb6b),
	.w3(32'hba25f085),
	.w4(32'hbaace623),
	.w5(32'hbb1030d0),
	.w6(32'hbacc1922),
	.w7(32'hbb1aab54),
	.w8(32'h3a883bde),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f5aaf),
	.w1(32'h3b072110),
	.w2(32'h38a4a6d8),
	.w3(32'h395ee414),
	.w4(32'h3a3d5847),
	.w5(32'hbb326af5),
	.w6(32'h3bd90064),
	.w7(32'h3b06da83),
	.w8(32'hbb2e32ed),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ba263),
	.w1(32'h3b1fe957),
	.w2(32'h3a5d7a03),
	.w3(32'hb902ae69),
	.w4(32'hb93a032d),
	.w5(32'h3b6fe1b1),
	.w6(32'h3b2de633),
	.w7(32'h3a448f3c),
	.w8(32'h3b2a665a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e4d45),
	.w1(32'h3bfc3888),
	.w2(32'h3b72873e),
	.w3(32'h3baebafa),
	.w4(32'h3a94e581),
	.w5(32'hbb42430d),
	.w6(32'h3baa33e0),
	.w7(32'h3b0c525d),
	.w8(32'hbac9159f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5121a0),
	.w1(32'hbb5a9e65),
	.w2(32'hbb431662),
	.w3(32'hbbbd6394),
	.w4(32'hbb582aaa),
	.w5(32'h3a425d8e),
	.w6(32'hbbc1d45b),
	.w7(32'hbb5f7473),
	.w8(32'h3b63b9c0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5233a0),
	.w1(32'hb9ad421f),
	.w2(32'hbae3f980),
	.w3(32'hb9a5fae2),
	.w4(32'hba35b1bb),
	.w5(32'h3a1eabac),
	.w6(32'hb9909f2a),
	.w7(32'hbb141f32),
	.w8(32'h376895b1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad283f3),
	.w1(32'h3bc9972f),
	.w2(32'h3bc27332),
	.w3(32'hbb2ba174),
	.w4(32'h3ad6a674),
	.w5(32'h3ae81e4d),
	.w6(32'h3b2364ff),
	.w7(32'h3b9e1316),
	.w8(32'hbb401620),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a62f06),
	.w1(32'hbb2821b3),
	.w2(32'h3b4b0017),
	.w3(32'h3b87a672),
	.w4(32'h3bc471c9),
	.w5(32'hbb1967ee),
	.w6(32'hba8953bc),
	.w7(32'h3af0bbe0),
	.w8(32'h3a80ad15),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdd0b5),
	.w1(32'h3b81b71b),
	.w2(32'h3b8c2982),
	.w3(32'hbb1922ca),
	.w4(32'hb85c52fb),
	.w5(32'hbbd35d45),
	.w6(32'h3af474ca),
	.w7(32'h3bb3a870),
	.w8(32'hbb8baa0b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb561e6e),
	.w1(32'hbb181184),
	.w2(32'hbb52091b),
	.w3(32'hbb51c881),
	.w4(32'hbb65299b),
	.w5(32'hbadf29e8),
	.w6(32'hbb4a4ba1),
	.w7(32'hbb57a959),
	.w8(32'hbab65f63),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3feee8),
	.w1(32'h39d1eaa9),
	.w2(32'hbab6f04e),
	.w3(32'hbaeb44e9),
	.w4(32'hbaf7c179),
	.w5(32'hbbabc252),
	.w6(32'h39dfb524),
	.w7(32'hba2d81c9),
	.w8(32'hba752da6),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3010a8),
	.w1(32'h3b62b6df),
	.w2(32'h3b931f44),
	.w3(32'hbae574e9),
	.w4(32'hbb6dd802),
	.w5(32'h3abb1ce1),
	.w6(32'h3a9c98d2),
	.w7(32'h3b277c6c),
	.w8(32'h3b4c7de8),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0407a6),
	.w1(32'h3ba6e571),
	.w2(32'h3ac041d5),
	.w3(32'h3a651e49),
	.w4(32'h3a845e0b),
	.w5(32'h3b4b6b18),
	.w6(32'h3b44a0e8),
	.w7(32'h3b64e025),
	.w8(32'h3b7bc387),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc5057),
	.w1(32'h3bf44e13),
	.w2(32'h3b99a135),
	.w3(32'h3a93c32a),
	.w4(32'hba836aba),
	.w5(32'h3b2003bc),
	.w6(32'h3b805834),
	.w7(32'h3b946a5b),
	.w8(32'h3aa95347),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64b93d),
	.w1(32'hbb9b09b7),
	.w2(32'hbb61b8c2),
	.w3(32'h3aec58b6),
	.w4(32'hba3afcb7),
	.w5(32'h3b01fb8e),
	.w6(32'hbb09077a),
	.w7(32'hbb10900c),
	.w8(32'h3bad256e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda6996),
	.w1(32'h3ab5513e),
	.w2(32'h3ad1c4b9),
	.w3(32'h3b34c03a),
	.w4(32'h3b22f798),
	.w5(32'h3bacc66b),
	.w6(32'h3b5c7525),
	.w7(32'h3b4dee49),
	.w8(32'h3b4ec895),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69d10c),
	.w1(32'hbb0eb35e),
	.w2(32'hb9837745),
	.w3(32'h3b4f5034),
	.w4(32'h3b37b17c),
	.w5(32'h3a0b115e),
	.w6(32'h397fa8a8),
	.w7(32'h3adefc7a),
	.w8(32'h3bf270be),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39966344),
	.w1(32'h3b6f400b),
	.w2(32'h3b522790),
	.w3(32'h3b93a6f6),
	.w4(32'h3bf13455),
	.w5(32'hb9df3ddb),
	.w6(32'h3c33fb9e),
	.w7(32'h3bf74407),
	.w8(32'hbae70b76),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bc1c7),
	.w1(32'h393aad29),
	.w2(32'hba5246bd),
	.w3(32'hbb4099d5),
	.w4(32'hbaaa9a79),
	.w5(32'hbbb25079),
	.w6(32'hbb1f43d8),
	.w7(32'h3904e793),
	.w8(32'hbb9f1dd4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46203c),
	.w1(32'h3a9b8780),
	.w2(32'h3a6cb863),
	.w3(32'hbb8df101),
	.w4(32'hbb11852b),
	.w5(32'hbbdb634c),
	.w6(32'hba3a7bef),
	.w7(32'h3a77c336),
	.w8(32'hbb97b1dd),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1819a2),
	.w1(32'hbbb3be1a),
	.w2(32'h3b006d86),
	.w3(32'hbbe13ee6),
	.w4(32'hb9b88eb1),
	.w5(32'h3c0784b9),
	.w6(32'hbb5202e9),
	.w7(32'h3b9275d9),
	.w8(32'h3c59c413),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4242f),
	.w1(32'h3b482f89),
	.w2(32'h3ad24012),
	.w3(32'h3c07e6bb),
	.w4(32'h3bdd627a),
	.w5(32'hbb3e8311),
	.w6(32'h3c1cc087),
	.w7(32'h3bee541f),
	.w8(32'hb9686ee3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b93996),
	.w1(32'h3a0d8223),
	.w2(32'hb8cf379f),
	.w3(32'hba9b7151),
	.w4(32'hb9c2bfca),
	.w5(32'h3ad40a15),
	.w6(32'h3ab449dc),
	.w7(32'h3b062489),
	.w8(32'h390880fb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26632c),
	.w1(32'hbb760d60),
	.w2(32'hbb912ca7),
	.w3(32'h39c455cf),
	.w4(32'hba939d88),
	.w5(32'hba174b92),
	.w6(32'hbb37abe5),
	.w7(32'hbb68c095),
	.w8(32'hbb0fbf4c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d6c03),
	.w1(32'hbb817a5d),
	.w2(32'hbb2c7d19),
	.w3(32'hbaeb3c8d),
	.w4(32'hbb3238b4),
	.w5(32'h3b2b3d27),
	.w6(32'hbb37f2dc),
	.w7(32'hbb258dd2),
	.w8(32'h3b85171d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acdf40),
	.w1(32'h3a16c393),
	.w2(32'hba60e321),
	.w3(32'h3b1fd6e5),
	.w4(32'h3a305866),
	.w5(32'hbc031968),
	.w6(32'h3b8ae027),
	.w7(32'h39a292d5),
	.w8(32'hbbc568e3),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3b986),
	.w1(32'hba1771d3),
	.w2(32'h3bcbcc89),
	.w3(32'hbb1eb257),
	.w4(32'h3b567126),
	.w5(32'hb9663de7),
	.w6(32'hbaf2a6a4),
	.w7(32'h3b8a4a9c),
	.w8(32'h38380701),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ab57e),
	.w1(32'h3ae82492),
	.w2(32'h3b4c5e87),
	.w3(32'hba576a61),
	.w4(32'hbaa7844d),
	.w5(32'hbaa21269),
	.w6(32'hb9a9462a),
	.w7(32'h3afd7021),
	.w8(32'hba46d1e7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e985e),
	.w1(32'hbb38e3c2),
	.w2(32'h3a84c9fd),
	.w3(32'hbb238b0a),
	.w4(32'h39a14424),
	.w5(32'h3b1bfe69),
	.w6(32'hba5c81be),
	.w7(32'hb8c572bb),
	.w8(32'h3ba5e6b7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b861bb3),
	.w1(32'h3b6303c5),
	.w2(32'hbb13ac1e),
	.w3(32'hbb3752c3),
	.w4(32'hba1b48f7),
	.w5(32'hbb70d0da),
	.w6(32'h3b1cfe98),
	.w7(32'h39528af7),
	.w8(32'hbabbdca4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39653bf0),
	.w1(32'hb9b81dc0),
	.w2(32'hbab5995f),
	.w3(32'hba9cb7d2),
	.w4(32'h398d76f7),
	.w5(32'hbab29e2c),
	.w6(32'hbb0b2325),
	.w7(32'hba086d30),
	.w8(32'hbb02271f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a2ca1),
	.w1(32'hba9053ca),
	.w2(32'hbb2ec59a),
	.w3(32'hbb21965b),
	.w4(32'hbadd2214),
	.w5(32'h3b912d8b),
	.w6(32'hbb3e15ad),
	.w7(32'hbb0c2bf5),
	.w8(32'h3ac72b06),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b111091),
	.w1(32'h3a32a4b1),
	.w2(32'h39dfd35d),
	.w3(32'h3b262bc4),
	.w4(32'h3b11f065),
	.w5(32'hbb4ec537),
	.w6(32'h3a1c844f),
	.w7(32'h3ae771c9),
	.w8(32'h3a9997eb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad01bc5),
	.w1(32'hbaac6e18),
	.w2(32'hbac03de7),
	.w3(32'hbb17ac8e),
	.w4(32'hbb32befb),
	.w5(32'h3a21a2c1),
	.w6(32'hb9b57085),
	.w7(32'hba7ff627),
	.w8(32'hb6e01490),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084799),
	.w1(32'h39735007),
	.w2(32'hba77b721),
	.w3(32'h39204a91),
	.w4(32'hba0c706d),
	.w5(32'hbb966ebb),
	.w6(32'h3b593cfa),
	.w7(32'hb8a7c87a),
	.w8(32'h3a5a2185),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90443ff),
	.w1(32'hbaaf9c71),
	.w2(32'hbb87ac54),
	.w3(32'h3b72bb53),
	.w4(32'h3b01166e),
	.w5(32'hbab8d3c1),
	.w6(32'h3bb80670),
	.w7(32'h3bbc713d),
	.w8(32'h3ac7bd07),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e4884),
	.w1(32'hbb0fd903),
	.w2(32'hbb9732f3),
	.w3(32'h389eab2c),
	.w4(32'hbb1860bb),
	.w5(32'h3b495d3b),
	.w6(32'hb9b6892d),
	.w7(32'hbb5bfb72),
	.w8(32'h3bbcee52),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d4fe22),
	.w1(32'hbae7d2c2),
	.w2(32'hbb44f587),
	.w3(32'h3b6f21ba),
	.w4(32'h3b141735),
	.w5(32'hba69a8f8),
	.w6(32'h3b885ba4),
	.w7(32'h3a511977),
	.w8(32'h3a82ecf7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21419b),
	.w1(32'hba9efe3e),
	.w2(32'hbaf5808d),
	.w3(32'hba0916f9),
	.w4(32'hbaad3dfc),
	.w5(32'h3abfb86e),
	.w6(32'h3a728d4d),
	.w7(32'hba02a73e),
	.w8(32'h39504e2f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07af99),
	.w1(32'hb99ee8fc),
	.w2(32'h39508522),
	.w3(32'hb9f73fc7),
	.w4(32'h3996df09),
	.w5(32'hbb277cde),
	.w6(32'hb8fb271e),
	.w7(32'h3a94f64e),
	.w8(32'hba3b819f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02ac76),
	.w1(32'hbb428947),
	.w2(32'hbac682cc),
	.w3(32'hbb90b7b2),
	.w4(32'hbad758bf),
	.w5(32'hba95a537),
	.w6(32'hbb875ae0),
	.w7(32'hbad968d3),
	.w8(32'hbab2672d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35357f),
	.w1(32'hbb69e1ba),
	.w2(32'hbb19b522),
	.w3(32'hba88a097),
	.w4(32'hbab14c04),
	.w5(32'h3b0cff49),
	.w6(32'hbb00ed12),
	.w7(32'hbb9a1197),
	.w8(32'h3b4205db),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c029f),
	.w1(32'hb981fd8b),
	.w2(32'hbb321e1c),
	.w3(32'h3ae9b51b),
	.w4(32'h3a58ecd6),
	.w5(32'h3ab4f1c4),
	.w6(32'h3b87d6ec),
	.w7(32'hb9a4113c),
	.w8(32'hb9968cb3),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae03f9e),
	.w1(32'hbb8b6d7f),
	.w2(32'hbbdf96af),
	.w3(32'h3ad9d59c),
	.w4(32'h3a9497db),
	.w5(32'hbbe17b0d),
	.w6(32'hbb193919),
	.w7(32'hbb759a86),
	.w8(32'hbb718b79),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77ab54),
	.w1(32'hb905a930),
	.w2(32'h3bbd8c4b),
	.w3(32'hbb9179e1),
	.w4(32'hba730d58),
	.w5(32'hbb9d39a1),
	.w6(32'hbb4ceb52),
	.w7(32'h3b64e185),
	.w8(32'hbb98a64c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb226ae0),
	.w1(32'h39022ee9),
	.w2(32'hbac4b03d),
	.w3(32'hbafd0efc),
	.w4(32'hbb4f8b6c),
	.w5(32'hbb0d567d),
	.w6(32'hbb202541),
	.w7(32'hb9732f12),
	.w8(32'hbaa7b047),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb403c39),
	.w1(32'hb95feb08),
	.w2(32'hba16ef20),
	.w3(32'hba3ed89f),
	.w4(32'h39c246d2),
	.w5(32'h3be09da1),
	.w6(32'h3aa807d4),
	.w7(32'h3b02d865),
	.w8(32'h3b9022b4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad88049),
	.w1(32'hbae6d098),
	.w2(32'h3a16f6e9),
	.w3(32'h3b72dfac),
	.w4(32'hb9b1eb35),
	.w5(32'h3bf4ce7c),
	.w6(32'hb97a3165),
	.w7(32'hbb0b4c6b),
	.w8(32'h3b41c21f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55006f),
	.w1(32'hbaf40787),
	.w2(32'hba3a63e0),
	.w3(32'h3baf806a),
	.w4(32'h3aff06de),
	.w5(32'hba813109),
	.w6(32'h3b7f3cc3),
	.w7(32'h3b875a7f),
	.w8(32'h3a68675a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51a3c5),
	.w1(32'hba6ee298),
	.w2(32'hb8f60730),
	.w3(32'hbad72107),
	.w4(32'hbaa2e22d),
	.w5(32'h3c0c09d0),
	.w6(32'hba331a38),
	.w7(32'hba8d6065),
	.w8(32'h3c04eb87),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8a207),
	.w1(32'h3b73b5ee),
	.w2(32'h39571ac2),
	.w3(32'h3b042a94),
	.w4(32'h3b012c2a),
	.w5(32'hba5f63f4),
	.w6(32'hb9ff2f4a),
	.w7(32'h3a7a9dd6),
	.w8(32'hbb42bff9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49d05c),
	.w1(32'hbb3c330c),
	.w2(32'h38e745db),
	.w3(32'hb9eb4882),
	.w4(32'hba78a10c),
	.w5(32'h3bb3d49c),
	.w6(32'hbb82fadc),
	.w7(32'hbb09edaf),
	.w8(32'h3b2f8b18),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad79af),
	.w1(32'hba81dd29),
	.w2(32'h3a116e73),
	.w3(32'h3bb1cf84),
	.w4(32'h3b7d9b27),
	.w5(32'hbb2d649d),
	.w6(32'h3b023df3),
	.w7(32'h3aa6388f),
	.w8(32'hbb566032),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28bc78),
	.w1(32'hbad7c118),
	.w2(32'hb8a7ad3e),
	.w3(32'hbaf49a13),
	.w4(32'hbb2a0166),
	.w5(32'hba9e9418),
	.w6(32'hbaf0b249),
	.w7(32'hb8914d4a),
	.w8(32'hbab83413),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c28e8),
	.w1(32'hbb1fb300),
	.w2(32'hba9dddc9),
	.w3(32'hbaa97154),
	.w4(32'hbb1c07e5),
	.w5(32'h3a9dc237),
	.w6(32'hbabe031e),
	.w7(32'hbaadbd56),
	.w8(32'h3a6e235a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10df67),
	.w1(32'hbb357579),
	.w2(32'hbb5531a8),
	.w3(32'h3aaa6a00),
	.w4(32'hb936c499),
	.w5(32'hbb3bc94e),
	.w6(32'hba234b9d),
	.w7(32'hbb0a918e),
	.w8(32'hbb7cac58),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0321f),
	.w1(32'hbbbcb3e0),
	.w2(32'hbbb3f9fb),
	.w3(32'hbb8a3c6e),
	.w4(32'hbad8e6e3),
	.w5(32'hbb21c907),
	.w6(32'hbb5fbd94),
	.w7(32'hbae39ca9),
	.w8(32'hb9ea151f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04d33f),
	.w1(32'hba96c7e7),
	.w2(32'h39a86849),
	.w3(32'hbaba1485),
	.w4(32'hbad8880b),
	.w5(32'hb8d57426),
	.w6(32'hba05579d),
	.w7(32'hb99c6ba9),
	.w8(32'hb81a5345),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78a432e),
	.w1(32'h3a42ac23),
	.w2(32'h3bb0006c),
	.w3(32'hb99e3c7e),
	.w4(32'hba44ef18),
	.w5(32'hba73fc0e),
	.w6(32'hbb110142),
	.w7(32'h3a841bc3),
	.w8(32'h3a6ceaf3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60ee94),
	.w1(32'h3a53b88c),
	.w2(32'hbb9853f1),
	.w3(32'hbad1d4ad),
	.w4(32'hba41a6b7),
	.w5(32'h3a4f9f3a),
	.w6(32'hba0f8232),
	.w7(32'hbb5626f0),
	.w8(32'h3a7f2836),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dafa9),
	.w1(32'h3a313b67),
	.w2(32'h3b181746),
	.w3(32'h3a4c62f8),
	.w4(32'hbac76ad5),
	.w5(32'hb9d535b0),
	.w6(32'hba42be3d),
	.w7(32'hb88156bb),
	.w8(32'h3a06e70d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf76499),
	.w1(32'h3a7bbe92),
	.w2(32'hb96776cc),
	.w3(32'h3a83db96),
	.w4(32'h3a892566),
	.w5(32'hbb97027c),
	.w6(32'h3b825c24),
	.w7(32'h3ad99758),
	.w8(32'hba9cc71f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba29ab7),
	.w1(32'h3b1afaef),
	.w2(32'h3b0c9307),
	.w3(32'hba1b052f),
	.w4(32'h39502927),
	.w5(32'h3982d519),
	.w6(32'h3b9cb1fd),
	.w7(32'h3b2509b3),
	.w8(32'h3b0683ea),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f3658),
	.w1(32'hb895bbf5),
	.w2(32'hba148f1f),
	.w3(32'h3ad18dbf),
	.w4(32'h3b0ef54c),
	.w5(32'hbb0415c6),
	.w6(32'h3a150706),
	.w7(32'hb978e92b),
	.w8(32'hbabfc1a9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c44cd),
	.w1(32'hb9e8b88c),
	.w2(32'hbabfdbf2),
	.w3(32'hb9826a25),
	.w4(32'hbabeff3f),
	.w5(32'h3a3ea4e2),
	.w6(32'h396c6987),
	.w7(32'hba96b85d),
	.w8(32'h39eeb7a1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34d356),
	.w1(32'h397a5f45),
	.w2(32'h3b0d9b83),
	.w3(32'h3b1eb13e),
	.w4(32'h3b6c0534),
	.w5(32'h3b8d71eb),
	.w6(32'h39df7042),
	.w7(32'h3a138ede),
	.w8(32'h3b9ba4d2),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacd101),
	.w1(32'hba53fa97),
	.w2(32'hbb6a03b8),
	.w3(32'hbafdd535),
	.w4(32'h3a5627ad),
	.w5(32'hbbc94a59),
	.w6(32'hbb6e8dd5),
	.w7(32'hbac23058),
	.w8(32'hbb1adf16),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d3e906),
	.w1(32'hbb218bf5),
	.w2(32'hbbc9de5c),
	.w3(32'hbb511315),
	.w4(32'hbb839f13),
	.w5(32'h3abb71d9),
	.w6(32'hba905717),
	.w7(32'hbba2594d),
	.w8(32'hb93b55ed),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb664dad),
	.w1(32'h3a87ab4d),
	.w2(32'h3a938e02),
	.w3(32'h39dd5ff4),
	.w4(32'h3a9d5679),
	.w5(32'hbb8a7d79),
	.w6(32'h3b16b41e),
	.w7(32'h3aa82a92),
	.w8(32'hba2f38e1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b5324),
	.w1(32'h3b822eef),
	.w2(32'h3b401de6),
	.w3(32'h3a6c85cd),
	.w4(32'h393204ff),
	.w5(32'h3c08d790),
	.w6(32'h3bb0fd94),
	.w7(32'h3b885134),
	.w8(32'h3bf59ac2),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc88850),
	.w1(32'h3bd5ebe5),
	.w2(32'h3b8f27d0),
	.w3(32'h3bc16f17),
	.w4(32'h3ac0f6e7),
	.w5(32'h3a821c0c),
	.w6(32'h3bbff999),
	.w7(32'h3b4725c2),
	.w8(32'hbac144cc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b348986),
	.w1(32'h3987dff7),
	.w2(32'h39b6857e),
	.w3(32'h3b92d192),
	.w4(32'h3b12ea44),
	.w5(32'h3a05e170),
	.w6(32'h3ad38ece),
	.w7(32'hba0e6abe),
	.w8(32'h3af3b559),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b285c7c),
	.w1(32'hba78c279),
	.w2(32'h3924b560),
	.w3(32'hba9cfc24),
	.w4(32'h38b81e7b),
	.w5(32'h3b0c562c),
	.w6(32'hbaa09a8b),
	.w7(32'hba379a0e),
	.w8(32'hba9705ef),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9af72),
	.w1(32'hba9128b7),
	.w2(32'h3b9b3c62),
	.w3(32'h3b2661e5),
	.w4(32'h3bb2951b),
	.w5(32'h3a85a4e1),
	.w6(32'h3a987d2c),
	.w7(32'h3ba7b320),
	.w8(32'h3a647f91),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ababce5),
	.w1(32'h3a3a20fa),
	.w2(32'h3a7744c0),
	.w3(32'h39410f3d),
	.w4(32'hb9a4e457),
	.w5(32'hbb5a66e1),
	.w6(32'h38e0e5ed),
	.w7(32'hb2b10190),
	.w8(32'hbb6569de),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94471e),
	.w1(32'hbbb98177),
	.w2(32'hbb6879e1),
	.w3(32'hbb81e92f),
	.w4(32'hbb56ea93),
	.w5(32'hbaacd50b),
	.w6(32'hbb33ced1),
	.w7(32'hbb8ba6d0),
	.w8(32'hba9a3a68),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb196e35),
	.w1(32'hba962d8e),
	.w2(32'hbb2f5a4d),
	.w3(32'h3a9eadd4),
	.w4(32'h39dcaf56),
	.w5(32'hbb0a5294),
	.w6(32'h3b0486aa),
	.w7(32'hbaa4e3b7),
	.w8(32'hbb3cb534),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb814639),
	.w1(32'hbb8d4c10),
	.w2(32'hbb6f34bc),
	.w3(32'hbb030c44),
	.w4(32'hb9866e25),
	.w5(32'hba6ea609),
	.w6(32'hba569b33),
	.w7(32'h3884ff92),
	.w8(32'hbaba77b7),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0005e7),
	.w1(32'hbb1460b9),
	.w2(32'hbaf99fe4),
	.w3(32'hba9cd3cb),
	.w4(32'hbadb1be8),
	.w5(32'hbb32758f),
	.w6(32'hbb0ee1cf),
	.w7(32'hbb04d7a5),
	.w8(32'hbb1be7fc),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a9127),
	.w1(32'hb9f9a3d9),
	.w2(32'hb96babb9),
	.w3(32'hba2cf985),
	.w4(32'hbaf9de12),
	.w5(32'hba87bf5d),
	.w6(32'hbaac116f),
	.w7(32'hbaac05c2),
	.w8(32'hbb203533),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71b57a1),
	.w1(32'hbac1b01f),
	.w2(32'hbaf17fdb),
	.w3(32'hba889d1d),
	.w4(32'hbb2855ac),
	.w5(32'hbb47908c),
	.w6(32'hbb7539e5),
	.w7(32'hbb890112),
	.w8(32'hbb1d8b7e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb376178),
	.w1(32'hbb5bebcb),
	.w2(32'hbb460809),
	.w3(32'hbafb7fd5),
	.w4(32'hbb137df0),
	.w5(32'hbb12e7f0),
	.w6(32'hbaee95a0),
	.w7(32'hbb5ffb8d),
	.w8(32'hbb17d990),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb062829),
	.w1(32'hbab1d805),
	.w2(32'hba86cafa),
	.w3(32'hbb136ae7),
	.w4(32'hbab2f963),
	.w5(32'h3ac7f599),
	.w6(32'hbacdf39a),
	.w7(32'hba20f28f),
	.w8(32'h3aea9f87),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1aa245),
	.w1(32'h3a4d8c55),
	.w2(32'h3adbe6ba),
	.w3(32'h3aaaf831),
	.w4(32'h3a66feff),
	.w5(32'h3b086f07),
	.w6(32'h3b49c508),
	.w7(32'h3b581e57),
	.w8(32'h3aed86d7),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13b7fe),
	.w1(32'hb8ad4f5a),
	.w2(32'h391ddcdd),
	.w3(32'h39b842e8),
	.w4(32'hba1ab134),
	.w5(32'h3bc50fd4),
	.w6(32'hb9c4f71f),
	.w7(32'hba540bf5),
	.w8(32'h3bd75bb0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb088cf),
	.w1(32'h3b9cda71),
	.w2(32'h3b4fc378),
	.w3(32'h3ba6713a),
	.w4(32'h3b5665f3),
	.w5(32'h3b031423),
	.w6(32'h3bb44150),
	.w7(32'h3b8dbd00),
	.w8(32'h3ae452c1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c309dd),
	.w1(32'hba67224d),
	.w2(32'hb8dfd364),
	.w3(32'h3b2dcd57),
	.w4(32'h3abcbd0c),
	.w5(32'hba60f803),
	.w6(32'h3afe83bd),
	.w7(32'h3acae19b),
	.w8(32'hbaefdb0c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb428799),
	.w1(32'hbaf4dff3),
	.w2(32'hba97a133),
	.w3(32'hbad0c98a),
	.w4(32'hbae0edfa),
	.w5(32'h3a8b8804),
	.w6(32'hbae6d0f5),
	.w7(32'hba8c6b44),
	.w8(32'h3a4d8d16),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7c8e7),
	.w1(32'h39082e97),
	.w2(32'hba2a28c4),
	.w3(32'h3a8225fb),
	.w4(32'h391a70f4),
	.w5(32'hba771cb3),
	.w6(32'h3a3745d7),
	.w7(32'hbafa3cf0),
	.w8(32'hba42bc48),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1793b),
	.w1(32'h3935e150),
	.w2(32'hbab7e5c5),
	.w3(32'h396a3ad9),
	.w4(32'hbad209df),
	.w5(32'hbb816c85),
	.w6(32'h39fbb800),
	.w7(32'h3845cca9),
	.w8(32'hbb58c0dd),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee741),
	.w1(32'hbb1f9c29),
	.w2(32'hbadffa6e),
	.w3(32'hbb51d5c7),
	.w4(32'hbb05d38f),
	.w5(32'hb9a249d6),
	.w6(32'h3a0ccb33),
	.w7(32'hbae5d44e),
	.w8(32'hbac62443),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fe26d),
	.w1(32'hbb2e0c0c),
	.w2(32'hb9e9c60a),
	.w3(32'hbb414e14),
	.w4(32'hbb0547aa),
	.w5(32'h3b3f5a3c),
	.w6(32'hbb21d367),
	.w7(32'h38021070),
	.w8(32'h3b7867e6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f060b),
	.w1(32'h3b521ab7),
	.w2(32'h3b480bb3),
	.w3(32'h3af46425),
	.w4(32'h3b329455),
	.w5(32'hbaa18837),
	.w6(32'h3b028d76),
	.w7(32'h3b39cf2e),
	.w8(32'hba06cf54),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8685ea),
	.w1(32'hb9ada47b),
	.w2(32'hba834f9f),
	.w3(32'h39f680bb),
	.w4(32'h38e09e47),
	.w5(32'hba956cf2),
	.w6(32'h3a42b2a4),
	.w7(32'h3b2d9ddb),
	.w8(32'hba0e6faa),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e345b1),
	.w1(32'hbad93451),
	.w2(32'hbaafabf8),
	.w3(32'hbaad17c7),
	.w4(32'hbb190b94),
	.w5(32'hbb0e1cd9),
	.w6(32'hbaa44654),
	.w7(32'hbb062f43),
	.w8(32'hb848c8e7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e57e1a),
	.w1(32'h3a868497),
	.w2(32'h3a535ea8),
	.w3(32'hbabafb67),
	.w4(32'hbabe9bd9),
	.w5(32'h3b1b6802),
	.w6(32'hbae7cfff),
	.w7(32'hbaaad135),
	.w8(32'h3b096057),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6e24b),
	.w1(32'h3a188f9a),
	.w2(32'hba7a5b55),
	.w3(32'h3ac92542),
	.w4(32'h3a0be9c2),
	.w5(32'hba8dea6f),
	.w6(32'h3b28d092),
	.w7(32'h3a7d79c9),
	.w8(32'hbacfee55),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03680b),
	.w1(32'hbaa74111),
	.w2(32'hbab183cc),
	.w3(32'h38973a8d),
	.w4(32'hba9c933d),
	.w5(32'h3af574c5),
	.w6(32'hbb09aaea),
	.w7(32'hbb2711e4),
	.w8(32'hbb3e2e10),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e3b6b),
	.w1(32'hbadba14a),
	.w2(32'hb881c633),
	.w3(32'h3a96a7ba),
	.w4(32'h3a198c9d),
	.w5(32'hb9316805),
	.w6(32'hbad7f94d),
	.w7(32'hbaf81a08),
	.w8(32'h3aee08c8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e4a74),
	.w1(32'h3aed75e6),
	.w2(32'h3afa74fa),
	.w3(32'h3a2c9080),
	.w4(32'hba52891c),
	.w5(32'h3b8fd325),
	.w6(32'h3a4e1b7a),
	.w7(32'h392bee7f),
	.w8(32'h3a4a45a1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5944a),
	.w1(32'hba21a6ed),
	.w2(32'hba88944d),
	.w3(32'h3b256e51),
	.w4(32'h3b2ceb58),
	.w5(32'hbaf6511d),
	.w6(32'h3a8c5880),
	.w7(32'h3a0f957f),
	.w8(32'hbab28d95),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1c032),
	.w1(32'hbadfcff1),
	.w2(32'hbb4ea289),
	.w3(32'hbae1b710),
	.w4(32'hbb17201e),
	.w5(32'hba78c672),
	.w6(32'hba0b07a7),
	.w7(32'hba71463f),
	.w8(32'h3a3ada5e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b144e3f),
	.w1(32'h3aec3dee),
	.w2(32'h399de299),
	.w3(32'hb8267475),
	.w4(32'hbb10663f),
	.w5(32'hbb612f41),
	.w6(32'h3b09630c),
	.w7(32'h3680d88c),
	.w8(32'hbb36875f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63b390),
	.w1(32'hbb00cb1a),
	.w2(32'hb8e9fa9f),
	.w3(32'hbafc91cc),
	.w4(32'hba74abf3),
	.w5(32'h3b8fb26a),
	.w6(32'hbacf2e87),
	.w7(32'hbaa0efb1),
	.w8(32'h3b34bb3f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule