module layer_10_featuremap_403(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbd0db),
	.w1(32'hba4ad76e),
	.w2(32'hb7b40ed9),
	.w3(32'hbae824ce),
	.w4(32'h3aeb33d0),
	.w5(32'hbaaf73a2),
	.w6(32'hba641a0c),
	.w7(32'h3b3298b6),
	.w8(32'h39a1f0a2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc7716),
	.w1(32'hbaedc30e),
	.w2(32'h3abb22d1),
	.w3(32'hba4880b0),
	.w4(32'hba166382),
	.w5(32'h3aebcb9a),
	.w6(32'hbb2bed62),
	.w7(32'hbb4f5230),
	.w8(32'hbb0ea421),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92030e7),
	.w1(32'hbb3298f4),
	.w2(32'hbb644d55),
	.w3(32'h3addc8e7),
	.w4(32'hbb50d329),
	.w5(32'h3a5eef4b),
	.w6(32'hbafd9b7c),
	.w7(32'h39992c61),
	.w8(32'hba3fed32),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69728b),
	.w1(32'h3a90f11f),
	.w2(32'hbb0aefac),
	.w3(32'h3ab2f44d),
	.w4(32'h3a0695ac),
	.w5(32'hba929dbb),
	.w6(32'hba5c8827),
	.w7(32'hb9bbe1e6),
	.w8(32'hbb5ad648),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5552c5),
	.w1(32'hbabee3de),
	.w2(32'hba3101f1),
	.w3(32'h3b4ea5aa),
	.w4(32'h3ad46465),
	.w5(32'h3a0ba5aa),
	.w6(32'hbb68952c),
	.w7(32'h3b7bc920),
	.w8(32'h3b1a8203),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9655b6),
	.w1(32'h3a9111a3),
	.w2(32'hbb8bdf3f),
	.w3(32'hb8949524),
	.w4(32'h3bcca289),
	.w5(32'hbac380d9),
	.w6(32'hbb250139),
	.w7(32'hbb5a1498),
	.w8(32'h3c291b0d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae4327),
	.w1(32'hbba9edb2),
	.w2(32'hba8a5a9a),
	.w3(32'hbad35662),
	.w4(32'hbbd32c3c),
	.w5(32'hbac88f55),
	.w6(32'h3b417e1d),
	.w7(32'h3a04b57c),
	.w8(32'hb9b2f767),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07832d),
	.w1(32'h3adf5f02),
	.w2(32'h387e1431),
	.w3(32'hba134328),
	.w4(32'h3b1ceecc),
	.w5(32'hbb9a746b),
	.w6(32'hba949320),
	.w7(32'hb88388b1),
	.w8(32'hbb006cd2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4037ac),
	.w1(32'hba95927a),
	.w2(32'h3ab9554b),
	.w3(32'h3b92a905),
	.w4(32'hb9cbbb33),
	.w5(32'hba5a1b60),
	.w6(32'h3b368b73),
	.w7(32'hbb578902),
	.w8(32'h3a2fe8e2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c2aa3),
	.w1(32'hbafd4881),
	.w2(32'h398ea5a8),
	.w3(32'hbb8b4a62),
	.w4(32'h3aea8c1e),
	.w5(32'h399d3c51),
	.w6(32'hbb166da1),
	.w7(32'h3a070a72),
	.w8(32'hbb613c91),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16d16f),
	.w1(32'h3a792fa0),
	.w2(32'h3abdf3aa),
	.w3(32'h3b05ed58),
	.w4(32'h3b1eecf2),
	.w5(32'h3b1528ac),
	.w6(32'h3b98a08c),
	.w7(32'hbb4da2ce),
	.w8(32'hbb1019f6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20cd4f),
	.w1(32'hbb1ea1e2),
	.w2(32'h3a9d1492),
	.w3(32'h3a8b7a32),
	.w4(32'hbb986fdc),
	.w5(32'hb9985ffd),
	.w6(32'hbac5ee94),
	.w7(32'hba9fa3bb),
	.w8(32'hbafb2ec7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb096405),
	.w1(32'hb8991fd3),
	.w2(32'h3a44dc06),
	.w3(32'h3aa2cf82),
	.w4(32'hba088fcb),
	.w5(32'hbae6c049),
	.w6(32'h391e7ad8),
	.w7(32'hbc01c48e),
	.w8(32'h3b068e1c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cdc4e),
	.w1(32'hbac3aeb5),
	.w2(32'h3a4d5b03),
	.w3(32'hbb73785f),
	.w4(32'hbbf2e147),
	.w5(32'hbadb3f41),
	.w6(32'hba64634c),
	.w7(32'h38b564af),
	.w8(32'hba1c668d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84a4f8),
	.w1(32'hb9cb38f9),
	.w2(32'h3a9fa94f),
	.w3(32'hbaa21902),
	.w4(32'hba11c560),
	.w5(32'hba963480),
	.w6(32'h3a1bd307),
	.w7(32'hbb85a158),
	.w8(32'hba7097e8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa856dc),
	.w1(32'hba92097d),
	.w2(32'h3982331b),
	.w3(32'h3ae4b1d7),
	.w4(32'hbb952b9e),
	.w5(32'hbb2104c3),
	.w6(32'h3a951b2a),
	.w7(32'hbba50b13),
	.w8(32'hbb3a07de),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12a2c2),
	.w1(32'h3a9ae66a),
	.w2(32'hba2c04b5),
	.w3(32'hbb2532a1),
	.w4(32'h3a53ae25),
	.w5(32'h3b9b1380),
	.w6(32'h3ae9602a),
	.w7(32'hbb168ddb),
	.w8(32'hbbaeb937),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d45d4),
	.w1(32'h3a61d03b),
	.w2(32'hbad76ae5),
	.w3(32'h3b627d0d),
	.w4(32'hb93be506),
	.w5(32'hba95b966),
	.w6(32'hbb48ce3a),
	.w7(32'hbaa719a2),
	.w8(32'hbb14ad29),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb417587),
	.w1(32'hba5d9ea8),
	.w2(32'h3ad10520),
	.w3(32'h3ac283e6),
	.w4(32'hbae199ea),
	.w5(32'h3aabe5f2),
	.w6(32'hb8aa266c),
	.w7(32'hbb734923),
	.w8(32'hbabd48be),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4d929),
	.w1(32'h3a4e505e),
	.w2(32'h3a1c407e),
	.w3(32'h3996c35c),
	.w4(32'h3befae78),
	.w5(32'h3cb68875),
	.w6(32'hbaca4b2f),
	.w7(32'hbb721f09),
	.w8(32'h3bbb5b15),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e175a),
	.w1(32'h3b0e1275),
	.w2(32'hb97f333c),
	.w3(32'hbb403242),
	.w4(32'h3b157c0d),
	.w5(32'hbb53f40d),
	.w6(32'h3aa398c0),
	.w7(32'hbb15260a),
	.w8(32'h3b3f5ada),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3725a),
	.w1(32'h3b9b9a20),
	.w2(32'h3b44f229),
	.w3(32'h39a80c4e),
	.w4(32'h3b81fff5),
	.w5(32'h3bb3a04b),
	.w6(32'h3a715ff0),
	.w7(32'hbae00e8b),
	.w8(32'h3c19904a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95b996),
	.w1(32'hbb7f895e),
	.w2(32'hbbc923b1),
	.w3(32'hb9457ce4),
	.w4(32'hbbe3722a),
	.w5(32'hbaae9e6c),
	.w6(32'hba58ca02),
	.w7(32'hba8a94bb),
	.w8(32'hba3b1d25),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1b511),
	.w1(32'hbb74d416),
	.w2(32'hba44d43f),
	.w3(32'h3c3ccc2a),
	.w4(32'h39844b9e),
	.w5(32'hbb0b38f1),
	.w6(32'h3b469c7c),
	.w7(32'hbb059fb2),
	.w8(32'hbace428d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be7b95),
	.w1(32'hba95a2c3),
	.w2(32'hb91138fd),
	.w3(32'hbab0ca8c),
	.w4(32'hbb931503),
	.w5(32'hbb5647d7),
	.w6(32'hba435467),
	.w7(32'hb9cdf9ef),
	.w8(32'hbb984ac6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea9b73),
	.w1(32'h3b0ff5d9),
	.w2(32'hb7b46d23),
	.w3(32'hba9e9d6b),
	.w4(32'h3c205f22),
	.w5(32'h3ba1ceaf),
	.w6(32'hbada82d4),
	.w7(32'h3c0e9596),
	.w8(32'h3c45e992),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba52d2),
	.w1(32'hbbae1535),
	.w2(32'h3b26a7d4),
	.w3(32'h3b042859),
	.w4(32'hbbe893b3),
	.w5(32'hbb436dde),
	.w6(32'h3c083130),
	.w7(32'h38e7f033),
	.w8(32'h3bb5919f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f332b),
	.w1(32'hbb3046ef),
	.w2(32'hbae9d2fa),
	.w3(32'h3ba082ad),
	.w4(32'hbb13c051),
	.w5(32'hbb271f3a),
	.w6(32'h3bc841d4),
	.w7(32'h3a1d3ea8),
	.w8(32'hbb082899),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b66dfd),
	.w1(32'hbb1c4ad1),
	.w2(32'hbaaa7ab7),
	.w3(32'h3b2486e2),
	.w4(32'hbae59220),
	.w5(32'h3b91787f),
	.w6(32'hbad9619c),
	.w7(32'hba8095b7),
	.w8(32'hb9c7448d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7bf1d),
	.w1(32'h3b51a222),
	.w2(32'hbab51ada),
	.w3(32'h3b9fda67),
	.w4(32'h3ae0916b),
	.w5(32'hbb8b4523),
	.w6(32'hb9e13ffd),
	.w7(32'hb800d446),
	.w8(32'h3978fcbd),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe4168),
	.w1(32'h39e1e536),
	.w2(32'hba9daf25),
	.w3(32'hbb185139),
	.w4(32'h3bc95758),
	.w5(32'h3c036405),
	.w6(32'hba3b40b6),
	.w7(32'hbae736cb),
	.w8(32'hb9a874ed),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53fae5),
	.w1(32'hba16362b),
	.w2(32'hbac2dcf8),
	.w3(32'h3bbe83e2),
	.w4(32'hbb216d4f),
	.w5(32'hb9f730c0),
	.w6(32'h3a7a7a16),
	.w7(32'hbb9b393d),
	.w8(32'hba8dfcbe),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e95fc),
	.w1(32'hbb9d1666),
	.w2(32'hbb30dab9),
	.w3(32'h3a4d236c),
	.w4(32'hbb01e340),
	.w5(32'h3b31dce6),
	.w6(32'h3a9a10a6),
	.w7(32'h3bce0de6),
	.w8(32'h3b1e4095),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6734ea),
	.w1(32'hb9fa4166),
	.w2(32'hbaaa88c1),
	.w3(32'h3a8e55fe),
	.w4(32'h3be7ecd0),
	.w5(32'h3b83ccb8),
	.w6(32'h3bb56b44),
	.w7(32'h3b9c1654),
	.w8(32'h3b81f7b1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984d0fc),
	.w1(32'h3aba4d53),
	.w2(32'h3b957119),
	.w3(32'h3b97678d),
	.w4(32'h3aa158dc),
	.w5(32'hbbb86d23),
	.w6(32'h3b79b8cd),
	.w7(32'h3acfcc3a),
	.w8(32'h39add5f0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05a449),
	.w1(32'h3a61ea49),
	.w2(32'hb996b792),
	.w3(32'h3b429908),
	.w4(32'h3ad20501),
	.w5(32'hb961f87f),
	.w6(32'h3aca9b83),
	.w7(32'h3a063add),
	.w8(32'hbb1418aa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d06da),
	.w1(32'hbb5f2932),
	.w2(32'hbbb749d8),
	.w3(32'h3a479e86),
	.w4(32'hbb434586),
	.w5(32'hb9c1275c),
	.w6(32'h38960e58),
	.w7(32'hb99565fd),
	.w8(32'hbb930139),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa8ba0),
	.w1(32'hbac8fb4a),
	.w2(32'hba893952),
	.w3(32'hbaaa707a),
	.w4(32'hbb9fbac8),
	.w5(32'hb9281e04),
	.w6(32'hbb5dd490),
	.w7(32'hbb97f628),
	.w8(32'hba768349),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39328784),
	.w1(32'hbb128541),
	.w2(32'hbab4791a),
	.w3(32'hb9a5ed04),
	.w4(32'hbb7d9a9b),
	.w5(32'hbb3b919d),
	.w6(32'hb91d75d3),
	.w7(32'h39544ea8),
	.w8(32'hbaf9b498),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892a69),
	.w1(32'h399e49c9),
	.w2(32'h39f980bf),
	.w3(32'h3ae13f01),
	.w4(32'hb9b85da8),
	.w5(32'hbaae010d),
	.w6(32'hbb8815c4),
	.w7(32'h3acc71bc),
	.w8(32'h3b555922),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b976aab),
	.w1(32'hbbcacd1d),
	.w2(32'h3ae48dcd),
	.w3(32'h3b9e2e9b),
	.w4(32'hbbd1c35e),
	.w5(32'hba2b83a0),
	.w6(32'h3b676f57),
	.w7(32'hbbc64646),
	.w8(32'hbb265924),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef1640),
	.w1(32'hba253602),
	.w2(32'hbb3ef464),
	.w3(32'h3a40bdfa),
	.w4(32'h39f442cc),
	.w5(32'hbb82922a),
	.w6(32'h3b4396c3),
	.w7(32'hbab2168f),
	.w8(32'hbb7ed4a9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbcdd5),
	.w1(32'hba2d5bae),
	.w2(32'h3a3a2c22),
	.w3(32'hbaf5f365),
	.w4(32'hbb7e5b55),
	.w5(32'hbb04722c),
	.w6(32'hbb26409e),
	.w7(32'hbb4944f4),
	.w8(32'h3a137287),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa86763),
	.w1(32'hbb2e89e6),
	.w2(32'h3a2e0c74),
	.w3(32'hbb0da8c4),
	.w4(32'hbba04e22),
	.w5(32'hba106ada),
	.w6(32'hbb08d1bb),
	.w7(32'hbb5584e7),
	.w8(32'hbb3c0491),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391067a5),
	.w1(32'hbadc8052),
	.w2(32'h39f5c8a1),
	.w3(32'h3ab86cb8),
	.w4(32'hba6bcaf2),
	.w5(32'hbb099513),
	.w6(32'hbb5c07b2),
	.w7(32'hbb3991ff),
	.w8(32'hba964e50),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dc319),
	.w1(32'h3b0daa1c),
	.w2(32'h3a9f290f),
	.w3(32'hba7eb24f),
	.w4(32'hbb4d7df3),
	.w5(32'hbb519a67),
	.w6(32'hbabb4394),
	.w7(32'hbbb5de5b),
	.w8(32'hbbd779ef),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada89fc),
	.w1(32'h39ef6c98),
	.w2(32'h3a8a8a76),
	.w3(32'hbaf06b50),
	.w4(32'hbb3f0518),
	.w5(32'hbb969ac6),
	.w6(32'h3b0520c4),
	.w7(32'hbba39fb1),
	.w8(32'hbae527a0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34fe25),
	.w1(32'hbbb64ed2),
	.w2(32'hbae8462f),
	.w3(32'hbbdaa5d7),
	.w4(32'hbb376e7a),
	.w5(32'hbaf9d611),
	.w6(32'hbb262046),
	.w7(32'h3b34c83d),
	.w8(32'hbb65b1c2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8b100),
	.w1(32'h3b9483f1),
	.w2(32'h3b068d59),
	.w3(32'h3a236127),
	.w4(32'hba479d85),
	.w5(32'hbbbef185),
	.w6(32'hbb185478),
	.w7(32'hbb45c4ea),
	.w8(32'hbb9431b4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d355c),
	.w1(32'hb8f42cde),
	.w2(32'hbb513130),
	.w3(32'h3b87eef7),
	.w4(32'hb99710b3),
	.w5(32'hbba938b2),
	.w6(32'hba1814ab),
	.w7(32'hba9c3443),
	.w8(32'hbb04b864),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40ec11),
	.w1(32'hbb25f958),
	.w2(32'h3b27997e),
	.w3(32'h396df030),
	.w4(32'hba0acfba),
	.w5(32'h3b0b05c9),
	.w6(32'h3a807d41),
	.w7(32'hbb3f4fd3),
	.w8(32'hbb803421),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3310fe),
	.w1(32'hbbae3208),
	.w2(32'hb9f81526),
	.w3(32'h389e545c),
	.w4(32'hbb519bb4),
	.w5(32'h3aea5ce8),
	.w6(32'hba1eac54),
	.w7(32'hbba0552e),
	.w8(32'h3a55322a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf26bf2),
	.w1(32'hbae8adc8),
	.w2(32'hbb71552e),
	.w3(32'h3969f5bb),
	.w4(32'hbb0e38fa),
	.w5(32'hbb59aaf8),
	.w6(32'h3b02b892),
	.w7(32'hbaea264a),
	.w8(32'h3a9f02b5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c4325),
	.w1(32'hbaa5e443),
	.w2(32'hba8ee13d),
	.w3(32'hba2e7c78),
	.w4(32'hbb31e606),
	.w5(32'hbb7eca60),
	.w6(32'h3b670827),
	.w7(32'hbb4a73f3),
	.w8(32'h3b6c2e06),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1ff40),
	.w1(32'h3bc30d8c),
	.w2(32'h3ba18a4d),
	.w3(32'h3b3b9352),
	.w4(32'hba747fbc),
	.w5(32'h39b26a55),
	.w6(32'h3b8df5b4),
	.w7(32'hbb68277b),
	.w8(32'h3aa43b12),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c55132),
	.w1(32'h3b1ac45b),
	.w2(32'h3b7af542),
	.w3(32'h3ab9f624),
	.w4(32'hbb329dbb),
	.w5(32'hbab7929f),
	.w6(32'hbb1868d3),
	.w7(32'hb8ea6493),
	.w8(32'h3b464ac3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88c61c),
	.w1(32'hbaf7db8c),
	.w2(32'h3a836edb),
	.w3(32'h3baf088b),
	.w4(32'hba486a6c),
	.w5(32'h3b215168),
	.w6(32'h3bc9a33e),
	.w7(32'hb98ca24c),
	.w8(32'h3b07d5ba),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a110f1f),
	.w1(32'h3b1472b4),
	.w2(32'hba7a600f),
	.w3(32'hb9c61abf),
	.w4(32'h3c7e0345),
	.w5(32'h3b7a150f),
	.w6(32'hb92f33b0),
	.w7(32'h3b8a07fe),
	.w8(32'h3c8286de),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5279f2),
	.w1(32'h3a9d1d84),
	.w2(32'hbb88658d),
	.w3(32'hbb5909d9),
	.w4(32'hb9af71e4),
	.w5(32'h3a34c484),
	.w6(32'h3bd771c4),
	.w7(32'hba92cbaa),
	.w8(32'hba5a25d8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81c741),
	.w1(32'hbb0e915f),
	.w2(32'hbc115e0f),
	.w3(32'h3aefc3d9),
	.w4(32'hbb5f6bf6),
	.w5(32'hbaadae1c),
	.w6(32'hbab53b42),
	.w7(32'h3784168a),
	.w8(32'hbb11396e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f6af9),
	.w1(32'h3b6d5197),
	.w2(32'h3b70a473),
	.w3(32'hbbca4bac),
	.w4(32'h3b4fdc79),
	.w5(32'h3b5c2705),
	.w6(32'hbb91b9d4),
	.w7(32'h3a215048),
	.w8(32'h3b11ee24),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109be7),
	.w1(32'h3ae543fc),
	.w2(32'h3b68cb1b),
	.w3(32'hba1a40f2),
	.w4(32'hba1fec72),
	.w5(32'hba0493b7),
	.w6(32'hba5bd026),
	.w7(32'h3a8a5405),
	.w8(32'h3a510691),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9672c),
	.w1(32'hbb306636),
	.w2(32'hbb353c98),
	.w3(32'h3ba7c70c),
	.w4(32'hbabc02fa),
	.w5(32'hb942cfbc),
	.w6(32'h38d1964c),
	.w7(32'hbaf22aeb),
	.w8(32'hbb97b900),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a9298),
	.w1(32'h3af7f881),
	.w2(32'h3b0da4f0),
	.w3(32'h39930d99),
	.w4(32'hbb11aa60),
	.w5(32'h3a37d1be),
	.w6(32'h394c0823),
	.w7(32'hb9bbce64),
	.w8(32'hba2c135a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a031664),
	.w1(32'h3aa517db),
	.w2(32'h3b39d0df),
	.w3(32'h3a37e4d5),
	.w4(32'h3aba4cfa),
	.w5(32'h3b227a8b),
	.w6(32'h3a968bc9),
	.w7(32'h3aa2afe1),
	.w8(32'h3b3ff34a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a9783),
	.w1(32'hbb3c001c),
	.w2(32'hbb474e84),
	.w3(32'h3b214f3c),
	.w4(32'hbba00db2),
	.w5(32'hbb168359),
	.w6(32'h3ae51520),
	.w7(32'hb9ce9c89),
	.w8(32'h3a0a2bcb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f9a63),
	.w1(32'h3bce58b2),
	.w2(32'h3aa7c365),
	.w3(32'hbaf4a6c9),
	.w4(32'hb95ab835),
	.w5(32'hbb7deead),
	.w6(32'hba14698d),
	.w7(32'hbae65244),
	.w8(32'hbb8b6af7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f09372),
	.w1(32'hbb406274),
	.w2(32'h3a9c8d54),
	.w3(32'h39606c32),
	.w4(32'h3bdd613a),
	.w5(32'hbb2ea4a1),
	.w6(32'hbba229b5),
	.w7(32'h3bcc4674),
	.w8(32'h3b480ebf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0d40e),
	.w1(32'hbb197a19),
	.w2(32'h3b7f15fb),
	.w3(32'hbad968b7),
	.w4(32'hbac6ad7e),
	.w5(32'hbab705d8),
	.w6(32'hbb76bcde),
	.w7(32'hbae65518),
	.w8(32'hbbd094ff),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb06cd5),
	.w1(32'hb926b6e2),
	.w2(32'h39691d26),
	.w3(32'h3b816bc7),
	.w4(32'hb89f8705),
	.w5(32'h390b0e93),
	.w6(32'hbb19f205),
	.w7(32'hba614545),
	.w8(32'hba67ebb9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb531e86f),
	.w1(32'hb507a74e),
	.w2(32'h351218db),
	.w3(32'h35d2dfbb),
	.w4(32'h36a00d2d),
	.w5(32'hb40d27f6),
	.w6(32'hb45ac164),
	.w7(32'h370a4a81),
	.w8(32'h369c111e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb625418d),
	.w1(32'hb5f4a93e),
	.w2(32'h351c0284),
	.w3(32'hb6909a92),
	.w4(32'hb5c9afee),
	.w5(32'h366df11e),
	.w6(32'h3636afaa),
	.w7(32'h36e1f38f),
	.w8(32'h371b1f6a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dc7dbe),
	.w1(32'h37274b3b),
	.w2(32'h371a3ec3),
	.w3(32'hb5f5f4ac),
	.w4(32'h371b18f5),
	.w5(32'h369b530a),
	.w6(32'h36fe3a4c),
	.w7(32'h36f5b99b),
	.w8(32'h378b020d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e32aa),
	.w1(32'hb8c095de),
	.w2(32'hb918ebfb),
	.w3(32'h38a5633f),
	.w4(32'h383c21ab),
	.w5(32'h37098ae1),
	.w6(32'h38fe3d59),
	.w7(32'h37ea12ce),
	.w8(32'hb8106fde),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36971c4c),
	.w1(32'hb3fa2f55),
	.w2(32'hb67aa765),
	.w3(32'h36c9e83a),
	.w4(32'h36ddf105),
	.w5(32'h3687abb1),
	.w6(32'h3790969a),
	.w7(32'h373c3730),
	.w8(32'h36ada410),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d9e35),
	.w1(32'hb9a0b3b9),
	.w2(32'hb97e4ab1),
	.w3(32'hb9ffdaba),
	.w4(32'hb97970dd),
	.w5(32'hb9883d8c),
	.w6(32'h397f7ee4),
	.w7(32'h36bdf439),
	.w8(32'hb95c7917),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43a137),
	.w1(32'hb9fb499a),
	.w2(32'hb50c6a2c),
	.w3(32'hba62e1c4),
	.w4(32'h39a13635),
	.w5(32'h394cbef4),
	.w6(32'hb9a4d584),
	.w7(32'hb8f9a494),
	.w8(32'h37dd5c23),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81b17f),
	.w1(32'hba108fd6),
	.w2(32'hba1cb0f3),
	.w3(32'hba8380bb),
	.w4(32'hba5d04c6),
	.w5(32'hba707831),
	.w6(32'hba143eaf),
	.w7(32'hba6e6ea3),
	.w8(32'hbaa38e8f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b8d77),
	.w1(32'hba049c51),
	.w2(32'hb95095ed),
	.w3(32'hb9ac457b),
	.w4(32'hb961ce8a),
	.w5(32'h390b4e37),
	.w6(32'hb8e93c6c),
	.w7(32'hb8d551b7),
	.w8(32'hb8f4f026),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2e8dc),
	.w1(32'hb8a50205),
	.w2(32'hb8119b1c),
	.w3(32'hba1c483a),
	.w4(32'hb9428118),
	.w5(32'hb9c99200),
	.w6(32'hb85e761b),
	.w7(32'hb960e366),
	.w8(32'hb9f60c21),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f0eba),
	.w1(32'h3737f984),
	.w2(32'h38c02754),
	.w3(32'hb90184cf),
	.w4(32'h385c65c8),
	.w5(32'h39076627),
	.w6(32'hb9d085b4),
	.w7(32'hb927a247),
	.w8(32'hb9044df7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba198f41),
	.w1(32'hb9f253bd),
	.w2(32'hba13cd07),
	.w3(32'hba027ca2),
	.w4(32'hb9f65a98),
	.w5(32'hba0a5c5f),
	.w6(32'hb93b1353),
	.w7(32'hb9e1fed0),
	.w8(32'hba2265cc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b0eeac),
	.w1(32'hb60c4061),
	.w2(32'hb4ca7f76),
	.w3(32'hb582b6e2),
	.w4(32'hb4eaf17c),
	.w5(32'h3520b392),
	.w6(32'h34ee980a),
	.w7(32'h35443e6e),
	.w8(32'h36353ba6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb700cbc0),
	.w1(32'hb72eb5a8),
	.w2(32'hb646e015),
	.w3(32'hb74e92f6),
	.w4(32'hb742593e),
	.w5(32'hb6a617ed),
	.w6(32'hb6cc7698),
	.w7(32'hb6dec36d),
	.w8(32'hb7103c3c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3669b046),
	.w1(32'h3684a8d1),
	.w2(32'h363e6f28),
	.w3(32'h368416c0),
	.w4(32'h3659f384),
	.w5(32'h3618c61a),
	.w6(32'h36a0c9ab),
	.w7(32'h36556eda),
	.w8(32'h35c8f0fd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372ff61a),
	.w1(32'h373a9c3b),
	.w2(32'h374283de),
	.w3(32'h3759e485),
	.w4(32'h3729fda0),
	.w5(32'h371291a2),
	.w6(32'hb6dbd373),
	.w7(32'hb70e37dc),
	.w8(32'hb7b2f318),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77c272),
	.w1(32'hba846625),
	.w2(32'hba8413c2),
	.w3(32'hba82837e),
	.w4(32'hba0c50a1),
	.w5(32'hba2e9f99),
	.w6(32'hbb011d44),
	.w7(32'hba739870),
	.w8(32'hb8139c19),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82db818),
	.w1(32'h37994a86),
	.w2(32'h38146216),
	.w3(32'h38374b43),
	.w4(32'h3911b03e),
	.w5(32'h37cd00c8),
	.w6(32'h371022c5),
	.w7(32'h3831a37f),
	.w8(32'h36865c5b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62cc79),
	.w1(32'hb98193cb),
	.w2(32'h382a2425),
	.w3(32'hba9fffd8),
	.w4(32'hba1df033),
	.w5(32'h390982c4),
	.w6(32'hba948ad0),
	.w7(32'hb9a94130),
	.w8(32'hb78546ea),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba704324),
	.w1(32'hb9b8b879),
	.w2(32'hba0c4425),
	.w3(32'hba51eaad),
	.w4(32'hb917544b),
	.w5(32'hba115d07),
	.w6(32'hb9d120ee),
	.w7(32'hb9c90027),
	.w8(32'hba21d743),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399059e1),
	.w1(32'h38d11599),
	.w2(32'h3894f5e7),
	.w3(32'h3995f885),
	.w4(32'h39010077),
	.w5(32'hb7fd09a0),
	.w6(32'h3958c485),
	.w7(32'h37788dce),
	.w8(32'hb91fbfe5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86d592e),
	.w1(32'h372477e7),
	.w2(32'h38fca47a),
	.w3(32'hb9e0b24c),
	.w4(32'h39aa9c43),
	.w5(32'h3998038c),
	.w6(32'hb8cad9ff),
	.w7(32'h3860ce15),
	.w8(32'h3938f69f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98928e5),
	.w1(32'hb8ea7583),
	.w2(32'hb93aa4eb),
	.w3(32'hb9e5006f),
	.w4(32'hb9160278),
	.w5(32'hb8df985d),
	.w6(32'hb9f55afc),
	.w7(32'hb9cdd84f),
	.w8(32'hb9b09013),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88da27),
	.w1(32'hba8a54c9),
	.w2(32'hba1590ed),
	.w3(32'hba870559),
	.w4(32'hb9f78a5d),
	.w5(32'h3875b3ef),
	.w6(32'hb9e96c8b),
	.w7(32'hb91d65b6),
	.w8(32'hb89a0820),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba029a92),
	.w1(32'hb9be0369),
	.w2(32'hb9ccff79),
	.w3(32'hbaae987c),
	.w4(32'hba34e2f4),
	.w5(32'hb9e03e9b),
	.w6(32'hba86a1a6),
	.w7(32'hba37da7d),
	.w8(32'hb9d90a04),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba191841),
	.w1(32'hb96ca457),
	.w2(32'h381e0a46),
	.w3(32'hb9e389f5),
	.w4(32'h3947f300),
	.w5(32'h3976a072),
	.w6(32'hb9b09096),
	.w7(32'hb91382b9),
	.w8(32'hb945821d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379abdfe),
	.w1(32'h37745d8a),
	.w2(32'hb7e67845),
	.w3(32'hb5c8efd0),
	.w4(32'hb7fa7f69),
	.w5(32'hb8812236),
	.w6(32'hb8dc7e92),
	.w7(32'hb84e3f2e),
	.w8(32'hb8891361),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc86ea),
	.w1(32'hba8b0e67),
	.w2(32'hba884ac6),
	.w3(32'hbac725a9),
	.w4(32'hba8e413f),
	.w5(32'hba1de438),
	.w6(32'hba909b43),
	.w7(32'hba925060),
	.w8(32'hba9a135f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38838f38),
	.w1(32'hba1672cb),
	.w2(32'hba8b6eb4),
	.w3(32'hba7ace00),
	.w4(32'hb922fd2d),
	.w5(32'hba9ad67b),
	.w6(32'hb9fc9333),
	.w7(32'hb9c28328),
	.w8(32'hba871de8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad465fd),
	.w1(32'hba8547cd),
	.w2(32'h39938cb1),
	.w3(32'hbaf26ee3),
	.w4(32'hba2eb4b1),
	.w5(32'hb8e34e68),
	.w6(32'hba019977),
	.w7(32'hba595bd5),
	.w8(32'hbaacd9de),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1a04b),
	.w1(32'hbad056b4),
	.w2(32'hbb245614),
	.w3(32'hbad11718),
	.w4(32'h396176af),
	.w5(32'hbabe4313),
	.w6(32'hbb1434ef),
	.w7(32'hb8909fc7),
	.w8(32'hba97c10c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc1b81),
	.w1(32'hba327bfe),
	.w2(32'hb9c42801),
	.w3(32'hbadb781a),
	.w4(32'hba6b217e),
	.w5(32'hb97f9b5a),
	.w6(32'hbaed39ab),
	.w7(32'hbab01caf),
	.w8(32'hba976c85),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b0935),
	.w1(32'hba7bda96),
	.w2(32'hba93b297),
	.w3(32'hbae3afbb),
	.w4(32'hb9f08eae),
	.w5(32'hb9bdf055),
	.w6(32'hba5eca4f),
	.w7(32'hba3b8ffd),
	.w8(32'hba8611ff),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78d4ce2),
	.w1(32'hb5d35bd3),
	.w2(32'hb6ba6230),
	.w3(32'hb6fdca6f),
	.w4(32'h364701ff),
	.w5(32'h37ff6cc9),
	.w6(32'hb6cfefea),
	.w7(32'h37cf02d1),
	.w8(32'h381c910c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad06b49),
	.w1(32'hba8d5820),
	.w2(32'hba147766),
	.w3(32'hba9ed203),
	.w4(32'hba17c92c),
	.w5(32'hb9948f83),
	.w6(32'hba57ffca),
	.w7(32'hb6db812e),
	.w8(32'hbaaa199a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e43b5f),
	.w1(32'hb8e4a91b),
	.w2(32'hb89ecc82),
	.w3(32'h39429bad),
	.w4(32'h37991815),
	.w5(32'hba47cd96),
	.w6(32'h3948dad1),
	.w7(32'h3851f8a0),
	.w8(32'hb89c8fa1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38153e0a),
	.w1(32'h35ef5caa),
	.w2(32'hb7000f45),
	.w3(32'h37ac4c69),
	.w4(32'hb6ce10cc),
	.w5(32'hb7029532),
	.w6(32'h37f785f6),
	.w7(32'h36de9040),
	.w8(32'h375ef1c4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884a913),
	.w1(32'hb786c3d4),
	.w2(32'h37137143),
	.w3(32'hb7ea2385),
	.w4(32'hb81190a5),
	.w5(32'hb6247106),
	.w6(32'hb94ae07f),
	.w7(32'hb91135d6),
	.w8(32'hb7a62ace),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9df0a2),
	.w1(32'hba4a55df),
	.w2(32'hba1700c9),
	.w3(32'hbaa09c2e),
	.w4(32'hba320f10),
	.w5(32'hb9ae0eb3),
	.w6(32'hba955202),
	.w7(32'hba640a6a),
	.w8(32'hba45579b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba368b64),
	.w1(32'hb941e4ad),
	.w2(32'h39458a64),
	.w3(32'hba683ff0),
	.w4(32'hb94463ce),
	.w5(32'h395bc094),
	.w6(32'hba9d632b),
	.w7(32'hba18e0eb),
	.w8(32'hb9d58356),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f79a60),
	.w1(32'hba0605e5),
	.w2(32'hba09e522),
	.w3(32'hba6f77f4),
	.w4(32'hba0df2c3),
	.w5(32'hb9d58597),
	.w6(32'hba25e8a3),
	.w7(32'hb9992697),
	.w8(32'hba235b73),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bc7fc),
	.w1(32'hba16d865),
	.w2(32'hb9e02cee),
	.w3(32'hb9e7f4ea),
	.w4(32'hb9b7f2d1),
	.w5(32'hb9e98e40),
	.w6(32'hba060937),
	.w7(32'hb9b5c109),
	.w8(32'hba178a05),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980a86b),
	.w1(32'h39a61d1e),
	.w2(32'h3993120a),
	.w3(32'h398d600d),
	.w4(32'h39941c74),
	.w5(32'h38937a2a),
	.w6(32'h383bd5f3),
	.w7(32'h3857e642),
	.w8(32'h37787ba8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bbdf1),
	.w1(32'hb9ace5a9),
	.w2(32'hb915351a),
	.w3(32'hba3f1f5b),
	.w4(32'hb9ce353d),
	.w5(32'h368972a5),
	.w6(32'hba15878a),
	.w7(32'hb9c62478),
	.w8(32'h38bfca8e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d691a2),
	.w1(32'hb8a90d75),
	.w2(32'h3905d6de),
	.w3(32'hba0b69ee),
	.w4(32'hb907bc51),
	.w5(32'h390a1d03),
	.w6(32'hba511b6c),
	.w7(32'hb9cf7cad),
	.w8(32'hb96b9c96),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb777fb8b),
	.w1(32'hb6d171f5),
	.w2(32'h329b2869),
	.w3(32'hb7890bfd),
	.w4(32'hb6d341dd),
	.w5(32'h3606001a),
	.w6(32'hb7653566),
	.w7(32'hb6d2c306),
	.w8(32'hb5ca9406),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e1372),
	.w1(32'hb7c92247),
	.w2(32'h377dfb42),
	.w3(32'hb84c25df),
	.w4(32'hb7f35025),
	.w5(32'h3776eb38),
	.w6(32'hb81f22b5),
	.w7(32'hb7f3176b),
	.w8(32'hb68fe714),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb793d169),
	.w1(32'hb874a0dd),
	.w2(32'hb8346778),
	.w3(32'h3825f1c7),
	.w4(32'h3829b85e),
	.w5(32'h38524f5b),
	.w6(32'hb6f49287),
	.w7(32'hb69a74c9),
	.w8(32'hb7aa3c3a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3781c05c),
	.w1(32'h3833fa7a),
	.w2(32'h383af80f),
	.w3(32'h366e6c1d),
	.w4(32'h378ddb89),
	.w5(32'h37fbe9b5),
	.w6(32'h375b602e),
	.w7(32'h38154bcb),
	.w8(32'h382250f3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0602af),
	.w1(32'hb9030519),
	.w2(32'h37da8f33),
	.w3(32'hba0c4df4),
	.w4(32'hb86ec4e6),
	.w5(32'h39013999),
	.w6(32'hba44a547),
	.w7(32'hb9d6e5d7),
	.w8(32'hb9a51e81),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ecf58),
	.w1(32'hb7b5ad3b),
	.w2(32'h39051c48),
	.w3(32'hb83926db),
	.w4(32'h384184c4),
	.w5(32'h3950cf23),
	.w6(32'h3810846c),
	.w7(32'h394c9207),
	.w8(32'h39473cb7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f04c4),
	.w1(32'hb9c35f38),
	.w2(32'hb9dcffbc),
	.w3(32'hb8daa342),
	.w4(32'hb9449fd8),
	.w5(32'hb9f64679),
	.w6(32'hba11d671),
	.w7(32'hb9553638),
	.w8(32'hb9bb7da2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9860c1f),
	.w1(32'hb88c2c94),
	.w2(32'hb9916975),
	.w3(32'hba212373),
	.w4(32'hb95f58a3),
	.w5(32'hb9d8931a),
	.w6(32'hb9ffbb04),
	.w7(32'hba0149de),
	.w8(32'hba575186),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369aee7a),
	.w1(32'hb60c0d07),
	.w2(32'hb5a4704d),
	.w3(32'h350a7a62),
	.w4(32'hb591f9dd),
	.w5(32'h30c6f070),
	.w6(32'h353a1d02),
	.w7(32'h35a5a87d),
	.w8(32'h35981528),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a37cb6),
	.w1(32'hb7ce4871),
	.w2(32'hb81d3e39),
	.w3(32'hb6e0f586),
	.w4(32'hb8043ba6),
	.w5(32'hb7cf5439),
	.w6(32'h37ebf386),
	.w7(32'hb669cca1),
	.w8(32'h3649a6cd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a4e52a),
	.w1(32'h365367f7),
	.w2(32'hb3f55cbe),
	.w3(32'h37107264),
	.w4(32'h361ac3db),
	.w5(32'hb5ac1e69),
	.w6(32'h36e550cb),
	.w7(32'h369bf70b),
	.w8(32'h369bb9ef),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f6f19),
	.w1(32'hb91e5f90),
	.w2(32'hb9912d7b),
	.w3(32'hba1467cf),
	.w4(32'hb9b29749),
	.w5(32'hb9ba4781),
	.w6(32'hb9331a43),
	.w7(32'hb9adaf5f),
	.w8(32'hb9f7775e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983de28),
	.w1(32'h3a0be967),
	.w2(32'hb951f80b),
	.w3(32'h3966bc84),
	.w4(32'hb8f5c0f7),
	.w5(32'hba1268cd),
	.w6(32'hb772d3f0),
	.w7(32'hb909dba7),
	.w8(32'hb5b0dc2e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba928c35),
	.w1(32'hba118638),
	.w2(32'hba25a159),
	.w3(32'hba9f54d7),
	.w4(32'hba40db8f),
	.w5(32'hb8f21406),
	.w6(32'hba15d7c6),
	.w7(32'hba5bd0a0),
	.w8(32'hba437e9f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b004cb),
	.w1(32'hb6d9fea2),
	.w2(32'hb85fd07d),
	.w3(32'h36a842cd),
	.w4(32'hb6ec9451),
	.w5(32'hb8236223),
	.w6(32'h382f4dcd),
	.w7(32'h3783dc32),
	.w8(32'hb7fc422b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3e44f41),
	.w1(32'h36eaa341),
	.w2(32'hb813c7e9),
	.w3(32'h38e6c3e4),
	.w4(32'hb85fbd02),
	.w5(32'hb888e022),
	.w6(32'h38ddb99a),
	.w7(32'h37e98283),
	.w8(32'hb9018e96),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d2d93b),
	.w1(32'hb96aa493),
	.w2(32'hb70c16c0),
	.w3(32'hb94f66a0),
	.w4(32'hb942e153),
	.w5(32'hb91b4641),
	.w6(32'hb996b891),
	.w7(32'hb9499f63),
	.w8(32'hb951f237),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcbc36),
	.w1(32'hb8e21d8b),
	.w2(32'hb8b38c11),
	.w3(32'hb9b1bda4),
	.w4(32'hb9341949),
	.w5(32'hb88bc6ec),
	.w6(32'hb9d054fb),
	.w7(32'hb9b3ef72),
	.w8(32'hb969ae92),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1714a7),
	.w1(32'hb8e2c4c3),
	.w2(32'h390ae71e),
	.w3(32'hba5fc33f),
	.w4(32'hb9b93edc),
	.w5(32'hb9b27d49),
	.w6(32'hba8421c5),
	.w7(32'hb9cf9981),
	.w8(32'hb93bf752),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78464f),
	.w1(32'hba2b6c4e),
	.w2(32'hba65d6f9),
	.w3(32'hba8ba2e8),
	.w4(32'hba2d5b27),
	.w5(32'hb9c107bf),
	.w6(32'hb8714327),
	.w7(32'hba355df7),
	.w8(32'hba340e05),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba211be2),
	.w1(32'hb9dc7e6e),
	.w2(32'hb97913e3),
	.w3(32'hba2ea460),
	.w4(32'hb9b2bb75),
	.w5(32'hb9727f9b),
	.w6(32'hba7da458),
	.w7(32'hb9e4bd6d),
	.w8(32'hba0439d9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3a9f6),
	.w1(32'hba3d1f28),
	.w2(32'hba1b0774),
	.w3(32'hbab84265),
	.w4(32'hb9bee1ea),
	.w5(32'hb9ff2fc9),
	.w6(32'hbad2df30),
	.w7(32'hbab4235c),
	.w8(32'hba1ac808),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aa2ed),
	.w1(32'hb9e20f40),
	.w2(32'hba0e1827),
	.w3(32'hba4fa058),
	.w4(32'hb9e5402e),
	.w5(32'hb9c7903c),
	.w6(32'hb8aa8883),
	.w7(32'hb984a52c),
	.w8(32'hba373e81),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c74d3e),
	.w1(32'hb89b9e59),
	.w2(32'h38470c71),
	.w3(32'hba19a574),
	.w4(32'hb8091ba3),
	.w5(32'h38cd3ce5),
	.w6(32'hba075583),
	.w7(32'hb9ddbc35),
	.w8(32'hb9b01656),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37f971),
	.w1(32'hba0d7bed),
	.w2(32'hb932821a),
	.w3(32'hba91a0a8),
	.w4(32'hb9e32847),
	.w5(32'h38a416f1),
	.w6(32'hba1e52d0),
	.w7(32'hb9ca229f),
	.w8(32'hb96f6af9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96429da),
	.w1(32'hb8924f2f),
	.w2(32'hb777ae53),
	.w3(32'hb95838db),
	.w4(32'hb86b8193),
	.w5(32'h37a45cbe),
	.w6(32'hb9959e48),
	.w7(32'hb9224516),
	.w8(32'hb910d191),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1260c7),
	.w1(32'hba0bd25f),
	.w2(32'hba49b84a),
	.w3(32'hba88bcea),
	.w4(32'hb9cf3058),
	.w5(32'hb995e57f),
	.w6(32'hbab9b255),
	.w7(32'hba279d8e),
	.w8(32'hba4e2424),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32c90d),
	.w1(32'hb9f55cab),
	.w2(32'hb8b99e6f),
	.w3(32'hba7339a3),
	.w4(32'hb96ae1cc),
	.w5(32'h3984942f),
	.w6(32'hba388376),
	.w7(32'hb9cdf68f),
	.w8(32'h393e9f35),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb628a5a1),
	.w1(32'hb62457ea),
	.w2(32'hb6a38a3a),
	.w3(32'hb6464dd7),
	.w4(32'hb6b7e080),
	.w5(32'hb6b931f6),
	.w6(32'h35170869),
	.w7(32'hb57b4dc9),
	.w8(32'hb6536e73),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37741e8d),
	.w1(32'h37c710a0),
	.w2(32'hb5ad52f4),
	.w3(32'h378f8520),
	.w4(32'h37b9f7a8),
	.w5(32'h37a32522),
	.w6(32'hb7a19c88),
	.w7(32'h37450e71),
	.w8(32'h37823145),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ae9fdd),
	.w1(32'h38c16018),
	.w2(32'h38646628),
	.w3(32'h3904a796),
	.w4(32'h39145fb5),
	.w5(32'h37b95601),
	.w6(32'h38f4e9ee),
	.w7(32'h38ba3dbf),
	.w8(32'h352b4a61),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94188f),
	.w1(32'hba6567f7),
	.w2(32'hb9f4710f),
	.w3(32'hba4a9f05),
	.w4(32'hb9c47beb),
	.w5(32'hb9402684),
	.w6(32'hba6fc2fb),
	.w7(32'hb9fafdf7),
	.w8(32'hb9a06d03),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac07de),
	.w1(32'hba335cb4),
	.w2(32'hba3a8c22),
	.w3(32'hb8cb1b19),
	.w4(32'hba514dd7),
	.w5(32'hb9964f04),
	.w6(32'hb8610517),
	.w7(32'hba020450),
	.w8(32'hba953251),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61ebc45),
	.w1(32'hb5becdda),
	.w2(32'h35e259b7),
	.w3(32'hb5e6b3c0),
	.w4(32'hb550d487),
	.w5(32'h350a6919),
	.w6(32'h35a71b67),
	.w7(32'h33e661be),
	.w8(32'h357f03b4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fffdf),
	.w1(32'hb9c4ddf5),
	.w2(32'hb9b81a36),
	.w3(32'hba8d44c4),
	.w4(32'hb9f18b5f),
	.w5(32'hb8fefc79),
	.w6(32'hba862b33),
	.w7(32'hba19c395),
	.w8(32'hba2939b0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22ca79),
	.w1(32'hb9d731de),
	.w2(32'hb9b27a38),
	.w3(32'hba45e059),
	.w4(32'hba14fddd),
	.w5(32'hb9f0f018),
	.w6(32'hba763c69),
	.w7(32'hba44d192),
	.w8(32'hba39d406),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99eb90),
	.w1(32'hb905d2b3),
	.w2(32'hba191f84),
	.w3(32'hbab5a0e6),
	.w4(32'hba6abef8),
	.w5(32'hba8fcd12),
	.w6(32'hba477e65),
	.w7(32'hba187aee),
	.w8(32'hba73e33d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a8f4e3),
	.w1(32'hb907785b),
	.w2(32'h386035da),
	.w3(32'hb9276f99),
	.w4(32'h378c8b1d),
	.w5(32'h39618ddf),
	.w6(32'hba04c6e9),
	.w7(32'hba0dd92c),
	.w8(32'hb9a5bcfa),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999493c),
	.w1(32'hb86592c6),
	.w2(32'h39a4a2a9),
	.w3(32'hba0ad2cb),
	.w4(32'hb948c5d7),
	.w5(32'h39de2295),
	.w6(32'h39a83677),
	.w7(32'h3988e6f6),
	.w8(32'h3991ac6c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386e15cf),
	.w1(32'h385b6b47),
	.w2(32'h38396500),
	.w3(32'h38c2b942),
	.w4(32'h389a5d45),
	.w5(32'h37abf680),
	.w6(32'h38a47cc5),
	.w7(32'h386c8645),
	.w8(32'h37ea676b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e0bcb),
	.w1(32'h39692365),
	.w2(32'h39c1f1bb),
	.w3(32'hb948020d),
	.w4(32'h398b3686),
	.w5(32'h39b1e0e1),
	.w6(32'hb9d5bd78),
	.w7(32'hb711be95),
	.w8(32'h3889d700),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82bdcb),
	.w1(32'hba6aaf85),
	.w2(32'hb961fa1e),
	.w3(32'hbabfc2c7),
	.w4(32'hb9621743),
	.w5(32'hb9049fef),
	.w6(32'hb9c88066),
	.w7(32'h39779fcf),
	.w8(32'hb90502fe),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f46d4),
	.w1(32'h395460b1),
	.w2(32'h392e8818),
	.w3(32'h397ef0cc),
	.w4(32'h39246b66),
	.w5(32'h38e4ca6c),
	.w6(32'h386ef67d),
	.w7(32'hb82887d0),
	.w8(32'hb80442a1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b685cc),
	.w1(32'hb8e3520d),
	.w2(32'hb8f61df8),
	.w3(32'hb94c1759),
	.w4(32'hb8cd5f0b),
	.w5(32'hb744a658),
	.w6(32'hb82d44e0),
	.w7(32'hb8d80432),
	.w8(32'hb95ea71d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72f440b),
	.w1(32'hb712b4a9),
	.w2(32'h35094e9b),
	.w3(32'hb780179b),
	.w4(32'hb67c2348),
	.w5(32'h35486089),
	.w6(32'hb727e3c9),
	.w7(32'hb79128f8),
	.w8(32'hb71b0cde),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e9b83),
	.w1(32'hb9fd4e65),
	.w2(32'hb9e6d707),
	.w3(32'hba5e1c76),
	.w4(32'hb9c3716f),
	.w5(32'hb9a7e101),
	.w6(32'hb93a5d70),
	.w7(32'hb9b87e7d),
	.w8(32'hba0663fa),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382367d2),
	.w1(32'h369a4931),
	.w2(32'hb79ed2ec),
	.w3(32'h387fe9df),
	.w4(32'h388860ed),
	.w5(32'hb7d7a408),
	.w6(32'h38a0cf85),
	.w7(32'h38374635),
	.w8(32'hb7b9755a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aaa71a),
	.w1(32'hb904abbe),
	.w2(32'h387ca5be),
	.w3(32'hb9d52124),
	.w4(32'hb93ebb60),
	.w5(32'h38b4891b),
	.w6(32'hba0cbb01),
	.w7(32'hb9b31b61),
	.w8(32'hb963daf2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d08919),
	.w1(32'h35e30865),
	.w2(32'hb6c285c1),
	.w3(32'hb752c37f),
	.w4(32'hb800dae2),
	.w5(32'hb735d65b),
	.w6(32'h3869ba3d),
	.w7(32'h379ae835),
	.w8(32'hb71d06e0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12629e),
	.w1(32'h39dc8a5a),
	.w2(32'hb56beb8e),
	.w3(32'h3a4569cb),
	.w4(32'h3a0591f0),
	.w5(32'h37271c47),
	.w6(32'h39e0f5a7),
	.w7(32'h396f327d),
	.w8(32'h380cde27),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367c786d),
	.w1(32'h369485a1),
	.w2(32'h3732cac3),
	.w3(32'h366fbf3e),
	.w4(32'h36810e2f),
	.w5(32'h37146b9f),
	.w6(32'h36e6219a),
	.w7(32'h371f4d92),
	.w8(32'h3794e79c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38429712),
	.w1(32'h37cc5022),
	.w2(32'hb7597c20),
	.w3(32'h38a09f52),
	.w4(32'h389477dd),
	.w5(32'h3775e768),
	.w6(32'h39169a95),
	.w7(32'h390b39f9),
	.w8(32'h38a0ee1d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d4759),
	.w1(32'hba29175e),
	.w2(32'hb97d504a),
	.w3(32'hba88328c),
	.w4(32'hb9ca26e0),
	.w5(32'h392626bb),
	.w6(32'hba274b45),
	.w7(32'hb9c7422c),
	.w8(32'hb94e991c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39c8f2),
	.w1(32'hb8b2d2cc),
	.w2(32'hb875248b),
	.w3(32'hba837ec7),
	.w4(32'hb90c74f9),
	.w5(32'h39a22793),
	.w6(32'hbaa9cfb0),
	.w7(32'hb9d2bf8a),
	.w8(32'hb9431c33),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944bf44),
	.w1(32'h390188ed),
	.w2(32'h3863dc82),
	.w3(32'h399f3f3a),
	.w4(32'h397a939f),
	.w5(32'h3936445c),
	.w6(32'h38977d12),
	.w7(32'h3854128c),
	.w8(32'h389063e0),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba433001),
	.w1(32'hb9865d13),
	.w2(32'hb80dab96),
	.w3(32'hba9e8b51),
	.w4(32'hba1d27e4),
	.w5(32'hb8c80a87),
	.w6(32'hbac9fd5b),
	.w7(32'hba852118),
	.w8(32'hba22046f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902bba8),
	.w1(32'hb8837119),
	.w2(32'hb68ee7b0),
	.w3(32'hb932f2c2),
	.w4(32'hb881125d),
	.w5(32'h380efce9),
	.w6(32'hb8d6eee3),
	.w7(32'hb88d8f4c),
	.w8(32'h383f7a46),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb026b8b),
	.w1(32'hbac7fa9c),
	.w2(32'hbaf827c4),
	.w3(32'hbb169e28),
	.w4(32'hbac56cdd),
	.w5(32'hba28b75a),
	.w6(32'hba5cc43c),
	.w7(32'hbac926c8),
	.w8(32'hba9e2371),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cce6ec),
	.w1(32'hb99968af),
	.w2(32'hb7f079ba),
	.w3(32'hb988369f),
	.w4(32'hb8243523),
	.w5(32'h3849eab2),
	.w6(32'hb99526c5),
	.w7(32'hb97db88f),
	.w8(32'hb974a7fa),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99ba63),
	.w1(32'hba259f9f),
	.w2(32'hb9f5865e),
	.w3(32'hba96536d),
	.w4(32'hba32d022),
	.w5(32'hb90d1b22),
	.w6(32'hba9783e5),
	.w7(32'hba58aa47),
	.w8(32'hba153c22),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb847f378),
	.w1(32'h37e2fc3a),
	.w2(32'h388b8c1f),
	.w3(32'hb80fc6af),
	.w4(32'h3815f7ee),
	.w5(32'h3852b7c5),
	.w6(32'h37eb28ac),
	.w7(32'h382a9208),
	.w8(32'h3890025e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cf242),
	.w1(32'hba016c39),
	.w2(32'hb979fd79),
	.w3(32'hba8233a5),
	.w4(32'hb9a0cc57),
	.w5(32'h397d6df4),
	.w6(32'hba0c23a6),
	.w7(32'hb95868d4),
	.w8(32'hb86e0c7a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a9bee0),
	.w1(32'hb56b363e),
	.w2(32'hb64fb8ab),
	.w3(32'hb4fe5adc),
	.w4(32'hb672c00c),
	.w5(32'hb64210c3),
	.w6(32'h36591792),
	.w7(32'h3609ebff),
	.w8(32'h3647141e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a74918),
	.w1(32'h38dd6689),
	.w2(32'h3904edb6),
	.w3(32'h38abdcc0),
	.w4(32'h38d72229),
	.w5(32'h387119ac),
	.w6(32'hb7534c0c),
	.w7(32'h382947c3),
	.w8(32'h38807e3f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383e27f9),
	.w1(32'h37f6c461),
	.w2(32'h3836a0d3),
	.w3(32'h3734d63c),
	.w4(32'hb75d8b37),
	.w5(32'h35d41d89),
	.w6(32'hb7f689ab),
	.w7(32'hb84c5531),
	.w8(32'hb823845b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba551e33),
	.w1(32'hba5ec188),
	.w2(32'hb9f7e802),
	.w3(32'hbaa548b6),
	.w4(32'hb9eb2a13),
	.w5(32'hba51bb28),
	.w6(32'hba3dc895),
	.w7(32'hba12ce7c),
	.w8(32'hb9f3230a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ae4fb7),
	.w1(32'hb499184b),
	.w2(32'h35a543a7),
	.w3(32'hb6087916),
	.w4(32'hb58c59f7),
	.w5(32'h35266a5e),
	.w6(32'h34f8f4d5),
	.w7(32'h3581756d),
	.w8(32'h35e60dca),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e1f602),
	.w1(32'hb7010b05),
	.w2(32'hb6693ac7),
	.w3(32'hb70b6225),
	.w4(32'h3656b224),
	.w5(32'h371edd40),
	.w6(32'h374971fe),
	.w7(32'h37527ee1),
	.w8(32'h36e75331),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b94e3b),
	.w1(32'h396d97b1),
	.w2(32'h3914726c),
	.w3(32'h38ea0e11),
	.w4(32'h39203986),
	.w5(32'h384f35ee),
	.w6(32'hb7feb638),
	.w7(32'hb85207c9),
	.w8(32'hb8db6802),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e933d),
	.w1(32'hba49cb50),
	.w2(32'hba84ae15),
	.w3(32'hba5b9d39),
	.w4(32'hb8f81f6a),
	.w5(32'hbabe42a6),
	.w6(32'hba1e9dd8),
	.w7(32'hba5d30a6),
	.w8(32'hbaca5b57),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9818540),
	.w1(32'hb8427d3f),
	.w2(32'h390a1052),
	.w3(32'hb95b14da),
	.w4(32'h38337d14),
	.w5(32'h37da39ae),
	.w6(32'hb81ab5f8),
	.w7(32'h382493ab),
	.w8(32'hb9429553),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38763212),
	.w1(32'h37c69954),
	.w2(32'h375c1fbb),
	.w3(32'h3836ba49),
	.w4(32'h373d7f24),
	.w5(32'hb7267fcc),
	.w6(32'h38932643),
	.w7(32'hb7127d23),
	.w8(32'h36c56b3a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb295d74),
	.w1(32'hba677524),
	.w2(32'hba594595),
	.w3(32'hbae4d899),
	.w4(32'hba6fa630),
	.w5(32'h37eff472),
	.w6(32'hba5f18c9),
	.w7(32'hba7c18cf),
	.w8(32'hbab329a3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d1e62),
	.w1(32'h391c54c0),
	.w2(32'h3a168ed5),
	.w3(32'hbae762f3),
	.w4(32'hb9ad4f1c),
	.w5(32'h3a7bd5fb),
	.w6(32'hbace83e2),
	.w7(32'hba513e6b),
	.w8(32'h3a2f9a68),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b26dc9),
	.w1(32'h387050d4),
	.w2(32'h3754e6b8),
	.w3(32'h3841098c),
	.w4(32'h38ea4109),
	.w5(32'hb71ce3c7),
	.w6(32'h393bc702),
	.w7(32'h385b48a3),
	.w8(32'hb8870ca0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4897c72),
	.w1(32'hb75b338c),
	.w2(32'hb751c840),
	.w3(32'h35c7e2bf),
	.w4(32'hb71965a8),
	.w5(32'hb79ea1ea),
	.w6(32'h36fac250),
	.w7(32'h3555aea4),
	.w8(32'hb6f3fbaf),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7118995),
	.w1(32'hb7503a59),
	.w2(32'hb678b86f),
	.w3(32'hb5ed62ef),
	.w4(32'h370d7857),
	.w5(32'h3758583b),
	.w6(32'h36badf2f),
	.w7(32'h3746a566),
	.w8(32'h374f6405),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3638f3b5),
	.w1(32'h349d3e08),
	.w2(32'hb5ed781f),
	.w3(32'h360c05f1),
	.w4(32'hb58bb56f),
	.w5(32'hb5b70dcc),
	.w6(32'h368a2149),
	.w7(32'h352c6b48),
	.w8(32'h357f6c31),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c40279),
	.w1(32'hb8f7d788),
	.w2(32'hb89b1901),
	.w3(32'hb9a3d1c8),
	.w4(32'hb91b48a8),
	.w5(32'hb9997fb4),
	.w6(32'hb96b5fe1),
	.w7(32'hb8710661),
	.w8(32'hb98eb714),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08f13a),
	.w1(32'hb941b6c9),
	.w2(32'hb9be71ab),
	.w3(32'hba9a2265),
	.w4(32'hba812085),
	.w5(32'hba477072),
	.w6(32'hba01d73f),
	.w7(32'hb8c5eb67),
	.w8(32'hb9ba790d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5d46c),
	.w1(32'hba31f93e),
	.w2(32'hb97c8034),
	.w3(32'hba9a361f),
	.w4(32'hb98cacde),
	.w5(32'h395ac803),
	.w6(32'hba81aceb),
	.w7(32'hba1fd31e),
	.w8(32'hba293273),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70afe6c),
	.w1(32'h38e9d26b),
	.w2(32'h3902bdb0),
	.w3(32'h3833050b),
	.w4(32'h38fb3048),
	.w5(32'h39012573),
	.w6(32'hb77bf2d0),
	.w7(32'h3922685e),
	.w8(32'h39442cdf),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe0354),
	.w1(32'hbb4c6501),
	.w2(32'hbc0e49eb),
	.w3(32'hbaaffd93),
	.w4(32'hba894a95),
	.w5(32'hbbe93288),
	.w6(32'hba2f6891),
	.w7(32'hb9b69ac0),
	.w8(32'hbc49fdb5),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44d5be),
	.w1(32'hbb36b4c5),
	.w2(32'hbb1789a7),
	.w3(32'h3a2c677e),
	.w4(32'hbbcbc52e),
	.w5(32'h3a869a3c),
	.w6(32'hbb9a60a2),
	.w7(32'hbbf59378),
	.w8(32'hbbb3dbb4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e1577),
	.w1(32'hb9af1a42),
	.w2(32'h3bc1941a),
	.w3(32'h3bf21c03),
	.w4(32'h3c01de41),
	.w5(32'h3b99362e),
	.w6(32'hbbe391c3),
	.w7(32'h3b2c8407),
	.w8(32'hbb678c0e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb295957),
	.w1(32'h3b36e7ce),
	.w2(32'h3b8c717c),
	.w3(32'hbc35162e),
	.w4(32'h3b21a188),
	.w5(32'hbb1a05ef),
	.w6(32'hbb9d279e),
	.w7(32'h3aea5f3b),
	.w8(32'hbc298fad),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4ec14),
	.w1(32'h3b5053db),
	.w2(32'h3b9ccda1),
	.w3(32'hbbfbaac2),
	.w4(32'h3b58e166),
	.w5(32'h3b13adb6),
	.w6(32'hbbc28a05),
	.w7(32'hba0bd807),
	.w8(32'hbad723af),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb70fe9),
	.w1(32'h3b9f0053),
	.w2(32'h3b0ee3d6),
	.w3(32'hba8e2eed),
	.w4(32'hba8cfb7b),
	.w5(32'hbba09193),
	.w6(32'hbb593c74),
	.w7(32'h3b8105af),
	.w8(32'hbaeaa216),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ecbdc),
	.w1(32'hbba4c4a4),
	.w2(32'hbad8c146),
	.w3(32'hbbfef294),
	.w4(32'hbbf4b4fe),
	.w5(32'hbb40f61c),
	.w6(32'hbb7a9310),
	.w7(32'hbb3b8afe),
	.w8(32'hbaa06e04),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03a1bb),
	.w1(32'h3b3905c4),
	.w2(32'h3bf232f2),
	.w3(32'hbbc85263),
	.w4(32'h3bd291e9),
	.w5(32'hbb7f0267),
	.w6(32'hbb089de8),
	.w7(32'h38c581e7),
	.w8(32'hba14a777),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7ebcc),
	.w1(32'hbc249726),
	.w2(32'hbb88c3a0),
	.w3(32'h3b2c6e0e),
	.w4(32'hbaef57b2),
	.w5(32'hbc513b2b),
	.w6(32'h3b1ec306),
	.w7(32'h39b7fcc5),
	.w8(32'h3b0fbf44),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af99150),
	.w1(32'hbb85ec3c),
	.w2(32'hbb821372),
	.w3(32'hbc00a4c2),
	.w4(32'h3a81418d),
	.w5(32'hbbb24080),
	.w6(32'h39412f52),
	.w7(32'hbaf71b1b),
	.w8(32'hbb24d8bc),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba3b6b),
	.w1(32'hbab37856),
	.w2(32'hbab24d3b),
	.w3(32'hbbb3c402),
	.w4(32'hbbbe3262),
	.w5(32'hbbe505e8),
	.w6(32'hbba1990a),
	.w7(32'h3b03adfc),
	.w8(32'h3a23cc61),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd17759),
	.w1(32'h3c1127f3),
	.w2(32'h3c1755ad),
	.w3(32'hbbd0841a),
	.w4(32'h3c70c25c),
	.w5(32'h3b736bb9),
	.w6(32'h390eeddb),
	.w7(32'h3b7fa9da),
	.w8(32'hb9f5c4bb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf768c7),
	.w1(32'hbb515c6b),
	.w2(32'hbc2d79fa),
	.w3(32'h3be18648),
	.w4(32'hbc0f08fc),
	.w5(32'hbc69d2c6),
	.w6(32'h3b996f75),
	.w7(32'h3b242aae),
	.w8(32'h3bf2c165),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae17f4b),
	.w1(32'hbb0fc9e4),
	.w2(32'h3ab656d2),
	.w3(32'h3c6be93e),
	.w4(32'hbb0484cd),
	.w5(32'hbad4e116),
	.w6(32'h3c254b49),
	.w7(32'hbbbe7995),
	.w8(32'h3a0be03e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9c25a),
	.w1(32'h3b09bbc1),
	.w2(32'hbb7122dc),
	.w3(32'h3b24b222),
	.w4(32'h3b4a459f),
	.w5(32'h3b0d0185),
	.w6(32'hbaa37fe8),
	.w7(32'hbb5d340e),
	.w8(32'hbbfea1a0),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3af094),
	.w1(32'hba82d97b),
	.w2(32'hbb978fac),
	.w3(32'h3b7cbd77),
	.w4(32'hba8bd285),
	.w5(32'hbbe3902b),
	.w6(32'hbb8c21bc),
	.w7(32'h3b9589c9),
	.w8(32'hba6c5a0f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee3122),
	.w1(32'hbb9ffb71),
	.w2(32'hbbc11592),
	.w3(32'hbb16a7a1),
	.w4(32'hbb56e430),
	.w5(32'h3ad2d4cd),
	.w6(32'hbbbde14d),
	.w7(32'hbbc40478),
	.w8(32'hbb202b7a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc140481),
	.w1(32'hbb23b58b),
	.w2(32'hb9c31ec6),
	.w3(32'hbc3d8b5d),
	.w4(32'h3ac03fa6),
	.w5(32'hbb967ddb),
	.w6(32'hbc21ae39),
	.w7(32'hbb894b50),
	.w8(32'hbc4c979e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0a1b1),
	.w1(32'hba0919cf),
	.w2(32'h3ac513ad),
	.w3(32'hbc356624),
	.w4(32'h3b852074),
	.w5(32'hbc31dfd8),
	.w6(32'hbbeac533),
	.w7(32'h3b297cb7),
	.w8(32'h3b6d6d81),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4fcbb),
	.w1(32'h3bdaafdc),
	.w2(32'h3b7695e1),
	.w3(32'hbbdc2973),
	.w4(32'h3a64b144),
	.w5(32'h39e26b13),
	.w6(32'h39e17fe2),
	.w7(32'hbba7b96e),
	.w8(32'h3a043970),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b3b95a),
	.w1(32'h3b065d09),
	.w2(32'h3b030ab5),
	.w3(32'h3c6718f7),
	.w4(32'hbb186026),
	.w5(32'h3bedfb47),
	.w6(32'hba97eb0f),
	.w7(32'hbb24f09e),
	.w8(32'h3b4fafbb),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99aa357),
	.w1(32'h3b63f0ba),
	.w2(32'h3b347ace),
	.w3(32'hb990dd86),
	.w4(32'h395dd39a),
	.w5(32'h39e6a4bc),
	.w6(32'h37669faa),
	.w7(32'h3b0658bd),
	.w8(32'hba31d104),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba935429),
	.w1(32'h3b77d0f2),
	.w2(32'hbb9a7fbd),
	.w3(32'hbb070b7c),
	.w4(32'h3b880cc0),
	.w5(32'h3c097ca7),
	.w6(32'hbb80e0f2),
	.w7(32'hbba78988),
	.w8(32'h3b0136ca),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92cfb79),
	.w1(32'h3b1fd5ad),
	.w2(32'h3a60bdbe),
	.w3(32'hbb496667),
	.w4(32'hba522bb8),
	.w5(32'hbad85dc0),
	.w6(32'hbbc30af8),
	.w7(32'h3b98cb03),
	.w8(32'h3a9737cd),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1c094),
	.w1(32'hba04cd54),
	.w2(32'h3b0658aa),
	.w3(32'hbae0325c),
	.w4(32'hbb4744ba),
	.w5(32'h39e224a2),
	.w6(32'hbbe622c3),
	.w7(32'hbb38a9fe),
	.w8(32'hbab53c40),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39014830),
	.w1(32'h3be5af77),
	.w2(32'h3af67093),
	.w3(32'hb9332ad8),
	.w4(32'h3add0c6e),
	.w5(32'hbb33a90a),
	.w6(32'hbb7278f0),
	.w7(32'h3abd7c34),
	.w8(32'hbbcd3e92),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c04cd),
	.w1(32'hbba332d2),
	.w2(32'h3b47bee7),
	.w3(32'hbb7b94cf),
	.w4(32'hbaadbcb2),
	.w5(32'h3cd0f826),
	.w6(32'hbbee0020),
	.w7(32'hbb870457),
	.w8(32'hbbbe1afa),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba89824),
	.w1(32'h3aa39805),
	.w2(32'hbc3e3cb9),
	.w3(32'hbbc85eee),
	.w4(32'hbbbbfb9c),
	.w5(32'hbb4573f3),
	.w6(32'hbc4463c8),
	.w7(32'hbba27ac2),
	.w8(32'h3abd5e84),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af23291),
	.w1(32'h3aa793ee),
	.w2(32'hbb4511ee),
	.w3(32'h3bd7ee0d),
	.w4(32'hba548091),
	.w5(32'hbba4200e),
	.w6(32'hbb17a1bc),
	.w7(32'hb95ad19e),
	.w8(32'hb9993a58),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b062c68),
	.w1(32'h3a9e65d3),
	.w2(32'h3c6b2cb2),
	.w3(32'hbae2881c),
	.w4(32'hbb19e32f),
	.w5(32'h3c9f1842),
	.w6(32'hb94f0a4f),
	.w7(32'h3c3bf840),
	.w8(32'h3c4ac1a4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf076c),
	.w1(32'h3b1aacef),
	.w2(32'h3af3d7fe),
	.w3(32'h3c2acd1d),
	.w4(32'h3b02cb45),
	.w5(32'hb8ee832e),
	.w6(32'h399d36e0),
	.w7(32'hbc040f37),
	.w8(32'hbb7c2427),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0cfb1),
	.w1(32'hb96f2747),
	.w2(32'hbab2c4fd),
	.w3(32'hbbbd74f7),
	.w4(32'hbb695b6c),
	.w5(32'hbbb1000a),
	.w6(32'h3b8f4416),
	.w7(32'hbb369761),
	.w8(32'h3b213881),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7f97a),
	.w1(32'h39c9eb08),
	.w2(32'hbb5eb36f),
	.w3(32'h3a92553a),
	.w4(32'h393c0e1a),
	.w5(32'h3b51e315),
	.w6(32'h3b025135),
	.w7(32'h3b7ad17b),
	.w8(32'hba57af2a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b2fe3),
	.w1(32'h3baa5d87),
	.w2(32'hbafd1cfa),
	.w3(32'h3b32fcbb),
	.w4(32'h3a6325aa),
	.w5(32'h3b8be6a1),
	.w6(32'hbb47ea49),
	.w7(32'h3af0cf45),
	.w8(32'hbb2ee24d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b1dcd),
	.w1(32'hbad00ef7),
	.w2(32'hbc2a0411),
	.w3(32'hbaa730aa),
	.w4(32'hb8c63840),
	.w5(32'hbc34e1ce),
	.w6(32'hbba23f9a),
	.w7(32'h3a4019ef),
	.w8(32'hbbbf5019),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6c807),
	.w1(32'h3a9d897b),
	.w2(32'h3ba42329),
	.w3(32'h3aabb038),
	.w4(32'hbbb861d4),
	.w5(32'hbbba072f),
	.w6(32'hbba7c73e),
	.w7(32'hbb531d0d),
	.w8(32'hbb0f4ced),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9a1b8),
	.w1(32'h3b343e90),
	.w2(32'hbb02ce78),
	.w3(32'h3bfbf9a4),
	.w4(32'hbb09665e),
	.w5(32'hbb0947b8),
	.w6(32'hbb25cf03),
	.w7(32'h3bccb4fc),
	.w8(32'h3baaac12),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc064c7),
	.w1(32'hbc09d08e),
	.w2(32'hbb7cf5e4),
	.w3(32'h3bc49840),
	.w4(32'hbc1d0fa8),
	.w5(32'hba52f051),
	.w6(32'h3b20eb1c),
	.w7(32'hbbbe7245),
	.w8(32'h3b757248),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee047b),
	.w1(32'hb988def6),
	.w2(32'h3c0e341f),
	.w3(32'h3c453bd1),
	.w4(32'h3b18d7fe),
	.w5(32'h3be054f7),
	.w6(32'h3bbc1f64),
	.w7(32'hb8902f81),
	.w8(32'h3b84a694),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6389fa),
	.w1(32'h3bae9dba),
	.w2(32'h3b272f7f),
	.w3(32'hbb88d492),
	.w4(32'h3ba4c68d),
	.w5(32'hbab6530f),
	.w6(32'h3b078673),
	.w7(32'h3b285a5d),
	.w8(32'hbab9e18a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39953121),
	.w1(32'hbb9d27d0),
	.w2(32'h3b9935c1),
	.w3(32'h3bc6e636),
	.w4(32'hbb7172d9),
	.w5(32'hbba2b9d5),
	.w6(32'h3b0772f4),
	.w7(32'hbad8c091),
	.w8(32'hbb80ec36),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb596254),
	.w1(32'hb8e7a143),
	.w2(32'hbc221bd1),
	.w3(32'hb9140464),
	.w4(32'hbbb83874),
	.w5(32'h3c65d7b5),
	.w6(32'h38d8adb1),
	.w7(32'hbb8eb985),
	.w8(32'hba60a800),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7811fc),
	.w1(32'hbb8f00cc),
	.w2(32'hb763b760),
	.w3(32'h3af128ce),
	.w4(32'hbc1908f8),
	.w5(32'h3c05915f),
	.w6(32'hbbb3729c),
	.w7(32'hbb58bb08),
	.w8(32'h3c576f28),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb69c0),
	.w1(32'h3b59208b),
	.w2(32'hbba86b55),
	.w3(32'hbbcef186),
	.w4(32'h39fc7b45),
	.w5(32'hbba2b327),
	.w6(32'hbbc13a2e),
	.w7(32'hba4ca0d6),
	.w8(32'h3b38ae69),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9fbc2),
	.w1(32'hb8a39fc0),
	.w2(32'h3ab2edff),
	.w3(32'h3a9fee81),
	.w4(32'hbb825fde),
	.w5(32'hbc3b1eea),
	.w6(32'h3a84ca59),
	.w7(32'hbc070381),
	.w8(32'hbc029a5c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e542d),
	.w1(32'h3a919eb3),
	.w2(32'h3b7ea719),
	.w3(32'h3ae8ae29),
	.w4(32'h3c2b5260),
	.w5(32'hbc2543da),
	.w6(32'hba110f7f),
	.w7(32'hba45742c),
	.w8(32'hbbaf49a1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3b6bd),
	.w1(32'h3b690dd3),
	.w2(32'h3a60bd3d),
	.w3(32'h3b3f254e),
	.w4(32'h3b788b6c),
	.w5(32'hbb479134),
	.w6(32'hb8e7adb6),
	.w7(32'h3a61ceed),
	.w8(32'hbabb5b13),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d7b49),
	.w1(32'hbb8557f3),
	.w2(32'hbc1161aa),
	.w3(32'hbbc426bc),
	.w4(32'hbbba0b76),
	.w5(32'hbc85384b),
	.w6(32'hbbeab778),
	.w7(32'h3b09f217),
	.w8(32'hbbb4421b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b601150),
	.w1(32'hbb1d1f3c),
	.w2(32'h3a9795d6),
	.w3(32'h3b395c23),
	.w4(32'h3b129ea2),
	.w5(32'hbb1746a2),
	.w6(32'hb9e21582),
	.w7(32'h3ba109b5),
	.w8(32'h3bbbf9b5),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb193aac),
	.w1(32'h3a43bf47),
	.w2(32'h3b44dfa1),
	.w3(32'h3b0a5888),
	.w4(32'h3b34c536),
	.w5(32'h3a1479a2),
	.w6(32'h3b223cf0),
	.w7(32'h39c80685),
	.w8(32'h3a8b20e9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7e883),
	.w1(32'hba2eacf5),
	.w2(32'hbbbddac0),
	.w3(32'hbbc5c3bc),
	.w4(32'h3949c527),
	.w5(32'hb9f4d3cd),
	.w6(32'hbbd57c40),
	.w7(32'hbb3aa79b),
	.w8(32'hbbbbd21c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29230c),
	.w1(32'h39cd3022),
	.w2(32'h3b37783a),
	.w3(32'hbbe60120),
	.w4(32'h3c22bba2),
	.w5(32'hbc0dcb23),
	.w6(32'hbb37f3c5),
	.w7(32'hbbcfb6b5),
	.w8(32'hbc0757e0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0608ec),
	.w1(32'hbb5a450d),
	.w2(32'h3b1973ef),
	.w3(32'h39622ec0),
	.w4(32'hbbaa75e7),
	.w5(32'h3af90fa7),
	.w6(32'hb9ae43a6),
	.w7(32'hbb89ccaa),
	.w8(32'hbc09d1a9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae07fc1),
	.w1(32'h3b0befcc),
	.w2(32'hbb9e0004),
	.w3(32'h3aec78a3),
	.w4(32'hbb8d07c2),
	.w5(32'hbba4393a),
	.w6(32'h3bb8e0ad),
	.w7(32'hbb996ccd),
	.w8(32'h3b941818),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef090d),
	.w1(32'hb90f1e19),
	.w2(32'hbb9bc575),
	.w3(32'h39ab6dcb),
	.w4(32'hbb3b8d59),
	.w5(32'h3a620845),
	.w6(32'hbbf78ee1),
	.w7(32'h3b9231aa),
	.w8(32'h3bfac2c3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd420a),
	.w1(32'hb983fbf0),
	.w2(32'h3929ac6e),
	.w3(32'h3b791781),
	.w4(32'hbae269b5),
	.w5(32'hbbfdf163),
	.w6(32'hbba20dba),
	.w7(32'h3b520cba),
	.w8(32'hbaf53dee),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2fd42),
	.w1(32'h39248aeb),
	.w2(32'hbac94ede),
	.w3(32'hbc3a5dd2),
	.w4(32'h3ba7cc0b),
	.w5(32'hbbcae062),
	.w6(32'hbb99e4bd),
	.w7(32'hbaddf97b),
	.w8(32'hbb9f52a2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd34d8c),
	.w1(32'hbc1f26df),
	.w2(32'hbc08e8e8),
	.w3(32'hbb41caa0),
	.w4(32'hbc6c1f71),
	.w5(32'hbb552af4),
	.w6(32'h3b8af873),
	.w7(32'h3ae8f718),
	.w8(32'h3b211112),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb061fb),
	.w1(32'h3b8c70ad),
	.w2(32'hba5ddb70),
	.w3(32'h3b0219c8),
	.w4(32'hbb975835),
	.w5(32'hba574775),
	.w6(32'h3b9a4a76),
	.w7(32'hbc018686),
	.w8(32'hbbc46c3d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule