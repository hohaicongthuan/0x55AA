module layer_6_featuremap_2(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3722ae16),
	.w1(32'hb77141a3),
	.w2(32'hb855732f),
	.w3(32'hb86c1e41),
	.w4(32'hb7f9256c),
	.w5(32'hb916e19c),
	.w6(32'hb91ec635),
	.w7(32'hb90f2a3c),
	.w8(32'hb95b23ed),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f3fddb),
	.w1(32'h36134139),
	.w2(32'h37796b6d),
	.w3(32'hb917cf96),
	.w4(32'hb5d09840),
	.w5(32'h388d93ec),
	.w6(32'hb99b62ba),
	.w7(32'hb91a1c5e),
	.w8(32'hb85a5a67),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89911d),
	.w1(32'hb9e0c3e7),
	.w2(32'h38d9ab57),
	.w3(32'hbaac75fe),
	.w4(32'hb9eb83db),
	.w5(32'hb96e5b69),
	.w6(32'hbaa5bd0d),
	.w7(32'hba108dc6),
	.w8(32'hba39e3bc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d59e78),
	.w1(32'hbb241b67),
	.w2(32'hbad80313),
	.w3(32'hb8df2dfa),
	.w4(32'hba81ae2a),
	.w5(32'h3bb89f60),
	.w6(32'hbb392e2d),
	.w7(32'h39ae3dc2),
	.w8(32'h3c028f48),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d981e8),
	.w1(32'hb98a2fb8),
	.w2(32'hbb1c00a0),
	.w3(32'h3aa895bf),
	.w4(32'h3ab5bf41),
	.w5(32'hb99f1ac2),
	.w6(32'hba1fe94b),
	.w7(32'hbb022bb8),
	.w8(32'hbb229aff),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a37c8),
	.w1(32'hb9447976),
	.w2(32'hb911488b),
	.w3(32'hb8efc2e1),
	.w4(32'hb9672e37),
	.w5(32'hb9360083),
	.w6(32'hb9561870),
	.w7(32'hb9b11d2d),
	.w8(32'hb9a1a349),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5928c8),
	.w1(32'hbb416a38),
	.w2(32'hbaed573d),
	.w3(32'hbb5de5d3),
	.w4(32'hbb5bd3ac),
	.w5(32'hbb5be213),
	.w6(32'hbaa40c8f),
	.w7(32'hbabdcbd8),
	.w8(32'hbaea1564),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d6d2b),
	.w1(32'hba42c813),
	.w2(32'hba86cd17),
	.w3(32'hba83dc13),
	.w4(32'hbab1a6a7),
	.w5(32'hbb13384f),
	.w6(32'hba1a5bf9),
	.w7(32'hbaa11d6f),
	.w8(32'hbb123321),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13f49f),
	.w1(32'hbafff9fb),
	.w2(32'hbaef3b09),
	.w3(32'hbb03a9fd),
	.w4(32'hbabc62c1),
	.w5(32'hb8e58f3e),
	.w6(32'hbb165158),
	.w7(32'hbadc93d2),
	.w8(32'h3891a7d3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58ce1f),
	.w1(32'h3a0cc088),
	.w2(32'h3a832117),
	.w3(32'h398ef011),
	.w4(32'h373a58ff),
	.w5(32'h394de8cd),
	.w6(32'h3a39d4d4),
	.w7(32'h399e603d),
	.w8(32'h3a130a7c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3f369),
	.w1(32'h3b1b60fb),
	.w2(32'hbb2a241e),
	.w3(32'h3b64b21d),
	.w4(32'h3b6f0ce9),
	.w5(32'h3b138dee),
	.w6(32'hbb135a87),
	.w7(32'hbaf9af5a),
	.w8(32'hbab41225),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09cf89),
	.w1(32'hba01c6cd),
	.w2(32'hb9d2d3b7),
	.w3(32'hb9b51d56),
	.w4(32'hb9e0e4b3),
	.w5(32'h3878adc7),
	.w6(32'hba2aeb6e),
	.w7(32'hb9e2eba2),
	.w8(32'hb86df4f2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f69bcf),
	.w1(32'hb6a980df),
	.w2(32'hb6a225fb),
	.w3(32'hb8561923),
	.w4(32'hb7f89879),
	.w5(32'hb852f3b6),
	.w6(32'hb87cc3e4),
	.w7(32'hb82984a9),
	.w8(32'hb864560c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc39b3e),
	.w1(32'h3ba22c20),
	.w2(32'h3a00a2eb),
	.w3(32'h3c09f764),
	.w4(32'h3bf4a065),
	.w5(32'h3b862f30),
	.w6(32'h3b0e8562),
	.w7(32'hbae69962),
	.w8(32'hbb4abfa6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab11fd0),
	.w1(32'hbb0faf04),
	.w2(32'hbb2b4d3d),
	.w3(32'hbac81597),
	.w4(32'hbb1c5f39),
	.w5(32'hba9bf316),
	.w6(32'hbb1f04fa),
	.w7(32'hbae3c262),
	.w8(32'hbaa3a3ed),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6106ea),
	.w1(32'hba3e4165),
	.w2(32'hbaf6663d),
	.w3(32'h3a30bbdb),
	.w4(32'hb91e260b),
	.w5(32'h3a1d09fc),
	.w6(32'hbb38877a),
	.w7(32'hbb6a065e),
	.w8(32'hba9c4e97),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb3304),
	.w1(32'h3c1e9054),
	.w2(32'h3c79c3bf),
	.w3(32'hbc521c2c),
	.w4(32'hbb31778a),
	.w5(32'h3c1bf5ed),
	.w6(32'hbba3d514),
	.w7(32'h3a00a5df),
	.w8(32'h3babe4ed),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f0ab87),
	.w1(32'h362eb541),
	.w2(32'h376d93a7),
	.w3(32'hb7977412),
	.w4(32'h378ba8c3),
	.w5(32'h37b3a7e9),
	.w6(32'hb811d4e1),
	.w7(32'hb76bdf27),
	.w8(32'hb68f1e4b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1ef4c),
	.w1(32'hbae9fd88),
	.w2(32'hbaefc928),
	.w3(32'hbb24b474),
	.w4(32'hbb16e2be),
	.w5(32'hbb885505),
	.w6(32'hba42a5a6),
	.w7(32'hbaabe100),
	.w8(32'hbade970e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399cf0c8),
	.w1(32'h3a047374),
	.w2(32'h3a9cd10e),
	.w3(32'h3b1b1398),
	.w4(32'h3b096bbf),
	.w5(32'h3b2fbb24),
	.w6(32'h3aa1b41d),
	.w7(32'h3a1cfe27),
	.w8(32'hb97b06aa),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba230fae),
	.w1(32'hbb3e4bb6),
	.w2(32'hb9e39b13),
	.w3(32'h3ab4fa3d),
	.w4(32'hb8d18daf),
	.w5(32'h3ba46d5f),
	.w6(32'h39b8e8b9),
	.w7(32'hb955d5d2),
	.w8(32'h3b0fb309),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbe6f2),
	.w1(32'h3b8e95f2),
	.w2(32'h3b1c1f53),
	.w3(32'h3c1d05d3),
	.w4(32'h3c175e65),
	.w5(32'h3c077c72),
	.w6(32'h3b9debe1),
	.w7(32'h3b154931),
	.w8(32'h3aa72577),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398da756),
	.w1(32'h37d60cc5),
	.w2(32'h39cd770e),
	.w3(32'h39971d3e),
	.w4(32'hb8821abb),
	.w5(32'hba07efd1),
	.w6(32'h3ae0f57a),
	.w7(32'h3ae5c96e),
	.w8(32'h3a7e615d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3a803),
	.w1(32'hba8eafd3),
	.w2(32'h3aa76b37),
	.w3(32'h3b471247),
	.w4(32'hb8b78e84),
	.w5(32'h39231c03),
	.w6(32'hba9336ea),
	.w7(32'hbbacfa54),
	.w8(32'hbaf88188),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42ec4b),
	.w1(32'hbc704211),
	.w2(32'hbc33d6f7),
	.w3(32'hbc0c1c0d),
	.w4(32'hbb508e47),
	.w5(32'h3c813bf1),
	.w6(32'hbc5dc588),
	.w7(32'hbc076b92),
	.w8(32'hba9c1f61),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45245a),
	.w1(32'hbab6f4a9),
	.w2(32'h3af5c6a4),
	.w3(32'hbb918a37),
	.w4(32'hba9bf4b7),
	.w5(32'h3c1956ad),
	.w6(32'hbbbcd736),
	.w7(32'h3a9a32de),
	.w8(32'h3c428e63),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95c728),
	.w1(32'h3ba2e00a),
	.w2(32'h3b8530bb),
	.w3(32'h3b4a5f58),
	.w4(32'h3a143965),
	.w5(32'h3a232626),
	.w6(32'h3a4d7ff5),
	.w7(32'hbb219a45),
	.w8(32'hba20e456),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9804f83),
	.w1(32'hb8a80377),
	.w2(32'h394cc137),
	.w3(32'hb96707dc),
	.w4(32'hb8fff170),
	.w5(32'h393bb6e1),
	.w6(32'hb946cd69),
	.w7(32'hb8bab8a0),
	.w8(32'h387f2647),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa646b5),
	.w1(32'h3a73f532),
	.w2(32'h39d24f20),
	.w3(32'h3ad6c544),
	.w4(32'h3aac7895),
	.w5(32'h3a9763c9),
	.w6(32'h3a2ee076),
	.w7(32'h38df1d7e),
	.w8(32'h35afa174),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89b16f),
	.w1(32'hbab1bf03),
	.w2(32'hbbf6748b),
	.w3(32'hbbb6e2e0),
	.w4(32'hbc2fdedf),
	.w5(32'hbbbbff82),
	.w6(32'hbc5508bf),
	.w7(32'hbc2a35ce),
	.w8(32'hbb03c576),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6eff1e4),
	.w1(32'hbcac5050),
	.w2(32'hbcfe707d),
	.w3(32'hb6bc9147),
	.w4(32'h3ad8c189),
	.w5(32'hbcebe7fa),
	.w6(32'hbc3540d4),
	.w7(32'h3ad11ee6),
	.w8(32'h3bf25d2d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29dd8d),
	.w1(32'hbbd63bc4),
	.w2(32'hbbf07570),
	.w3(32'hbbdaf33a),
	.w4(32'hbb1c6229),
	.w5(32'h3c3fdf1b),
	.w6(32'hbc3e758d),
	.w7(32'hbcadb4fc),
	.w8(32'hbc2ead66),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05b2b9),
	.w1(32'h3c500fda),
	.w2(32'h3c849041),
	.w3(32'hbacd8d63),
	.w4(32'hbd4177b0),
	.w5(32'hbdea42f6),
	.w6(32'h3d058e7f),
	.w7(32'h3dae3aae),
	.w8(32'h3d47d84d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2233b0),
	.w1(32'h3d334dde),
	.w2(32'h3d1a5d39),
	.w3(32'hbd72af29),
	.w4(32'hbbb26e15),
	.w5(32'h3c3b9d19),
	.w6(32'h3c5c3d06),
	.w7(32'h3d0d4a7c),
	.w8(32'h3cc1ccb0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d76fd77),
	.w1(32'h3c7ec11e),
	.w2(32'hbbdee4f1),
	.w3(32'h3bb5303d),
	.w4(32'hbb9706c0),
	.w5(32'hbc66ef23),
	.w6(32'h3b408374),
	.w7(32'h3c0c232f),
	.w8(32'h3c0dbf82),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf794f1),
	.w1(32'hbcb5c9ba),
	.w2(32'hbd8042f0),
	.w3(32'h3c45d2f9),
	.w4(32'h3cbf89a9),
	.w5(32'h3d0a4f97),
	.w6(32'h3c4c4556),
	.w7(32'h3c9d58e5),
	.w8(32'hbbfb95c0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda9b7e),
	.w1(32'h3ac4d8f6),
	.w2(32'hbd0a4474),
	.w3(32'hbb52ce45),
	.w4(32'h3c50335e),
	.w5(32'h3aa518d9),
	.w6(32'h3c982b86),
	.w7(32'hba297850),
	.w8(32'h391712e5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d622a),
	.w1(32'hbd53c27c),
	.w2(32'hbcbd9084),
	.w3(32'h3bb5a221),
	.w4(32'hbbf05ff5),
	.w5(32'h3aa690ec),
	.w6(32'hbd4bb9be),
	.w7(32'hbd3d51e0),
	.w8(32'hbcd74673),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01c52e),
	.w1(32'h3b329fa6),
	.w2(32'h3c1084d2),
	.w3(32'hbba64bbf),
	.w4(32'h3c335cb5),
	.w5(32'h3c6a254a),
	.w6(32'h3c1cf576),
	.w7(32'h3c4fc90b),
	.w8(32'h3c35d52a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e63f2),
	.w1(32'h3b858918),
	.w2(32'hbbedd78d),
	.w3(32'h3d0c4cd8),
	.w4(32'h3d0621e5),
	.w5(32'h3d58f116),
	.w6(32'hbb9c7c81),
	.w7(32'hbc17ee52),
	.w8(32'hbca35166),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01909d),
	.w1(32'h3b873188),
	.w2(32'hbb9f902d),
	.w3(32'h3b591451),
	.w4(32'h3aac117f),
	.w5(32'h3c5ef861),
	.w6(32'hba22fc6c),
	.w7(32'hba5ce9db),
	.w8(32'hbbefe4bb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5b251),
	.w1(32'h3c1da389),
	.w2(32'h3c12472b),
	.w3(32'h3b89ffd8),
	.w4(32'h3c67c9e3),
	.w5(32'h3c6efff7),
	.w6(32'h3c2b6a58),
	.w7(32'h3c0d7e47),
	.w8(32'h3c23d46c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbae90c),
	.w1(32'hbcd16e36),
	.w2(32'hbd67dc94),
	.w3(32'h3c58dfdf),
	.w4(32'hbc3fca0f),
	.w5(32'h3ba39a70),
	.w6(32'hbb6b5e59),
	.w7(32'hbab869e3),
	.w8(32'hbc1926f0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5fceb),
	.w1(32'hbbe9a0d7),
	.w2(32'hbbeb4c27),
	.w3(32'hbb3adceb),
	.w4(32'h3a9e94ea),
	.w5(32'h38314951),
	.w6(32'hbbfb2226),
	.w7(32'h3a31361a),
	.w8(32'h3c0e1a14),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebe1b7),
	.w1(32'h3bba6c07),
	.w2(32'h3ce34cfa),
	.w3(32'h3bc93b9f),
	.w4(32'h3c1959d6),
	.w5(32'hbce2deac),
	.w6(32'h3b6ac9e6),
	.w7(32'hbbe15706),
	.w8(32'hbc046aa3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a137603),
	.w1(32'h3c89d073),
	.w2(32'h3cf13437),
	.w3(32'hbb99f516),
	.w4(32'h3b9b1860),
	.w5(32'h3b66b717),
	.w6(32'hbc381e97),
	.w7(32'h38a9e3da),
	.w8(32'h39c7cb6b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5725b9),
	.w1(32'hbc9e1347),
	.w2(32'hbd1cc6d8),
	.w3(32'hbb7572f6),
	.w4(32'hbd2711aa),
	.w5(32'h3cfd8f18),
	.w6(32'hbc743050),
	.w7(32'hbd85f69e),
	.w8(32'h3b75fe46),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc717f40),
	.w1(32'hbcb1a075),
	.w2(32'hbcf30829),
	.w3(32'h3bdab6c9),
	.w4(32'hbcd685df),
	.w5(32'hbc553355),
	.w6(32'hbc87d163),
	.w7(32'hbca3f6a9),
	.w8(32'h3c076dd6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca035b),
	.w1(32'h3d54bf63),
	.w2(32'hbd136756),
	.w3(32'h3cffa0e2),
	.w4(32'h3c8ed01c),
	.w5(32'h3caf0427),
	.w6(32'h3c65bf38),
	.w7(32'hbc2b82db),
	.w8(32'hbcfc25a5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca66513),
	.w1(32'hbcc69495),
	.w2(32'hbcbba720),
	.w3(32'hbcf9caa3),
	.w4(32'hbcbebd6b),
	.w5(32'hbcbe0a9f),
	.w6(32'h3b3346ae),
	.w7(32'h3c3d0715),
	.w8(32'h3c428121),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0d761),
	.w1(32'hbc4fd1df),
	.w2(32'hbca99558),
	.w3(32'hbc823b15),
	.w4(32'h3b3613a9),
	.w5(32'h3c53ec13),
	.w6(32'hbb164b85),
	.w7(32'hbc0774ca),
	.w8(32'hbb97789b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bdc86),
	.w1(32'h3ccac5e2),
	.w2(32'h3d98bc9d),
	.w3(32'h3c03a665),
	.w4(32'hbccab151),
	.w5(32'hbb08f8bb),
	.w6(32'hbbb13ec3),
	.w7(32'h3c8fd942),
	.w8(32'hba4f11c0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe9405),
	.w1(32'h3bc4d447),
	.w2(32'hbcd2fd4a),
	.w3(32'hbc0e808b),
	.w4(32'hba26ff2c),
	.w5(32'h3c00a803),
	.w6(32'h3cbcab37),
	.w7(32'hbc23caf6),
	.w8(32'hbc2888fb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6e4d2),
	.w1(32'hbcaf80cb),
	.w2(32'hbd40b73f),
	.w3(32'hbc1a584f),
	.w4(32'hbc1426d9),
	.w5(32'h3aa09002),
	.w6(32'hbc2861ce),
	.w7(32'hbc6efe10),
	.w8(32'hbcd1bd39),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc018e89),
	.w1(32'hbb050d11),
	.w2(32'h3bc192a7),
	.w3(32'hbac1ed5d),
	.w4(32'hbd270b65),
	.w5(32'hbd36625e),
	.w6(32'hbc5a4f19),
	.w7(32'hbc92f3c9),
	.w8(32'h3b81e8fb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07563b),
	.w1(32'hbc9508f4),
	.w2(32'hbd05bcf0),
	.w3(32'hbb179174),
	.w4(32'h3ca13aef),
	.w5(32'hbcb57f78),
	.w6(32'h3ad12f3b),
	.w7(32'hbcfdb84b),
	.w8(32'hbb29f34b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1b17e),
	.w1(32'hbc20b1f5),
	.w2(32'hbd57aed2),
	.w3(32'h3bb0a7fc),
	.w4(32'h3ca2e22e),
	.w5(32'h3c4e1746),
	.w6(32'hbb7507e1),
	.w7(32'h3c7bfb68),
	.w8(32'hbb4ed834),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4cbc9),
	.w1(32'h39cf0edb),
	.w2(32'hbb08bec3),
	.w3(32'hbcbf520a),
	.w4(32'hbb65e662),
	.w5(32'hbba990d0),
	.w6(32'h3c5e5147),
	.w7(32'hbbb083ef),
	.w8(32'hbb341f4f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf7276),
	.w1(32'h3c3307aa),
	.w2(32'h3cc5068d),
	.w3(32'hbb3c9063),
	.w4(32'hbcc55252),
	.w5(32'h3cdea1f1),
	.w6(32'hbce2586a),
	.w7(32'h3c2da9ce),
	.w8(32'hbd08d7f1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a2cb9),
	.w1(32'hbaea1b36),
	.w2(32'hbc072a43),
	.w3(32'hbb5caf96),
	.w4(32'hbc0f6b4e),
	.w5(32'hbbdbb30c),
	.w6(32'hbd4d2709),
	.w7(32'hbd52c93c),
	.w8(32'hbc919986),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8d726),
	.w1(32'hbbb9ddbb),
	.w2(32'hbc940a58),
	.w3(32'h3b15b0ff),
	.w4(32'hbba07491),
	.w5(32'h3b1884ec),
	.w6(32'hbc671188),
	.w7(32'hbc62211d),
	.w8(32'hbc990e25),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59cb72),
	.w1(32'h3c4882cd),
	.w2(32'hbb55ab1b),
	.w3(32'hbb1f2d6f),
	.w4(32'h3cb8d729),
	.w5(32'h3c678f3a),
	.w6(32'hbc4cfd4d),
	.w7(32'hbbf3a9b6),
	.w8(32'hbc40612f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4273f),
	.w1(32'hbc6b6f23),
	.w2(32'hbca39844),
	.w3(32'hbc7eaec4),
	.w4(32'hbc86c451),
	.w5(32'hbc80652a),
	.w6(32'hbce5987c),
	.w7(32'hbccc0e4d),
	.w8(32'hbca5be12),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ce0e3),
	.w1(32'h3b2202fb),
	.w2(32'h3b49d940),
	.w3(32'h3b3321ae),
	.w4(32'h3b0f7f09),
	.w5(32'h3b948c2e),
	.w6(32'h3a67a9c4),
	.w7(32'h39ba34b1),
	.w8(32'h3b375942),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule