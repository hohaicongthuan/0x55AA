module layer_10_featuremap_73(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52d8b5),
	.w1(32'hbb82f050),
	.w2(32'h3b46d632),
	.w3(32'h3c152112),
	.w4(32'hba051532),
	.w5(32'hbc2e63a7),
	.w6(32'h3c16ac77),
	.w7(32'h3ab3c5db),
	.w8(32'hbca2edd4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f801a),
	.w1(32'h3cd3a6f9),
	.w2(32'h3ba33857),
	.w3(32'h3b95fb74),
	.w4(32'h3cde5b4b),
	.w5(32'h3ca08a9f),
	.w6(32'hbb535276),
	.w7(32'h3c39ef77),
	.w8(32'h3bcbc238),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2ea10),
	.w1(32'h3cc76447),
	.w2(32'hbbcadf86),
	.w3(32'h3d235ee3),
	.w4(32'h3d034251),
	.w5(32'hbb20442e),
	.w6(32'h3c5ad5f4),
	.w7(32'h3c157b61),
	.w8(32'h3a8bb74e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb02fed),
	.w1(32'h3c0cbd98),
	.w2(32'h3a58d131),
	.w3(32'h3934ad3f),
	.w4(32'h3a855b70),
	.w5(32'hbba75259),
	.w6(32'h3c05a25f),
	.w7(32'hbb950a22),
	.w8(32'h3c249864),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956b821),
	.w1(32'h3bca87ae),
	.w2(32'h3cbade98),
	.w3(32'h3c5f2fc3),
	.w4(32'h3bec54fc),
	.w5(32'h3d136bb7),
	.w6(32'h3c432b4f),
	.w7(32'h3b5b7ca0),
	.w8(32'h3cd0a682),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdef194),
	.w1(32'h3bb85d52),
	.w2(32'hbca6d7a1),
	.w3(32'h3cfff22c),
	.w4(32'h3c89030c),
	.w5(32'hbcaeaf3f),
	.w6(32'h3c8d7103),
	.w7(32'h3b4902b2),
	.w8(32'hbcb56780),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d13dcc9),
	.w1(32'hbc675b75),
	.w2(32'h3bdfdf1f),
	.w3(32'h3d0ef16a),
	.w4(32'hbc7ee6e0),
	.w5(32'h3abcdc75),
	.w6(32'h3cfdb908),
	.w7(32'hbca5f641),
	.w8(32'h3bbcd9df),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68b292),
	.w1(32'hbbcacd84),
	.w2(32'h3ba6a325),
	.w3(32'h3bade269),
	.w4(32'hbbeb70f1),
	.w5(32'h3bd96e64),
	.w6(32'h3c54a263),
	.w7(32'h3b25a4d5),
	.w8(32'h3bdcdb5f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc51324),
	.w1(32'hbb4fd339),
	.w2(32'hbbd7dbe1),
	.w3(32'h3b3a6395),
	.w4(32'hbba5c44a),
	.w5(32'h3c1bcfef),
	.w6(32'h3a897a66),
	.w7(32'hbc0f0c1d),
	.w8(32'h3c11e861),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82937e),
	.w1(32'h3c8724e1),
	.w2(32'hbc84db33),
	.w3(32'h3d110fd8),
	.w4(32'h3cf82bdd),
	.w5(32'hbc9817f4),
	.w6(32'h3d10cbd3),
	.w7(32'h3cfefcb0),
	.w8(32'hbc7faab3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c5079),
	.w1(32'hbc816617),
	.w2(32'hb9c2ab14),
	.w3(32'hbc541685),
	.w4(32'hbc96c1ca),
	.w5(32'h3c136800),
	.w6(32'hbc476348),
	.w7(32'hbc78ad9b),
	.w8(32'h3c0d40bc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ce609),
	.w1(32'h3afc5447),
	.w2(32'hbbeafbf0),
	.w3(32'h3c43e4fd),
	.w4(32'h3c166220),
	.w5(32'hbc36ac74),
	.w6(32'h3c528490),
	.w7(32'h3bc680a6),
	.w8(32'hbc1df76a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56c6b4),
	.w1(32'hbaaef796),
	.w2(32'hbdedf624),
	.w3(32'hb95244f4),
	.w4(32'hbb3944ae),
	.w5(32'hbe2724ce),
	.w6(32'hb7101d52),
	.w7(32'h39edc9b9),
	.w8(32'hbe002a1e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe28704d),
	.w1(32'hbdab9f58),
	.w2(32'h3c338922),
	.w3(32'hbe64a960),
	.w4(32'hbe0f08c8),
	.w5(32'h3c2bf889),
	.w6(32'hbe2f8c09),
	.w7(32'hbdc0b810),
	.w8(32'h3b9370b1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c087b08),
	.w1(32'h3c94475a),
	.w2(32'hbbe90d3c),
	.w3(32'h3c988099),
	.w4(32'h3c9add81),
	.w5(32'hbbb5dbd8),
	.w6(32'h3c24eea9),
	.w7(32'h3c37b927),
	.w8(32'hbc36e4ca),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bf5a1),
	.w1(32'hbadb2c6f),
	.w2(32'hbc21b8b5),
	.w3(32'hba4d1f87),
	.w4(32'hbb8c2478),
	.w5(32'hbc09cfd9),
	.w6(32'hbbf2538d),
	.w7(32'hbc05829f),
	.w8(32'hbbf84888),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fc876),
	.w1(32'hbbf2692a),
	.w2(32'h3a2d0ced),
	.w3(32'h3acd6b10),
	.w4(32'hbc0fa563),
	.w5(32'h3b458466),
	.w6(32'h3a58339c),
	.w7(32'hbbdf5dc6),
	.w8(32'hb921c052),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66a9fd),
	.w1(32'h3c1355fb),
	.w2(32'hbda09596),
	.w3(32'h3c94c93f),
	.w4(32'h3c0c5193),
	.w5(32'hbdd21db3),
	.w6(32'h3c8e7e24),
	.w7(32'h3c32b358),
	.w8(32'hbdaccef8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdcf6db6),
	.w1(32'hbd88421c),
	.w2(32'h3b230606),
	.w3(32'hbe004634),
	.w4(32'hbdb36b0b),
	.w5(32'hbbd14e74),
	.w6(32'hbddb7b0e),
	.w7(32'hbd7a5b25),
	.w8(32'hbad0afc3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb962e99),
	.w1(32'hbabe1b0c),
	.w2(32'h3c413c85),
	.w3(32'hbb9073a9),
	.w4(32'hbb9b0989),
	.w5(32'h3b9e5e5a),
	.w6(32'hbb1c8374),
	.w7(32'hbb98a97f),
	.w8(32'h3ae818b9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b050695),
	.w1(32'hbbaaabc9),
	.w2(32'h3beaa99c),
	.w3(32'h3b34c9e4),
	.w4(32'hba5c050b),
	.w5(32'h3ca1436b),
	.w6(32'hbbb4837b),
	.w7(32'hbb5972cb),
	.w8(32'h3c048997),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87295e),
	.w1(32'h3c2c6eeb),
	.w2(32'hbcd9cff3),
	.w3(32'h3c55ff51),
	.w4(32'h3c720a05),
	.w5(32'hbce39b7b),
	.w6(32'h3c1d98f9),
	.w7(32'h3bdb20a6),
	.w8(32'hbc8baa69),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cc475),
	.w1(32'hbb937754),
	.w2(32'hbaed07ba),
	.w3(32'hbc22d292),
	.w4(32'hbb897ced),
	.w5(32'hbb1bb630),
	.w6(32'h38a2d796),
	.w7(32'h3ba642b7),
	.w8(32'h3ae65173),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0f8fa),
	.w1(32'h3b57d332),
	.w2(32'hbdacc2d7),
	.w3(32'h3b128c0d),
	.w4(32'h39804f56),
	.w5(32'hbdf986e5),
	.w6(32'h3bfcaaa4),
	.w7(32'h3bcda162),
	.w8(32'hbdc2a49b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdfe0fd1),
	.w1(32'hbd9981ee),
	.w2(32'h3c163907),
	.w3(32'hbe3505f6),
	.w4(32'hbdd3cbca),
	.w5(32'h3b9f031f),
	.w6(32'hbe06c676),
	.w7(32'hbd71d556),
	.w8(32'hbc32fb0d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e8240),
	.w1(32'h3c073632),
	.w2(32'h3c4cf897),
	.w3(32'h3c145206),
	.w4(32'h3b9bf842),
	.w5(32'hbb32f873),
	.w6(32'hbbaf964a),
	.w7(32'h39b81ac5),
	.w8(32'hbbd77057),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25b8ce),
	.w1(32'h398a7696),
	.w2(32'h39d24aa7),
	.w3(32'hbc4130fc),
	.w4(32'hbb07c773),
	.w5(32'h3a69db7c),
	.w6(32'hb80fbc7e),
	.w7(32'h3bb23ebc),
	.w8(32'h3a122483),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ace32c),
	.w1(32'hba08cb6c),
	.w2(32'hbc0aee6f),
	.w3(32'h3a95aced),
	.w4(32'hba2739fd),
	.w5(32'hbbac1ab6),
	.w6(32'h3a1a7243),
	.w7(32'hba11df65),
	.w8(32'hbbcb53db),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75d01c),
	.w1(32'hbb317552),
	.w2(32'h3b1109f0),
	.w3(32'hba688518),
	.w4(32'hba400a28),
	.w5(32'h3bbdfed6),
	.w6(32'hbbbc6d58),
	.w7(32'hba92c44b),
	.w8(32'h3a8d0db5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85f06c),
	.w1(32'hb98a9f19),
	.w2(32'h3a1ea98b),
	.w3(32'hbaeba73a),
	.w4(32'h3b1658b7),
	.w5(32'hbac1bbed),
	.w6(32'hbada257e),
	.w7(32'h3b8a88bb),
	.w8(32'hb9deec70),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e7908),
	.w1(32'hb99ba78d),
	.w2(32'h3b74da1b),
	.w3(32'hba9a18be),
	.w4(32'hbadc0a9c),
	.w5(32'hbb7179b7),
	.w6(32'h39268715),
	.w7(32'hba263c47),
	.w8(32'h3bae5cb9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b25be),
	.w1(32'h3a3e342d),
	.w2(32'h3b6e6d0e),
	.w3(32'hbbbc58af),
	.w4(32'hbbb06c6c),
	.w5(32'h3b438a02),
	.w6(32'h3bac7a18),
	.w7(32'h3bedad70),
	.w8(32'hb99c904b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cd259),
	.w1(32'h3b244e36),
	.w2(32'h3a10aa2f),
	.w3(32'h3b265ea0),
	.w4(32'hb9b781f6),
	.w5(32'hbb282465),
	.w6(32'h3b521d90),
	.w7(32'h3b2aa533),
	.w8(32'hbb1f1320),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab59ee8),
	.w1(32'hba603d65),
	.w2(32'h3a06d876),
	.w3(32'hbb5f971d),
	.w4(32'hbb4e710c),
	.w5(32'h3b874004),
	.w6(32'hbb540bc7),
	.w7(32'hbb0e9a07),
	.w8(32'h3b29f7bc),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34bcce),
	.w1(32'hbb33e2aa),
	.w2(32'hbb50feea),
	.w3(32'h39dc4ad1),
	.w4(32'hbb684c7d),
	.w5(32'hbb359c6f),
	.w6(32'h3bd7a77c),
	.w7(32'hbba1a0f7),
	.w8(32'hbb7a1e87),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85297c),
	.w1(32'h3b0539c9),
	.w2(32'hbb40a13d),
	.w3(32'hba71d4c0),
	.w4(32'h3af9c486),
	.w5(32'hbb38c05c),
	.w6(32'hbab67169),
	.w7(32'h3b006611),
	.w8(32'hbb92362f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fe695),
	.w1(32'h3a6f1c62),
	.w2(32'hbbc782db),
	.w3(32'hbb038b9a),
	.w4(32'h3aabe145),
	.w5(32'hbc043615),
	.w6(32'h39a52047),
	.w7(32'h3bce0a0e),
	.w8(32'hbc0f153d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9e89a),
	.w1(32'h397ac631),
	.w2(32'hba53795a),
	.w3(32'h38a24968),
	.w4(32'h39dce49e),
	.w5(32'h3b458aa1),
	.w6(32'h3ae73d37),
	.w7(32'h3af2ad8b),
	.w8(32'h3bf91793),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f46e4b),
	.w1(32'hbab43edd),
	.w2(32'hbadae995),
	.w3(32'h3b734813),
	.w4(32'h3b0d8d50),
	.w5(32'hbbd631f9),
	.w6(32'h3bf58fb1),
	.w7(32'h3bbf2ec9),
	.w8(32'hbc24f29d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce7a81),
	.w1(32'h3bb0038a),
	.w2(32'h3b2db5dc),
	.w3(32'h3bccea0b),
	.w4(32'h3bd8dcee),
	.w5(32'h3b2af225),
	.w6(32'hbb34e7fc),
	.w7(32'h3b5204d6),
	.w8(32'h39c718b2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1faa3b),
	.w1(32'h3b04612c),
	.w2(32'hbb821d33),
	.w3(32'h3af62e36),
	.w4(32'h3b95d3c9),
	.w5(32'h3a06c2c7),
	.w6(32'h3b2d6027),
	.w7(32'h3bd395f5),
	.w8(32'hb98bd511),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaad397),
	.w1(32'hb9b9b0a7),
	.w2(32'hbc04a282),
	.w3(32'h3bd73250),
	.w4(32'h3beeaa9b),
	.w5(32'hbbc1a642),
	.w6(32'h3b52d2fb),
	.w7(32'h3b0638f0),
	.w8(32'h3bb208bd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc105eb0),
	.w1(32'hbc250c67),
	.w2(32'hbc0c6b86),
	.w3(32'hbc3fbee0),
	.w4(32'hbc1fa31b),
	.w5(32'hbbb15887),
	.w6(32'hbb4a2af0),
	.w7(32'hb92d3a02),
	.w8(32'hbbc2c6b6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a7fc9),
	.w1(32'hbb11c755),
	.w2(32'hbbeeb5c7),
	.w3(32'h3abbfed9),
	.w4(32'h3b0f0849),
	.w5(32'hbbbec9da),
	.w6(32'h3ae5d5a2),
	.w7(32'h3b27d4ba),
	.w8(32'hbb7565ad),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54d848),
	.w1(32'hbb378bf1),
	.w2(32'h3ab23962),
	.w3(32'hbb6d2396),
	.w4(32'h39b5a9d0),
	.w5(32'h3b51f6bb),
	.w6(32'hbb60a890),
	.w7(32'h3a1123a8),
	.w8(32'hbb619c98),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97a017),
	.w1(32'hbb1e9852),
	.w2(32'hbb29b508),
	.w3(32'h3b2d0e0f),
	.w4(32'hba2f33f2),
	.w5(32'hbb5e940f),
	.w6(32'h3a80a389),
	.w7(32'h3b0ed5e8),
	.w8(32'h3a0bef03),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2606ff),
	.w1(32'hbb9b3f78),
	.w2(32'h3ac6b184),
	.w3(32'hbbedcb6f),
	.w4(32'hbb97117b),
	.w5(32'h3bc59bf6),
	.w6(32'hbb923d2e),
	.w7(32'hbbafc4aa),
	.w8(32'h3be3b2ca),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6e5cc),
	.w1(32'hbae61e90),
	.w2(32'hbc03260e),
	.w3(32'hba37a8e5),
	.w4(32'hbab17329),
	.w5(32'hbba4a34b),
	.w6(32'h3bed0810),
	.w7(32'hb936f33c),
	.w8(32'hbb923533),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb374042),
	.w1(32'hbab0071e),
	.w2(32'hbb52a793),
	.w3(32'h3a31aa97),
	.w4(32'h3b1cab71),
	.w5(32'hbb81f63c),
	.w6(32'h3a45c69d),
	.w7(32'h3b35abbd),
	.w8(32'hbb45b545),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70e89e),
	.w1(32'hbb233b7a),
	.w2(32'hba5f17a7),
	.w3(32'hbbe3f741),
	.w4(32'hbbfc5048),
	.w5(32'hbbb6d341),
	.w6(32'hbb1afc56),
	.w7(32'hbad361f3),
	.w8(32'h3abcde27),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a5916),
	.w1(32'hbc3dd484),
	.w2(32'hbabf09fd),
	.w3(32'hbc844556),
	.w4(32'hbc606bab),
	.w5(32'h3b0d29a2),
	.w6(32'hbc587894),
	.w7(32'hbc4a49b8),
	.w8(32'h3bd35c1d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19bff5),
	.w1(32'hba38fd20),
	.w2(32'hbc09d434),
	.w3(32'h3b8d3fc1),
	.w4(32'h3b5ba5e8),
	.w5(32'hbc5c08e0),
	.w6(32'h3c18c325),
	.w7(32'h3acd9998),
	.w8(32'hbc30dcdf),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e3fa7),
	.w1(32'hbc5cbff2),
	.w2(32'hb9d428a1),
	.w3(32'hbc9abd9e),
	.w4(32'hbc8b5bbc),
	.w5(32'h39b9a5d5),
	.w6(32'hbc9192e4),
	.w7(32'hbc41b361),
	.w8(32'hbadfa6ca),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29779e),
	.w1(32'hba5de4de),
	.w2(32'hbbacc18d),
	.w3(32'h3b20777e),
	.w4(32'h3983029a),
	.w5(32'hbb37e7f0),
	.w6(32'hbacd288c),
	.w7(32'hbb91cbce),
	.w8(32'hba92e816),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9a5b6),
	.w1(32'hbc060744),
	.w2(32'h3bf656a2),
	.w3(32'hbc02b7dc),
	.w4(32'h3a5294a2),
	.w5(32'hbb4f13ce),
	.w6(32'hbbbb656c),
	.w7(32'hbb1fb7de),
	.w8(32'hbbda8013),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6d128),
	.w1(32'h3b6f4e74),
	.w2(32'h3b1a76be),
	.w3(32'h3a629434),
	.w4(32'h3abda02c),
	.w5(32'hbbc2fafe),
	.w6(32'hba62aa57),
	.w7(32'h3abc8b5d),
	.w8(32'hbbd5a56d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0268e),
	.w1(32'hbad83d56),
	.w2(32'hbb0cc229),
	.w3(32'hbb2e1b0c),
	.w4(32'hbb6f43f9),
	.w5(32'hbb19c5b2),
	.w6(32'hbb0755e4),
	.w7(32'h3bb7119f),
	.w8(32'hbb0141fc),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32c6fd),
	.w1(32'h3b584df5),
	.w2(32'hb8e63373),
	.w3(32'hbb436487),
	.w4(32'h3b2b4398),
	.w5(32'hbb162014),
	.w6(32'hbbaae690),
	.w7(32'h3b0efb21),
	.w8(32'hbbaaacf1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23c329),
	.w1(32'hb9fbb790),
	.w2(32'hbb8e9d78),
	.w3(32'hba30b576),
	.w4(32'h3a285b6b),
	.w5(32'hbb43be57),
	.w6(32'h3b848b58),
	.w7(32'h3bec979f),
	.w8(32'hbb411a0a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53451b),
	.w1(32'h3a72db1b),
	.w2(32'hbbe5e2b8),
	.w3(32'h39ab6243),
	.w4(32'hbaee2c43),
	.w5(32'hbb773034),
	.w6(32'hbab86379),
	.w7(32'hbb787515),
	.w8(32'hbb332c1e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd176e),
	.w1(32'h3a60f804),
	.w2(32'h3a4a6b8a),
	.w3(32'h39642f30),
	.w4(32'hba8ef69b),
	.w5(32'h3b2030ca),
	.w6(32'h3b339671),
	.w7(32'hbacaf09b),
	.w8(32'h3b9c2259),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae45168),
	.w1(32'hbbed3bca),
	.w2(32'h3a3e3a72),
	.w3(32'h3b3a8bd9),
	.w4(32'hba196c77),
	.w5(32'h3a51bcc3),
	.w6(32'h3b2c381a),
	.w7(32'h3a5bb32d),
	.w8(32'h3b08fa91),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb932a2),
	.w1(32'h3c079804),
	.w2(32'h3b0609f1),
	.w3(32'hba3afda3),
	.w4(32'h3bb8264e),
	.w5(32'h3b9f042d),
	.w6(32'h3983619b),
	.w7(32'h3bb9aff0),
	.w8(32'h3bb70a4f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacea935),
	.w1(32'h3b52572b),
	.w2(32'hbb56502d),
	.w3(32'h3b82cc90),
	.w4(32'h3badbced),
	.w5(32'hbbd39717),
	.w6(32'h3a97cf65),
	.w7(32'h3b092f5e),
	.w8(32'hbba3ae35),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84c04b),
	.w1(32'h3af9e5bf),
	.w2(32'h3a28e3cc),
	.w3(32'hbbe663b7),
	.w4(32'hbae9b6ca),
	.w5(32'h3a41c598),
	.w6(32'hbb3a17d7),
	.w7(32'hba2812f8),
	.w8(32'h3a38aa67),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fbcce),
	.w1(32'hbb2f8188),
	.w2(32'hbb3d6653),
	.w3(32'hba32e909),
	.w4(32'hbaafab3f),
	.w5(32'hbafb10f7),
	.w6(32'hba4d6544),
	.w7(32'hbad2cb2f),
	.w8(32'hbb62cbc6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48078c),
	.w1(32'hbb570d61),
	.w2(32'hbae9dfd4),
	.w3(32'h3b43b080),
	.w4(32'hbabfbcec),
	.w5(32'hbb29c2f6),
	.w6(32'h3b323f83),
	.w7(32'hbb13ec30),
	.w8(32'h3981cda8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d294a),
	.w1(32'hbb055d82),
	.w2(32'hb967529c),
	.w3(32'hbb721096),
	.w4(32'hbb7328dd),
	.w5(32'hba2ee2d7),
	.w6(32'hba9fb7c8),
	.w7(32'hbb49371d),
	.w8(32'h39e7a61a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cefe5),
	.w1(32'h3b3f714b),
	.w2(32'h39a66b4c),
	.w3(32'hb987d964),
	.w4(32'h3b170731),
	.w5(32'h3b9412ab),
	.w6(32'h3943f1bc),
	.w7(32'h3b6fad9c),
	.w8(32'h3b1809d9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd50583),
	.w1(32'hbad23f29),
	.w2(32'hbc6e8ebd),
	.w3(32'h3c153ba8),
	.w4(32'h3acaa0d5),
	.w5(32'hbc8a94e5),
	.w6(32'h3c0d3303),
	.w7(32'h3a9244a2),
	.w8(32'hbc526bd3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8d60c),
	.w1(32'hbb4227e9),
	.w2(32'h3b2bb82e),
	.w3(32'h3af31361),
	.w4(32'hbb8e8b0e),
	.w5(32'hb81e7f88),
	.w6(32'h3b904f99),
	.w7(32'hbb86a0b6),
	.w8(32'hba3f5aea),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b633646),
	.w1(32'h3a7cec7f),
	.w2(32'h3a208b87),
	.w3(32'h3b01e8db),
	.w4(32'h3a0d3cdf),
	.w5(32'hb8afadf1),
	.w6(32'hba2ef4d8),
	.w7(32'hbb07ce71),
	.w8(32'hb95e37a7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca059),
	.w1(32'hbb8a26bf),
	.w2(32'h3abc89ef),
	.w3(32'hbbc9e321),
	.w4(32'hbc06bde1),
	.w5(32'hb95c0436),
	.w6(32'hbb90de15),
	.w7(32'hbb6e4bb0),
	.w8(32'h3ad6176c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad88fb5),
	.w1(32'hbaa91983),
	.w2(32'hbb7397d3),
	.w3(32'h3ab25744),
	.w4(32'h3b411dce),
	.w5(32'hbad23805),
	.w6(32'h3af96b97),
	.w7(32'h3baaaba9),
	.w8(32'hbb2872e0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383dc8d3),
	.w1(32'h39ca958f),
	.w2(32'hbb826617),
	.w3(32'h3b2da809),
	.w4(32'h3b72c30f),
	.w5(32'hbbd59ae8),
	.w6(32'h3b0acbaf),
	.w7(32'h3b96f726),
	.w8(32'hbb7221e1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a252d04),
	.w1(32'h3b3b8ee9),
	.w2(32'hbc0cad39),
	.w3(32'hbb32ba78),
	.w4(32'h394d18af),
	.w5(32'hbc819231),
	.w6(32'hbb171f6b),
	.w7(32'h3a9a8f3d),
	.w8(32'hbbfb12d3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7885bd),
	.w1(32'hbc3ac264),
	.w2(32'hbc0786b9),
	.w3(32'hbc90b745),
	.w4(32'hbc8d7960),
	.w5(32'hbc448dc4),
	.w6(32'hbc4badb6),
	.w7(32'hbc133e33),
	.w8(32'hbae6f3be),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6126e4),
	.w1(32'hbc055496),
	.w2(32'h3b69aa84),
	.w3(32'hbc74f6e7),
	.w4(32'hbc25740a),
	.w5(32'h3b11d9ff),
	.w6(32'hbc09a890),
	.w7(32'hbbc86284),
	.w8(32'h3bdf93ce),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b602ffc),
	.w1(32'hbb0720c1),
	.w2(32'h3a93761a),
	.w3(32'h3b3e7dff),
	.w4(32'hba58a97e),
	.w5(32'h3b85131b),
	.w6(32'h3ba8c31c),
	.w7(32'h3b4c9444),
	.w8(32'h3af5717b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b803f2a),
	.w1(32'hba03fb88),
	.w2(32'hbb1f03e3),
	.w3(32'h3b9dd986),
	.w4(32'hba4f8910),
	.w5(32'hbb383cdf),
	.w6(32'h3b10af72),
	.w7(32'hb9d02f82),
	.w8(32'hbaca3842),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5c2d9),
	.w1(32'hbab739f1),
	.w2(32'h3a149073),
	.w3(32'h39e82e52),
	.w4(32'hbb132313),
	.w5(32'hba9273dd),
	.w6(32'h3a9f33e0),
	.w7(32'hbb8ffecb),
	.w8(32'hbac26ca4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75bfb6),
	.w1(32'hba8aee7e),
	.w2(32'hbacfde21),
	.w3(32'h3b68b39c),
	.w4(32'hbad9dcf3),
	.w5(32'h38f4c0bd),
	.w6(32'h3b3116b0),
	.w7(32'hbb1f0147),
	.w8(32'hb8d7538c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be8ee5),
	.w1(32'hbac32044),
	.w2(32'h3c0dd568),
	.w3(32'hbb5d8865),
	.w4(32'hbaf080b2),
	.w5(32'h3be6d22d),
	.w6(32'hba9493b7),
	.w7(32'hbb250a45),
	.w8(32'h3bf8896d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29e0ba),
	.w1(32'hbbad0713),
	.w2(32'h39d6f1e7),
	.w3(32'h3b4e80cc),
	.w4(32'hbb25d8bb),
	.w5(32'hbb087911),
	.w6(32'h3c00a61a),
	.w7(32'h38b14d90),
	.w8(32'hbb7874ec),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb699ad3),
	.w1(32'hbc0402f9),
	.w2(32'h38f5cbd2),
	.w3(32'hbc205cac),
	.w4(32'hbbd87af3),
	.w5(32'hba953949),
	.w6(32'hbbb39ea2),
	.w7(32'hbc1bf347),
	.w8(32'h3a69ffdd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d2d9f),
	.w1(32'hbab790a7),
	.w2(32'h3b3b8877),
	.w3(32'hbbc2138a),
	.w4(32'hbb0c77f9),
	.w5(32'h3b4d0d4e),
	.w6(32'hbb74f382),
	.w7(32'hbb1d2269),
	.w8(32'h3b6766b4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c5080),
	.w1(32'h3ac742ab),
	.w2(32'hb9d8cdc1),
	.w3(32'h3b9aeaad),
	.w4(32'h3b31d1a0),
	.w5(32'h39887ede),
	.w6(32'h3bad62b4),
	.w7(32'h3b6fb4d8),
	.w8(32'h3aa131ea),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c4fcb),
	.w1(32'h3a0ff619),
	.w2(32'hba30b547),
	.w3(32'h3a8c75ca),
	.w4(32'h3a85deba),
	.w5(32'hbb0dd5c5),
	.w6(32'h3ad0d8ac),
	.w7(32'h3b0125b9),
	.w8(32'hbb0257e5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc315519),
	.w1(32'hbc1c3887),
	.w2(32'hbac62eed),
	.w3(32'hbc7e0680),
	.w4(32'hbc3288a2),
	.w5(32'hbab23c3f),
	.w6(32'hbc11523a),
	.w7(32'hbc36ca2d),
	.w8(32'hbbfe9582),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b056d47),
	.w1(32'hbb482d6f),
	.w2(32'hbb64a700),
	.w3(32'h3b6c43b4),
	.w4(32'h3a918220),
	.w5(32'hbc31bc55),
	.w6(32'h3ace7325),
	.w7(32'hba8f72c7),
	.w8(32'hbc11cbff),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b180475),
	.w1(32'h3a90fcf1),
	.w2(32'hba8f8414),
	.w3(32'hbb5ccbaa),
	.w4(32'hbafe67aa),
	.w5(32'hbb2a30be),
	.w6(32'hbb12dced),
	.w7(32'h39b418d2),
	.w8(32'hbbaa95a6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58546b),
	.w1(32'h3a0b64c6),
	.w2(32'hba59dadc),
	.w3(32'h3b655472),
	.w4(32'hb9b4cb28),
	.w5(32'h3b2e8ed5),
	.w6(32'h3b089403),
	.w7(32'hbb448476),
	.w8(32'h3b151ac7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a329d),
	.w1(32'hb9b7b190),
	.w2(32'hbad72397),
	.w3(32'h3b94b567),
	.w4(32'h3b3bb3c8),
	.w5(32'hb8f2ddb7),
	.w6(32'h3b941a71),
	.w7(32'h3b44ea6b),
	.w8(32'h388231ff),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19547a),
	.w1(32'h3a862193),
	.w2(32'h3b41c957),
	.w3(32'h3b537b78),
	.w4(32'h3aaf2664),
	.w5(32'hb9d2a0b9),
	.w6(32'h3b5eab63),
	.w7(32'h3a969a50),
	.w8(32'h3a5ac459),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7720f3),
	.w1(32'h3b21f5a5),
	.w2(32'hb96be3ce),
	.w3(32'h3a8e23f2),
	.w4(32'h3b1cb7d1),
	.w5(32'hb9b8d686),
	.w6(32'hbaad68d2),
	.w7(32'hbaba27d7),
	.w8(32'hbac2a65c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b2d14),
	.w1(32'h3bc35e71),
	.w2(32'h3adc51e1),
	.w3(32'hbbeccf76),
	.w4(32'hbb2f9e2c),
	.w5(32'h3a8c1a5d),
	.w6(32'hbc20cc97),
	.w7(32'hbb06b6b6),
	.w8(32'h3928d277),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65e2bd),
	.w1(32'h3b17e2fb),
	.w2(32'hbc6069af),
	.w3(32'h3ad758e3),
	.w4(32'h3bc24476),
	.w5(32'hbc484a3c),
	.w6(32'hbaf32833),
	.w7(32'h3be9e0c2),
	.w8(32'hbb386a56),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc834132),
	.w1(32'hbc854464),
	.w2(32'h3b1b6917),
	.w3(32'hbc8c5d09),
	.w4(32'hbc6acabe),
	.w5(32'h3ba73390),
	.w6(32'hbc6e7b74),
	.w7(32'hbc47d769),
	.w8(32'h3b9ac73d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52dbf7),
	.w1(32'hbaddc2b6),
	.w2(32'hbaf0a50d),
	.w3(32'hbab3d538),
	.w4(32'hbbcc97e5),
	.w5(32'hb9fa1e90),
	.w6(32'hb91006de),
	.w7(32'hbb1380c0),
	.w8(32'hbb8efbba),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b8aff),
	.w1(32'h3b4a7942),
	.w2(32'hbbb48276),
	.w3(32'hbb0462d1),
	.w4(32'h3b7e9e99),
	.w5(32'hbc218794),
	.w6(32'hbb2d5b84),
	.w7(32'h3ab2c9d7),
	.w8(32'hbb0c5f6c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfcdd9),
	.w1(32'hbb23191d),
	.w2(32'hbbd62bed),
	.w3(32'hbc201520),
	.w4(32'hbbfab1bb),
	.w5(32'hbbfee065),
	.w6(32'hbb1f6547),
	.w7(32'h3afd3fd9),
	.w8(32'hbb16c5f2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcd2d5),
	.w1(32'hbbfae653),
	.w2(32'hbb49675a),
	.w3(32'hbc0ea263),
	.w4(32'hbbcbd574),
	.w5(32'hbb34c7cc),
	.w6(32'hbaf41225),
	.w7(32'h3a951896),
	.w8(32'h3a498558),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f013cd),
	.w1(32'h3a8befac),
	.w2(32'hbafe604b),
	.w3(32'h3b7c6bc4),
	.w4(32'hba92ce6d),
	.w5(32'h38c177a3),
	.w6(32'h3b98b656),
	.w7(32'hbab5e93d),
	.w8(32'h3b1cde7e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24df87),
	.w1(32'h3b5c727d),
	.w2(32'h3c033dc4),
	.w3(32'hbaa22f5c),
	.w4(32'h3a680991),
	.w5(32'h3c21098d),
	.w6(32'hbae8c681),
	.w7(32'hba23bf73),
	.w8(32'h3c4ecb6b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd5e71),
	.w1(32'hba837cbb),
	.w2(32'hbb071d11),
	.w3(32'hba5bee6a),
	.w4(32'hbba8fedd),
	.w5(32'hb9b3321a),
	.w6(32'h3a711b65),
	.w7(32'hbb5c63a9),
	.w8(32'h390a0280),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacecba3),
	.w1(32'h3a641222),
	.w2(32'hbb9f38ce),
	.w3(32'hbadc1db8),
	.w4(32'h39a89065),
	.w5(32'hbb8076d3),
	.w6(32'hbae7736d),
	.w7(32'hbb012bdd),
	.w8(32'hbb0a6d0b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e9065),
	.w1(32'hba4f104f),
	.w2(32'h3b32b200),
	.w3(32'hbb744212),
	.w4(32'hba664b74),
	.w5(32'h3bac7c8f),
	.w6(32'hbb87bdd5),
	.w7(32'hba7f970e),
	.w8(32'h3b2abc62),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1d1dd),
	.w1(32'h3b21f28e),
	.w2(32'hba6ebfe1),
	.w3(32'h3b72ce09),
	.w4(32'h3c082f4f),
	.w5(32'hbb9a88c6),
	.w6(32'h3b54daeb),
	.w7(32'h3c06b04c),
	.w8(32'hbb97f9ca),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb471240),
	.w1(32'h38ec1f99),
	.w2(32'hba9dae0b),
	.w3(32'hbbd2b21d),
	.w4(32'h38beda01),
	.w5(32'h3a472060),
	.w6(32'hbc2bfb2f),
	.w7(32'h3ae5260e),
	.w8(32'h3b95e020),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa19db),
	.w1(32'hbb87c2b7),
	.w2(32'hbc5c1b7f),
	.w3(32'h3a46128f),
	.w4(32'hbb7a0e5c),
	.w5(32'hbc7f64e3),
	.w6(32'h3b3cec68),
	.w7(32'h3b2bdb8a),
	.w8(32'hbc364a32),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc909883),
	.w1(32'hbc8d598d),
	.w2(32'h3a1f6ce5),
	.w3(32'hbcafdb49),
	.w4(32'hbc9020bd),
	.w5(32'h3a2f0fa4),
	.w6(32'hbc7b2e36),
	.w7(32'hbc628b01),
	.w8(32'h3b24fbb1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe65e42),
	.w1(32'h3a64bcf1),
	.w2(32'h3bed113e),
	.w3(32'hbb184f1d),
	.w4(32'h3aed5df8),
	.w5(32'h3ba11789),
	.w6(32'h3a716761),
	.w7(32'h3b01c2c2),
	.w8(32'h3b49d47c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbefbd3),
	.w1(32'h3b8a04b7),
	.w2(32'hbac3b53b),
	.w3(32'h3b926ec8),
	.w4(32'hb932ff0a),
	.w5(32'hbb39d242),
	.w6(32'h3b91170c),
	.w7(32'hbaf4c150),
	.w8(32'hbb06f104),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb800796b),
	.w1(32'hbbd7385f),
	.w2(32'hba3ea255),
	.w3(32'hbb8b1a21),
	.w4(32'hbb9bb0df),
	.w5(32'hbbfeee4d),
	.w6(32'hbb7d842a),
	.w7(32'hbb86b2c4),
	.w8(32'hbc2d877d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc0f31),
	.w1(32'h3a123535),
	.w2(32'hbbb23751),
	.w3(32'hba464c02),
	.w4(32'h3b2dacc8),
	.w5(32'hbaf11427),
	.w6(32'hbb80b30d),
	.w7(32'hbadc2e8e),
	.w8(32'hb95f3e56),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96bc79),
	.w1(32'hbabf2436),
	.w2(32'hbc50a99c),
	.w3(32'hbaf26b5c),
	.w4(32'hb9c33e17),
	.w5(32'hbbca730d),
	.w6(32'h3aa38ccc),
	.w7(32'h3adea34c),
	.w8(32'hbbe4d5d8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bc6c3),
	.w1(32'hbba70e93),
	.w2(32'hbb8fca40),
	.w3(32'h3b163775),
	.w4(32'h3b28a964),
	.w5(32'h3a2c2ae8),
	.w6(32'h39cdec69),
	.w7(32'h3a96d94a),
	.w8(32'hba7a5317),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d0f85),
	.w1(32'hbb4b402b),
	.w2(32'hbb34aa4b),
	.w3(32'h3b34df0b),
	.w4(32'h3ac082c5),
	.w5(32'hbaf795ca),
	.w6(32'h3b04ddd4),
	.w7(32'h3a7da9e2),
	.w8(32'h3c25f168),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92ba64),
	.w1(32'hba14c558),
	.w2(32'hbbd981e0),
	.w3(32'hbbe4e370),
	.w4(32'hbbce4d1d),
	.w5(32'hbbb237db),
	.w6(32'h3c0953d1),
	.w7(32'h3c169394),
	.w8(32'hba17cd10),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd074ee),
	.w1(32'hbb930a39),
	.w2(32'h3ac39d62),
	.w3(32'hbbdeaede),
	.w4(32'hbb8b9938),
	.w5(32'h39f0e78c),
	.w6(32'h383ae507),
	.w7(32'h3bdaaf02),
	.w8(32'h3a6da329),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb04211),
	.w1(32'h3b9561b7),
	.w2(32'h3afca9d3),
	.w3(32'hba855f4f),
	.w4(32'h3b8d8302),
	.w5(32'h3a2225b6),
	.w6(32'hba1171da),
	.w7(32'h3a9a28af),
	.w8(32'h38c1573e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb1b80),
	.w1(32'h3aa514ce),
	.w2(32'hbb1f156c),
	.w3(32'h39c64847),
	.w4(32'h3a89f2b2),
	.w5(32'hbb74a4f6),
	.w6(32'h3a21d13f),
	.w7(32'h3aa27aff),
	.w8(32'hbafce767),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bbcb8),
	.w1(32'hb9cc12d3),
	.w2(32'h3bc2d0b9),
	.w3(32'hbb90f8be),
	.w4(32'hbb3174f0),
	.w5(32'h3c109f81),
	.w6(32'hbb58d2c8),
	.w7(32'hba32d7a1),
	.w8(32'h3c7403e7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86a644),
	.w1(32'hbb09efba),
	.w2(32'hbabcbbd8),
	.w3(32'h3bc6c4b3),
	.w4(32'hbb366091),
	.w5(32'h3a3763e0),
	.w6(32'h3becf482),
	.w7(32'hbaacdfdb),
	.w8(32'hb90528cb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e96f4),
	.w1(32'h3a9f88f7),
	.w2(32'hb9e65b16),
	.w3(32'hb82f012e),
	.w4(32'h3aa49adf),
	.w5(32'h3b0b54e5),
	.w6(32'hbae88375),
	.w7(32'h3a4698cd),
	.w8(32'h3c042379),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a147c),
	.w1(32'hbb3cb35b),
	.w2(32'h3bc0729b),
	.w3(32'hbb650eb7),
	.w4(32'hbbcaa561),
	.w5(32'h3bdbaf47),
	.w6(32'hbacfe2ab),
	.w7(32'hbbb2b2df),
	.w8(32'h3b7fa48f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae30845),
	.w1(32'hbb71a24a),
	.w2(32'hbb7e4ce4),
	.w3(32'hbb55250d),
	.w4(32'hbbcee4df),
	.w5(32'hbbaad2f2),
	.w6(32'h3809da09),
	.w7(32'hbb6fee0e),
	.w8(32'hbac85c3d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc505f),
	.w1(32'hbba2c27a),
	.w2(32'h3af698fb),
	.w3(32'hbc28d2e0),
	.w4(32'hbb9c8799),
	.w5(32'h3aea3853),
	.w6(32'hbbfea160),
	.w7(32'hbb4581fa),
	.w8(32'hba60f760),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0157f),
	.w1(32'h3bc02036),
	.w2(32'h3be62db3),
	.w3(32'h3b6feecf),
	.w4(32'h3be80b22),
	.w5(32'h3a097095),
	.w6(32'h3b17ee72),
	.w7(32'h3bbdb3cc),
	.w8(32'h3ab7f999),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b469b0d),
	.w1(32'h3bb75aad),
	.w2(32'h3b0ea7f2),
	.w3(32'hbaa317f8),
	.w4(32'h3b5c2a4d),
	.w5(32'h3ba96946),
	.w6(32'h3724ddd6),
	.w7(32'h3ae68668),
	.w8(32'h3aaef6e1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8764f4),
	.w1(32'hbb8820dd),
	.w2(32'hbbf8aa38),
	.w3(32'h3b8857b6),
	.w4(32'h3b11acef),
	.w5(32'hbc22d6e4),
	.w6(32'h3a9e00e9),
	.w7(32'h3ae5f138),
	.w8(32'hbbbf94f1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c7dcc),
	.w1(32'hbc35232f),
	.w2(32'hbba5cde7),
	.w3(32'hbc5b35f7),
	.w4(32'hbc278e20),
	.w5(32'h3b0d19d2),
	.w6(32'hbc6e7f57),
	.w7(32'hbc2509b8),
	.w8(32'hbba93b37),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc241b85),
	.w1(32'hbbf63177),
	.w2(32'hbb71f395),
	.w3(32'hbade229b),
	.w4(32'hbaf84e17),
	.w5(32'hbb8e8485),
	.w6(32'hbb90a363),
	.w7(32'hbbdb9e4a),
	.w8(32'hbb855064),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7072e),
	.w1(32'h3b7c98c1),
	.w2(32'hbbd07e96),
	.w3(32'h3b06271b),
	.w4(32'h3bc908cb),
	.w5(32'hbbbeb2da),
	.w6(32'hbb803929),
	.w7(32'h3bc520c5),
	.w8(32'hbbbc1e37),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8b639),
	.w1(32'hba5572e2),
	.w2(32'hbbb28466),
	.w3(32'h3a8fafef),
	.w4(32'h390de673),
	.w5(32'h3b888d9f),
	.w6(32'h39f25fea),
	.w7(32'h3aaeea19),
	.w8(32'h3b6df525),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac04035),
	.w1(32'hbb1a3cad),
	.w2(32'h3b059f46),
	.w3(32'h3b9a71ce),
	.w4(32'h3952c047),
	.w5(32'h3a3d6a23),
	.w6(32'h3b7e663f),
	.w7(32'hbb5caafe),
	.w8(32'h3abc8f57),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe60fe),
	.w1(32'hbbb49935),
	.w2(32'h3a3e0b98),
	.w3(32'h3b42534d),
	.w4(32'hba973098),
	.w5(32'hbb965edc),
	.w6(32'h3b4ad43f),
	.w7(32'h3a677cb6),
	.w8(32'hbb9dfe4c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b236120),
	.w1(32'h3bcb0c7e),
	.w2(32'h3a36cee4),
	.w3(32'hba9ccbb4),
	.w4(32'h3b4eafcb),
	.w5(32'hbaeff2f3),
	.w6(32'hbb2bb4b4),
	.w7(32'h3b3efe0b),
	.w8(32'hbaaba884),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a843c34),
	.w1(32'h3a084768),
	.w2(32'hbb7d94b8),
	.w3(32'hba9a6f68),
	.w4(32'hbaf1392d),
	.w5(32'hbc3810d9),
	.w6(32'hbaa5e23f),
	.w7(32'hbad9a71c),
	.w8(32'hbbd4499e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdf290),
	.w1(32'hbb948766),
	.w2(32'hbafc70fc),
	.w3(32'hbbf59910),
	.w4(32'hbb8efaea),
	.w5(32'hba9b139a),
	.w6(32'hbc346b94),
	.w7(32'hbbcb1028),
	.w8(32'h388bcb11),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a266090),
	.w1(32'h39aad1e5),
	.w2(32'hbc25c363),
	.w3(32'h3a51ac8f),
	.w4(32'h39ce4f2b),
	.w5(32'hbc5b9aa8),
	.w6(32'h3aa2d985),
	.w7(32'h3a556974),
	.w8(32'hbc462c48),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa82206),
	.w1(32'hb8afa554),
	.w2(32'hbb8e32d4),
	.w3(32'hbb14a616),
	.w4(32'h3a77387e),
	.w5(32'h3a81b240),
	.w6(32'hbbc7443d),
	.w7(32'hbaed83dd),
	.w8(32'h3bef7f4e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ed4f1),
	.w1(32'hba7b7f19),
	.w2(32'hbaf03f1d),
	.w3(32'h39dd8dd0),
	.w4(32'h3b92ad16),
	.w5(32'hba3ff6ee),
	.w6(32'h3b8b3f17),
	.w7(32'h3b97426e),
	.w8(32'hbb7dbd77),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a268c36),
	.w1(32'hbb39fec5),
	.w2(32'h3a02f710),
	.w3(32'h3af75fa3),
	.w4(32'hb9b43618),
	.w5(32'h39c0ee94),
	.w6(32'h3ac24aca),
	.w7(32'hbafbe924),
	.w8(32'h3a44529c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa008c),
	.w1(32'h39f6edef),
	.w2(32'h3b72d128),
	.w3(32'h3a9eaabb),
	.w4(32'hba167feb),
	.w5(32'h3bc104bf),
	.w6(32'h3a6690ff),
	.w7(32'hbaa919c5),
	.w8(32'hbae0ce84),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac45848),
	.w1(32'h3b8d439d),
	.w2(32'hbb5a9a6a),
	.w3(32'h3ba6ee85),
	.w4(32'h3c13ed2d),
	.w5(32'hbb4e4fb2),
	.w6(32'h3a836980),
	.w7(32'h3baa655f),
	.w8(32'hba825821),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1375e6),
	.w1(32'h3b9aadf4),
	.w2(32'h3b9a33dc),
	.w3(32'h3ac69d0e),
	.w4(32'h3b5d571c),
	.w5(32'h3b78732c),
	.w6(32'hbb5e4c36),
	.w7(32'h3b2c165a),
	.w8(32'h3bfa3704),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383bd2ae),
	.w1(32'hbb2ba605),
	.w2(32'hba5efef0),
	.w3(32'h3b14a274),
	.w4(32'hb986c906),
	.w5(32'hba737daf),
	.w6(32'h3bd20416),
	.w7(32'h3b9ae535),
	.w8(32'hb9838bd4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39371a69),
	.w1(32'h3ab2a272),
	.w2(32'hbc1e55f3),
	.w3(32'hb916114c),
	.w4(32'hb91b9018),
	.w5(32'hbc469751),
	.w6(32'hb913b9aa),
	.w7(32'hb962d6f0),
	.w8(32'hbc00ac0c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28427c),
	.w1(32'hbc34f621),
	.w2(32'hbb449934),
	.w3(32'hbcaba9ed),
	.w4(32'hbc864850),
	.w5(32'h3b044aa0),
	.w6(32'hbc807019),
	.w7(32'hbc6af823),
	.w8(32'h3ba4028a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac033f1),
	.w1(32'hb9f2c5c1),
	.w2(32'h3a26af5f),
	.w3(32'h3b75cda6),
	.w4(32'h3b0401e1),
	.w5(32'hbb20609a),
	.w6(32'h3b44266e),
	.w7(32'h3b734afd),
	.w8(32'hb769b3fe),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b4803),
	.w1(32'h3b07aaf4),
	.w2(32'hbc262910),
	.w3(32'hba0f2164),
	.w4(32'hb993e952),
	.w5(32'hbc03e693),
	.w6(32'h3ac1c4fc),
	.w7(32'h3ac3bf2c),
	.w8(32'hbc291095),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78228d),
	.w1(32'hbbcb8aa7),
	.w2(32'hbaba6a75),
	.w3(32'hbacb02d6),
	.w4(32'hbbf67ef5),
	.w5(32'h3b9d2ab6),
	.w6(32'hbbe799ac),
	.w7(32'hbc11460b),
	.w8(32'h3c0db247),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8556ea),
	.w1(32'hb8c730d0),
	.w2(32'hbc311afa),
	.w3(32'hbb000571),
	.w4(32'hba8dc344),
	.w5(32'hbc5c522f),
	.w6(32'h3b6102cf),
	.w7(32'h39f8a40c),
	.w8(32'hbc0ad467),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc619401),
	.w1(32'hbc2c9187),
	.w2(32'h3ac91284),
	.w3(32'hbc90adc4),
	.w4(32'hbc450dd5),
	.w5(32'h38a9d029),
	.w6(32'hbc6c873d),
	.w7(32'hbc1ab2fb),
	.w8(32'h3a86377a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3df5d9),
	.w1(32'h3a410d84),
	.w2(32'hbc738184),
	.w3(32'h3b809085),
	.w4(32'h3a11dddc),
	.w5(32'hbb04f341),
	.w6(32'h3b45da64),
	.w7(32'h3ad9e960),
	.w8(32'hbbedb3a3),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8c9fe),
	.w1(32'h3b986a51),
	.w2(32'hbbba7ab4),
	.w3(32'h3c74feb4),
	.w4(32'h3c0dd504),
	.w5(32'hb98a8aa7),
	.w6(32'h3c099309),
	.w7(32'h3be0bcde),
	.w8(32'h3c466fee),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c0386),
	.w1(32'hbbff5df3),
	.w2(32'h3ac4fe66),
	.w3(32'hbbef52e1),
	.w4(32'hbc4030e8),
	.w5(32'h3b8ca4d9),
	.w6(32'h3c200108),
	.w7(32'h3b8ffd5a),
	.w8(32'h3b5bbb8d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a465277),
	.w1(32'hb9bfa583),
	.w2(32'h3870c098),
	.w3(32'h3b6639b7),
	.w4(32'h3b18d89c),
	.w5(32'hbc772ece),
	.w6(32'h3b290125),
	.w7(32'h3b285695),
	.w8(32'hbc38ec0b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8f09d),
	.w1(32'hbb3bca97),
	.w2(32'h3af610f3),
	.w3(32'hbc9f8efe),
	.w4(32'hbc1a93fc),
	.w5(32'hbb24c1b5),
	.w6(32'hbc486b3b),
	.w7(32'hbc0a468c),
	.w8(32'hbca1d0dd),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c267de8),
	.w1(32'h3c123b6c),
	.w2(32'hba592af5),
	.w3(32'hbc2c755a),
	.w4(32'h3a22e44d),
	.w5(32'h3b23dd7d),
	.w6(32'hbc8e6ffa),
	.w7(32'hbc16f438),
	.w8(32'hbb06e2a2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6ffdf),
	.w1(32'hbb588aa5),
	.w2(32'h3c31319c),
	.w3(32'h397907db),
	.w4(32'h3ac1a8de),
	.w5(32'h3b90cd15),
	.w6(32'hbb6840af),
	.w7(32'hbb1c539b),
	.w8(32'hbb58f5af),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beca552),
	.w1(32'hbc143fb3),
	.w2(32'h3b6e2082),
	.w3(32'hbc64f6e7),
	.w4(32'hbceb7128),
	.w5(32'h3c204bd6),
	.w6(32'hbcbf5cf5),
	.w7(32'hbcc4c289),
	.w8(32'h3bdd9450),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be83bb2),
	.w1(32'h3bf04955),
	.w2(32'hbc382000),
	.w3(32'h3c3d5163),
	.w4(32'h3c1271ab),
	.w5(32'h3bd1166b),
	.w6(32'h3c168aee),
	.w7(32'h3c1053ab),
	.w8(32'h3c3c214d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad834f6),
	.w1(32'h3ae28383),
	.w2(32'hbbb0a1d3),
	.w3(32'h3c42744b),
	.w4(32'h3c1517b0),
	.w5(32'h3b012fda),
	.w6(32'h3c62d22a),
	.w7(32'h3bf8015a),
	.w8(32'hbb89253e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a818b58),
	.w1(32'hbb51a9a7),
	.w2(32'hbc12b00e),
	.w3(32'h3bcd9fd2),
	.w4(32'h3a7008cf),
	.w5(32'hbb928142),
	.w6(32'hba92013d),
	.w7(32'hbb05f042),
	.w8(32'h3c863fd1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef6e3f),
	.w1(32'hb8c8a514),
	.w2(32'hbbeffe5a),
	.w3(32'hbaa34cc1),
	.w4(32'hbbf47e1f),
	.w5(32'hbc3e4b25),
	.w6(32'h3c4b1b0b),
	.w7(32'hba38f0d0),
	.w8(32'hbbd5e7f4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19bb21),
	.w1(32'h3c8ca627),
	.w2(32'h3bb9f61f),
	.w3(32'h3bed1776),
	.w4(32'h3cb9dae4),
	.w5(32'h3b95ae97),
	.w6(32'h3bcf3f5f),
	.w7(32'h3c59887f),
	.w8(32'h3bbabf02),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e53cb),
	.w1(32'h3910a48e),
	.w2(32'hbb4d327a),
	.w3(32'h3b9f793a),
	.w4(32'h3b3b3faa),
	.w5(32'h3c0a66d9),
	.w6(32'h3aa22b56),
	.w7(32'h3a7e2c2c),
	.w8(32'h3b3c026f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae9232),
	.w1(32'hbbd8a283),
	.w2(32'hbbcb1990),
	.w3(32'h3bb4dc74),
	.w4(32'hbb377771),
	.w5(32'hbc92439d),
	.w6(32'h3afbe8b4),
	.w7(32'hbb73f1b4),
	.w8(32'h3bf5e4b9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d95eb),
	.w1(32'hba70b0e9),
	.w2(32'hbb3e1b12),
	.w3(32'hbce71f29),
	.w4(32'hbb9e44f1),
	.w5(32'hb96c1fe3),
	.w6(32'hb78576e9),
	.w7(32'h3a3eb57e),
	.w8(32'hb9b1263d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aba71),
	.w1(32'h3b6c76a5),
	.w2(32'h3bb8eb7f),
	.w3(32'h3bf1f85a),
	.w4(32'h3bc3e06f),
	.w5(32'hba266891),
	.w6(32'h3be362b5),
	.w7(32'h3bfcc8e4),
	.w8(32'h3b830a4e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82523e),
	.w1(32'hbc49d922),
	.w2(32'h3bab19cc),
	.w3(32'hbc8da328),
	.w4(32'hbcc6cbcb),
	.w5(32'h3b9434ad),
	.w6(32'hbc34cf80),
	.w7(32'hbad53ff5),
	.w8(32'h3bed59c7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ba222),
	.w1(32'h3b27be7a),
	.w2(32'hbc83122b),
	.w3(32'h3bdddf48),
	.w4(32'h3bb5084c),
	.w5(32'hbcb20a85),
	.w6(32'h3c11b82e),
	.w7(32'h3c84fdf3),
	.w8(32'hbbb2a080),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc278cc8),
	.w1(32'hbb9793ec),
	.w2(32'hba07575b),
	.w3(32'hbd008e31),
	.w4(32'hbc2ea8e8),
	.w5(32'h3c5d8ef9),
	.w6(32'hbc9e473e),
	.w7(32'hbb8b6911),
	.w8(32'h3c768e6a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc864ddf),
	.w1(32'hbc091655),
	.w2(32'hbb212a7f),
	.w3(32'hbcc632e9),
	.w4(32'hbcaadc3f),
	.w5(32'hbb7009e3),
	.w6(32'hbbce7f9c),
	.w7(32'hbc3c2d29),
	.w8(32'hbb63339c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfcc43),
	.w1(32'h3a90e6e8),
	.w2(32'hb9e21ad0),
	.w3(32'h3a1342ab),
	.w4(32'hbaa848df),
	.w5(32'hbba5795b),
	.w6(32'hba4dc578),
	.w7(32'h3ace24e1),
	.w8(32'hbad4ba82),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7df973),
	.w1(32'h3b860d0a),
	.w2(32'h3c25433a),
	.w3(32'hbc427a98),
	.w4(32'hbc375949),
	.w5(32'h3ba57eb1),
	.w6(32'hbc04ac2a),
	.w7(32'hbbb74148),
	.w8(32'h3a3fba80),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaf2c1),
	.w1(32'hbbbfd0ef),
	.w2(32'hbc00aa1e),
	.w3(32'hbc3484d0),
	.w4(32'hbc8258be),
	.w5(32'hbcc13d16),
	.w6(32'h3acd9146),
	.w7(32'h3a9987a7),
	.w8(32'hbc3329f4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d7f87),
	.w1(32'hbaf41b89),
	.w2(32'h3bacf24b),
	.w3(32'hbc2cdfa0),
	.w4(32'h3bf271d4),
	.w5(32'h3a66d15c),
	.w6(32'h3bc257dd),
	.w7(32'h3c954014),
	.w8(32'hbbfaa9d9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94858e8),
	.w1(32'hbb89cb1a),
	.w2(32'hbaa96761),
	.w3(32'hbc0f63bb),
	.w4(32'hbc271571),
	.w5(32'hba830472),
	.w6(32'hbb163c7f),
	.w7(32'hbbfc11e4),
	.w8(32'hbc31bc6e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e4da1),
	.w1(32'hbb4d0d7a),
	.w2(32'hbc55c65f),
	.w3(32'hbbf8a1f6),
	.w4(32'hba5f92db),
	.w5(32'h3b415f72),
	.w6(32'hbbf6fb45),
	.w7(32'hbb692de6),
	.w8(32'h3c89f4b0),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbbd4b),
	.w1(32'hbbc3bc64),
	.w2(32'h3c72fc57),
	.w3(32'h3b2f583b),
	.w4(32'h3a854843),
	.w5(32'h3ca0870e),
	.w6(32'h3c931d0b),
	.w7(32'hbc1dd470),
	.w8(32'hbb46fb27),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c756578),
	.w1(32'h3b8de786),
	.w2(32'hbc25653c),
	.w3(32'h3c40a320),
	.w4(32'hbbd3f1c4),
	.w5(32'hbcaffccf),
	.w6(32'hbc57d15a),
	.w7(32'hbc19d6f1),
	.w8(32'hbc649c52),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bbed18),
	.w1(32'h3c9304b7),
	.w2(32'h3bacb2f9),
	.w3(32'hbc23aae2),
	.w4(32'h3bb35507),
	.w5(32'h3aad234e),
	.w6(32'hbc6e08ab),
	.w7(32'hbaabb5ae),
	.w8(32'h3b3b3f51),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b548108),
	.w1(32'hbb6ce63c),
	.w2(32'h3b5c46dc),
	.w3(32'h38dc62bf),
	.w4(32'hbba9e581),
	.w5(32'h3b898f74),
	.w6(32'h3b290fab),
	.w7(32'hbb938f63),
	.w8(32'hbb9c4047),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea8655),
	.w1(32'hbc1b0f4c),
	.w2(32'hbc027a4b),
	.w3(32'h3c22e64c),
	.w4(32'hbbbf6778),
	.w5(32'hbb2060f6),
	.w6(32'h3ad0d4ea),
	.w7(32'hbc89a5eb),
	.w8(32'hbb8d0b54),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02f0cd),
	.w1(32'hbbe3854a),
	.w2(32'hbb79006f),
	.w3(32'h3a5de429),
	.w4(32'hbaf0bff9),
	.w5(32'h39f9659a),
	.w6(32'h3ab63aa2),
	.w7(32'h3b2ad455),
	.w8(32'h3c26245b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb417b8c),
	.w1(32'hba8ed58c),
	.w2(32'hbc6b3ec8),
	.w3(32'hb829a17e),
	.w4(32'h3966f41d),
	.w5(32'hbc263d14),
	.w6(32'h3bd6c935),
	.w7(32'h3b8564da),
	.w8(32'h3ae5148f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fac13),
	.w1(32'hbbb3974e),
	.w2(32'hbb9fa622),
	.w3(32'hbc8d188c),
	.w4(32'hbbfe1417),
	.w5(32'h3ab4592e),
	.w6(32'hbbce37c1),
	.w7(32'hbb92dd4f),
	.w8(32'hbbc92898),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389544cf),
	.w1(32'hbc05a4fd),
	.w2(32'hb986ad49),
	.w3(32'h3bcb6151),
	.w4(32'hbc005753),
	.w5(32'h3a8d3cab),
	.w6(32'h3be7d84c),
	.w7(32'h38f49007),
	.w8(32'hbae00d14),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c84dd),
	.w1(32'hb9c56071),
	.w2(32'h3b3ff570),
	.w3(32'h3bf63d50),
	.w4(32'h3b4c0c9a),
	.w5(32'h3c332739),
	.w6(32'h3bbbcf30),
	.w7(32'h393f7aaa),
	.w8(32'h3a0e33f0),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6b70b),
	.w1(32'h3ba1feda),
	.w2(32'hbb585ddc),
	.w3(32'h3c391da5),
	.w4(32'h3b7d7ccb),
	.w5(32'hbb5d0421),
	.w6(32'h3bd4a99d),
	.w7(32'h3b81b2e8),
	.w8(32'hbbb78858),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7cd01),
	.w1(32'hbab7d670),
	.w2(32'hbc229a14),
	.w3(32'h37667ccc),
	.w4(32'hbb5dba12),
	.w5(32'hbbde6b7d),
	.w6(32'hbba45ac2),
	.w7(32'hbbd202cc),
	.w8(32'hbbf93503),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb449d0),
	.w1(32'hba38a8d0),
	.w2(32'hba907d39),
	.w3(32'h3a74ec5f),
	.w4(32'h3b85d9dc),
	.w5(32'hbbc5f98e),
	.w6(32'h3a909a64),
	.w7(32'h3b637538),
	.w8(32'hbbb6496f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a246a),
	.w1(32'hbbf6fda5),
	.w2(32'hbb12596b),
	.w3(32'hbc7d1df0),
	.w4(32'hbb7e0a64),
	.w5(32'hbb917ff8),
	.w6(32'hbbdcdb44),
	.w7(32'hbb119676),
	.w8(32'hb97fafdd),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70e68e),
	.w1(32'h3b381a9b),
	.w2(32'hbb130f02),
	.w3(32'hbbe89273),
	.w4(32'hbc2ebadd),
	.w5(32'hb9c6d911),
	.w6(32'h37338bfb),
	.w7(32'hbc47052f),
	.w8(32'hbaab5ab3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb19a50),
	.w1(32'hba86b991),
	.w2(32'hbc01ae6e),
	.w3(32'h3c110b16),
	.w4(32'h3aabeb72),
	.w5(32'hbbec5fc3),
	.w6(32'h3bc9598a),
	.w7(32'h389a56d6),
	.w8(32'hbb87271b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd0f5b),
	.w1(32'h3a20e9f8),
	.w2(32'hba808e91),
	.w3(32'hbb8240de),
	.w4(32'h3b79913f),
	.w5(32'hbb449557),
	.w6(32'h3b089aae),
	.w7(32'h3bcdfb1b),
	.w8(32'hbb04f43c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60748a),
	.w1(32'h3b34c6f8),
	.w2(32'hbbdb4b8d),
	.w3(32'hbbc140a6),
	.w4(32'hbad650dc),
	.w5(32'hbbb56382),
	.w6(32'hbb62ba10),
	.w7(32'hbb825220),
	.w8(32'hbb0335e0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e4e04),
	.w1(32'hbc0df11c),
	.w2(32'h3bbe328e),
	.w3(32'hbc6ef69a),
	.w4(32'hbbb7098d),
	.w5(32'hbbf3955c),
	.w6(32'hbb58a334),
	.w7(32'h3b376e66),
	.w8(32'hbc84b797),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ea538),
	.w1(32'h3b8b67f4),
	.w2(32'hbbb6b6f9),
	.w3(32'hbb2ed3dc),
	.w4(32'hba9cf111),
	.w5(32'hba893544),
	.w6(32'hbc337b78),
	.w7(32'hbc3b0bf8),
	.w8(32'hbb14d9c4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61f6f1),
	.w1(32'hba837e65),
	.w2(32'h3c33a29a),
	.w3(32'h3c06cae4),
	.w4(32'h3b0feb4d),
	.w5(32'h3c2fedda),
	.w6(32'h3be66e97),
	.w7(32'h3af06442),
	.w8(32'h3c2b49ed),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bf01f),
	.w1(32'h3bbded4e),
	.w2(32'h3c2dc3ed),
	.w3(32'h3bd3c2eb),
	.w4(32'h3c2cfe3a),
	.w5(32'h394e3c26),
	.w6(32'h3ba07eb7),
	.w7(32'h3c193754),
	.w8(32'hba8f9a2a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c8212),
	.w1(32'h3bbbbc15),
	.w2(32'h3bc8b765),
	.w3(32'hbbbdacce),
	.w4(32'hbc0b2a5e),
	.w5(32'hbc43d52c),
	.w6(32'hba8cf972),
	.w7(32'hbb67f59b),
	.w8(32'hbb79d3e4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12e436),
	.w1(32'hbbc9708b),
	.w2(32'hbc687a2c),
	.w3(32'hbc79ff6c),
	.w4(32'hbc0fa877),
	.w5(32'hbc6a0d1d),
	.w6(32'hbc0ec955),
	.w7(32'h3b6b8c2a),
	.w8(32'hbb39e60d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca95e32),
	.w1(32'hbbe5d306),
	.w2(32'hb8800ba2),
	.w3(32'hbcb01ed7),
	.w4(32'hbca68b84),
	.w5(32'h3abd576e),
	.w6(32'hbc4ee8ca),
	.w7(32'hbc882b49),
	.w8(32'h3aa8c71f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e5955),
	.w1(32'hba035b55),
	.w2(32'hb82cede4),
	.w3(32'h3c6eb84b),
	.w4(32'h3a914364),
	.w5(32'hba411bca),
	.w6(32'h3c24fed6),
	.w7(32'h3b44de44),
	.w8(32'hbb6a2584),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c9cc5),
	.w1(32'h3a08ddba),
	.w2(32'hbb4259cc),
	.w3(32'hbb665585),
	.w4(32'hbb69d0e8),
	.w5(32'hba5177b2),
	.w6(32'hbacb7289),
	.w7(32'h39cc658b),
	.w8(32'hbaebcff6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fbdfb),
	.w1(32'hbafea884),
	.w2(32'h38863edf),
	.w3(32'h3c215c69),
	.w4(32'h3bb0561e),
	.w5(32'h3b3b3edf),
	.w6(32'h3bf297ed),
	.w7(32'h3b81c4f4),
	.w8(32'h3c37f5f2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884a008),
	.w1(32'hbacd0ed0),
	.w2(32'hbc0c11f2),
	.w3(32'h3a1e8e23),
	.w4(32'hbc17ae08),
	.w5(32'hbb893b93),
	.w6(32'h3bfaddd8),
	.w7(32'hbc50425a),
	.w8(32'h3c1c5b82),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfed7fc),
	.w1(32'hbc432205),
	.w2(32'hbbcb4ee4),
	.w3(32'hbcbd9887),
	.w4(32'hbcb4ce81),
	.w5(32'hbc3e86f8),
	.w6(32'hbc07d290),
	.w7(32'hbb654260),
	.w8(32'h3abc7ca4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc233ca0),
	.w1(32'h3a83971c),
	.w2(32'hbbdc848e),
	.w3(32'hbc40b160),
	.w4(32'hbad70417),
	.w5(32'hbc99c4a5),
	.w6(32'hba9d6b7e),
	.w7(32'hba8a13a4),
	.w8(32'hbbc4526d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc573573),
	.w1(32'h3a9128da),
	.w2(32'hbb119085),
	.w3(32'hbc8f20aa),
	.w4(32'h3b8fdc3b),
	.w5(32'hbb9cbe48),
	.w6(32'hbc246dd2),
	.w7(32'h3c14211b),
	.w8(32'hbb0b41b8),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397625cb),
	.w1(32'hbbf64edc),
	.w2(32'h3b80616f),
	.w3(32'h399fed2d),
	.w4(32'hbc2b21a2),
	.w5(32'h3b4431c6),
	.w6(32'hbb122878),
	.w7(32'hbc25b468),
	.w8(32'h3b5527b9),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc609e),
	.w1(32'h3b178366),
	.w2(32'h3c2b1c98),
	.w3(32'h3b810b91),
	.w4(32'h3b33af9d),
	.w5(32'hbad81eb3),
	.w6(32'h3b509d4d),
	.w7(32'h3b02c5e4),
	.w8(32'hbad55590),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9b6b1),
	.w1(32'hbb28ef3b),
	.w2(32'h3ae34750),
	.w3(32'hbc701d0e),
	.w4(32'hbbe64458),
	.w5(32'hbaf7e355),
	.w6(32'hbb8624b4),
	.w7(32'hbbf62a19),
	.w8(32'hbbc6e012),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11f480),
	.w1(32'hbb7e5eb4),
	.w2(32'hba758978),
	.w3(32'hbbf880f1),
	.w4(32'hbc569ac0),
	.w5(32'hb8ba2baf),
	.w6(32'hbc16c758),
	.w7(32'hbbb8c2bd),
	.w8(32'hba12e769),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc41420),
	.w1(32'h3abe2a76),
	.w2(32'hbb48d320),
	.w3(32'h3bdb52b4),
	.w4(32'h3be1b0cb),
	.w5(32'h3b3fbe52),
	.w6(32'h3c168bc5),
	.w7(32'h3baa739b),
	.w8(32'h3950cb95),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22c643),
	.w1(32'h3b4ef55b),
	.w2(32'hbaaac528),
	.w3(32'h3c99761e),
	.w4(32'h3c31ff69),
	.w5(32'h39b65792),
	.w6(32'h3c564596),
	.w7(32'h3a447a75),
	.w8(32'h39886dd8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ebdcd),
	.w1(32'hbad7bc8d),
	.w2(32'hbbac3382),
	.w3(32'hba1586fb),
	.w4(32'hba9a52c9),
	.w5(32'hbb8ef7e7),
	.w6(32'hba1f171d),
	.w7(32'hbb314f66),
	.w8(32'hba397b38),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb096558),
	.w1(32'hbb21f77a),
	.w2(32'hb9903f64),
	.w3(32'h3a7015f1),
	.w4(32'hba08253a),
	.w5(32'hbaa932b8),
	.w6(32'h3b9aed74),
	.w7(32'h3ae3a42e),
	.w8(32'hbb262c5b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af37974),
	.w1(32'hbb54c61f),
	.w2(32'h3c614a8f),
	.w3(32'hbb363495),
	.w4(32'hbbb9f5e7),
	.w5(32'hbc6f98c9),
	.w6(32'hbb19e2bd),
	.w7(32'hbc018207),
	.w8(32'hbcbd72a4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ef336),
	.w1(32'hbbb3a6cf),
	.w2(32'h3bc09304),
	.w3(32'hbcf582fe),
	.w4(32'hbcc76ac4),
	.w5(32'h3b07f5a8),
	.w6(32'hbcafa0d0),
	.w7(32'hbca8b465),
	.w8(32'h3a88b0ae),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1085fa),
	.w1(32'h3ae28ba1),
	.w2(32'hbbbf8741),
	.w3(32'h3b29e62d),
	.w4(32'h394506a4),
	.w5(32'hbbc522bf),
	.w6(32'hb9a133dd),
	.w7(32'h3a92d310),
	.w8(32'h3c388b81),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca3234),
	.w1(32'h3b354019),
	.w2(32'h3956e06e),
	.w3(32'hbc491344),
	.w4(32'hb9c0a6ec),
	.w5(32'hbc8a684c),
	.w6(32'hbb4033d6),
	.w7(32'hbb924215),
	.w8(32'hbc98c472),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a271b),
	.w1(32'hbc6b7b0d),
	.w2(32'hbbc43176),
	.w3(32'hbd05643c),
	.w4(32'hbcb43a0f),
	.w5(32'h3ba9b211),
	.w6(32'hbcb85bb4),
	.w7(32'hbc5e3260),
	.w8(32'h3a7eb010),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb612118),
	.w1(32'h3a95569b),
	.w2(32'h3a70b406),
	.w3(32'h3bb3c309),
	.w4(32'h3bc13780),
	.w5(32'hbc2eacd4),
	.w6(32'h3bd6dffb),
	.w7(32'h3bd719f2),
	.w8(32'h3be339ff),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b606d6e),
	.w1(32'h3c1e4fd1),
	.w2(32'h3bdeaa1e),
	.w3(32'hbb68424a),
	.w4(32'h3b3c7afc),
	.w5(32'hbb1e6e7d),
	.w6(32'h3bbc4420),
	.w7(32'h3be9a655),
	.w8(32'h3a90ad60),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9323d0),
	.w1(32'h3c2fc9c8),
	.w2(32'hbb2142d9),
	.w3(32'hbc165435),
	.w4(32'hbb63ffe6),
	.w5(32'hbc0e3087),
	.w6(32'hbae44977),
	.w7(32'h3b2a6367),
	.w8(32'hbbf8e8eb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92b6a4),
	.w1(32'h398f6af5),
	.w2(32'h3b31eae4),
	.w3(32'hbbb6eea6),
	.w4(32'hbbf0510b),
	.w5(32'hbb41c19b),
	.w6(32'hbb80e8ae),
	.w7(32'hbb160039),
	.w8(32'hbc1fb537),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b8441),
	.w1(32'hbba57cfe),
	.w2(32'hbc8d9941),
	.w3(32'hbc10ad12),
	.w4(32'hbbf56fe4),
	.w5(32'hbcd8ccb8),
	.w6(32'hbbaa3627),
	.w7(32'h3ad54568),
	.w8(32'hbca1d0ea),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99a016),
	.w1(32'hbbb263be),
	.w2(32'hbae7a0ef),
	.w3(32'hbd137356),
	.w4(32'hbc3930fe),
	.w5(32'hbbd541ff),
	.w6(32'hbcd8191e),
	.w7(32'hb9c28bfa),
	.w8(32'hbbe33125),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c833),
	.w1(32'hba480afe),
	.w2(32'hbbad4278),
	.w3(32'hbbcca27e),
	.w4(32'hbb88fdd9),
	.w5(32'hbc21f622),
	.w6(32'hbb1468ea),
	.w7(32'hbb9a572d),
	.w8(32'hbc134446),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb688346),
	.w1(32'hbb04c9b7),
	.w2(32'hbc12ad35),
	.w3(32'hbbe259f1),
	.w4(32'hbbc3da2e),
	.w5(32'h3b015f48),
	.w6(32'hbbe0dd0b),
	.w7(32'hbbae02f4),
	.w8(32'hbb205877),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56e13),
	.w1(32'h3a54bfa4),
	.w2(32'hbc3bd9ae),
	.w3(32'hbab0d8d9),
	.w4(32'hbb7e37be),
	.w5(32'hbc8589dc),
	.w6(32'hbb6b9260),
	.w7(32'hbb798b24),
	.w8(32'hbb27d3ea),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55c358),
	.w1(32'h3be8f0b5),
	.w2(32'hbc686a61),
	.w3(32'hbc381f4e),
	.w4(32'h3b0c3730),
	.w5(32'hbc81303f),
	.w6(32'hbbf17117),
	.w7(32'h3baaa942),
	.w8(32'h3a9aec6a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc875f4e),
	.w1(32'hbbc2d465),
	.w2(32'hbb53516e),
	.w3(32'hbc97448f),
	.w4(32'hbbf1ef50),
	.w5(32'hbbeb4eb1),
	.w6(32'hbb36ac9f),
	.w7(32'hbac2220f),
	.w8(32'hb890bd17),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39304e),
	.w1(32'h3b98bd6d),
	.w2(32'hbc682a47),
	.w3(32'hbb4d0408),
	.w4(32'hba57dc67),
	.w5(32'hbc940b61),
	.w6(32'h3b68e112),
	.w7(32'h3b189a31),
	.w8(32'hbc92707f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09907c),
	.w1(32'hbb896a76),
	.w2(32'h3c70c507),
	.w3(32'hbc854fe9),
	.w4(32'hbc2d83d3),
	.w5(32'h3c48cafd),
	.w6(32'hbc8183e0),
	.w7(32'hbaa83993),
	.w8(32'h3a9f1811),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04dedb),
	.w1(32'h3abb283d),
	.w2(32'hbc5ea25b),
	.w3(32'hbbf17e1a),
	.w4(32'hbc4e5896),
	.w5(32'hbce6f1d6),
	.w6(32'hbc7be352),
	.w7(32'hbc33ae74),
	.w8(32'hbbd83eab),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13c00b),
	.w1(32'hbbabdb3d),
	.w2(32'h3c4760b5),
	.w3(32'hbcc99abc),
	.w4(32'hbc46a7bb),
	.w5(32'h3bcb9a16),
	.w6(32'hbc4c0e08),
	.w7(32'hbc0e0e35),
	.w8(32'hbb55a578),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06b183),
	.w1(32'h382723a0),
	.w2(32'h39bf4c0d),
	.w3(32'hba33a1bf),
	.w4(32'hbc2739be),
	.w5(32'h3bc6c485),
	.w6(32'hbc5d1b89),
	.w7(32'hbc54f6e9),
	.w8(32'h3adf739e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d1bca),
	.w1(32'h3b971b8f),
	.w2(32'hbae4a470),
	.w3(32'h3c2d2ef4),
	.w4(32'h3c10597b),
	.w5(32'hba414e0c),
	.w6(32'h3b5b40f8),
	.w7(32'h3aada677),
	.w8(32'h3bcdf051),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa0541),
	.w1(32'h3bf8b78c),
	.w2(32'h3a8ec3ad),
	.w3(32'h3a942c75),
	.w4(32'h3b98e15e),
	.w5(32'h3b8f267b),
	.w6(32'h3c0a1a69),
	.w7(32'h3b86a75a),
	.w8(32'h385afdb7),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae30963),
	.w1(32'hba8114e0),
	.w2(32'hbbdd5020),
	.w3(32'h3b87bf2d),
	.w4(32'h3b165b99),
	.w5(32'hbcc13bf0),
	.w6(32'hbaa8e28f),
	.w7(32'hbaa6d5d7),
	.w8(32'hbbe5d21d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eb307),
	.w1(32'hbbd03893),
	.w2(32'h3bc4c41a),
	.w3(32'hbcf82d10),
	.w4(32'hbc5ed897),
	.w5(32'hbb751163),
	.w6(32'hbc25b859),
	.w7(32'hba4f109e),
	.w8(32'h3b166c68),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be78d1b),
	.w1(32'h3c16b781),
	.w2(32'h3a66285f),
	.w3(32'h3a1355f8),
	.w4(32'h3bed66f9),
	.w5(32'h3bb59939),
	.w6(32'h3c0c9ac7),
	.w7(32'h3b83d66a),
	.w8(32'h3b01b0b6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24a890),
	.w1(32'hbbc98e75),
	.w2(32'hb92b6c04),
	.w3(32'h3bf06ec7),
	.w4(32'hb959444e),
	.w5(32'h3b2ac072),
	.w6(32'h3ba29458),
	.w7(32'h3c102cf2),
	.w8(32'h3b445539),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f6e4e),
	.w1(32'h3adc7440),
	.w2(32'h3bdacf84),
	.w3(32'h3b922bcb),
	.w4(32'h3b128f8e),
	.w5(32'h3bc3295a),
	.w6(32'h3b471550),
	.w7(32'h3b034285),
	.w8(32'h3be746ce),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e746),
	.w1(32'h3b24c9ed),
	.w2(32'h3ae66f26),
	.w3(32'h3b71e184),
	.w4(32'h3b9eb595),
	.w5(32'h3c0f3ba2),
	.w6(32'h3b9887dc),
	.w7(32'h3baf97f0),
	.w8(32'h3bcbf51b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f80d3),
	.w1(32'hbcecd084),
	.w2(32'hbb4b925e),
	.w3(32'hbc8b2cdd),
	.w4(32'hbd129001),
	.w5(32'hbb195f9f),
	.w6(32'hbc5555f0),
	.w7(32'hbcd44cbc),
	.w8(32'hbb9d5e91),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7e87c),
	.w1(32'hbab63732),
	.w2(32'hbbd7e265),
	.w3(32'h3a5dc868),
	.w4(32'h39bb9df2),
	.w5(32'hbcaf8a80),
	.w6(32'hba69c406),
	.w7(32'hba58390f),
	.w8(32'hbc3e3d8b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46b188),
	.w1(32'hbc3640a4),
	.w2(32'hbb91daeb),
	.w3(32'hbcf2919a),
	.w4(32'hbc3c382d),
	.w5(32'hbc51c0a4),
	.w6(32'hbca6b253),
	.w7(32'h3b6282db),
	.w8(32'hbaf43e7c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88d76c),
	.w1(32'hbb026eb7),
	.w2(32'hbbc8271c),
	.w3(32'hbce4d38b),
	.w4(32'hbc4c6f24),
	.w5(32'hbb218965),
	.w6(32'hbc22dbbf),
	.w7(32'h39a71ee1),
	.w8(32'h3acbebca),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58999d),
	.w1(32'hbb4038d8),
	.w2(32'hbbdfd0dd),
	.w3(32'hbc8c2088),
	.w4(32'hbb64b54e),
	.w5(32'hbc65e8fc),
	.w6(32'hbc745b53),
	.w7(32'hba930ff5),
	.w8(32'hbc2d3cb5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule