module layer_10_featuremap_189(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ce1a0f),
	.w1(32'hb754277c),
	.w2(32'hb6ac3db4),
	.w3(32'hb5dd3326),
	.w4(32'hb7840bc0),
	.w5(32'h3612c68f),
	.w6(32'hb702129e),
	.w7(32'hb784c4f6),
	.w8(32'hb7142ed9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae34d5d),
	.w1(32'hbb0f6a23),
	.w2(32'hbb04d35b),
	.w3(32'hbaee80b9),
	.w4(32'hba64e80e),
	.w5(32'hba01b773),
	.w6(32'hbaa6bea3),
	.w7(32'hb95064c5),
	.w8(32'hb9f6bec0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6995e65),
	.w1(32'hb6a7b660),
	.w2(32'hb69aff2b),
	.w3(32'hb658d4bb),
	.w4(32'hb65109cc),
	.w5(32'hb68215d5),
	.w6(32'hb6fa766f),
	.w7(32'hb675611f),
	.w8(32'hb6e645a8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cc9ae0),
	.w1(32'h39271304),
	.w2(32'h39b77808),
	.w3(32'hb880125a),
	.w4(32'h38ac9f65),
	.w5(32'hb9035887),
	.w6(32'h3817e771),
	.w7(32'hb883c16c),
	.w8(32'hb86822da),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9295730),
	.w1(32'h371668af),
	.w2(32'h39af29f4),
	.w3(32'hb9d7c16c),
	.w4(32'hb9a7455a),
	.w5(32'h38c51b8a),
	.w6(32'hb9ef5b4c),
	.w7(32'hb9e52136),
	.w8(32'hb88ccd81),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361b9e45),
	.w1(32'h361eebe5),
	.w2(32'hb6b70b85),
	.w3(32'hb437b25e),
	.w4(32'h36a970f0),
	.w5(32'hb70c9055),
	.w6(32'hb50800e9),
	.w7(32'h3497c059),
	.w8(32'hb7619463),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a2713),
	.w1(32'hb8a18c88),
	.w2(32'h383fe604),
	.w3(32'hb90934ba),
	.w4(32'hb90aca65),
	.w5(32'h3956283d),
	.w6(32'hb91821ae),
	.w7(32'hb9188bf2),
	.w8(32'h39e50ef3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b625e8e),
	.w1(32'h3b6326c7),
	.w2(32'h3b9596b5),
	.w3(32'h3b28e5f9),
	.w4(32'h3aa77355),
	.w5(32'h39fed2e5),
	.w6(32'h3b3d3007),
	.w7(32'h3ae97b52),
	.w8(32'h3ab94c25),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393faa0b),
	.w1(32'h3a662978),
	.w2(32'h3ab1aad0),
	.w3(32'hb919baa4),
	.w4(32'h3a12222c),
	.w5(32'h3a85d213),
	.w6(32'hb9d2f005),
	.w7(32'hb9647976),
	.w8(32'h3a01ebb2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a39ee9),
	.w1(32'h3951981d),
	.w2(32'hb9dc0c6e),
	.w3(32'hba615e2c),
	.w4(32'h39768d8b),
	.w5(32'h3a2fd8a0),
	.w6(32'h3a8a0935),
	.w7(32'h3a87da9a),
	.w8(32'h3a8f31ec),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eb368),
	.w1(32'h387d8111),
	.w2(32'h3a89f08b),
	.w3(32'h397f5871),
	.w4(32'h39285679),
	.w5(32'h3a5d5791),
	.w6(32'h398eb2d2),
	.w7(32'h35c69005),
	.w8(32'h3a463fdb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba007b63),
	.w1(32'hb8e9b60b),
	.w2(32'h39c53133),
	.w3(32'h3820e4a6),
	.w4(32'hb9be2dcd),
	.w5(32'hb8907362),
	.w6(32'h359088d3),
	.w7(32'hb5dc5d2d),
	.w8(32'h38f7c663),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c00b1d),
	.w1(32'h3a6db01b),
	.w2(32'h3b016c6f),
	.w3(32'hba464380),
	.w4(32'h3a0e8563),
	.w5(32'h3aff6662),
	.w6(32'h38c817a8),
	.w7(32'h3a232b31),
	.w8(32'h3aa207e6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b91ce6),
	.w1(32'h3a349f0b),
	.w2(32'h3a6d7100),
	.w3(32'h39fff6b8),
	.w4(32'h3a33ccf6),
	.w5(32'h3a2b235d),
	.w6(32'h3a69a4eb),
	.w7(32'h3a1762a9),
	.w8(32'h39897fe8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa18008),
	.w1(32'hba87e950),
	.w2(32'h39ce0b4e),
	.w3(32'hbadee226),
	.w4(32'hb9b58f3a),
	.w5(32'h391ec652),
	.w6(32'hba7857db),
	.w7(32'hb9429334),
	.w8(32'h3988e1ec),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a7fde),
	.w1(32'h3a2a763f),
	.w2(32'h3aaee05a),
	.w3(32'hba9c8af7),
	.w4(32'h3a0eaf7a),
	.w5(32'h38a434a7),
	.w6(32'h39d7e60a),
	.w7(32'h3a6a525c),
	.w8(32'h3ad44e26),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b287af),
	.w1(32'hb9bd56ee),
	.w2(32'hb9a592ed),
	.w3(32'hb8087846),
	.w4(32'h38a0792c),
	.w5(32'h38ce3d89),
	.w6(32'hb8e83af5),
	.w7(32'h38a5b800),
	.w8(32'h38ae2eeb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb3f5b),
	.w1(32'h3c096533),
	.w2(32'h3c1bc085),
	.w3(32'h3be83e4d),
	.w4(32'h3bb7506b),
	.w5(32'h3bad3fa7),
	.w6(32'h3bb0a860),
	.w7(32'h3b6f863a),
	.w8(32'h3b3bfadb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acaf7bd),
	.w1(32'h3b269c19),
	.w2(32'h3b15ee45),
	.w3(32'h3b0a02b7),
	.w4(32'h3af3fe35),
	.w5(32'h3acf41c5),
	.w6(32'h3af81288),
	.w7(32'h3a995d46),
	.w8(32'h3a45b113),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7259ff2),
	.w1(32'hb76ea1fa),
	.w2(32'hb7f3fa34),
	.w3(32'hb705ab30),
	.w4(32'hb6532d70),
	.w5(32'hb70b4af0),
	.w6(32'hb740737c),
	.w7(32'hb710b7ea),
	.w8(32'hb78c176a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f1c9aa),
	.w1(32'h365bda11),
	.w2(32'hb7eef49d),
	.w3(32'h36aa1478),
	.w4(32'h36e9a94b),
	.w5(32'hb7d9a73c),
	.w6(32'hb69b3aaf),
	.w7(32'hb6c5e306),
	.w8(32'hb7f02c44),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad154e8),
	.w1(32'hbaa7e785),
	.w2(32'hba891a25),
	.w3(32'hbac9dc05),
	.w4(32'hba8ca672),
	.w5(32'hba607df2),
	.w6(32'hba98d49e),
	.w7(32'hba15dde0),
	.w8(32'hba158475),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4d41c),
	.w1(32'h3c20401a),
	.w2(32'h3bdad78d),
	.w3(32'h3bdde998),
	.w4(32'h3b21d833),
	.w5(32'h3bcc5779),
	.w6(32'h3bed7ff8),
	.w7(32'h3b1f6b1b),
	.w8(32'h3b8d7c87),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9939e23),
	.w1(32'hba3a4d89),
	.w2(32'hba98bc60),
	.w3(32'hbb11996d),
	.w4(32'hba9b2998),
	.w5(32'hba200174),
	.w6(32'hb9ac016f),
	.w7(32'h3a07b227),
	.w8(32'h3a46aed1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8145af),
	.w1(32'hbabfaf63),
	.w2(32'hbb060290),
	.w3(32'hbb5bc7cc),
	.w4(32'hbafb07a1),
	.w5(32'hbac4b557),
	.w6(32'hba90275c),
	.w7(32'h3a5fd1c8),
	.w8(32'h3a7dde5d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad9bbb),
	.w1(32'hb874c8a1),
	.w2(32'hb8c25174),
	.w3(32'hb954595b),
	.w4(32'hb894549e),
	.w5(32'h38c8110c),
	.w6(32'h386865aa),
	.w7(32'hb8a41a3a),
	.w8(32'hb885af7b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82fe4ce),
	.w1(32'hb83a59f0),
	.w2(32'hb8abf99c),
	.w3(32'hb81f2165),
	.w4(32'hb7f5a0f1),
	.w5(32'hb85b94c8),
	.w6(32'hb8477a7b),
	.w7(32'hb73521c1),
	.w8(32'hb81c6895),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0161d2),
	.w1(32'hba9c8a5d),
	.w2(32'hba0daa5e),
	.w3(32'hbb0e463d),
	.w4(32'hba516212),
	.w5(32'h39a669cb),
	.w6(32'hbafd3e16),
	.w7(32'hba21a20c),
	.w8(32'h390b28dd),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf7d5a),
	.w1(32'hb990300b),
	.w2(32'h37f67279),
	.w3(32'hba01facd),
	.w4(32'hba20e023),
	.w5(32'hba313154),
	.w6(32'hb98038b6),
	.w7(32'hb715fda3),
	.w8(32'hb982e4f6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6bca9),
	.w1(32'hbab9b85c),
	.w2(32'hbaa2f198),
	.w3(32'hbb3d35f8),
	.w4(32'hbaac9d85),
	.w5(32'hba44148a),
	.w6(32'hbac3856a),
	.w7(32'hb9e1a939),
	.w8(32'hb9e66e2f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d10116),
	.w1(32'hb79d1655),
	.w2(32'hb7f251f4),
	.w3(32'hb77e2805),
	.w4(32'hb722a7cd),
	.w5(32'hb7b18a19),
	.w6(32'hb7efa41b),
	.w7(32'hb774778f),
	.w8(32'hb7b65740),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7870d7c),
	.w1(32'hb77a6d86),
	.w2(32'hb88bc5b5),
	.w3(32'h361497f7),
	.w4(32'hb76e5f6f),
	.w5(32'hb8a02a50),
	.w6(32'hb6e6c7e7),
	.w7(32'hb8209e3f),
	.w8(32'hb8cf4288),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93264cd),
	.w1(32'hb7ff879e),
	.w2(32'h37d8a1ca),
	.w3(32'hb9ea7b13),
	.w4(32'hba06b540),
	.w5(32'hb9aad5a3),
	.w6(32'h39137ad4),
	.w7(32'hb94b2c27),
	.w8(32'hb91875e4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39788b62),
	.w1(32'hb9fd3027),
	.w2(32'hba4cab45),
	.w3(32'hb999bf0e),
	.w4(32'hb9848c8e),
	.w5(32'hb9ccc53f),
	.w6(32'h38cc4995),
	.w7(32'h38bcaa88),
	.w8(32'h378d8a3e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83fd916),
	.w1(32'hb71589aa),
	.w2(32'hb70bd37a),
	.w3(32'hb6cfeff2),
	.w4(32'hb75b9218),
	.w5(32'hb68f93de),
	.w6(32'h38d621ea),
	.w7(32'h391b3a13),
	.w8(32'h39048a1b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2ea28),
	.w1(32'h391968ee),
	.w2(32'h39307710),
	.w3(32'h3988f40a),
	.w4(32'hb8848f77),
	.w5(32'hb927d77e),
	.w6(32'h39fdd0a4),
	.w7(32'h383504c4),
	.w8(32'h38cd9821),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b005ebf),
	.w1(32'h3b25fbf8),
	.w2(32'h3af4110d),
	.w3(32'h3b19c981),
	.w4(32'h3aa07f2c),
	.w5(32'h3a08a42f),
	.w6(32'h3b407f9c),
	.w7(32'hb9d7f1e3),
	.w8(32'h3985382f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f0935),
	.w1(32'hbbc717d8),
	.w2(32'hbbab7e43),
	.w3(32'hbbe2fae3),
	.w4(32'hbb92ca68),
	.w5(32'hbb30b24f),
	.w6(32'hbb8107fd),
	.w7(32'hba9fc938),
	.w8(32'hbacc72c4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac41d9),
	.w1(32'hbba6e55f),
	.w2(32'hbb73a72f),
	.w3(32'hbbd6cea3),
	.w4(32'hbb2f1036),
	.w5(32'hb9ddd94b),
	.w6(32'hbbbbc394),
	.w7(32'hba49600c),
	.w8(32'h3996a1af),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f894b),
	.w1(32'hba840a45),
	.w2(32'hba55a2f1),
	.w3(32'hbac16a55),
	.w4(32'hb9a94fec),
	.w5(32'hb9da64c6),
	.w6(32'hba7014c2),
	.w7(32'hb94425f3),
	.w8(32'hb957e51f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38802c06),
	.w1(32'h3874dc8a),
	.w2(32'h37c7a230),
	.w3(32'h38a3bfa7),
	.w4(32'h389e17d6),
	.w5(32'h37f06476),
	.w6(32'h38b7a871),
	.w7(32'h381c2372),
	.w8(32'hb876da34),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81446d7),
	.w1(32'hb8a36780),
	.w2(32'hb92a6081),
	.w3(32'hb8b3e362),
	.w4(32'hb8bd3d70),
	.w5(32'hb8fa1771),
	.w6(32'hb91f9c54),
	.w7(32'hb8d6a1ad),
	.w8(32'hb8ff4e3b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39097bc5),
	.w1(32'hb8aa1c6d),
	.w2(32'h36d89dc0),
	.w3(32'h36dd39ee),
	.w4(32'hb99a9e26),
	.w5(32'h3888ddac),
	.w6(32'h391d5d5e),
	.w7(32'hb8fc494d),
	.w8(32'h3914556e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5f5db),
	.w1(32'h3abe8f26),
	.w2(32'h3a7ef2b9),
	.w3(32'h3a20180a),
	.w4(32'h39e5c7b1),
	.w5(32'h38b783eb),
	.w6(32'h3b02199d),
	.w7(32'h3a8c4451),
	.w8(32'h3a0049ca),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d52a17),
	.w1(32'hb9a79a00),
	.w2(32'hb923cc94),
	.w3(32'hbafe221d),
	.w4(32'hba9434f3),
	.w5(32'hb990737a),
	.w6(32'hba3f5018),
	.w7(32'hb90e91d9),
	.w8(32'h38fabbfb),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b405b8),
	.w1(32'hba1e34cb),
	.w2(32'hba9e003d),
	.w3(32'hbb13c470),
	.w4(32'hba47bb52),
	.w5(32'hba3c999c),
	.w6(32'hb9357c0c),
	.w7(32'h3a10a6b6),
	.w8(32'h39e7df60),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ba86e),
	.w1(32'h3ab1801a),
	.w2(32'h3a48628f),
	.w3(32'hb93692fa),
	.w4(32'h39c7c8bc),
	.w5(32'hba7a91a3),
	.w6(32'h3b221301),
	.w7(32'h3a870b31),
	.w8(32'h39585ed2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd72fca),
	.w1(32'h3c21b1ab),
	.w2(32'h3c2a5915),
	.w3(32'h3bfa203d),
	.w4(32'h3bde12f9),
	.w5(32'h3bd4cdd0),
	.w6(32'h3bcca63e),
	.w7(32'h3b553704),
	.w8(32'h3b4765dc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84b546a),
	.w1(32'h38930e03),
	.w2(32'hb64c6f25),
	.w3(32'hb69aa51b),
	.w4(32'hb6b6da5f),
	.w5(32'hb8f8bb48),
	.w6(32'hb7006463),
	.w7(32'hb8b51d42),
	.w8(32'hb981dfe2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a588a13),
	.w1(32'h3a0c5ac8),
	.w2(32'h39f97b84),
	.w3(32'h3a365cac),
	.w4(32'h3a00cfc5),
	.w5(32'h3a5e29f0),
	.w6(32'h39aed421),
	.w7(32'h39b62a38),
	.w8(32'h3a617208),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60ae96e),
	.w1(32'hb841510d),
	.w2(32'hb8581e84),
	.w3(32'hb912d586),
	.w4(32'hb95756db),
	.w5(32'hb7a1ce9d),
	.w6(32'hb942f1cd),
	.w7(32'hb9995717),
	.w8(32'hb8e40e2e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c276b3),
	.w1(32'hb919c47a),
	.w2(32'hb8fb737c),
	.w3(32'hba0f22a3),
	.w4(32'hb9f65665),
	.w5(32'h38039d74),
	.w6(32'hb7b748c4),
	.w7(32'h39c9f8e6),
	.w8(32'h3a1c034f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bb7a0),
	.w1(32'h3a7aefb1),
	.w2(32'h3a8fc111),
	.w3(32'h3a48721e),
	.w4(32'h39ba9822),
	.w5(32'h394876af),
	.w6(32'h3a7270ef),
	.w7(32'h397a4305),
	.w8(32'h39a8d1e6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840d62),
	.w1(32'h3bad214c),
	.w2(32'h3b974ab3),
	.w3(32'h3ba677d0),
	.w4(32'h3b3e9a19),
	.w5(32'h3af53676),
	.w6(32'h3b63b4f4),
	.w7(32'h39a01e36),
	.w8(32'h3a9ab420),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e9651),
	.w1(32'h3a1bb1d3),
	.w2(32'h3a8df2fb),
	.w3(32'h39395761),
	.w4(32'hb712187a),
	.w5(32'h39b4aa66),
	.w6(32'h393dcf90),
	.w7(32'h391f656d),
	.w8(32'h39e235c6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f7bf59),
	.w1(32'h373d02a3),
	.w2(32'h3819576f),
	.w3(32'hb791b9f5),
	.w4(32'h3786df67),
	.w5(32'h383598cf),
	.w6(32'hb728980b),
	.w7(32'h3706ad7b),
	.w8(32'h376ded97),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77081c2),
	.w1(32'hb77db736),
	.w2(32'hb7934638),
	.w3(32'hb7934feb),
	.w4(32'hb76bb455),
	.w5(32'hb7667a7b),
	.w6(32'hb7b8cd71),
	.w7(32'hb751822c),
	.w8(32'hb78c5d7b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6924f4b),
	.w1(32'hb54e750c),
	.w2(32'hb7f6d1a3),
	.w3(32'hb8762355),
	.w4(32'hb858728f),
	.w5(32'h37d7c94b),
	.w6(32'hb8afbafb),
	.w7(32'hb80bc7e7),
	.w8(32'hb53bfebb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b9675),
	.w1(32'hb8ba3eb2),
	.w2(32'h36c4616f),
	.w3(32'hb99a56b2),
	.w4(32'hb96a2a8c),
	.w5(32'h3839f719),
	.w6(32'hb93ad031),
	.w7(32'hb8f6f3aa),
	.w8(32'h38c5fc3d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980681e),
	.w1(32'h37047a27),
	.w2(32'h39835309),
	.w3(32'hb98ecb89),
	.w4(32'h382fa5e3),
	.w5(32'h38dcb083),
	.w6(32'hb98c81e0),
	.w7(32'h38f3a28c),
	.w8(32'h394d8e1b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af81a12),
	.w1(32'h3b1f385c),
	.w2(32'h3b15193e),
	.w3(32'h3ae1a53c),
	.w4(32'h3ab49228),
	.w5(32'h3a9a7c92),
	.w6(32'h3aa6b120),
	.w7(32'h3a86dfb3),
	.w8(32'h3aa5c033),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b155aff),
	.w1(32'h3b1d0afe),
	.w2(32'h3ab1ac40),
	.w3(32'h3b21d3a7),
	.w4(32'h3a58dc1d),
	.w5(32'h3b21ff4c),
	.w6(32'h3ab683cd),
	.w7(32'h3a91bdd9),
	.w8(32'h3acb979d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bac771),
	.w1(32'hb6258a32),
	.w2(32'hb8184001),
	.w3(32'h38146b46),
	.w4(32'hb7e57f12),
	.w5(32'hb86ce9e7),
	.w6(32'h3823c402),
	.w7(32'hb8291138),
	.w8(32'hb89ea025),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ce376d),
	.w1(32'h359e9a1f),
	.w2(32'hb732986e),
	.w3(32'h36db9509),
	.w4(32'h36e238a5),
	.w5(32'hb6590f25),
	.w6(32'h363afeda),
	.w7(32'h34e43048),
	.w8(32'hb768bb28),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91049d7),
	.w1(32'hb8c16209),
	.w2(32'hb8382639),
	.w3(32'hb8ef17cc),
	.w4(32'hb8667ec3),
	.w5(32'hb7aba2e6),
	.w6(32'hb8c2b041),
	.w7(32'hb89303be),
	.w8(32'hb8c367fe),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d71dfd),
	.w1(32'h366dff6d),
	.w2(32'hb7c86cce),
	.w3(32'hb6c92b3e),
	.w4(32'hb62c6c27),
	.w5(32'hb808746a),
	.w6(32'hb7fa67e0),
	.w7(32'hb7898516),
	.w8(32'hb85a71ca),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08ef05),
	.w1(32'h3a55f92b),
	.w2(32'h3a2ff968),
	.w3(32'h39a0a301),
	.w4(32'h384eb878),
	.w5(32'h370b83ba),
	.w6(32'h3a483622),
	.w7(32'h3a15f2f4),
	.w8(32'h3a035b11),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4680c8),
	.w1(32'hba0098be),
	.w2(32'h3a0e0558),
	.w3(32'hbb1e8b5c),
	.w4(32'hba83c7e1),
	.w5(32'hba4cafb2),
	.w6(32'h3882401b),
	.w7(32'h3a6ba350),
	.w8(32'h3ada3e7e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7314dc),
	.w1(32'h3b3af0f4),
	.w2(32'h3b695d7a),
	.w3(32'h3ae71bad),
	.w4(32'hb8bc5561),
	.w5(32'h3b2d7dfa),
	.w6(32'h3b31ac4d),
	.w7(32'h3af41f69),
	.w8(32'h3b35bfa7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c1f81),
	.w1(32'hbb0bd28d),
	.w2(32'hbb3d8352),
	.w3(32'hbb8b7a47),
	.w4(32'hbb09a6cd),
	.w5(32'hba49ecc8),
	.w6(32'hbac5b176),
	.w7(32'h39ca10b8),
	.w8(32'h39cd5a49),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb695d0dd),
	.w1(32'hb5519a34),
	.w2(32'hb78d042d),
	.w3(32'h36abc4ce),
	.w4(32'h3769fbe2),
	.w5(32'hb7056827),
	.w6(32'h36301a18),
	.w7(32'hb6e59f10),
	.w8(32'hb7e020bb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6db42b8),
	.w1(32'hb7ab8943),
	.w2(32'hb891944d),
	.w3(32'h369af96b),
	.w4(32'h35953c65),
	.w5(32'hb7f678e9),
	.w6(32'hb7c29009),
	.w7(32'hb7d235a4),
	.w8(32'hb87c2dbc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c35e93),
	.w1(32'h37b3729f),
	.w2(32'hb81d2f64),
	.w3(32'hb5475b6c),
	.w4(32'h3735388b),
	.w5(32'hb8036855),
	.w6(32'hb855e68b),
	.w7(32'hb76af180),
	.w8(32'hb8808940),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5c281),
	.w1(32'h3a8685e8),
	.w2(32'h3a9d526b),
	.w3(32'h39e79824),
	.w4(32'h3a462fc9),
	.w5(32'h3a318eac),
	.w6(32'h3a1d98ee),
	.w7(32'h3a274c05),
	.w8(32'h3a161210),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bf2808),
	.w1(32'h36e057f8),
	.w2(32'hb7aa5304),
	.w3(32'hb7280f5f),
	.w4(32'hb727094c),
	.w5(32'hb83a21f5),
	.w6(32'hb7bb6fa2),
	.w7(32'hb807d021),
	.w8(32'hb87db9e3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab80393),
	.w1(32'h3b801fb4),
	.w2(32'h3b4b911b),
	.w3(32'h3b5fbca4),
	.w4(32'h3b4b7ac6),
	.w5(32'h3a82e30f),
	.w6(32'h3b5dd955),
	.w7(32'h3a54efa2),
	.w8(32'h39b11bbd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0db55d),
	.w1(32'h3b8c6712),
	.w2(32'h3bd842ba),
	.w3(32'h3b6497cd),
	.w4(32'h3b9fb0b1),
	.w5(32'h3a833074),
	.w6(32'h3be80f9a),
	.w7(32'h3b8ebca5),
	.w8(32'h3b6a281a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8286b6),
	.w1(32'hba903c26),
	.w2(32'hb90ffa2e),
	.w3(32'hbb197cd5),
	.w4(32'hba4e6e53),
	.w5(32'h3a2b028e),
	.w6(32'hbaba2071),
	.w7(32'h38201132),
	.w8(32'h39ee9867),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe4993),
	.w1(32'h3ab8a66f),
	.w2(32'h3ad29506),
	.w3(32'h3a91d508),
	.w4(32'h3a567013),
	.w5(32'h3a7ecdce),
	.w6(32'h3b02a334),
	.w7(32'h3aa3205a),
	.w8(32'h3aab601f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96daa6d),
	.w1(32'h39590b67),
	.w2(32'h395bdcc5),
	.w3(32'hb9b3ddb0),
	.w4(32'hb9606f6c),
	.w5(32'hb9ce1f1c),
	.w6(32'h3a1e3079),
	.w7(32'h39b31910),
	.w8(32'h3a39a1dd),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ccb75a),
	.w1(32'h391d693e),
	.w2(32'h399b2680),
	.w3(32'hb9d6dfb7),
	.w4(32'hb96de09f),
	.w5(32'h39e089db),
	.w6(32'hb8b8f664),
	.w7(32'h3932037e),
	.w8(32'h3a0a5ccd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeee10a),
	.w1(32'h3b626410),
	.w2(32'h3b339951),
	.w3(32'h3b303f12),
	.w4(32'h3b0d0ed3),
	.w5(32'h3acf631a),
	.w6(32'h3afec882),
	.w7(32'h3a898f82),
	.w8(32'h3a20d882),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3780e4ca),
	.w1(32'h377dbddf),
	.w2(32'h36439953),
	.w3(32'h36d41223),
	.w4(32'h370fb3cd),
	.w5(32'hb6f8d305),
	.w6(32'hb65a1884),
	.w7(32'hb74a61a1),
	.w8(32'hb8097d3f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85aa133),
	.w1(32'hb8107137),
	.w2(32'hb82ad03e),
	.w3(32'hb845e02a),
	.w4(32'hb8285734),
	.w5(32'hb73f671c),
	.w6(32'hb7cb5ecc),
	.w7(32'hb7f4930c),
	.w8(32'hb7cd1044),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e39f45),
	.w1(32'hb924f210),
	.w2(32'hb989f14e),
	.w3(32'hb9daf7ce),
	.w4(32'hb9396905),
	.w5(32'hb8a88958),
	.w6(32'hb9bf4799),
	.w7(32'hb8d61c4d),
	.w8(32'hb905a179),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b13417),
	.w1(32'hb7f854cd),
	.w2(32'hb6ccdf0c),
	.w3(32'hb7f2f6e8),
	.w4(32'hb7cc4c53),
	.w5(32'h3717a587),
	.w6(32'hb52da1ad),
	.w7(32'h36fde33a),
	.w8(32'h37cd3d0d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab33365),
	.w1(32'hbad87420),
	.w2(32'hbb4f39c8),
	.w3(32'hbb2dda7c),
	.w4(32'hba9aabf1),
	.w5(32'hbab7642c),
	.w6(32'hbac1fc79),
	.w7(32'hb9e86aa2),
	.w8(32'hba6a2b47),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8491917),
	.w1(32'hb88c92ef),
	.w2(32'h3650911b),
	.w3(32'hb8f0d9bf),
	.w4(32'hb909a886),
	.w5(32'hb935f9b7),
	.w6(32'h3914764a),
	.w7(32'h383d8963),
	.w8(32'hb8a2a7b3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d3253),
	.w1(32'h39a1e402),
	.w2(32'h3958705a),
	.w3(32'hba0a1f2c),
	.w4(32'h39d1a741),
	.w5(32'h3a2d13fd),
	.w6(32'h394404b6),
	.w7(32'h3a409019),
	.w8(32'h3a22b135),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb92c75),
	.w1(32'h3bbaedee),
	.w2(32'h3b880993),
	.w3(32'h3c04e842),
	.w4(32'h3b645e0a),
	.w5(32'h3aa5e6d8),
	.w6(32'h3c04ceed),
	.w7(32'h3b7793b4),
	.w8(32'h3b1fba0d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a0c7e),
	.w1(32'hba529242),
	.w2(32'h38840df5),
	.w3(32'hbae4178a),
	.w4(32'hb9b6bcf3),
	.w5(32'hb93e661f),
	.w6(32'hba7a1c27),
	.w7(32'hb7f74b48),
	.w8(32'h392d8a3a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1dc44),
	.w1(32'h3b0469b9),
	.w2(32'h3b28cb04),
	.w3(32'h3a63e908),
	.w4(32'h38cfd006),
	.w5(32'h3b4a9853),
	.w6(32'h39a701e1),
	.w7(32'hba9f1ede),
	.w8(32'h3ab1c67e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3420f),
	.w1(32'hbaeebc75),
	.w2(32'hbac9196f),
	.w3(32'hbad87019),
	.w4(32'hbaa19a81),
	.w5(32'hba1da9ee),
	.w6(32'hbacaa78a),
	.w7(32'hba9a08c5),
	.w8(32'hb9e44732),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a835af3),
	.w1(32'h3a9455fb),
	.w2(32'h3ab7a7a5),
	.w3(32'h3a4a81b7),
	.w4(32'h3a0eb914),
	.w5(32'h3a7e3b47),
	.w6(32'h3ac643d4),
	.w7(32'h3ab7b4cd),
	.w8(32'h3ad49f8e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9974f7),
	.w1(32'hba8a990f),
	.w2(32'hbacff679),
	.w3(32'hbaf97685),
	.w4(32'hbabfc784),
	.w5(32'hba7ba14c),
	.w6(32'hbabacb57),
	.w7(32'hba9659dd),
	.w8(32'hba456b39),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0acaf),
	.w1(32'hbadbc331),
	.w2(32'hba800f1a),
	.w3(32'hbb0eb306),
	.w4(32'hba57c9f2),
	.w5(32'hb9d13f23),
	.w6(32'hbabea4e6),
	.w7(32'hb98a29c2),
	.w8(32'hb9b7bc1d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951dde2),
	.w1(32'hb9cff770),
	.w2(32'hb979b7f9),
	.w3(32'hb95ec0fd),
	.w4(32'hb9eb01dd),
	.w5(32'h389807b6),
	.w6(32'hb9adaeb9),
	.w7(32'hba4d59ad),
	.w8(32'hb89e374f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a556bf3),
	.w1(32'h3a85ba85),
	.w2(32'h3adc7e4f),
	.w3(32'h3872d925),
	.w4(32'hb9a6f3c3),
	.w5(32'h3a499dbd),
	.w6(32'h3a932a39),
	.w7(32'h391c7dd3),
	.w8(32'h3a4b5fa9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9204bd4),
	.w1(32'hb96f0f2e),
	.w2(32'hba747ecb),
	.w3(32'hba341649),
	.w4(32'hba82c5bf),
	.w5(32'hb832865b),
	.w6(32'hba7040ad),
	.w7(32'hba239466),
	.w8(32'h3a1496c7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81cb43),
	.w1(32'h3c010666),
	.w2(32'h3bac401c),
	.w3(32'h3bebb6c8),
	.w4(32'h3bb51311),
	.w5(32'h3b1196b8),
	.w6(32'h3bea5dea),
	.w7(32'h3b5d1d64),
	.w8(32'h3b1996fd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60d6e5),
	.w1(32'hbb93462d),
	.w2(32'hbb11efcf),
	.w3(32'hbbb03439),
	.w4(32'hbb6f0fa5),
	.w5(32'h3b2905d9),
	.w6(32'hbba0b174),
	.w7(32'hbb8781dc),
	.w8(32'h38398fc0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba835a25),
	.w1(32'hbb0a757d),
	.w2(32'hbb0a72c9),
	.w3(32'hbb6ff1ce),
	.w4(32'hbad94e0d),
	.w5(32'hba7c671e),
	.w6(32'hbaadcf58),
	.w7(32'hb986d8f9),
	.w8(32'hba2574ed),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b052526),
	.w1(32'h3b46bdda),
	.w2(32'h3b7b82d0),
	.w3(32'h3a9bc3a7),
	.w4(32'h3a25c1bb),
	.w5(32'h3b5664a3),
	.w6(32'h3aa51bf8),
	.w7(32'hbaaa84f5),
	.w8(32'h3a964734),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d40de),
	.w1(32'hba02cb7c),
	.w2(32'hba4bd70e),
	.w3(32'h38a39e59),
	.w4(32'hba412930),
	.w5(32'hba5ee7fb),
	.w6(32'h3819eec9),
	.w7(32'hba382718),
	.w8(32'hba8ac66a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ea4e),
	.w1(32'h3c257c0d),
	.w2(32'h3c139a59),
	.w3(32'h3be3af29),
	.w4(32'h3c0dd8c6),
	.w5(32'h3b9d8ff2),
	.w6(32'h3c18babf),
	.w7(32'h3b8a2bc8),
	.w8(32'h3b5fbfc8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab8b13),
	.w1(32'hb8f637a4),
	.w2(32'h39b6bb55),
	.w3(32'hba935689),
	.w4(32'h3a91994e),
	.w5(32'h3a7ae8b3),
	.w6(32'hba4d2695),
	.w7(32'h39ce8a57),
	.w8(32'h3a1f0d22),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9558568),
	.w1(32'hb8f9f325),
	.w2(32'hb891d1a0),
	.w3(32'hb8cbf49d),
	.w4(32'h37e891a9),
	.w5(32'h392e508a),
	.w6(32'hb955cb84),
	.w7(32'hb5811b0c),
	.w8(32'h3817eb5c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397fa89b),
	.w1(32'h39663967),
	.w2(32'hba116eb1),
	.w3(32'h398c5f85),
	.w4(32'hb6ef2366),
	.w5(32'h39ad135f),
	.w6(32'h3985ccf3),
	.w7(32'h3959117f),
	.w8(32'hb95600a2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d1801),
	.w1(32'hb8fdcee6),
	.w2(32'h39de7c60),
	.w3(32'hbaadaf3f),
	.w4(32'hb926e27d),
	.w5(32'h399aee7e),
	.w6(32'h37836c4b),
	.w7(32'h3a103ce2),
	.w8(32'h398b8d8a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e82a4),
	.w1(32'hba698a58),
	.w2(32'hba869d1f),
	.w3(32'hbb411112),
	.w4(32'hbac77c07),
	.w5(32'hba44b887),
	.w6(32'hba892b82),
	.w7(32'hb9d3fa73),
	.w8(32'hb99402d2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c31e5),
	.w1(32'hba04ccd8),
	.w2(32'h3abd055f),
	.w3(32'hbae5b843),
	.w4(32'hba474c9a),
	.w5(32'h3a979905),
	.w6(32'hba158226),
	.w7(32'hb84e2e27),
	.w8(32'h39dd04a3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2a49b),
	.w1(32'h39088c91),
	.w2(32'h37667cc0),
	.w3(32'hb8cc24e5),
	.w4(32'h3964cdc6),
	.w5(32'h3a6b4433),
	.w6(32'h3990b4c8),
	.w7(32'h39f6f57b),
	.w8(32'h39f2367a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83b0d4),
	.w1(32'h3a383772),
	.w2(32'h3a7b2478),
	.w3(32'h39c2aefa),
	.w4(32'h38275914),
	.w5(32'hb9ffd230),
	.w6(32'h3a3d2fd1),
	.w7(32'h39dedfe0),
	.w8(32'h3a1738df),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab478f3),
	.w1(32'h3ae83f73),
	.w2(32'h3a7bb93e),
	.w3(32'h3aa37ee4),
	.w4(32'h3aa53ac9),
	.w5(32'h3a9b9034),
	.w6(32'h3ab016a1),
	.w7(32'h3a60d689),
	.w8(32'h3a840597),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80158e4),
	.w1(32'h380307a3),
	.w2(32'hb7cac838),
	.w3(32'hba890e18),
	.w4(32'hb9a4070c),
	.w5(32'h38de4205),
	.w6(32'hba4265a6),
	.w7(32'h39762b6d),
	.w8(32'h3a2158cd),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8e841),
	.w1(32'h383d09da),
	.w2(32'h3852cc0c),
	.w3(32'h38d8c238),
	.w4(32'h387488f3),
	.w5(32'hb67d8556),
	.w6(32'h38ab91d5),
	.w7(32'h38271cbc),
	.w8(32'h3730d57f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3801e316),
	.w1(32'h37bcac5d),
	.w2(32'h3613fc62),
	.w3(32'hb6d429e8),
	.w4(32'h37266137),
	.w5(32'hb75cf7e9),
	.w6(32'hb7f4be4e),
	.w7(32'hb78cb89e),
	.w8(32'hb7c98265),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ace60c),
	.w1(32'h371ed3b6),
	.w2(32'hb72801e7),
	.w3(32'hb7f4fc83),
	.w4(32'hb7a1f92c),
	.w5(32'hb7fa15f9),
	.w6(32'hb790f4d6),
	.w7(32'hb7d9b5fb),
	.w8(32'hb807ea01),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ffe0ec),
	.w1(32'h38bee7b1),
	.w2(32'hb85c45e9),
	.w3(32'hb9a2d7cc),
	.w4(32'hb9de2036),
	.w5(32'hb9c58cd6),
	.w6(32'hb8b38e15),
	.w7(32'hb984faf2),
	.w8(32'h390fd7ad),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d1ef5),
	.w1(32'hbad1f16a),
	.w2(32'hba9cd1af),
	.w3(32'hbb1590cf),
	.w4(32'hbaaa8906),
	.w5(32'hba0063b4),
	.w6(32'hbb0059cc),
	.w7(32'hba8576c6),
	.w8(32'hb9e29323),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b79195),
	.w1(32'h399f4a1b),
	.w2(32'h3a89f12a),
	.w3(32'hb9dd6c39),
	.w4(32'hb9a4a0e8),
	.w5(32'h39e5541c),
	.w6(32'hba2323d0),
	.w7(32'hba1aa3e5),
	.w8(32'h39207a5f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa046b9),
	.w1(32'h3ae9a624),
	.w2(32'h3b095518),
	.w3(32'h3a79d374),
	.w4(32'h3a3f7624),
	.w5(32'h3a18e298),
	.w6(32'h3ac56c3a),
	.w7(32'h39ee6c6b),
	.w8(32'h3a1bddae),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0011a8),
	.w1(32'hbb44d56c),
	.w2(32'hbb391b0a),
	.w3(32'hbb37b0c6),
	.w4(32'hba7b069c),
	.w5(32'hba0097af),
	.w6(32'hbb186903),
	.w7(32'hb95381ae),
	.w8(32'hb972488e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90308c5),
	.w1(32'hb8cea69d),
	.w2(32'hb8bf2350),
	.w3(32'hb88a415f),
	.w4(32'h3614f115),
	.w5(32'h3870d148),
	.w6(32'h3717951c),
	.w7(32'h383ca5fd),
	.w8(32'h37ad54dc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dd6164),
	.w1(32'h38e5ef84),
	.w2(32'h3963e147),
	.w3(32'hb692c67c),
	.w4(32'h3861356b),
	.w5(32'h3949497a),
	.w6(32'hb801488d),
	.w7(32'h38a73346),
	.w8(32'h395fb322),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80bf133),
	.w1(32'hb76e98ae),
	.w2(32'hb7a64d4c),
	.w3(32'hb7454ee4),
	.w4(32'h3484112a),
	.w5(32'hb79f7dd7),
	.w6(32'hb7fdee38),
	.w7(32'hb73680bd),
	.w8(32'hb7b45dc2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3a3f1),
	.w1(32'hba8ae92b),
	.w2(32'hb9057868),
	.w3(32'hba6094c8),
	.w4(32'hba8a1ba8),
	.w5(32'h3a521110),
	.w6(32'hba07e872),
	.w7(32'hba8185d6),
	.w8(32'hbb1fc450),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46c44e),
	.w1(32'h3aff348f),
	.w2(32'h39c6c10d),
	.w3(32'hba8ca028),
	.w4(32'h3a1e6293),
	.w5(32'h39e21be6),
	.w6(32'h3a57321b),
	.w7(32'h3a32d9d9),
	.w8(32'h3ac8639d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00b36d),
	.w1(32'h39490276),
	.w2(32'h3bb1ba6d),
	.w3(32'h3b2318c1),
	.w4(32'hb9a66c36),
	.w5(32'h3b36b507),
	.w6(32'hba2e4d67),
	.w7(32'h3b0839a3),
	.w8(32'h3aa78fd7),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4b3ec),
	.w1(32'h3abd1f10),
	.w2(32'h3ad38a39),
	.w3(32'h3b7c8960),
	.w4(32'h3ae3e085),
	.w5(32'h3b49d1c0),
	.w6(32'h3a652965),
	.w7(32'h3ace0482),
	.w8(32'h3af1a7c4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08cc1f),
	.w1(32'h3ae47c79),
	.w2(32'h3aa0727d),
	.w3(32'h3b0800c8),
	.w4(32'h3a299923),
	.w5(32'h3a179c4d),
	.w6(32'hb9ea7a44),
	.w7(32'hba910889),
	.w8(32'hba6336ba),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce828c),
	.w1(32'h3aba5b93),
	.w2(32'hbb92e006),
	.w3(32'hba9682f1),
	.w4(32'hbae8b312),
	.w5(32'hbba866f1),
	.w6(32'hb9670927),
	.w7(32'hbbcd1cf1),
	.w8(32'hbacc50d5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5122b4),
	.w1(32'hb9d87817),
	.w2(32'hb96f3bf6),
	.w3(32'hbaeab737),
	.w4(32'hb865803a),
	.w5(32'hb93ec114),
	.w6(32'h3acaac45),
	.w7(32'h3b06fae9),
	.w8(32'h3b4a618b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97ef0c),
	.w1(32'hba91bdd7),
	.w2(32'hbb816a09),
	.w3(32'h3b048e00),
	.w4(32'hba673487),
	.w5(32'hbb1a584d),
	.w6(32'hbb0a566e),
	.w7(32'hbb75e42a),
	.w8(32'hba13febf),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87adba),
	.w1(32'h3b872bce),
	.w2(32'h3b432c28),
	.w3(32'h3bdbb6e5),
	.w4(32'h3aea951b),
	.w5(32'h3b274abf),
	.w6(32'h3ae7764b),
	.w7(32'h3a8317b5),
	.w8(32'h3b47c378),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa43f1c),
	.w1(32'hba4f993d),
	.w2(32'hb9b263c2),
	.w3(32'hba99c03c),
	.w4(32'hb8e7ae46),
	.w5(32'h3a45719d),
	.w6(32'hbb01f043),
	.w7(32'hba689204),
	.w8(32'hb99ac87b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b260844),
	.w1(32'h39290a1f),
	.w2(32'h3ac290ec),
	.w3(32'h3b251eda),
	.w4(32'h3a164265),
	.w5(32'h3b09bc3b),
	.w6(32'h3a7764f3),
	.w7(32'h3a78ca2e),
	.w8(32'h3ad9c561),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c376f),
	.w1(32'hb9fa85eb),
	.w2(32'h3b01786a),
	.w3(32'h3b84851d),
	.w4(32'hba9f4745),
	.w5(32'h3af5d403),
	.w6(32'hba26812d),
	.w7(32'hbab72ce7),
	.w8(32'h3b14d7d5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21b439),
	.w1(32'hb802d93b),
	.w2(32'hbb156034),
	.w3(32'h3a5118e6),
	.w4(32'hbaccdc63),
	.w5(32'hba914fda),
	.w6(32'hbb8b7704),
	.w7(32'hbbafd1e0),
	.w8(32'hbbac6554),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cbe4b),
	.w1(32'h37d0cad5),
	.w2(32'hbb134b42),
	.w3(32'hb956e375),
	.w4(32'hbae7c4c2),
	.w5(32'hbb28c88a),
	.w6(32'hbafb5db3),
	.w7(32'hbb970ca1),
	.w8(32'hbad4170b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a504e53),
	.w1(32'hb9908fb1),
	.w2(32'hba9ed058),
	.w3(32'h39c7dca0),
	.w4(32'hb97978ec),
	.w5(32'hb7ea1e58),
	.w6(32'hb9a4a366),
	.w7(32'hba95283a),
	.w8(32'hbab21c8d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8abfc7),
	.w1(32'hbb872357),
	.w2(32'hba9cc25d),
	.w3(32'hbb93c514),
	.w4(32'hbb32a4b4),
	.w5(32'h3acc858a),
	.w6(32'hbbdefa81),
	.w7(32'hbb854351),
	.w8(32'hba42e904),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b529470),
	.w1(32'h3b239e79),
	.w2(32'hbac50def),
	.w3(32'h3b6ad9d5),
	.w4(32'h3a6966c3),
	.w5(32'hb864a52e),
	.w6(32'h3b6ed907),
	.w7(32'hbb38fb47),
	.w8(32'h3a0ad581),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b585834),
	.w1(32'h3a044232),
	.w2(32'h39e1a124),
	.w3(32'h3bb6357c),
	.w4(32'h3a42a351),
	.w5(32'h39dd05ee),
	.w6(32'h3a69da8e),
	.w7(32'h3a24bc1c),
	.w8(32'h3acf1bce),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd278e),
	.w1(32'h3b090bc1),
	.w2(32'h3affd7b8),
	.w3(32'h3af1ba02),
	.w4(32'h3abeb285),
	.w5(32'h3b14226e),
	.w6(32'h39cbab6c),
	.w7(32'hba66ea9c),
	.w8(32'h3a0eb8d2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b256937),
	.w1(32'hb9f78f49),
	.w2(32'hb98d32d6),
	.w3(32'h3af70f0f),
	.w4(32'h3a23aed2),
	.w5(32'h3b23c1d9),
	.w6(32'hba458d80),
	.w7(32'h3a21623b),
	.w8(32'h3ad58749),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba954cdb),
	.w1(32'hba920578),
	.w2(32'h3a3bc6d7),
	.w3(32'hbb036331),
	.w4(32'hb9039e1a),
	.w5(32'h3a9d9c02),
	.w6(32'hba8985d1),
	.w7(32'h3923e932),
	.w8(32'h3a34becf),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5451f8),
	.w1(32'h3a8675cd),
	.w2(32'h3ac39274),
	.w3(32'hba16cdd5),
	.w4(32'h3a821fd2),
	.w5(32'h3ad9af3f),
	.w6(32'h3a0c1a52),
	.w7(32'h3aec5449),
	.w8(32'h3a32b281),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13db72),
	.w1(32'hb8d30c11),
	.w2(32'hb8d1620f),
	.w3(32'h3a050160),
	.w4(32'hbb0dbbf1),
	.w5(32'hbb18f597),
	.w6(32'hbaa83271),
	.w7(32'hbba8c2b7),
	.w8(32'hbb5421a2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a924168),
	.w1(32'hba0dfcdb),
	.w2(32'hbb790c8c),
	.w3(32'hbb1f144c),
	.w4(32'hbb115864),
	.w5(32'hbb861cb3),
	.w6(32'hbb70d061),
	.w7(32'hbbb64369),
	.w8(32'hbb32da50),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbee305),
	.w1(32'h3ba62304),
	.w2(32'h3c448c91),
	.w3(32'hbbc6b0e1),
	.w4(32'hbb15538c),
	.w5(32'h3c16c645),
	.w6(32'h3b85a69b),
	.w7(32'h3c4542f5),
	.w8(32'h3b0ee0ae),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05d1c4),
	.w1(32'h3b48e473),
	.w2(32'h3b8bcd9f),
	.w3(32'hbaa7085c),
	.w4(32'h3b02acd8),
	.w5(32'h3b5b8cd7),
	.w6(32'h3a69dc37),
	.w7(32'h38c4238f),
	.w8(32'h3ab4741c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a474d),
	.w1(32'h39f38372),
	.w2(32'h3aa1ab84),
	.w3(32'h393e8e67),
	.w4(32'hbb0d7171),
	.w5(32'hb9d64a45),
	.w6(32'hbb532431),
	.w7(32'hbb6951d6),
	.w8(32'hb99d5c1d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adadc46),
	.w1(32'h3a3ef178),
	.w2(32'hbab7f04c),
	.w3(32'hb906c129),
	.w4(32'hbabe9e11),
	.w5(32'hba374596),
	.w6(32'hbb316efc),
	.w7(32'hbb345dd8),
	.w8(32'h3ad44a5f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cd2b6),
	.w1(32'h399fae6b),
	.w2(32'h3a6a477a),
	.w3(32'hbb03b4eb),
	.w4(32'hb908d506),
	.w5(32'h37fc2050),
	.w6(32'hba6983e7),
	.w7(32'hba0a511b),
	.w8(32'hba912789),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b6a640),
	.w1(32'h3b095250),
	.w2(32'h3acc23cc),
	.w3(32'hbac31b16),
	.w4(32'hbab60a22),
	.w5(32'hb9b2d35a),
	.w6(32'hba9c9cec),
	.w7(32'hbab26ce0),
	.w8(32'hbaa99722),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8573c47),
	.w1(32'hb9435dee),
	.w2(32'h3c646f2b),
	.w3(32'hbb3ada00),
	.w4(32'hbb39e798),
	.w5(32'h3c5d2601),
	.w6(32'hbba6792b),
	.w7(32'h3b605c85),
	.w8(32'hbb02a42b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4aebe),
	.w1(32'hbb619fd7),
	.w2(32'hbab8e500),
	.w3(32'h3b2a3bb6),
	.w4(32'h38547576),
	.w5(32'h3a8f3e75),
	.w6(32'h392c6ee1),
	.w7(32'h3a2dedf2),
	.w8(32'h3b85ff98),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fd530),
	.w1(32'h3b077da0),
	.w2(32'h3b083d7c),
	.w3(32'h3be4d73d),
	.w4(32'h3a238489),
	.w5(32'h3a0c7bb6),
	.w6(32'h3a800842),
	.w7(32'hba5b7d26),
	.w8(32'hba9348fe),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bf25e),
	.w1(32'h3a733b2c),
	.w2(32'h38e1ad9f),
	.w3(32'hba361eaf),
	.w4(32'hb91b61c5),
	.w5(32'hb8c50516),
	.w6(32'hb9ab3b93),
	.w7(32'hbae60fed),
	.w8(32'hbaa0fa43),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab563a4),
	.w1(32'hbb18c93f),
	.w2(32'hbb0c5dfa),
	.w3(32'h39858da0),
	.w4(32'hbb2364cc),
	.w5(32'hbb1df121),
	.w6(32'hbb2658aa),
	.w7(32'hbb222bc8),
	.w8(32'hba987e94),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb427fbf),
	.w1(32'hba1bb07e),
	.w2(32'hbb00b21a),
	.w3(32'hba8bb5d4),
	.w4(32'hba4dfd0a),
	.w5(32'h39f3535b),
	.w6(32'hba43a59b),
	.w7(32'h3b13c4f4),
	.w8(32'hbb2eaa86),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb369503),
	.w1(32'hba0c019c),
	.w2(32'h3a02ceae),
	.w3(32'hba08929d),
	.w4(32'hbb0f090e),
	.w5(32'h3aeb1039),
	.w6(32'hbaa104dc),
	.w7(32'hb90306d0),
	.w8(32'h3a933ed8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85d860),
	.w1(32'h3ac17f1f),
	.w2(32'h3a9fbc41),
	.w3(32'h3a0e0ac1),
	.w4(32'hb8bb5dfa),
	.w5(32'hb94326b5),
	.w6(32'hb9c18eb4),
	.w7(32'hbb0646b0),
	.w8(32'hbad99a85),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a085672),
	.w1(32'h3ad9e30d),
	.w2(32'h3a057be4),
	.w3(32'hbae64aed),
	.w4(32'h3b038464),
	.w5(32'h3b5789bd),
	.w6(32'h3a513945),
	.w7(32'h3b23ce95),
	.w8(32'h3b7938fb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5d32b),
	.w1(32'h3a18b266),
	.w2(32'h3a489d9a),
	.w3(32'h3b43daf8),
	.w4(32'h3a45b506),
	.w5(32'h3ad21e5e),
	.w6(32'hb9ce0be7),
	.w7(32'h3a36bc90),
	.w8(32'h3a9d6dec),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12e7d1),
	.w1(32'h3ab33fce),
	.w2(32'h3ae0d697),
	.w3(32'h3a4ce255),
	.w4(32'h3aa020c7),
	.w5(32'h3ad998a0),
	.w6(32'h393729e0),
	.w7(32'h39f606e9),
	.w8(32'h3a888a15),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfdf4a),
	.w1(32'h3a2f291f),
	.w2(32'h3a85c567),
	.w3(32'h3a60b142),
	.w4(32'h38f93bb6),
	.w5(32'h3ac72353),
	.w6(32'hb9fc762c),
	.w7(32'hba0dd481),
	.w8(32'h3ac453b4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbb442),
	.w1(32'h3b0c3cee),
	.w2(32'hb8577d2b),
	.w3(32'h3b44120b),
	.w4(32'h3be48ded),
	.w5(32'h3b4163b5),
	.w6(32'h3c3a60f6),
	.w7(32'h3b5f685d),
	.w8(32'h3c02bfbd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac96d07),
	.w1(32'hba674f70),
	.w2(32'hbab91f6a),
	.w3(32'h3bc74778),
	.w4(32'hb9f5bf4e),
	.w5(32'hb9f614c7),
	.w6(32'h3a1163ff),
	.w7(32'hb9e1ce38),
	.w8(32'hb9631842),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e99229),
	.w1(32'hba902b53),
	.w2(32'hbae644d2),
	.w3(32'hb9e8e9e0),
	.w4(32'h3a562666),
	.w5(32'h3aaa4d68),
	.w6(32'hbadfdf24),
	.w7(32'hbaaa962b),
	.w8(32'hb9d35c87),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e29d0),
	.w1(32'hbbc64be1),
	.w2(32'hbb1ae653),
	.w3(32'hba8988aa),
	.w4(32'hbacb9db0),
	.w5(32'h3b2dad26),
	.w6(32'hbbb7139e),
	.w7(32'hbab9d9f3),
	.w8(32'h3b615e12),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16567a),
	.w1(32'hbaca2f41),
	.w2(32'h3a9618b6),
	.w3(32'h3b7f8f66),
	.w4(32'hbb5b1593),
	.w5(32'hba66a750),
	.w6(32'hbb1046dc),
	.w7(32'hbb07d0e1),
	.w8(32'hbac2d0da),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8545f4a),
	.w1(32'h3a5e60b9),
	.w2(32'h3afc7441),
	.w3(32'h382586d2),
	.w4(32'hba1e1157),
	.w5(32'h3a843bb4),
	.w6(32'hb9acbd1c),
	.w7(32'h3a27085e),
	.w8(32'h393a6614),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b173fee),
	.w1(32'h3a9c753a),
	.w2(32'hbb15f2d1),
	.w3(32'h3a9e8c58),
	.w4(32'h3922c433),
	.w5(32'hba951d85),
	.w6(32'h3b4f0f99),
	.w7(32'hbb0f95d1),
	.w8(32'h3aa59dbc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39443413),
	.w1(32'h3bd5c6f9),
	.w2(32'h3c8d107d),
	.w3(32'hbab8fa9e),
	.w4(32'h3a057834),
	.w5(32'h3c73f959),
	.w6(32'h39d502d9),
	.w7(32'h3c084513),
	.w8(32'h3a8501d3),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c431f94),
	.w1(32'hb9ab8e79),
	.w2(32'hba9f3145),
	.w3(32'h3bc3c4ba),
	.w4(32'hb98ef376),
	.w5(32'hb9f906f5),
	.w6(32'hba856100),
	.w7(32'hbb1353bc),
	.w8(32'hba708a4f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d00162),
	.w1(32'h3945d22e),
	.w2(32'h3a431b24),
	.w3(32'hb9fd70e3),
	.w4(32'h39ea474f),
	.w5(32'h3a90b2e2),
	.w6(32'hba53b374),
	.w7(32'hba22b1f3),
	.w8(32'h39a9e4fb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad42135),
	.w1(32'h395dc9a9),
	.w2(32'h3aabe65d),
	.w3(32'h3b11cd37),
	.w4(32'h3a8d593f),
	.w5(32'h3b149753),
	.w6(32'hb9562042),
	.w7(32'h3abc3dae),
	.w8(32'h3a9d9026),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf8958),
	.w1(32'h3ad8d3ca),
	.w2(32'h3b22bca8),
	.w3(32'h3a37a565),
	.w4(32'h3a86f4f1),
	.w5(32'h3a136fa1),
	.w6(32'h39c10f4b),
	.w7(32'h3ba0cb38),
	.w8(32'h3b1c4e91),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18e622),
	.w1(32'h39f0871a),
	.w2(32'hba8934e4),
	.w3(32'h3a520430),
	.w4(32'hb88604c0),
	.w5(32'hb9e21804),
	.w6(32'hb98f75be),
	.w7(32'hbaf40371),
	.w8(32'h3b21b116),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2188ab),
	.w1(32'hb9200011),
	.w2(32'hba650e32),
	.w3(32'h3b482359),
	.w4(32'h393e6fbd),
	.w5(32'hb9cb0b57),
	.w6(32'hba26b391),
	.w7(32'hba67756c),
	.w8(32'h3aceb1c9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0132d2),
	.w1(32'hbac13c72),
	.w2(32'hbb1c4dd5),
	.w3(32'h3b1436f3),
	.w4(32'hba1fbc55),
	.w5(32'hba33db86),
	.w6(32'hba4016fa),
	.w7(32'hbab4fea7),
	.w8(32'h3a03f4ec),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ec909),
	.w1(32'hbb4c966f),
	.w2(32'h3a665b68),
	.w3(32'hbad12894),
	.w4(32'h3ac4f20f),
	.w5(32'h3b7fa6e8),
	.w6(32'h3b462cf6),
	.w7(32'h3b71932b),
	.w8(32'h3b8c16da),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c40e6),
	.w1(32'h3b0115f6),
	.w2(32'hba15f47e),
	.w3(32'h3a8dfdb8),
	.w4(32'h39caec5f),
	.w5(32'h38e48b43),
	.w6(32'h3a9005fc),
	.w7(32'h38400b11),
	.w8(32'h38975228),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44f57c),
	.w1(32'hb781380b),
	.w2(32'h3a488459),
	.w3(32'hbaa8871d),
	.w4(32'h39fc0d5a),
	.w5(32'h3b503ba1),
	.w6(32'h3858e201),
	.w7(32'h3b184fdc),
	.w8(32'hbae7835f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafe506),
	.w1(32'h3ae6b78f),
	.w2(32'h3ac4fddc),
	.w3(32'h39ada943),
	.w4(32'h3a9dbda9),
	.w5(32'h3b6c1bd2),
	.w6(32'h39734bc7),
	.w7(32'h3abdc0bd),
	.w8(32'h3a8a3a34),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b880e49),
	.w1(32'h3bbb7e72),
	.w2(32'h3ba33dcc),
	.w3(32'h3b2a7dee),
	.w4(32'h3b1f27ac),
	.w5(32'h3b4e6883),
	.w6(32'h3b51bc2a),
	.w7(32'h3aee4b7e),
	.w8(32'h3afc1b90),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7da8e2),
	.w1(32'hbaff7e6f),
	.w2(32'hbaabbef6),
	.w3(32'hbb3f9801),
	.w4(32'hbb410cb0),
	.w5(32'hb9e08e9e),
	.w6(32'hbb7c1217),
	.w7(32'hbabde77b),
	.w8(32'h3952797a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c08f89),
	.w1(32'hba7499af),
	.w2(32'h388ec0be),
	.w3(32'hb8c97a02),
	.w4(32'hbaa0feda),
	.w5(32'hba8b9d2e),
	.w6(32'hba53c1fc),
	.w7(32'hbabb37d8),
	.w8(32'hba3e0d51),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c3f906),
	.w1(32'hbb509688),
	.w2(32'hbaa6ca0d),
	.w3(32'h3a194a90),
	.w4(32'hbb0969da),
	.w5(32'hbabbd4d3),
	.w6(32'hbb406602),
	.w7(32'hbb0b1e31),
	.w8(32'hbba724ff),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc606db),
	.w1(32'hbb5f15e3),
	.w2(32'hba9addf0),
	.w3(32'hbaf9961b),
	.w4(32'hba39f0a0),
	.w5(32'h3b03b766),
	.w6(32'hbb5ec927),
	.w7(32'hba72188d),
	.w8(32'h3b0b9221),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7d8eb),
	.w1(32'hba8d21c7),
	.w2(32'hb93f4401),
	.w3(32'h3b59602a),
	.w4(32'hba978a34),
	.w5(32'h39bac978),
	.w6(32'hba9b4196),
	.w7(32'hba5f9cd0),
	.w8(32'hb989b432),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb94c4),
	.w1(32'hba62c824),
	.w2(32'hbac7878b),
	.w3(32'hb9e08e87),
	.w4(32'hba216e6d),
	.w5(32'h3abcda1d),
	.w6(32'hbaa81c54),
	.w7(32'h3a80adce),
	.w8(32'hba02a15a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45e5ad),
	.w1(32'h3b484ccd),
	.w2(32'h3a667eef),
	.w3(32'hbaf413a8),
	.w4(32'h3b569069),
	.w5(32'h3ac7f62c),
	.w6(32'h3baf3ff2),
	.w7(32'h3b5c581d),
	.w8(32'h3bcc074f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39868bee),
	.w1(32'h3b384aaa),
	.w2(32'h3ad9e451),
	.w3(32'h3b1a6d44),
	.w4(32'h3b1d3f40),
	.w5(32'h3ba04cd9),
	.w6(32'h3bc55dc3),
	.w7(32'h3bc0438e),
	.w8(32'h3b065415),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4436a),
	.w1(32'h3ae27cdc),
	.w2(32'h39826404),
	.w3(32'h3b0e3227),
	.w4(32'h3a78cb71),
	.w5(32'h3a0e833b),
	.w6(32'h3a7075e6),
	.w7(32'h38a66333),
	.w8(32'h3aed9a97),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b132a19),
	.w1(32'hbac4b61f),
	.w2(32'h3b52edd5),
	.w3(32'h3ae31e47),
	.w4(32'hbae2ea04),
	.w5(32'h3b73cf93),
	.w6(32'hbb2e0481),
	.w7(32'h3a243058),
	.w8(32'h3953f60e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0027b),
	.w1(32'h3a873ae2),
	.w2(32'h3a88fd52),
	.w3(32'hb9cc684f),
	.w4(32'h3adb7ebc),
	.w5(32'h3b4410d3),
	.w6(32'h3a243796),
	.w7(32'h3ac11878),
	.w8(32'h3a1e8701),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38015f54),
	.w1(32'h3a53cbbe),
	.w2(32'h3a7884e0),
	.w3(32'h3a51a214),
	.w4(32'h3a0ac883),
	.w5(32'h3a81328c),
	.w6(32'hb8f7b7d0),
	.w7(32'hb982b8e5),
	.w8(32'hb80a6091),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b6507),
	.w1(32'h3affca2f),
	.w2(32'h3afd4281),
	.w3(32'h3aecf7bd),
	.w4(32'h3ac3713f),
	.w5(32'h3a8f1474),
	.w6(32'h3a2d3be6),
	.w7(32'h39c941b2),
	.w8(32'h39f48b3a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8d976),
	.w1(32'h3b1e4088),
	.w2(32'h3ab6e665),
	.w3(32'h3ae420d0),
	.w4(32'h37da6af9),
	.w5(32'hb971f999),
	.w6(32'hb9fe4770),
	.w7(32'hbb24f660),
	.w8(32'hbaffd2c1),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7501c6),
	.w1(32'h39c49681),
	.w2(32'h3b23f351),
	.w3(32'h39a1ce0d),
	.w4(32'hb68c51f7),
	.w5(32'h3b058193),
	.w6(32'h3af2f1cb),
	.w7(32'h3ae114a3),
	.w8(32'h3ad3b63b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba950b96),
	.w1(32'hbb8910e3),
	.w2(32'hbbb3f625),
	.w3(32'hbafe3e84),
	.w4(32'hbb662254),
	.w5(32'hbb0f0b37),
	.w6(32'hbb8d3a06),
	.w7(32'hbb1a02f9),
	.w8(32'hbab097aa),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf77d9),
	.w1(32'hbb038f6a),
	.w2(32'h39a85274),
	.w3(32'hbb97caa1),
	.w4(32'hbaba7122),
	.w5(32'h3ae730e2),
	.w6(32'hbb7f0a70),
	.w7(32'hbb0e08c1),
	.w8(32'h39b61e94),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2b1ab),
	.w1(32'hba037cba),
	.w2(32'h3b5b3b08),
	.w3(32'h3b3dd861),
	.w4(32'hba41617d),
	.w5(32'h3b47b3f5),
	.w6(32'hba0f84eb),
	.w7(32'h3b26024b),
	.w8(32'hb8219eab),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b94f0),
	.w1(32'hbbd52254),
	.w2(32'hbbf3958d),
	.w3(32'hbbaf8f92),
	.w4(32'hbb51a582),
	.w5(32'hbb1d0dbc),
	.w6(32'hbbcfa9ff),
	.w7(32'hbbc5659c),
	.w8(32'hba9b94b2),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98b908),
	.w1(32'h3ad49f8d),
	.w2(32'h3b15bfea),
	.w3(32'hbb922197),
	.w4(32'hb9bace3b),
	.w5(32'h37b73d8b),
	.w6(32'h3a21ffe9),
	.w7(32'hbae635dc),
	.w8(32'hbabd8484),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac286e7),
	.w1(32'h3ac08430),
	.w2(32'h3b86cd51),
	.w3(32'hba9e9304),
	.w4(32'h3b8cde12),
	.w5(32'h3beeb9a7),
	.w6(32'h3be04c62),
	.w7(32'h3bfc3f27),
	.w8(32'h3b90c17c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a4568),
	.w1(32'hb95b0e18),
	.w2(32'hba563dc6),
	.w3(32'h3b95a6a2),
	.w4(32'hbaaebea0),
	.w5(32'hbae401ce),
	.w6(32'hb8c47abe),
	.w7(32'hba2981d0),
	.w8(32'h39e5feff),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1be893),
	.w1(32'h398d386b),
	.w2(32'h3adb50c0),
	.w3(32'hb9e81fa8),
	.w4(32'hb9014daa),
	.w5(32'h3aa2ec65),
	.w6(32'hbaab5c9a),
	.w7(32'hbaf0fa27),
	.w8(32'hba8df5c2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a494dcb),
	.w1(32'hbad4f1eb),
	.w2(32'hb9aaddbc),
	.w3(32'hba7097d9),
	.w4(32'hba13faae),
	.w5(32'hba8dcdcc),
	.w6(32'hba009dba),
	.w7(32'h3a9151bf),
	.w8(32'h3af1930d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40fdaf),
	.w1(32'h3c39988e),
	.w2(32'h3c88f60c),
	.w3(32'h3aa39174),
	.w4(32'hb9a4d932),
	.w5(32'h3c5ca8cb),
	.w6(32'h3b58e02e),
	.w7(32'h3bfd4c12),
	.w8(32'hbaab61e7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a8408),
	.w1(32'hba45295d),
	.w2(32'hbb166fa1),
	.w3(32'h3b02200b),
	.w4(32'hba7d22e7),
	.w5(32'hba631c28),
	.w6(32'h392a0bb7),
	.w7(32'hb947f522),
	.w8(32'h3af0fe96),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07a21d),
	.w1(32'h3a68afc9),
	.w2(32'h3ab646ce),
	.w3(32'h3a907919),
	.w4(32'hb9db78f9),
	.w5(32'h3a9b9e8d),
	.w6(32'hba859e60),
	.w7(32'h39883478),
	.w8(32'h39b953e5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf4fb4),
	.w1(32'h3a8367fb),
	.w2(32'h3aa95708),
	.w3(32'hbad31d4a),
	.w4(32'hb9f8a487),
	.w5(32'hb9cacedd),
	.w6(32'hb9443b8f),
	.w7(32'hbae7ef38),
	.w8(32'hbac0e29a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae58815),
	.w1(32'h3986957a),
	.w2(32'hba5c2fa4),
	.w3(32'hb83f6934),
	.w4(32'h3a355e08),
	.w5(32'h39b68966),
	.w6(32'h3a60fe13),
	.w7(32'hb94fb680),
	.w8(32'h3ae19ad2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb0bc7),
	.w1(32'h3a88dd9b),
	.w2(32'h3a9b31c5),
	.w3(32'h3abda22f),
	.w4(32'h38b1fe4f),
	.w5(32'hba3692d4),
	.w6(32'h3ac66c87),
	.w7(32'hbb0e481f),
	.w8(32'hbaecc83e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba10a2f),
	.w1(32'h3bdf1160),
	.w2(32'h3bb1816b),
	.w3(32'h3b00a7ed),
	.w4(32'h3b0e4dbd),
	.w5(32'h3a8fa97f),
	.w6(32'h3b2cb04e),
	.w7(32'hbab08467),
	.w8(32'hba1edd61),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bcd6e),
	.w1(32'h3ad3daf4),
	.w2(32'h3ac5591a),
	.w3(32'h3b38c498),
	.w4(32'h3b564211),
	.w5(32'h3af1286e),
	.w6(32'h3b4dd2dc),
	.w7(32'h394fb5f9),
	.w8(32'h3a746edf),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcbe02),
	.w1(32'hb848d8b0),
	.w2(32'h3aaa8dad),
	.w3(32'hbaa78335),
	.w4(32'hba01be62),
	.w5(32'h3ac1f9dc),
	.w6(32'h39886544),
	.w7(32'h3ae62786),
	.w8(32'h3af17102),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cafa4),
	.w1(32'hbb102e1b),
	.w2(32'h3b5a36e4),
	.w3(32'h3a9f8c50),
	.w4(32'h398d2340),
	.w5(32'h3b746d87),
	.w6(32'h3b833a09),
	.w7(32'h3b41b2e5),
	.w8(32'h3b6693ee),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f37ae),
	.w1(32'h3ac09f9f),
	.w2(32'h3ab2fdc2),
	.w3(32'h3b50d42a),
	.w4(32'h3992606a),
	.w5(32'h39ca5494),
	.w6(32'h3a2598fb),
	.w7(32'h39efd965),
	.w8(32'h39ead9cf),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc7171),
	.w1(32'h39f3c139),
	.w2(32'hba65b895),
	.w3(32'hb9451842),
	.w4(32'h3a7d2882),
	.w5(32'hb9fdf89d),
	.w6(32'hbad8f623),
	.w7(32'hbb559826),
	.w8(32'h3a185bea),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9f641),
	.w1(32'h3b018771),
	.w2(32'h3c199311),
	.w3(32'h3aa519c5),
	.w4(32'h399cfc87),
	.w5(32'h3c2c6f93),
	.w6(32'h3bc4504f),
	.w7(32'h3c895d48),
	.w8(32'hb92bba29),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c118d),
	.w1(32'hba274dfe),
	.w2(32'hbb2eee1e),
	.w3(32'hbb20939b),
	.w4(32'hbac67498),
	.w5(32'hbb2d2cdc),
	.w6(32'hbae44a68),
	.w7(32'hbae06019),
	.w8(32'hbb81b9d1),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb966143),
	.w1(32'h3a4e23a0),
	.w2(32'h396b189b),
	.w3(32'hbb1fd2b2),
	.w4(32'hb8ee423e),
	.w5(32'h393bf93e),
	.w6(32'h3a4d4dca),
	.w7(32'h3a19328d),
	.w8(32'h3add39c1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a81e6),
	.w1(32'h3920a588),
	.w2(32'h39df5eaa),
	.w3(32'h3a94876d),
	.w4(32'hba3d4fe8),
	.w5(32'h3a791f38),
	.w6(32'h3a29498b),
	.w7(32'hba694c94),
	.w8(32'h3b379ee0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab13d3f),
	.w1(32'hbab397da),
	.w2(32'hb9e5b6d1),
	.w3(32'hb9df62ad),
	.w4(32'hba596de7),
	.w5(32'h39fc992c),
	.w6(32'hbaef6ab9),
	.w7(32'h3aed058c),
	.w8(32'hbb4a7927),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4c46d),
	.w1(32'hba31330e),
	.w2(32'hbba38196),
	.w3(32'hbb7812b2),
	.w4(32'h39855137),
	.w5(32'hbb4e5f7f),
	.w6(32'h3a850203),
	.w7(32'hba81893f),
	.w8(32'h3ac356e6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47bba5),
	.w1(32'h3b27012d),
	.w2(32'h3bb7298f),
	.w3(32'h3b206156),
	.w4(32'h3af89a79),
	.w5(32'h3b82ac54),
	.w6(32'h37f333b9),
	.w7(32'hbad86ab3),
	.w8(32'h3ac50260),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d9289),
	.w1(32'h3afa62b2),
	.w2(32'h3ac047c3),
	.w3(32'h3b97d28a),
	.w4(32'h376a2ced),
	.w5(32'h3a016458),
	.w6(32'h39bca8c4),
	.w7(32'hb9bb91e9),
	.w8(32'h39ae8ae1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf4f5f),
	.w1(32'hba724a23),
	.w2(32'h39bffab4),
	.w3(32'h3aa04260),
	.w4(32'hb980be59),
	.w5(32'h3ab078c1),
	.w6(32'hbafa7234),
	.w7(32'hbab65711),
	.w8(32'hb8a962f6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55bec4),
	.w1(32'h3b09dc43),
	.w2(32'h3b35e005),
	.w3(32'h3b903de7),
	.w4(32'h3ab99f46),
	.w5(32'h3b03b2d2),
	.w6(32'h3aafd04e),
	.w7(32'h3a906e79),
	.w8(32'h3a0437e5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c2fda6),
	.w1(32'h3aa74db8),
	.w2(32'h3a92a873),
	.w3(32'hb9d806d5),
	.w4(32'hba03ac70),
	.w5(32'hb9a1f4f3),
	.w6(32'hba221cdd),
	.w7(32'hbac288ed),
	.w8(32'hba4cc88f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7faee),
	.w1(32'h3b061d13),
	.w2(32'h3b210a46),
	.w3(32'hba32c6e5),
	.w4(32'hba8a5854),
	.w5(32'hba2489aa),
	.w6(32'hbade5ebe),
	.w7(32'hbb87f814),
	.w8(32'hbb4a40a9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bb84f),
	.w1(32'hba948b98),
	.w2(32'h383dacd1),
	.w3(32'hba5fb038),
	.w4(32'hb9e41c99),
	.w5(32'h3a84c5fe),
	.w6(32'hbb07a3f6),
	.w7(32'hbad3d14a),
	.w8(32'hb90edf0e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5a6ea),
	.w1(32'hba78e97b),
	.w2(32'hba7bd9bd),
	.w3(32'h3b102a6b),
	.w4(32'hbadd5670),
	.w5(32'hbaa69efe),
	.w6(32'hba89ddae),
	.w7(32'hba7e5763),
	.w8(32'hb7e5e798),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964e0f4),
	.w1(32'h3b44bc08),
	.w2(32'h3b528700),
	.w3(32'hba811da2),
	.w4(32'h3a96ba76),
	.w5(32'h3aa01815),
	.w6(32'h3a75f7b6),
	.w7(32'h3a5cd123),
	.w8(32'h3aad11c5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a690c),
	.w1(32'hbaf88e5e),
	.w2(32'h3b55e9d5),
	.w3(32'h3b311fcd),
	.w4(32'hbb25fed4),
	.w5(32'h3a779d7e),
	.w6(32'hbaff0955),
	.w7(32'h3b42ee02),
	.w8(32'h3aca3b45),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b881d31),
	.w1(32'h3b85a08a),
	.w2(32'h3b7474a1),
	.w3(32'h3b4ad2eb),
	.w4(32'h3afc9c14),
	.w5(32'h3aecca64),
	.w6(32'h3af4bc3c),
	.w7(32'h3a89013d),
	.w8(32'h3b12e793),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9001db),
	.w1(32'h3a21ad95),
	.w2(32'hba1c9550),
	.w3(32'h3b76ef5b),
	.w4(32'h3958afe0),
	.w5(32'hba1156ea),
	.w6(32'h3ab24c2e),
	.w7(32'h391fcccb),
	.w8(32'hb9edf31a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980d0c7),
	.w1(32'h3a19f787),
	.w2(32'hbaadeecd),
	.w3(32'hba657cc0),
	.w4(32'h3a0884f0),
	.w5(32'hba0c5a54),
	.w6(32'hb93705b7),
	.w7(32'hbb2892f8),
	.w8(32'hba068c8b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b953e),
	.w1(32'hbada6a9d),
	.w2(32'h3942bb74),
	.w3(32'h38efb31d),
	.w4(32'hba10bedc),
	.w5(32'h3ad77cd7),
	.w6(32'hbb45a57b),
	.w7(32'hbb113660),
	.w8(32'hb9276657),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fb6ce),
	.w1(32'hb955287f),
	.w2(32'h397d81b2),
	.w3(32'h3b5ac5f3),
	.w4(32'h39100af9),
	.w5(32'h3a853c36),
	.w6(32'hba9b3738),
	.w7(32'hba9e81e2),
	.w8(32'hb9e1a5f5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a577b98),
	.w1(32'hb9a029bd),
	.w2(32'h39ee953c),
	.w3(32'h3ac8bd6f),
	.w4(32'hb893a359),
	.w5(32'h3a97e378),
	.w6(32'hbacbf6f2),
	.w7(32'hbabb8ef8),
	.w8(32'hb96f7472),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada79f8),
	.w1(32'h3a90aaae),
	.w2(32'h3a2f48c2),
	.w3(32'h3b13e05f),
	.w4(32'hbacca8f5),
	.w5(32'hbb0d23b9),
	.w6(32'hba8c482f),
	.w7(32'hbb260015),
	.w8(32'hbab06dba),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980b71a),
	.w1(32'h3a4a3474),
	.w2(32'h3bb36179),
	.w3(32'h3a13d2b7),
	.w4(32'h3a6326c3),
	.w5(32'h3bf21de8),
	.w6(32'hb8a77b26),
	.w7(32'h3bd7bcc3),
	.w8(32'hba1e343e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdfbd8),
	.w1(32'h3b6515a1),
	.w2(32'h3b4fde9b),
	.w3(32'hbaf29946),
	.w4(32'h392f600f),
	.w5(32'h3a9381f3),
	.w6(32'h39729c57),
	.w7(32'hb94f6f08),
	.w8(32'h3a0a4f4f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b434344),
	.w1(32'h3aafc08d),
	.w2(32'h3b391a63),
	.w3(32'h3a868e29),
	.w4(32'hb8b486ec),
	.w5(32'h3ab98ee2),
	.w6(32'h38973635),
	.w7(32'h3abf667c),
	.w8(32'h3a62aa57),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb9d73),
	.w1(32'h3999e537),
	.w2(32'h3a19de2f),
	.w3(32'h3aaa75ec),
	.w4(32'h39bdf9d8),
	.w5(32'h3a50424c),
	.w6(32'hba221f11),
	.w7(32'hba228772),
	.w8(32'h3910216a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8ca4a),
	.w1(32'h3acaccdd),
	.w2(32'h3a0b40ba),
	.w3(32'h3acef1e5),
	.w4(32'hbaa2ba3f),
	.w5(32'hbb7b8c22),
	.w6(32'h382ad9d7),
	.w7(32'hbaa366cf),
	.w8(32'hb9b046c1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45a719),
	.w1(32'h39bb37d8),
	.w2(32'hbb225e0a),
	.w3(32'hbb5e6e29),
	.w4(32'hb858833d),
	.w5(32'hbab013f0),
	.w6(32'hba55f911),
	.w7(32'hbb48915d),
	.w8(32'h3afd10a0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d85e1),
	.w1(32'h3bc3c7ec),
	.w2(32'h3bafc0e0),
	.w3(32'h3bade369),
	.w4(32'h3ae00e97),
	.w5(32'h3b8e217d),
	.w6(32'h3b27b56f),
	.w7(32'h3a3e8421),
	.w8(32'hb9c7bdc0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21059f),
	.w1(32'h39606b12),
	.w2(32'hb7e6c5cc),
	.w3(32'hba257f27),
	.w4(32'h39a9c88d),
	.w5(32'h39652c98),
	.w6(32'h3968f0f4),
	.w7(32'h393ea7b0),
	.w8(32'hb92dbb8c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa349fa),
	.w1(32'h3a035c5c),
	.w2(32'h39d7ecf7),
	.w3(32'hb9d42285),
	.w4(32'hba28b4e7),
	.w5(32'hbad06954),
	.w6(32'h3a7433e5),
	.w7(32'hb9a1926f),
	.w8(32'h3a712117),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule