module layer_6_featuremap_111(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21cdf8),
	.w1(32'hb8a5d7ae),
	.w2(32'h3afbb7ed),
	.w3(32'hbb44e4c6),
	.w4(32'h3b6429a9),
	.w5(32'hba9681f4),
	.w6(32'hba3e85ef),
	.w7(32'h3b7404d9),
	.w8(32'hb9cee4bf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395783c8),
	.w1(32'hbc0751fa),
	.w2(32'hbbe95a5b),
	.w3(32'hbbe9ef4e),
	.w4(32'hbc08bf19),
	.w5(32'hbc0d5cf1),
	.w6(32'hbba5cb70),
	.w7(32'h3a8a1c98),
	.w8(32'hbada20b0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55af01),
	.w1(32'hbc87ef48),
	.w2(32'h3a92ead9),
	.w3(32'h3bf71f9a),
	.w4(32'h3b7f39b5),
	.w5(32'hbbeb63a5),
	.w6(32'hbb9cb795),
	.w7(32'hbb76174c),
	.w8(32'h39cd65a5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcd6ae),
	.w1(32'hb9588a8f),
	.w2(32'h3a8bae77),
	.w3(32'h3acde152),
	.w4(32'h3b029e25),
	.w5(32'h3a93e867),
	.w6(32'h3ac9d7b4),
	.w7(32'h3bb70599),
	.w8(32'h3bb9efed),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f7f72),
	.w1(32'hbc134b64),
	.w2(32'hbca64bf0),
	.w3(32'h3c7033c5),
	.w4(32'h3cb7a646),
	.w5(32'h3cd5d608),
	.w6(32'hbd21e2a3),
	.w7(32'hbd6a319b),
	.w8(32'hbce46e31),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf2452),
	.w1(32'hbb573393),
	.w2(32'hba9027d4),
	.w3(32'hbb3d6a24),
	.w4(32'h3b10a957),
	.w5(32'h3b26c019),
	.w6(32'hbb89efe9),
	.w7(32'hbab90fc8),
	.w8(32'h3abadcae),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5c234),
	.w1(32'hbc411432),
	.w2(32'hbb90178f),
	.w3(32'hbb418c4f),
	.w4(32'hbb96cb14),
	.w5(32'hbab36486),
	.w6(32'hbaf839b7),
	.w7(32'h3a9cfa9b),
	.w8(32'hbb0c6bcb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cef60),
	.w1(32'hbd4be258),
	.w2(32'hbd604c2e),
	.w3(32'h3c44aa29),
	.w4(32'h3c9d7361),
	.w5(32'h3b7e6ed3),
	.w6(32'h3bae546d),
	.w7(32'hba819a08),
	.w8(32'hbbcac150),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd16a354),
	.w1(32'h3c6fc3b7),
	.w2(32'h3cdda41c),
	.w3(32'hbb3865e8),
	.w4(32'h3b46708f),
	.w5(32'h3c953c6f),
	.w6(32'hbca11766),
	.w7(32'hbc8d8779),
	.w8(32'hbc88a9df),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b330efa),
	.w1(32'hb9ec8a43),
	.w2(32'h3b69bd8a),
	.w3(32'hbb46ac18),
	.w4(32'h3ac5475c),
	.w5(32'h3a80af9f),
	.w6(32'hbbd86068),
	.w7(32'hbbdc7fde),
	.w8(32'hbbfa1aee),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cb047),
	.w1(32'h3a7ac96e),
	.w2(32'h3c4256c5),
	.w3(32'hbab2301e),
	.w4(32'hbb253438),
	.w5(32'hbc1f6c0d),
	.w6(32'h3c1154cb),
	.w7(32'h3c43cf55),
	.w8(32'hbc0d62ac),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d0b70),
	.w1(32'h3c02aa0c),
	.w2(32'h3c18fca6),
	.w3(32'h3bac5c62),
	.w4(32'h3bb24884),
	.w5(32'h3aae8b4e),
	.w6(32'h3b040435),
	.w7(32'h3b5aa0dc),
	.w8(32'hbb395e45),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf87b),
	.w1(32'h3a0a52a2),
	.w2(32'h3c2de4d9),
	.w3(32'hbb42e469),
	.w4(32'h3ba91145),
	.w5(32'hbaf0e0fa),
	.w6(32'hbafc258d),
	.w7(32'h3c0ba7fa),
	.w8(32'hbb101839),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc110eff),
	.w1(32'hbb7ecd5c),
	.w2(32'hbbe79c77),
	.w3(32'h3b578a27),
	.w4(32'h3c50de06),
	.w5(32'h3c9424c1),
	.w6(32'hbca20d6f),
	.w7(32'hbcabccc0),
	.w8(32'hbc2ad35d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6931af),
	.w1(32'hbc64c74c),
	.w2(32'hbc318150),
	.w3(32'hbc1282c9),
	.w4(32'hbc1eb410),
	.w5(32'hbc564011),
	.w6(32'h396a6a55),
	.w7(32'h3bca4f8e),
	.w8(32'h3b828b1c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57499c),
	.w1(32'hbb83414d),
	.w2(32'hbaeb6a4a),
	.w3(32'hbb28f217),
	.w4(32'hbb46e65a),
	.w5(32'hbb7c3bac),
	.w6(32'h3b783fbd),
	.w7(32'h3b937106),
	.w8(32'h3b9fc909),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac39afb),
	.w1(32'hb9bf8508),
	.w2(32'hbc6015b2),
	.w3(32'h3c2fc13f),
	.w4(32'h3aadf248),
	.w5(32'h3c1ac9d3),
	.w6(32'h3c107d3d),
	.w7(32'h3c366043),
	.w8(32'h3ca38c42),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bb17b),
	.w1(32'h3b25e890),
	.w2(32'h3bf904ff),
	.w3(32'hba809888),
	.w4(32'h3b662c60),
	.w5(32'h3b35d8d0),
	.w6(32'hbb0a7a26),
	.w7(32'h3a851de2),
	.w8(32'hbaabacc1),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b747ea4),
	.w1(32'hbb30244b),
	.w2(32'hbb5f472c),
	.w3(32'hba1d07a6),
	.w4(32'hbb23e3cb),
	.w5(32'hbba220d6),
	.w6(32'h3a3df24e),
	.w7(32'hbb0fc0ea),
	.w8(32'hbb82895b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2c761),
	.w1(32'h38ed300d),
	.w2(32'h3c018aea),
	.w3(32'hbc926d12),
	.w4(32'hbc7ede4f),
	.w5(32'hbbc7bdb0),
	.w6(32'h39427d8b),
	.w7(32'h3a358e5e),
	.w8(32'hba787868),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba864b5f),
	.w1(32'hba1d61bb),
	.w2(32'hba9f896a),
	.w3(32'h3b1f838f),
	.w4(32'h3a3f44c1),
	.w5(32'h3a0e18eb),
	.w6(32'h3b5d923e),
	.w7(32'h3bc8c925),
	.w8(32'h3b19b09e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a301f),
	.w1(32'h3c4a44bb),
	.w2(32'h3cb5ce83),
	.w3(32'h3bd7ded8),
	.w4(32'h3bd79e01),
	.w5(32'h3b9f23d3),
	.w6(32'h3c6dc3be),
	.w7(32'h3ca99602),
	.w8(32'h3c038440),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34c172),
	.w1(32'hbc0c927d),
	.w2(32'h3a9609ac),
	.w3(32'hbbf2c787),
	.w4(32'hbb4b0bea),
	.w5(32'hbc69281d),
	.w6(32'h3b84d8c2),
	.w7(32'h3c94621d),
	.w8(32'hbc03d3d2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf84b4a),
	.w1(32'h3ced8e73),
	.w2(32'h3d70a68d),
	.w3(32'hbd41603d),
	.w4(32'hbd59aa31),
	.w5(32'hbd320083),
	.w6(32'h3c681b5d),
	.w7(32'h3b007af1),
	.w8(32'hbb42403e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cea4e1a),
	.w1(32'hbb947642),
	.w2(32'hbb81d47d),
	.w3(32'h3a81aae0),
	.w4(32'h3c2210f8),
	.w5(32'h3c63c714),
	.w6(32'h3bba3c32),
	.w7(32'h3c8a5063),
	.w8(32'h3c80825d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca97164),
	.w1(32'h3aa690ec),
	.w2(32'h3a86f0a6),
	.w3(32'hbbf8c439),
	.w4(32'hbbec2277),
	.w5(32'hbbf61bf5),
	.w6(32'hbb6e9a41),
	.w7(32'hbbedfe6b),
	.w8(32'h3a661683),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b706),
	.w1(32'h3bc366cb),
	.w2(32'h3c201675),
	.w3(32'h3bbc76f9),
	.w4(32'h39d0cc4f),
	.w5(32'hb98abb80),
	.w6(32'h3bfe047f),
	.w7(32'hb9402181),
	.w8(32'hbb4e416b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c419d9e),
	.w1(32'hbb4a69e6),
	.w2(32'hb9d92cdb),
	.w3(32'hba5c2d46),
	.w4(32'h3a4fdfb7),
	.w5(32'h3aeffa4b),
	.w6(32'hb9804518),
	.w7(32'h3b441ad4),
	.w8(32'h3b0bfc57),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1993b4),
	.w1(32'h389c094b),
	.w2(32'hbad98c0c),
	.w3(32'hbb2f6f4a),
	.w4(32'hbb8c9ce6),
	.w5(32'hbb91a55b),
	.w6(32'h3a63fc49),
	.w7(32'hbab65e2c),
	.w8(32'hba4a677f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba98841),
	.w1(32'hbcbf8c17),
	.w2(32'hbcaed79b),
	.w3(32'hbd1b13ab),
	.w4(32'hbce606f2),
	.w5(32'h3b80206f),
	.w6(32'hbcc359f7),
	.w7(32'hbb10d7bb),
	.w8(32'h3c0ddf3b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44026a),
	.w1(32'hbcb6ea46),
	.w2(32'hbcc076a6),
	.w3(32'h3cde1bfe),
	.w4(32'h3d0896d2),
	.w5(32'h3c2659a6),
	.w6(32'h3ccee488),
	.w7(32'h3d6a4272),
	.w8(32'h3d76897f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32c53b),
	.w1(32'hbca0d664),
	.w2(32'hbc040ce0),
	.w3(32'hbc0196f9),
	.w4(32'h3b80c30e),
	.w5(32'h3bc378c0),
	.w6(32'hbc80546a),
	.w7(32'hbc40e9a8),
	.w8(32'hbbe71ea7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02b9c3),
	.w1(32'hbb76bc56),
	.w2(32'h3bfb971a),
	.w3(32'hbc1e03e0),
	.w4(32'hbd077139),
	.w5(32'hbcce3b62),
	.w6(32'h3ba9e610),
	.w7(32'h3ce66ab4),
	.w8(32'h3cc9ddbe),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06d111),
	.w1(32'hb921406c),
	.w2(32'hbc5afe07),
	.w3(32'hbc78b5f2),
	.w4(32'hbb55552b),
	.w5(32'hbbad19f7),
	.w6(32'hbc806cb0),
	.w7(32'hbc48737d),
	.w8(32'hbb3ff8f1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bec29),
	.w1(32'hbaa7c672),
	.w2(32'hbb3eb2a0),
	.w3(32'h3a1a3bb5),
	.w4(32'hba41de7f),
	.w5(32'h3aab631d),
	.w6(32'hbbc81db9),
	.w7(32'hbbcfb649),
	.w8(32'hbad80418),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff46eb),
	.w1(32'hbb3c9c7c),
	.w2(32'h3acfa844),
	.w3(32'hbbc54918),
	.w4(32'hb9e184cd),
	.w5(32'h3ac63550),
	.w6(32'hbbb99e63),
	.w7(32'h3a3a3c88),
	.w8(32'h3b912c8f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ffed),
	.w1(32'h3adc2062),
	.w2(32'hb9140148),
	.w3(32'h3ad3384d),
	.w4(32'h3ba1add3),
	.w5(32'h3addbec5),
	.w6(32'hba157b08),
	.w7(32'h3ab001c6),
	.w8(32'h3a49f13b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e8500),
	.w1(32'h3adeb72a),
	.w2(32'h3aa56883),
	.w3(32'hb8c10e5f),
	.w4(32'hba39e80e),
	.w5(32'h3ae94c87),
	.w6(32'h3bc1de7c),
	.w7(32'h3bd5a9fc),
	.w8(32'h3c104b90),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2a394),
	.w1(32'hbbdf7715),
	.w2(32'hbc13ac84),
	.w3(32'h3b7e56c0),
	.w4(32'hbb486338),
	.w5(32'hbbed7214),
	.w6(32'hbb50b14a),
	.w7(32'hbb9923e1),
	.w8(32'hbc8b4531),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c7832),
	.w1(32'hbc777fd7),
	.w2(32'h3bdca27a),
	.w3(32'hbc883130),
	.w4(32'hbcf2b611),
	.w5(32'hbc6a8682),
	.w6(32'hbc8a490c),
	.w7(32'hbac14f4f),
	.w8(32'h3b98a618),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb823262),
	.w1(32'h3c01395b),
	.w2(32'h3cc5e8fd),
	.w3(32'h3b59ce11),
	.w4(32'hbc0e0e92),
	.w5(32'hbc8cd3f3),
	.w6(32'hbc3c800f),
	.w7(32'h3b7ba191),
	.w8(32'hbc20c4e9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4a536),
	.w1(32'hbb45ca59),
	.w2(32'hbaeaaf6e),
	.w3(32'hba5274be),
	.w4(32'hbb2089ba),
	.w5(32'hbb90c238),
	.w6(32'h3a824b8d),
	.w7(32'h3b4c328d),
	.w8(32'h390ed27f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e1dcd),
	.w1(32'h3b2f0e72),
	.w2(32'hbaec9d22),
	.w3(32'h3b5288c6),
	.w4(32'h3bcc53fd),
	.w5(32'hbb23f80e),
	.w6(32'h3b8bcbd3),
	.w7(32'h3b0aca40),
	.w8(32'hba4eba43),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ec554),
	.w1(32'hbcaa6499),
	.w2(32'hbcb68db6),
	.w3(32'hbca122d7),
	.w4(32'hbc02999e),
	.w5(32'hb9e71b56),
	.w6(32'hbc30b64a),
	.w7(32'h3cc31c8c),
	.w8(32'h3cf81d8e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03f715),
	.w1(32'h3bd4c7da),
	.w2(32'h3c1fb428),
	.w3(32'hbbbd8191),
	.w4(32'hbab80ab6),
	.w5(32'hbb5728f4),
	.w6(32'hbb2d21a5),
	.w7(32'hbbae309e),
	.w8(32'hbc145ee8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a247847),
	.w1(32'hbcaeeacc),
	.w2(32'hbc21009e),
	.w3(32'hbb7d2794),
	.w4(32'hbcbc4689),
	.w5(32'hbcf62e5c),
	.w6(32'hbb44ca85),
	.w7(32'hbc643059),
	.w8(32'hbcd9cdf4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04ac79),
	.w1(32'hbcd3ef7f),
	.w2(32'hbca062f9),
	.w3(32'hbb923270),
	.w4(32'hbc043f7f),
	.w5(32'hbb947c22),
	.w6(32'hbb927f06),
	.w7(32'hb8779ee0),
	.w8(32'h3c42618b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76227c),
	.w1(32'hbbbf45e5),
	.w2(32'h3c537574),
	.w3(32'hbc5fcc33),
	.w4(32'hbcac4d88),
	.w5(32'hbc8e6797),
	.w6(32'h3c885e6e),
	.w7(32'h3d1438c4),
	.w8(32'h3cf76fbf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2be0c),
	.w1(32'hbb8757be),
	.w2(32'hbb5dfeb2),
	.w3(32'hbb917ae1),
	.w4(32'hbbe9436b),
	.w5(32'hbbe2fba4),
	.w6(32'hbb2347a9),
	.w7(32'hbba4421b),
	.w8(32'hbbde3c98),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb01f66),
	.w1(32'hbcb6999e),
	.w2(32'hbca94c39),
	.w3(32'h3cbc1d98),
	.w4(32'h3d0c324b),
	.w5(32'h3c39a315),
	.w6(32'h3c1efd90),
	.w7(32'h3c83f14a),
	.w8(32'h3c7d9f26),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb00e79),
	.w1(32'h3bbccaee),
	.w2(32'h3c1c9601),
	.w3(32'h3b74aad3),
	.w4(32'hb82151d8),
	.w5(32'h39c53a2a),
	.w6(32'h3bd50694),
	.w7(32'h3c3044fc),
	.w8(32'h3bd81d5f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf9e0f),
	.w1(32'hbc08d525),
	.w2(32'hbb8c43a2),
	.w3(32'hbbfce670),
	.w4(32'hbbf731cc),
	.w5(32'hbb707d77),
	.w6(32'hbb1f7611),
	.w7(32'hbab61984),
	.w8(32'hbabb29f8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ab0de),
	.w1(32'hbb1d6f2f),
	.w2(32'h3c0d3cf0),
	.w3(32'hbaf74e8c),
	.w4(32'hbb0de56a),
	.w5(32'h3af08448),
	.w6(32'h3bd89ec4),
	.w7(32'h3c29e9c7),
	.w8(32'h3c3996fa),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc48ce1),
	.w1(32'hbbf19171),
	.w2(32'h3aab683f),
	.w3(32'hbb3539a1),
	.w4(32'hbc021dcf),
	.w5(32'hbbf71409),
	.w6(32'h3bc73af1),
	.w7(32'h3c7566ee),
	.w8(32'h3c7850de),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b0ee4),
	.w1(32'h3b626a1a),
	.w2(32'h3be580a9),
	.w3(32'hbc0d94ca),
	.w4(32'hbc2b3f84),
	.w5(32'hbc1ddcc5),
	.w6(32'hbab40f63),
	.w7(32'h3b460e8e),
	.w8(32'hbb58c08a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28bba8),
	.w1(32'hbc370def),
	.w2(32'hb9b431aa),
	.w3(32'h3a82c097),
	.w4(32'hbb2b0278),
	.w5(32'hbbaac044),
	.w6(32'hbaa73e7c),
	.w7(32'hbcaba5bc),
	.w8(32'hbbdc0a3d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcebefc3),
	.w1(32'hba99b192),
	.w2(32'hba587bd0),
	.w3(32'hba2a4f1c),
	.w4(32'hbb7148dc),
	.w5(32'hbbe5c901),
	.w6(32'hba67d393),
	.w7(32'h3b26b007),
	.w8(32'hbb8a442f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd007a0),
	.w1(32'hbb7c9c5c),
	.w2(32'h3c39fbac),
	.w3(32'h3b9e5474),
	.w4(32'hbb2ac35e),
	.w5(32'h3b82c8f4),
	.w6(32'h3b46c45a),
	.w7(32'hbbbf2f37),
	.w8(32'hbca6b07e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4156ec),
	.w1(32'h38cd8151),
	.w2(32'hb9279ca0),
	.w3(32'hba951d29),
	.w4(32'h3947fbe5),
	.w5(32'h3af8301b),
	.w6(32'hba8be591),
	.w7(32'hbb104c9b),
	.w8(32'hb9d152e1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ab8fc),
	.w1(32'h3b7112a5),
	.w2(32'h3c46cd2b),
	.w3(32'h3c48ee93),
	.w4(32'hb9e118e1),
	.w5(32'h3c4348fb),
	.w6(32'h3cd16c1a),
	.w7(32'h3d20fd42),
	.w8(32'h3bcbd0f4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be51af5),
	.w1(32'hbabb7706),
	.w2(32'hbbac983b),
	.w3(32'hbb3f4b52),
	.w4(32'hbba8a5a1),
	.w5(32'hba81f6a4),
	.w6(32'hbb1fc1dc),
	.w7(32'hbb8d3536),
	.w8(32'h3a2dff0a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8df86c),
	.w1(32'h3bcdb835),
	.w2(32'h3bc97096),
	.w3(32'hbc0218cf),
	.w4(32'hbc49d61c),
	.w5(32'hbb1c7e6d),
	.w6(32'h3be6a54d),
	.w7(32'h3c1b5581),
	.w8(32'h3b95d13c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58a65e),
	.w1(32'hbc586fc1),
	.w2(32'hbd241cec),
	.w3(32'hbc50aac2),
	.w4(32'hbcbce8e9),
	.w5(32'hbc4ac671),
	.w6(32'h3ca1e49b),
	.w7(32'h3d347f2d),
	.w8(32'h3c8c91d7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5190a9),
	.w1(32'hbbcb5488),
	.w2(32'hb9d24f45),
	.w3(32'hbbc4aa52),
	.w4(32'hbab76af1),
	.w5(32'h3aa122d6),
	.w6(32'hbb8646c1),
	.w7(32'hbb203cad),
	.w8(32'h3b877a05),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule