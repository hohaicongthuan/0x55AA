module layer_10_featuremap_173(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb683cd3a),
	.w1(32'hb66fd694),
	.w2(32'hb71f563a),
	.w3(32'hb6230d79),
	.w4(32'hb63da5c6),
	.w5(32'hb78beac5),
	.w6(32'hb6b81f44),
	.w7(32'hb72be878),
	.w8(32'hb69edc32),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b79aec),
	.w1(32'h358c387f),
	.w2(32'h38c70759),
	.w3(32'h366345c8),
	.w4(32'h38f086b1),
	.w5(32'h390c399c),
	.w6(32'h390ee44b),
	.w7(32'h3911c6bb),
	.w8(32'h3981ef2b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5839e49),
	.w1(32'hb62d9402),
	.w2(32'hb6239a66),
	.w3(32'h35243601),
	.w4(32'hb49840ee),
	.w5(32'hb5a5fdcf),
	.w6(32'hb65d52b0),
	.w7(32'hb68d01fa),
	.w8(32'hb6c8c602),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6467dfc),
	.w1(32'hb7a9f4a3),
	.w2(32'hb827b665),
	.w3(32'h37511a0f),
	.w4(32'h37b9c022),
	.w5(32'hb765b0a1),
	.w6(32'h375ca568),
	.w7(32'h37a74af4),
	.w8(32'hb72b3ccd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b5c7cc),
	.w1(32'h3600d4d3),
	.w2(32'hb6a7666b),
	.w3(32'h370a4c93),
	.w4(32'h3630e55f),
	.w5(32'h3584658e),
	.w6(32'h37044073),
	.w7(32'h34efaf66),
	.w8(32'hb6f9f621),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c99ba0),
	.w1(32'h375641f7),
	.w2(32'hb4ebbd0b),
	.w3(32'h374a277e),
	.w4(32'h35c83159),
	.w5(32'hb74162d7),
	.w6(32'h33494cba),
	.w7(32'hb7215c28),
	.w8(32'hb793c109),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39306090),
	.w1(32'h394a2132),
	.w2(32'hb8ac72ea),
	.w3(32'h395b8dfc),
	.w4(32'h3969cb79),
	.w5(32'h39367c13),
	.w6(32'h38c6afda),
	.w7(32'h38a36c85),
	.w8(32'hb80191b8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7efb0c7),
	.w1(32'hb89d325b),
	.w2(32'hb994ba9e),
	.w3(32'hba082e1d),
	.w4(32'hb9fd52d0),
	.w5(32'hba451bde),
	.w6(32'hba21d125),
	.w7(32'hb9bd9f11),
	.w8(32'hb97defe7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2aa3a),
	.w1(32'hb7307a8f),
	.w2(32'h361834dc),
	.w3(32'h375eb1bd),
	.w4(32'h383ba441),
	.w5(32'h38a38839),
	.w6(32'hb79a8590),
	.w7(32'h381c041d),
	.w8(32'h3838c390),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eac339),
	.w1(32'h3a1f21d5),
	.w2(32'h3a240834),
	.w3(32'hba345bcd),
	.w4(32'h382bad82),
	.w5(32'h39190220),
	.w6(32'hbaafd9bf),
	.w7(32'hba5069d7),
	.w8(32'hba0e3fa3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a7159c),
	.w1(32'h35bd3e4f),
	.w2(32'hb72a6344),
	.w3(32'h3788ddcb),
	.w4(32'hb6d0b0b8),
	.w5(32'hb728f715),
	.w6(32'h3614e96e),
	.w7(32'hb70f8c64),
	.w8(32'hb790f939),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efb6f2),
	.w1(32'h383a5780),
	.w2(32'h3a25e5aa),
	.w3(32'hb99f3ea4),
	.w4(32'h395202f3),
	.w5(32'h3a7beb0e),
	.w6(32'hb876e9fe),
	.w7(32'h3a1afc28),
	.w8(32'h3a8c49ef),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03326a),
	.w1(32'h3a17cdae),
	.w2(32'h3a2ed67a),
	.w3(32'hba80adcd),
	.w4(32'hb914d7e1),
	.w5(32'hb93647fe),
	.w6(32'hbac7c5fe),
	.w7(32'hba360886),
	.w8(32'hb9e663f7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb841df4e),
	.w1(32'h395310b5),
	.w2(32'h3990839f),
	.w3(32'hb7c43c70),
	.w4(32'h37b156cc),
	.w5(32'h39443952),
	.w6(32'hb8a83eda),
	.w7(32'h3834e17b),
	.w8(32'h3928470e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388596eb),
	.w1(32'h3988334a),
	.w2(32'h39a4f605),
	.w3(32'hb9c734e9),
	.w4(32'hb96cca46),
	.w5(32'hb86c1b7f),
	.w6(32'hb984f982),
	.w7(32'hb80dcdfe),
	.w8(32'h396c947e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888a328),
	.w1(32'h38b7cee4),
	.w2(32'h3906892f),
	.w3(32'hb9c1afa8),
	.w4(32'hb98e20cb),
	.w5(32'hb9bcd3cc),
	.w6(32'hba31e7b3),
	.w7(32'hb9eaa69f),
	.w8(32'hb9faf022),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371381f9),
	.w1(32'h35625fce),
	.w2(32'hb6d08380),
	.w3(32'hb696d7d6),
	.w4(32'hb61e8c08),
	.w5(32'hb70ecd3f),
	.w6(32'hb585d105),
	.w7(32'hb6a6ecd7),
	.w8(32'hb7346588),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34a3d075),
	.w1(32'h3964f3be),
	.w2(32'h36b841cf),
	.w3(32'hba07c8a5),
	.w4(32'hb90270c5),
	.w5(32'hb985ded1),
	.w6(32'hba71681d),
	.w7(32'hb9b1d443),
	.w8(32'hba164f24),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d3224),
	.w1(32'hb8a8d14c),
	.w2(32'hb8c4204b),
	.w3(32'hba1b49f8),
	.w4(32'hb9adf913),
	.w5(32'hb9ababfa),
	.w6(32'hba3fc380),
	.w7(32'hb9ca9be3),
	.w8(32'hb9cc1e42),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364872cc),
	.w1(32'h3342475e),
	.w2(32'hb68755c4),
	.w3(32'h367f563b),
	.w4(32'h34e7632a),
	.w5(32'hb6993799),
	.w6(32'h35d60c30),
	.w7(32'hb619e764),
	.w8(32'hb6d25c7a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f3504f),
	.w1(32'h36505b17),
	.w2(32'h3568334e),
	.w3(32'h36e4fa11),
	.w4(32'h3607e67d),
	.w5(32'hb655b740),
	.w6(32'h35da3e15),
	.w7(32'hb5f6eb99),
	.w8(32'hb725170e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a31d94),
	.w1(32'h36aa48e3),
	.w2(32'hb79c1a27),
	.w3(32'h385bd178),
	.w4(32'h38e9fbcc),
	.w5(32'h389c6aa6),
	.w6(32'h386bc553),
	.w7(32'h38d13779),
	.w8(32'h38f5863d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02f18d),
	.w1(32'h3999445f),
	.w2(32'hb99ec0c4),
	.w3(32'hb9a01e5c),
	.w4(32'hb93032fd),
	.w5(32'hba2b5d43),
	.w6(32'hb9885d98),
	.w7(32'hb8b314e7),
	.w8(32'h3a07e3ed),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909f032),
	.w1(32'h3a232b4f),
	.w2(32'h39fe80c4),
	.w3(32'hba0e4a64),
	.w4(32'hb83ef337),
	.w5(32'hb81f2659),
	.w6(32'hba82c159),
	.w7(32'hba20384f),
	.w8(32'hb99f511d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f86caf),
	.w1(32'h39931d1e),
	.w2(32'h3a3bc5a4),
	.w3(32'hba3dfef8),
	.w4(32'hb925c3b6),
	.w5(32'h395afbf3),
	.w6(32'hba48237a),
	.w7(32'hb954be24),
	.w8(32'h39f35a07),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e5ab0a),
	.w1(32'h3772a565),
	.w2(32'hb56535ce),
	.w3(32'h377bec11),
	.w4(32'h37972f5d),
	.w5(32'h3685826a),
	.w6(32'h3782c984),
	.w7(32'h362d80ef),
	.w8(32'hb66a0420),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb736e146),
	.w1(32'hb6989f8d),
	.w2(32'hb680004d),
	.w3(32'h35eb598c),
	.w4(32'h371e4364),
	.w5(32'h372e1d90),
	.w6(32'h3707947c),
	.w7(32'h35ee720f),
	.w8(32'hb59066b8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb973895b),
	.w1(32'h39020e49),
	.w2(32'h399c0b27),
	.w3(32'hb95ec9d4),
	.w4(32'h394bb070),
	.w5(32'h39935ce2),
	.w6(32'hb99e9833),
	.w7(32'hb8401bbd),
	.w8(32'h397b9d15),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba009ee8),
	.w1(32'hb8f6e887),
	.w2(32'hb8d82508),
	.w3(32'hb9992d14),
	.w4(32'hb7b74134),
	.w5(32'h38e93de5),
	.w6(32'hb812b1da),
	.w7(32'h39560727),
	.w8(32'h39b41412),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3747e90b),
	.w1(32'h39ea457d),
	.w2(32'h3a0070f2),
	.w3(32'hb9c4564d),
	.w4(32'h3755342a),
	.w5(32'h390e4135),
	.w6(32'hba064d1d),
	.w7(32'hb9158205),
	.w8(32'h38fe3c89),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72d094d),
	.w1(32'hb66b924a),
	.w2(32'hb658d9ec),
	.w3(32'hb6ed0dd8),
	.w4(32'hb600a9f8),
	.w5(32'hb5d51337),
	.w6(32'hb49b466d),
	.w7(32'h3467a9bc),
	.w8(32'h34941105),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3465d167),
	.w1(32'hb675b73e),
	.w2(32'hb66e7cfc),
	.w3(32'h33c782f0),
	.w4(32'hb66360e4),
	.w5(32'hb686c7c9),
	.w6(32'hb67ae408),
	.w7(32'hb710dc5b),
	.w8(32'hb7453e89),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974848d),
	.w1(32'h39a92f50),
	.w2(32'h38e49808),
	.w3(32'hb99e2249),
	.w4(32'hb95ea0b6),
	.w5(32'hb9b35c81),
	.w6(32'hb9a9ef56),
	.w7(32'hb991e526),
	.w8(32'hb980e224),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a47a4),
	.w1(32'h383156c6),
	.w2(32'h39562eb6),
	.w3(32'hb9113a17),
	.w4(32'hb775a952),
	.w5(32'h38c1dff9),
	.w6(32'hb76f8652),
	.w7(32'h38e5b77c),
	.w8(32'h396ea387),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81238d3),
	.w1(32'h36a15681),
	.w2(32'h386c5918),
	.w3(32'hb86b6ace),
	.w4(32'hb80da558),
	.w5(32'hb719d991),
	.w6(32'hb7b2e43e),
	.w7(32'h35b76b2c),
	.w8(32'h37a0f24e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89dbdc7),
	.w1(32'h39146785),
	.w2(32'hb7aad35e),
	.w3(32'hb90bddfe),
	.w4(32'h38a7cccb),
	.w5(32'hb7519676),
	.w6(32'hb93691fb),
	.w7(32'hb7701352),
	.w8(32'hb8452890),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9829299),
	.w1(32'h382d28a1),
	.w2(32'hb98719f2),
	.w3(32'h39783ae6),
	.w4(32'h37227479),
	.w5(32'hba9af7b6),
	.w6(32'hb94d0daa),
	.w7(32'hb9cf6935),
	.w8(32'hba244aa4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba0ea7),
	.w1(32'hb9cae5b0),
	.w2(32'h39b698f2),
	.w3(32'hb85a2b85),
	.w4(32'h3a889545),
	.w5(32'h3ae4bf2d),
	.w6(32'h39935878),
	.w7(32'h3a867f00),
	.w8(32'h3b05aa17),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67c8d6),
	.w1(32'hb9e63ba3),
	.w2(32'hb7dc50cd),
	.w3(32'h3713f766),
	.w4(32'h3a57b1bc),
	.w5(32'h3a893a94),
	.w6(32'h3a4c7a7b),
	.w7(32'h3aa4e72e),
	.w8(32'h3ae11c2b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382d8423),
	.w1(32'h38eff646),
	.w2(32'h39b469e7),
	.w3(32'hb9761d26),
	.w4(32'hb8cca836),
	.w5(32'h3931c899),
	.w6(32'hb9a56e3b),
	.w7(32'hb8cd0801),
	.w8(32'h39545561),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3795f4e0),
	.w1(32'h3711e3af),
	.w2(32'hb6c4361b),
	.w3(32'h36cf9d56),
	.w4(32'hb53743bc),
	.w5(32'hb74b719d),
	.w6(32'h352f3a59),
	.w7(32'hb717ba33),
	.w8(32'hb8002927),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79a5649),
	.w1(32'h358b6a7e),
	.w2(32'hb701e08e),
	.w3(32'h379ea9ef),
	.w4(32'h37f29430),
	.w5(32'h37f3815b),
	.w6(32'h37d2e8b3),
	.w7(32'h37b7c72a),
	.w8(32'h37b9c8f3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad3fe8),
	.w1(32'hb9868dcc),
	.w2(32'hb93a75c7),
	.w3(32'hb9963e32),
	.w4(32'hb90fa13a),
	.w5(32'hb89d25af),
	.w6(32'hb7920809),
	.w7(32'h38b646f3),
	.w8(32'h38ac8905),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a7cf3),
	.w1(32'h39ae66e0),
	.w2(32'h39f57cbe),
	.w3(32'hba59fe59),
	.w4(32'hb9f67a92),
	.w5(32'hb96d6c6f),
	.w6(32'hbaaa1e65),
	.w7(32'hba36b0b6),
	.w8(32'hb9fb933f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e666c1),
	.w1(32'h3a2ab8bd),
	.w2(32'h3a1d4c66),
	.w3(32'hb9f76973),
	.w4(32'h38e0b00f),
	.w5(32'h39428c8b),
	.w6(32'hba15d104),
	.w7(32'hb8a1b437),
	.w8(32'h3981d46e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f75c4),
	.w1(32'h3a40b79a),
	.w2(32'h3a1480ab),
	.w3(32'hba0e122f),
	.w4(32'h3889d044),
	.w5(32'h37fe719b),
	.w6(32'hba879040),
	.w7(32'hba18e8c0),
	.w8(32'hb99037ba),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d7abb),
	.w1(32'h3997d3ef),
	.w2(32'h3a09c2b9),
	.w3(32'hb9cf401f),
	.w4(32'h361762ad),
	.w5(32'h399626a5),
	.w6(32'hb9fb8ce4),
	.w7(32'h38f127f9),
	.w8(32'h3a0c0fdc),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ae5a2),
	.w1(32'hb92636eb),
	.w2(32'hba1ea679),
	.w3(32'hba281dd7),
	.w4(32'hba274352),
	.w5(32'hba844d73),
	.w6(32'hbab1a8f7),
	.w7(32'hba896496),
	.w8(32'hba96ad02),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37431e77),
	.w1(32'h37a4f03c),
	.w2(32'h37952860),
	.w3(32'h3752d785),
	.w4(32'h37869fb9),
	.w5(32'h372fedef),
	.w6(32'h372bbc81),
	.w7(32'h375ce47f),
	.w8(32'h351e4e14),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380e1855),
	.w1(32'h3884236f),
	.w2(32'h38623a9b),
	.w3(32'h37ff29a0),
	.w4(32'h3844fe0d),
	.w5(32'h3829903a),
	.w6(32'h370acb28),
	.w7(32'h37cff336),
	.w8(32'h37fd1bb4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372bef8c),
	.w1(32'h37c8b4e8),
	.w2(32'h36a92a6e),
	.w3(32'h3752cb89),
	.w4(32'h37cf3a94),
	.w5(32'h3686769b),
	.w6(32'h3658ec06),
	.w7(32'h3739154f),
	.w8(32'hb6a907d5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bf00bd),
	.w1(32'h39ab8588),
	.w2(32'h380f1b8a),
	.w3(32'hb9bb7e75),
	.w4(32'h3896eee8),
	.w5(32'h371f39ad),
	.w6(32'hb9c51277),
	.w7(32'hb9bab072),
	.w8(32'hb968eac3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bef609),
	.w1(32'h38f4cfe3),
	.w2(32'h3859b6de),
	.w3(32'h3771de19),
	.w4(32'h388140e4),
	.w5(32'h379ffb84),
	.w6(32'hb70de1f2),
	.w7(32'h37de1f23),
	.w8(32'h37c3ea82),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a924b),
	.w1(32'h3a13468d),
	.w2(32'h399d1b5c),
	.w3(32'hb9b1c913),
	.w4(32'h38a203e4),
	.w5(32'hb99beb48),
	.w6(32'hba70fb8b),
	.w7(32'hba0f74bb),
	.w8(32'hba2fdbb3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc698f),
	.w1(32'h3843f370),
	.w2(32'h38abdc11),
	.w3(32'hb88325eb),
	.w4(32'h38522e8b),
	.w5(32'h38bd93e7),
	.w6(32'hb8270384),
	.w7(32'h389b1d89),
	.w8(32'h3918a115),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5eaedb1),
	.w1(32'h361ea79a),
	.w2(32'hb5b7466e),
	.w3(32'hb5db4910),
	.w4(32'h362a8ac3),
	.w5(32'hb58d9f81),
	.w6(32'h36d960a5),
	.w7(32'h359fd5c4),
	.w8(32'h33ac047c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c0761e),
	.w1(32'h36b1c1ee),
	.w2(32'h3645f77e),
	.w3(32'h3687954a),
	.w4(32'h36c879f6),
	.w5(32'h37042e70),
	.w6(32'h37082399),
	.w7(32'h36a5f142),
	.w8(32'h35f5966c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ab02b8),
	.w1(32'hb68b53b6),
	.w2(32'h36786acb),
	.w3(32'hb6b5be28),
	.w4(32'hb6cc844d),
	.w5(32'h369cdcc0),
	.w6(32'hb742d9bf),
	.w7(32'hb6f1dd54),
	.w8(32'hb6940736),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bbefb),
	.w1(32'hb919e053),
	.w2(32'hb8d7aa46),
	.w3(32'hb92f4797),
	.w4(32'hb8ad7f80),
	.w5(32'hb8056e49),
	.w6(32'h383d471d),
	.w7(32'h3892eac2),
	.w8(32'h38a1d09f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f516f5),
	.w1(32'h3904f5bf),
	.w2(32'h38592b0a),
	.w3(32'h3827f198),
	.w4(32'h3890b023),
	.w5(32'hb801a845),
	.w6(32'hb66df786),
	.w7(32'h37b4ae3d),
	.w8(32'hb7a8d458),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f151e1),
	.w1(32'h39632eca),
	.w2(32'h39def0d1),
	.w3(32'hba148fd2),
	.w4(32'h37cf87e6),
	.w5(32'h38513139),
	.w6(32'hba3aca90),
	.w7(32'hb91ac7f4),
	.w8(32'hb88aa739),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939ab4c),
	.w1(32'hb8b0004d),
	.w2(32'hb87aeeaf),
	.w3(32'hb8b583a3),
	.w4(32'hb7f13637),
	.w5(32'hb8a6f36b),
	.w6(32'hb904efc1),
	.w7(32'hb705d1c7),
	.w8(32'hb87dadc9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36999a03),
	.w1(32'h368696b1),
	.w2(32'hb69028cc),
	.w3(32'h34ac5ce8),
	.w4(32'h364c65bb),
	.w5(32'hb71606e1),
	.w6(32'h35bb9476),
	.w7(32'hb67b19b2),
	.w8(32'hb6b32b2a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3669fef1),
	.w1(32'hb5ea1e2d),
	.w2(32'hb6c66b47),
	.w3(32'h3581c05a),
	.w4(32'hb642ca6d),
	.w5(32'hb6ede3e0),
	.w6(32'h35195fbd),
	.w7(32'hb692f70b),
	.w8(32'hb72dd682),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b1ff4e),
	.w1(32'h371b4e7a),
	.w2(32'h37d38231),
	.w3(32'h363aca6f),
	.w4(32'h364a5f47),
	.w5(32'h3713c94b),
	.w6(32'hb6f1dffd),
	.w7(32'hb70f3fe4),
	.w8(32'hb72becd0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a5435b),
	.w1(32'hb68d2cf9),
	.w2(32'hb668f7db),
	.w3(32'h36145ef6),
	.w4(32'hb5d975b3),
	.w5(32'hb5eceb54),
	.w6(32'hb5b894c6),
	.w7(32'hb52e225f),
	.w8(32'hb706780b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9186b5f),
	.w1(32'hb9267cdc),
	.w2(32'h39711477),
	.w3(32'hb8e9a118),
	.w4(32'hb9126c2d),
	.w5(32'hb91c4bc2),
	.w6(32'hba2ae9ef),
	.w7(32'hb9e48259),
	.w8(32'hb9df3b50),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4e374),
	.w1(32'h3a1fbc4e),
	.w2(32'h39a51dda),
	.w3(32'h388aaec1),
	.w4(32'h39d44ef8),
	.w5(32'h396d1e23),
	.w6(32'hb920d97d),
	.w7(32'hb7c98abb),
	.w8(32'hb8c80366),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db4957),
	.w1(32'h3939053e),
	.w2(32'h3a18e5c9),
	.w3(32'hb9a05c29),
	.w4(32'h38eced47),
	.w5(32'h39fa266d),
	.w6(32'hb985d52f),
	.w7(32'h3921cbf6),
	.w8(32'h3a17c9e2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eff59f),
	.w1(32'h3a8455eb),
	.w2(32'h3b0ead0c),
	.w3(32'hba5cf755),
	.w4(32'hb99fa529),
	.w5(32'h3a12b483),
	.w6(32'hb998215f),
	.w7(32'h3a07c3e4),
	.w8(32'h3aca80ae),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37105c13),
	.w1(32'h3625620c),
	.w2(32'hb75ebed9),
	.w3(32'h372c0d54),
	.w4(32'hb2b8c31b),
	.w5(32'hb75b78d2),
	.w6(32'h35bb51c4),
	.w7(32'hb735b7ed),
	.w8(32'hb7aa04ff),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37276b9e),
	.w1(32'hb5b0abb7),
	.w2(32'hb75ba017),
	.w3(32'h374382a2),
	.w4(32'h34a33a7c),
	.w5(32'hb74d42bc),
	.w6(32'h3645ec2b),
	.w7(32'hb7128633),
	.w8(32'hb7c3c084),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3708ae72),
	.w1(32'hb59f4103),
	.w2(32'hb780975b),
	.w3(32'h3736b3d7),
	.w4(32'hb6284c73),
	.w5(32'hb791b578),
	.w6(32'hb6a8d84e),
	.w7(32'hb77423f7),
	.w8(32'hb800126d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9757331),
	.w1(32'h3863efa0),
	.w2(32'h38092dc5),
	.w3(32'hb90c7065),
	.w4(32'hb64aabad),
	.w5(32'h37520026),
	.w6(32'hb91b9005),
	.w7(32'hb86e39da),
	.w8(32'hb86ed54f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37495e2f),
	.w1(32'h371e3312),
	.w2(32'h36327bf0),
	.w3(32'h378e16a9),
	.w4(32'h3777acb6),
	.w5(32'h361b739f),
	.w6(32'h368269d4),
	.w7(32'h350707ba),
	.w8(32'hb70b5d0f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b8faf),
	.w1(32'h391b358b),
	.w2(32'hb80e7c24),
	.w3(32'h3799bd28),
	.w4(32'hb8e719eb),
	.w5(32'hb9547e0a),
	.w6(32'hb996d119),
	.w7(32'hb9b17879),
	.w8(32'hb9d621c3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba315b51),
	.w1(32'hb99ce656),
	.w2(32'h38e5f0c0),
	.w3(32'hba0c2d9b),
	.w4(32'hba508513),
	.w5(32'hb9f0d0ca),
	.w6(32'hba54fe5f),
	.w7(32'hba29f110),
	.w8(32'hb9610a0e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993fee7),
	.w1(32'h39724ce6),
	.w2(32'h383a1cfe),
	.w3(32'hba40d933),
	.w4(32'hba02e300),
	.w5(32'hba005971),
	.w6(32'hba51aed3),
	.w7(32'hba413f5f),
	.w8(32'hba11e3a4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c627e),
	.w1(32'h3959ca10),
	.w2(32'h39192d01),
	.w3(32'hb981be52),
	.w4(32'hb87e3c54),
	.w5(32'hb89fde6b),
	.w6(32'hb9edd5e4),
	.w7(32'hb985cfc7),
	.w8(32'hb8cbf2be),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395757a9),
	.w1(32'h39a13e31),
	.w2(32'hb81cfe6d),
	.w3(32'hb8201453),
	.w4(32'h39483271),
	.w5(32'hb8c33206),
	.w6(32'hb9b23e67),
	.w7(32'hb990ede4),
	.w8(32'hb9ba83a9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2991f),
	.w1(32'h39408950),
	.w2(32'h3915c64f),
	.w3(32'hb8953783),
	.w4(32'h3846dfbc),
	.w5(32'h372f7eae),
	.w6(32'hb880a63d),
	.w7(32'h37ab6c9e),
	.w8(32'h37fa75b1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a36ba),
	.w1(32'h378f0046),
	.w2(32'hb9d93d1f),
	.w3(32'hb915d433),
	.w4(32'h389f098c),
	.w5(32'hb963f0fd),
	.w6(32'hb9e31310),
	.w7(32'hb9c654e8),
	.w8(32'hba02835c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34a49875),
	.w1(32'hb61090f1),
	.w2(32'hb629640d),
	.w3(32'h354e1453),
	.w4(32'hb5c7c863),
	.w5(32'hb619d6e9),
	.w6(32'hb57730ec),
	.w7(32'hb5f90c72),
	.w8(32'hb68044ea),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36930fcb),
	.w1(32'h362b7bec),
	.w2(32'hb63c4a8c),
	.w3(32'h3642046d),
	.w4(32'h35f230b3),
	.w5(32'hb6c75dd4),
	.w6(32'h3660a1b7),
	.w7(32'hb5ed4400),
	.w8(32'hb69e62be),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b354b5),
	.w1(32'h36655af5),
	.w2(32'h36c1ab93),
	.w3(32'h36804c50),
	.w4(32'hb629fe16),
	.w5(32'hb54d7d68),
	.w6(32'h36aa4e35),
	.w7(32'hb5b64eb1),
	.w8(32'hb7545611),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74d74ff),
	.w1(32'hb696d24e),
	.w2(32'hb67e081e),
	.w3(32'hb7932a48),
	.w4(32'hb6866c80),
	.w5(32'hb528d84c),
	.w6(32'hb6868218),
	.w7(32'hb5b27579),
	.w8(32'hb3862439),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8445d7c),
	.w1(32'h39f8d41c),
	.w2(32'h39e371d1),
	.w3(32'h37628a5e),
	.w4(32'h38917571),
	.w5(32'h3a311799),
	.w6(32'hb9852047),
	.w7(32'hb6dec956),
	.w8(32'h3a287678),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e208d),
	.w1(32'h37923c74),
	.w2(32'h36dba8e6),
	.w3(32'hb882c2cf),
	.w4(32'hb9428c41),
	.w5(32'hb9440729),
	.w6(32'h38dd928c),
	.w7(32'h386fc2fb),
	.w8(32'h37c6fbbf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a238ed9),
	.w1(32'h3a385f48),
	.w2(32'h38944efe),
	.w3(32'hb8c4ba1f),
	.w4(32'h37c8308f),
	.w5(32'hb998983e),
	.w6(32'hba1e9b4d),
	.w7(32'hb9b397fa),
	.w8(32'hba056132),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6e6cc),
	.w1(32'hb857156d),
	.w2(32'hb8100a2f),
	.w3(32'hba2847e0),
	.w4(32'hba0e2640),
	.w5(32'hb9e24fcb),
	.w6(32'hba7efc96),
	.w7(32'hba65ed0c),
	.w8(32'hba57771e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98113a0),
	.w1(32'hb7f9bc02),
	.w2(32'h397ce3fc),
	.w3(32'hb8eba5b8),
	.w4(32'h3958ec9f),
	.w5(32'h39a90bb6),
	.w6(32'h39937b90),
	.w7(32'h39fb7f33),
	.w8(32'h3a476212),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb2ab37bd),
	.w1(32'h3794bf04),
	.w2(32'hb8cc567a),
	.w3(32'h38f7b817),
	.w4(32'h3940b817),
	.w5(32'hb806d5a8),
	.w6(32'hb8056e80),
	.w7(32'h39085996),
	.w8(32'h374f4202),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec6631),
	.w1(32'h3a0c2aa7),
	.w2(32'h3a069ddb),
	.w3(32'h39c8f837),
	.w4(32'h3a42c224),
	.w5(32'h3a29185b),
	.w6(32'h39c574bc),
	.w7(32'h3a1a0f0f),
	.w8(32'h3a2a1022),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a77ae1),
	.w1(32'h3a39b51d),
	.w2(32'h3a6f71f1),
	.w3(32'hb9f01af9),
	.w4(32'hb76b0028),
	.w5(32'h39c09327),
	.w6(32'hba3fa16f),
	.w7(32'hb805db0d),
	.w8(32'h39f36e6e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39835f01),
	.w1(32'h3a05c2bc),
	.w2(32'h39ead70f),
	.w3(32'hb8ae1205),
	.w4(32'hb8875fa5),
	.w5(32'hb99c23f6),
	.w6(32'hba108772),
	.w7(32'hb95a5e8d),
	.w8(32'hba0e0b88),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cf9ea9),
	.w1(32'h39622605),
	.w2(32'hb99d7399),
	.w3(32'hba07deb6),
	.w4(32'hb9750db2),
	.w5(32'h39527e07),
	.w6(32'hb9e0e2fc),
	.w7(32'hb88e463e),
	.w8(32'h39b0219b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb627cd36),
	.w1(32'h373dde4a),
	.w2(32'h37b9a749),
	.w3(32'hb68e0ecb),
	.w4(32'h36e4e960),
	.w5(32'h37ec88b1),
	.w6(32'h36b0d8ca),
	.w7(32'h3787f163),
	.w8(32'hb66e7147),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3697c46c),
	.w1(32'h3a1bb9b1),
	.w2(32'h39becde3),
	.w3(32'hba3cf964),
	.w4(32'hb972f5e3),
	.w5(32'hb94a1b59),
	.w6(32'hba47e839),
	.w7(32'hb9ad0840),
	.w8(32'hb87786ea),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925b361),
	.w1(32'h39e4c102),
	.w2(32'h39f34af1),
	.w3(32'h39f06394),
	.w4(32'h39ac6b0f),
	.w5(32'h390478f2),
	.w6(32'h38bfdce4),
	.w7(32'hb71cde8c),
	.w8(32'h395e9d79),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a060da7),
	.w1(32'h3a21ba29),
	.w2(32'h39034f67),
	.w3(32'h38830588),
	.w4(32'hb85052f1),
	.w5(32'hba4052f4),
	.w6(32'h37b763a3),
	.w7(32'hb9516fba),
	.w8(32'hba1fd2ca),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e56157),
	.w1(32'h39edee7a),
	.w2(32'h3a06eb40),
	.w3(32'h398d7341),
	.w4(32'h3ac3ffce),
	.w5(32'h3b15ec00),
	.w6(32'h3a0a05e2),
	.w7(32'h3abfb65a),
	.w8(32'h3b1531d5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2b30c),
	.w1(32'h3a3bde4b),
	.w2(32'h39e3ae73),
	.w3(32'hb9ba267f),
	.w4(32'hb93bba6e),
	.w5(32'hb98225df),
	.w6(32'hba6db763),
	.w7(32'hba35e881),
	.w8(32'hba04bfc3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a270b21),
	.w1(32'h3a591cf3),
	.w2(32'h3976bbe8),
	.w3(32'h3998122a),
	.w4(32'h39cbe5ff),
	.w5(32'h39814358),
	.w6(32'hb93be02a),
	.w7(32'h38ad99b6),
	.w8(32'h399492b5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787a04e),
	.w1(32'h370f2243),
	.w2(32'h36ec98b3),
	.w3(32'h3739bff8),
	.w4(32'h3735109f),
	.w5(32'h3565fb2c),
	.w6(32'hb61700ec),
	.w7(32'hb69d23c4),
	.w8(32'hb68aae17),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b96736),
	.w1(32'h39ba107b),
	.w2(32'hb8d96a46),
	.w3(32'hba5567c1),
	.w4(32'hba00ee21),
	.w5(32'hba459c69),
	.w6(32'hba767b93),
	.w7(32'hba7dd752),
	.w8(32'hba2dc3ba),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99809fa),
	.w1(32'h3892bf1e),
	.w2(32'h3a4c3d4c),
	.w3(32'hb883dad3),
	.w4(32'hb7f18ad5),
	.w5(32'h39ffb9c4),
	.w6(32'h38884b5d),
	.w7(32'hb88b78fc),
	.w8(32'h39d9a029),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6948d1b),
	.w1(32'hb681750b),
	.w2(32'hb6f3f50b),
	.w3(32'hb6247f3b),
	.w4(32'hb50a13c2),
	.w5(32'hb655cc52),
	.w6(32'hb6e3cb5e),
	.w7(32'hb64f2d35),
	.w8(32'hb69843ae),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f927f2),
	.w1(32'h3814f44e),
	.w2(32'hb8ad120d),
	.w3(32'h37c1eaaf),
	.w4(32'h38c3b9d8),
	.w5(32'hb8732e84),
	.w6(32'h378d9f65),
	.w7(32'h3790f02c),
	.w8(32'hb87bcd5c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb975c673),
	.w1(32'h37ef1b8b),
	.w2(32'h38de8bf0),
	.w3(32'hba2f7eb0),
	.w4(32'hba0e1c87),
	.w5(32'hb9d6a340),
	.w6(32'hba6314da),
	.w7(32'hba1ce83d),
	.w8(32'hb9f4565b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fac695),
	.w1(32'h39be37e6),
	.w2(32'h3998a61b),
	.w3(32'hb993e3b5),
	.w4(32'hb81c8c59),
	.w5(32'hb5035603),
	.w6(32'hb9ec56b9),
	.w7(32'hb9bdc9d2),
	.w8(32'hb90eb7ec),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e139c8),
	.w1(32'hb913dd2b),
	.w2(32'hb86a347d),
	.w3(32'hb97e7dc8),
	.w4(32'hb96ccae1),
	.w5(32'hb958ef09),
	.w6(32'hb9336f29),
	.w7(32'h387b965f),
	.w8(32'h3934f4e1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39458cb0),
	.w1(32'h39ada14f),
	.w2(32'hb91ce27f),
	.w3(32'h3871d2a4),
	.w4(32'h3741c2bc),
	.w5(32'hb9e87e3e),
	.w6(32'h38975d90),
	.w7(32'hb8dbbc12),
	.w8(32'hb8cc540a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e15f63),
	.w1(32'h391a3122),
	.w2(32'h3912680a),
	.w3(32'h38d0f8a2),
	.w4(32'h3979ba71),
	.w5(32'h39baaeb7),
	.w6(32'h38646e66),
	.w7(32'h39a03a6f),
	.w8(32'h39eda200),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397338c3),
	.w1(32'h3966913a),
	.w2(32'h384cae89),
	.w3(32'h389fea02),
	.w4(32'h374cd564),
	.w5(32'hb8aae5e6),
	.w6(32'hb9b7caca),
	.w7(32'hb9c0b848),
	.w8(32'hb9ef09ae),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e45b22),
	.w1(32'h3943644e),
	.w2(32'h3973d5cd),
	.w3(32'hb93765d6),
	.w4(32'hb6e25cb4),
	.w5(32'h38accf6a),
	.w6(32'hb9650c54),
	.w7(32'hb90a1185),
	.w8(32'h38333256),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367cf7d2),
	.w1(32'h33df4651),
	.w2(32'h341ff2fc),
	.w3(32'h36a2af65),
	.w4(32'h31c94071),
	.w5(32'h362fe11f),
	.w6(32'hb595147b),
	.w7(32'h3535d730),
	.w8(32'hb50a6739),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5eca2f5),
	.w1(32'hb6a0460d),
	.w2(32'hb71f9eb3),
	.w3(32'hb63a2c35),
	.w4(32'hb60b7ff1),
	.w5(32'hb70e9b87),
	.w6(32'hb52f17e1),
	.w7(32'hb6327986),
	.w8(32'hb737a49c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38153a71),
	.w1(32'h37b4251c),
	.w2(32'h3737345d),
	.w3(32'h37a53ff8),
	.w4(32'h37a6cca7),
	.w5(32'h37697a19),
	.w6(32'h373e6efd),
	.w7(32'h37946cbd),
	.w8(32'h376b9d57),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37212f3f),
	.w1(32'h36d294ca),
	.w2(32'hb6981e5b),
	.w3(32'h36e35c00),
	.w4(32'h363f7f65),
	.w5(32'hb7043207),
	.w6(32'hb65c01a6),
	.w7(32'hb724e9f7),
	.w8(32'hb78e6070),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a6699),
	.w1(32'h39e4f8a9),
	.w2(32'h39b432fa),
	.w3(32'hb9a7fa1c),
	.w4(32'h36e715c9),
	.w5(32'h3792a349),
	.w6(32'hba0884e4),
	.w7(32'hb9abbf22),
	.w8(32'hb919b85b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e137a5),
	.w1(32'h36fd5f4b),
	.w2(32'h36356714),
	.w3(32'h373a7e13),
	.w4(32'h373afd68),
	.w5(32'h369a7896),
	.w6(32'h36e092a5),
	.w7(32'h368b4347),
	.w8(32'h35c31c85),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82e1c0a),
	.w1(32'h3855aa55),
	.w2(32'h389ab49c),
	.w3(32'hb963a162),
	.w4(32'hb922fb46),
	.w5(32'h37a6e8a3),
	.w6(32'hb9b853eb),
	.w7(32'hb9a63641),
	.w8(32'hb93c696b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d4587f),
	.w1(32'h38f96b93),
	.w2(32'hba31778d),
	.w3(32'hb958c1cd),
	.w4(32'h381f1248),
	.w5(32'hba04f086),
	.w6(32'hb8d91c68),
	.w7(32'hb8e74044),
	.w8(32'h3827ae57),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h355124bb),
	.w1(32'h37534334),
	.w2(32'h378c978e),
	.w3(32'h36dbb5c5),
	.w4(32'h37865675),
	.w5(32'hb7591e3f),
	.w6(32'h370a0df8),
	.w7(32'h372a3896),
	.w8(32'hb716ef0a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb796ce24),
	.w1(32'hb7b8706f),
	.w2(32'hb81e7f1c),
	.w3(32'h37eb5113),
	.w4(32'h37fab0f0),
	.w5(32'h37df73c7),
	.w6(32'h37ba7c6a),
	.w7(32'h3780063a),
	.w8(32'h370c5d9d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34cc5087),
	.w1(32'hb685175f),
	.w2(32'hb6744e76),
	.w3(32'h3663b9da),
	.w4(32'hb5895ae0),
	.w5(32'hb61684cf),
	.w6(32'h36035264),
	.w7(32'hb462321d),
	.w8(32'hb64b85ad),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d141d8),
	.w1(32'hb8a7da3d),
	.w2(32'hb91ab314),
	.w3(32'hb7ce8e4b),
	.w4(32'hb9b28068),
	.w5(32'hb9dee2fe),
	.w6(32'hb90cd536),
	.w7(32'hb92138a3),
	.w8(32'hb8bca7d5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974be8b),
	.w1(32'h37fad199),
	.w2(32'hb9fb522b),
	.w3(32'h3846ecdb),
	.w4(32'h3982d8df),
	.w5(32'h3835f095),
	.w6(32'hb91492b8),
	.w7(32'hb9bbf51d),
	.w8(32'hb9b43ed7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b096c),
	.w1(32'h393f48e3),
	.w2(32'hb9bd6eb7),
	.w3(32'hb9eb7c40),
	.w4(32'h39b7a971),
	.w5(32'h39209436),
	.w6(32'hba8aa610),
	.w7(32'hba3a9c4f),
	.w8(32'hba58c833),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8179d07),
	.w1(32'hb9d13e4b),
	.w2(32'hb99c92d0),
	.w3(32'h3a650d41),
	.w4(32'hb97eaba5),
	.w5(32'hb988916c),
	.w6(32'hb9ea922a),
	.w7(32'hb9df7de7),
	.w8(32'hb9eaf60d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00b5d1),
	.w1(32'hb8f14bf7),
	.w2(32'h371462d6),
	.w3(32'hba2c673c),
	.w4(32'hb8e14f85),
	.w5(32'hb97b28ff),
	.w6(32'hb93b5f3c),
	.w7(32'hb900f5db),
	.w8(32'hb9910835),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9306320),
	.w1(32'hb9aba1e2),
	.w2(32'hba340d26),
	.w3(32'hba0a2629),
	.w4(32'hb963624e),
	.w5(32'h399dd694),
	.w6(32'h385d8d16),
	.w7(32'hb5b39ad8),
	.w8(32'hb9b53ca1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8c277),
	.w1(32'h3950a177),
	.w2(32'hb878dfc8),
	.w3(32'hba1cb83e),
	.w4(32'hb686dde2),
	.w5(32'hb96201c8),
	.w6(32'hb97c6e66),
	.w7(32'hb9f8686e),
	.w8(32'hb9d223ae),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e2802),
	.w1(32'h3a3d6d36),
	.w2(32'h3953dabc),
	.w3(32'h39127081),
	.w4(32'h39d92408),
	.w5(32'hb9636069),
	.w6(32'h39c26562),
	.w7(32'h3921053f),
	.w8(32'hb9db3c3b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a97a0),
	.w1(32'h38b7eb95),
	.w2(32'hba1430b4),
	.w3(32'hba1442d7),
	.w4(32'hb9e8f69e),
	.w5(32'hba609e06),
	.w6(32'hba53b590),
	.w7(32'hba816692),
	.w8(32'hba8533c5),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23e68e),
	.w1(32'h3957008a),
	.w2(32'h3944686f),
	.w3(32'hba937754),
	.w4(32'hb93faaaf),
	.w5(32'hb925b3c7),
	.w6(32'hb9cc29c6),
	.w7(32'hb958dd3c),
	.w8(32'h393be85b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3872c55a),
	.w1(32'h39c786ae),
	.w2(32'h397e2a0a),
	.w3(32'hb922fdae),
	.w4(32'hb93bc772),
	.w5(32'hb8bce46d),
	.w6(32'hba5c8883),
	.w7(32'hba1c0da4),
	.w8(32'hb9ba8352),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918ed75),
	.w1(32'h3a36115c),
	.w2(32'hb9415c0d),
	.w3(32'hb9a445d3),
	.w4(32'h399adbb9),
	.w5(32'hb9a4bde3),
	.w6(32'hb9d95df9),
	.w7(32'hb8b7c2e5),
	.w8(32'hba20e911),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be39f8),
	.w1(32'h39d6940f),
	.w2(32'h3a014787),
	.w3(32'hba26f6cc),
	.w4(32'hb91132f1),
	.w5(32'h39a8346e),
	.w6(32'hb99e8368),
	.w7(32'h383a2e02),
	.w8(32'h395d7817),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14c958),
	.w1(32'h3a0a1621),
	.w2(32'hb8540b07),
	.w3(32'hb8be4b8c),
	.w4(32'hb9825153),
	.w5(32'hb937db8c),
	.w6(32'hb7fa69b8),
	.w7(32'hb978f44b),
	.w8(32'hb82c730f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39835919),
	.w1(32'h38cfe492),
	.w2(32'h388f5ba6),
	.w3(32'hb8f7cdb6),
	.w4(32'hb77fb687),
	.w5(32'h390b3e5b),
	.w6(32'hb99233b1),
	.w7(32'hb8e6f0b5),
	.w8(32'hb752874f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398215e2),
	.w1(32'h3a26df4a),
	.w2(32'h39914b62),
	.w3(32'hb93700f6),
	.w4(32'hb89b3432),
	.w5(32'h37aa0a64),
	.w6(32'hb92e709d),
	.w7(32'h38197984),
	.w8(32'h3a39775c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59acb6),
	.w1(32'h38f055a4),
	.w2(32'hb995b9e6),
	.w3(32'h39cf5b65),
	.w4(32'h3897bd98),
	.w5(32'h39cf3339),
	.w6(32'h39aedb3d),
	.w7(32'hb8b94239),
	.w8(32'h399ccc9e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a024d50),
	.w1(32'h3944b3d4),
	.w2(32'h371f632a),
	.w3(32'hb8f0fd76),
	.w4(32'h389c447b),
	.w5(32'hb8f6b358),
	.w6(32'h38bd5b58),
	.w7(32'hb90f5793),
	.w8(32'hb8fe88f2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920066f),
	.w1(32'h39635b16),
	.w2(32'h39cc82c6),
	.w3(32'hb8e4cf1d),
	.w4(32'hb930ac32),
	.w5(32'hb9c2c6a2),
	.w6(32'h38076123),
	.w7(32'h38df2523),
	.w8(32'hb95401ea),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994a94e),
	.w1(32'hb8c13626),
	.w2(32'h38a3a666),
	.w3(32'hba184a68),
	.w4(32'hb954a47d),
	.w5(32'hb9519414),
	.w6(32'hb9273cef),
	.w7(32'hb992aaf8),
	.w8(32'hb98491c8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381de05a),
	.w1(32'hb8841420),
	.w2(32'h38305dba),
	.w3(32'hba83e92f),
	.w4(32'hb9fb9b8b),
	.w5(32'hb94891d4),
	.w6(32'hba45f9cb),
	.w7(32'hb9a5c41f),
	.w8(32'hb930c9c5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c0209),
	.w1(32'h3996bd1e),
	.w2(32'h3a19291d),
	.w3(32'hbacbc514),
	.w4(32'hb9a0bcac),
	.w5(32'hb9892df4),
	.w6(32'hba8479a9),
	.w7(32'hba0e76db),
	.w8(32'hb9a57013),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37341444),
	.w1(32'hb925d043),
	.w2(32'hb994d410),
	.w3(32'h389b5540),
	.w4(32'hb983b6a8),
	.w5(32'hb9c9ab16),
	.w6(32'h3843aaf1),
	.w7(32'hb90da830),
	.w8(32'h382e9a93),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88af575),
	.w1(32'h384f3777),
	.w2(32'hb9f92144),
	.w3(32'hba448aaa),
	.w4(32'h36f7e0cc),
	.w5(32'h39872ef2),
	.w6(32'hba30aac6),
	.w7(32'hb9bd8df0),
	.w8(32'hba5a23dc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87b2cd1),
	.w1(32'h3a0a313c),
	.w2(32'h39d1aee9),
	.w3(32'h3897675b),
	.w4(32'hb7a5002d),
	.w5(32'hb953538e),
	.w6(32'h385d4416),
	.w7(32'h39a28971),
	.w8(32'h3946489f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d1764d),
	.w1(32'h3928ff4b),
	.w2(32'h36ac0da8),
	.w3(32'hb981d0c5),
	.w4(32'hb7c4cc49),
	.w5(32'hb8b191cd),
	.w6(32'hba13dd44),
	.w7(32'hba244afa),
	.w8(32'hb9ce8a85),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a29189),
	.w1(32'h39dcb173),
	.w2(32'h3972c054),
	.w3(32'hb7e7e727),
	.w4(32'hb893de5f),
	.w5(32'hb9d7a5c6),
	.w6(32'hb99e0e50),
	.w7(32'hb9127cab),
	.w8(32'hb9396c6a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dadeb1),
	.w1(32'h39efa842),
	.w2(32'h39c011a0),
	.w3(32'hb9b7ce69),
	.w4(32'h3827b652),
	.w5(32'hb8c1d734),
	.w6(32'h39b406b2),
	.w7(32'h3a119f5d),
	.w8(32'h39dfeb42),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8076ec7),
	.w1(32'h37248951),
	.w2(32'hb8c283d5),
	.w3(32'hba1b1c07),
	.w4(32'hb8c9eb65),
	.w5(32'hb929a360),
	.w6(32'h38b4265e),
	.w7(32'h37a5493d),
	.w8(32'h391be8c1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d7904d),
	.w1(32'hb967de1f),
	.w2(32'hb8e2b7a7),
	.w3(32'hb9da5d3e),
	.w4(32'hb9852e14),
	.w5(32'h389aa28f),
	.w6(32'hba65a1c0),
	.w7(32'hb8e325bc),
	.w8(32'h39c678db),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947ff04),
	.w1(32'h38d5f5aa),
	.w2(32'h3a91b4d7),
	.w3(32'hb476f600),
	.w4(32'h39aa529a),
	.w5(32'h3a81aa57),
	.w6(32'hb7da3ecb),
	.w7(32'h3a3ee7b4),
	.w8(32'h3a98dad6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb846c1c4),
	.w1(32'hb89ae773),
	.w2(32'h397e508f),
	.w3(32'hb96861f5),
	.w4(32'hb9389b78),
	.w5(32'h37adb519),
	.w6(32'hb88f8e36),
	.w7(32'h38a1969f),
	.w8(32'h38fa2b50),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2302a),
	.w1(32'hb93995ff),
	.w2(32'hb9ad7bb6),
	.w3(32'hb95b93e3),
	.w4(32'hb922ed9a),
	.w5(32'hb9a37277),
	.w6(32'hb45a4be9),
	.w7(32'hb9654c5c),
	.w8(32'hb91a8f90),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924c3a0),
	.w1(32'h38eb9e86),
	.w2(32'hb55fc580),
	.w3(32'hb8a2db92),
	.w4(32'h370bc4fb),
	.w5(32'hb8b2cfa9),
	.w6(32'h398de4e3),
	.w7(32'h392ff65d),
	.w8(32'h391a967d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f86d78),
	.w1(32'h383aa19d),
	.w2(32'h39ec27cf),
	.w3(32'hb9765926),
	.w4(32'hb9138c06),
	.w5(32'hb9f88e37),
	.w6(32'hb9b2bf7d),
	.w7(32'hb8ccba0c),
	.w8(32'hb93c6897),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3764da80),
	.w1(32'h3a09b8b4),
	.w2(32'h3a1814c3),
	.w3(32'h38ebff9e),
	.w4(32'h399b155f),
	.w5(32'h3a1cf322),
	.w6(32'h39bb9e78),
	.w7(32'h3a2c5dd2),
	.w8(32'h389b9aa0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c73bf0),
	.w1(32'h38e3a74a),
	.w2(32'hb984ed25),
	.w3(32'hb973ea85),
	.w4(32'hb9048901),
	.w5(32'hb91a90d9),
	.w6(32'hb9fd8059),
	.w7(32'hb9eaf8e5),
	.w8(32'hb9c80173),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c690c),
	.w1(32'hb7f237dd),
	.w2(32'hb9159634),
	.w3(32'hba17601d),
	.w4(32'hb8e5820d),
	.w5(32'hb961c95f),
	.w6(32'h3916db09),
	.w7(32'h38a7087e),
	.w8(32'h3901c368),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3829b796),
	.w1(32'hb9cb8dda),
	.w2(32'hb97491d5),
	.w3(32'h39c0340e),
	.w4(32'hb93caaf9),
	.w5(32'hba3c4be1),
	.w6(32'h38d1d228),
	.w7(32'hb8e5f450),
	.w8(32'hb934eab8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f3ea7),
	.w1(32'hb951212e),
	.w2(32'hb91d4b6d),
	.w3(32'hb9b745d6),
	.w4(32'hb9559dd7),
	.w5(32'hb9c11a5c),
	.w6(32'hb968464d),
	.w7(32'hb9991a07),
	.w8(32'hb9fbb377),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03773c),
	.w1(32'hb923fb54),
	.w2(32'hb905097c),
	.w3(32'hba26ca90),
	.w4(32'hb9136ffa),
	.w5(32'hb948b54e),
	.w6(32'hb9094aa7),
	.w7(32'hb987712a),
	.w8(32'hb9194d0f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d3648),
	.w1(32'hb9b4b899),
	.w2(32'hb9887266),
	.w3(32'hba35188f),
	.w4(32'hba1cd9dd),
	.w5(32'hb9b68381),
	.w6(32'hba4f303f),
	.w7(32'hba0e81f9),
	.w8(32'hb8bdc645),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e6e534),
	.w1(32'h39dcd200),
	.w2(32'hb82e59cb),
	.w3(32'hb9f67e25),
	.w4(32'h39abc6cd),
	.w5(32'hb985678b),
	.w6(32'hb9e6175c),
	.w7(32'hb9ebc00c),
	.w8(32'hba3cb5da),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa0901),
	.w1(32'hb9589f7d),
	.w2(32'hb92b785b),
	.w3(32'hb98a3a74),
	.w4(32'hb8bfd2b4),
	.w5(32'hb797e726),
	.w6(32'h394797b5),
	.w7(32'h38e27309),
	.w8(32'h38a8e9b8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397eecc5),
	.w1(32'h3a1ee65c),
	.w2(32'h3a123a92),
	.w3(32'hb9db6c4f),
	.w4(32'h382db1dd),
	.w5(32'h387d8c8b),
	.w6(32'hb9248faf),
	.w7(32'h38adde6c),
	.w8(32'h3904da38),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6c2fa),
	.w1(32'h399413a9),
	.w2(32'hb7f687c9),
	.w3(32'hb9359533),
	.w4(32'h39c25857),
	.w5(32'h388c5321),
	.w6(32'h39a23dbb),
	.w7(32'h39185e83),
	.w8(32'hb92b3cd2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b5e03),
	.w1(32'h3a718e32),
	.w2(32'h3aa76f87),
	.w3(32'hba0cd3fb),
	.w4(32'h39c87909),
	.w5(32'h3a3c8fd5),
	.w6(32'hbab84e9e),
	.w7(32'h37d78652),
	.w8(32'h399bf27d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a71a7c),
	.w1(32'h390f7078),
	.w2(32'hb8ceec1a),
	.w3(32'hb7f89cd0),
	.w4(32'h39916a76),
	.w5(32'h398e19d4),
	.w6(32'hba0410b5),
	.w7(32'hb8e6ad68),
	.w8(32'h38fbe901),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f2d1a),
	.w1(32'hb91a4cc0),
	.w2(32'hba7a20d0),
	.w3(32'hb967abd2),
	.w4(32'hb9ea9be9),
	.w5(32'hb9811191),
	.w6(32'hba55ed38),
	.w7(32'hba7732e2),
	.w8(32'hba6ad410),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986051b),
	.w1(32'h399b5d82),
	.w2(32'h3a467753),
	.w3(32'hb98b0887),
	.w4(32'h379cc63f),
	.w5(32'h3963c442),
	.w6(32'h39295f90),
	.w7(32'h39e8c5f5),
	.w8(32'h390b6a8a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6368d6),
	.w1(32'h3a294c76),
	.w2(32'h39c8c4a4),
	.w3(32'h390af5c9),
	.w4(32'h39669bed),
	.w5(32'h38f2a7c5),
	.w6(32'h36ee1e69),
	.w7(32'h38cb7cc4),
	.w8(32'hb833b62e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a22a8),
	.w1(32'hb936cb6c),
	.w2(32'hb7e16e78),
	.w3(32'hb8c6774b),
	.w4(32'hb8acfb66),
	.w5(32'hb8a09e7a),
	.w6(32'hb96fca03),
	.w7(32'hb96250c8),
	.w8(32'h35f43b1f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a8732d),
	.w1(32'h389a0c18),
	.w2(32'hb939da66),
	.w3(32'hb690dc21),
	.w4(32'h376b7ef4),
	.w5(32'hba1a79f6),
	.w6(32'h398c806f),
	.w7(32'hb8cae501),
	.w8(32'hb98433d6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382d0d23),
	.w1(32'h38bf28e1),
	.w2(32'hb98a763c),
	.w3(32'h38fd422c),
	.w4(32'hb909090f),
	.w5(32'h396844c0),
	.w6(32'hb8ae5410),
	.w7(32'hb7d8fd34),
	.w8(32'hb9854146),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381a791b),
	.w1(32'h3a045552),
	.w2(32'h398e54c5),
	.w3(32'h3a25690c),
	.w4(32'h3a09199d),
	.w5(32'h38f2ca93),
	.w6(32'hb928c765),
	.w7(32'hb9b80ace),
	.w8(32'hb9274f6f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971219b),
	.w1(32'hb9626c3e),
	.w2(32'hb79a8cca),
	.w3(32'hb9bdd2ad),
	.w4(32'hb8d51ed5),
	.w5(32'hb8f55f42),
	.w6(32'hb86e549a),
	.w7(32'hb97f0eda),
	.w8(32'hb9b32182),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98256a1),
	.w1(32'hb9a38de8),
	.w2(32'hb9a888ac),
	.w3(32'hb7d4b919),
	.w4(32'hb947283f),
	.w5(32'hb995f856),
	.w6(32'hb99a11bb),
	.w7(32'hb99d1cf5),
	.w8(32'hb98c10ab),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e22ebc),
	.w1(32'h38aee462),
	.w2(32'h39521791),
	.w3(32'hba174370),
	.w4(32'h3928bf4f),
	.w5(32'h39319c49),
	.w6(32'h3895b372),
	.w7(32'h387f3447),
	.w8(32'h3985bd6e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92438ed),
	.w1(32'h3a946eb3),
	.w2(32'h3a13cfe7),
	.w3(32'h3874e2a0),
	.w4(32'h3a2b12f7),
	.w5(32'h386f3141),
	.w6(32'h3806b62a),
	.w7(32'h39b31635),
	.w8(32'h39c0736c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2de24),
	.w1(32'h39f97496),
	.w2(32'hb9945399),
	.w3(32'h398bf63d),
	.w4(32'h38ae5cf8),
	.w5(32'hb973edb3),
	.w6(32'h39828c21),
	.w7(32'hb93ebfef),
	.w8(32'hb9c4c528),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d39571),
	.w1(32'hba0d1bb7),
	.w2(32'hb9e8511d),
	.w3(32'hb956a2c7),
	.w4(32'hb9cf8904),
	.w5(32'hb9f37164),
	.w6(32'hba037f43),
	.w7(32'hb9a5e211),
	.w8(32'hb9f0842c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eefa9),
	.w1(32'h3a7fcb1f),
	.w2(32'h3afd29c9),
	.w3(32'hbb1eca97),
	.w4(32'hba59c605),
	.w5(32'hba3fa626),
	.w6(32'hbb2f5308),
	.w7(32'hbaa99b97),
	.w8(32'hba263c99),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0d60d),
	.w1(32'hb895c65a),
	.w2(32'h3a0b3ed9),
	.w3(32'hba105c86),
	.w4(32'hb8a6c7ec),
	.w5(32'h399effa1),
	.w6(32'hba63e16d),
	.w7(32'hb95d3244),
	.w8(32'h38bebd30),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17e3db),
	.w1(32'hb976f844),
	.w2(32'hb8f79684),
	.w3(32'hba4dc6de),
	.w4(32'hb9073999),
	.w5(32'hb7f69370),
	.w6(32'hb96f4ee4),
	.w7(32'hb90a5c3a),
	.w8(32'h38425da8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379fa177),
	.w1(32'hb90b86c5),
	.w2(32'h391e84e9),
	.w3(32'h391b4ad6),
	.w4(32'hb947fb7a),
	.w5(32'hb9ba840b),
	.w6(32'h3892f066),
	.w7(32'h391b895b),
	.w8(32'hb9c1a370),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8296093),
	.w1(32'h38beee89),
	.w2(32'hb8fb31a2),
	.w3(32'h39355e68),
	.w4(32'h3968b9af),
	.w5(32'h38121d23),
	.w6(32'h394dd646),
	.w7(32'h388eb0ee),
	.w8(32'hb900a9ff),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93243e7),
	.w1(32'hb9ef9330),
	.w2(32'hb982dea3),
	.w3(32'hb8dff5c5),
	.w4(32'hb9a29cfb),
	.w5(32'hb93ac0e4),
	.w6(32'hb9afc77b),
	.w7(32'hb91da7fc),
	.w8(32'hb9794e50),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cd41a8),
	.w1(32'h39a0d6b1),
	.w2(32'hb92ea456),
	.w3(32'hb998d51f),
	.w4(32'hb6e1b474),
	.w5(32'hb9187edb),
	.w6(32'hb85c225c),
	.w7(32'hb8e1e7c6),
	.w8(32'hb99dc370),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae0764),
	.w1(32'h3a8132f9),
	.w2(32'h3a4a7ae7),
	.w3(32'h39b093ae),
	.w4(32'h39a310ab),
	.w5(32'h3923379b),
	.w6(32'hba1fa85a),
	.w7(32'hb9d44605),
	.w8(32'hb9d6fd57),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8c65c),
	.w1(32'h3a09a496),
	.w2(32'h3a3a99e9),
	.w3(32'hba96c36a),
	.w4(32'hb9ceafd3),
	.w5(32'hb99acbff),
	.w6(32'hba2eb8e8),
	.w7(32'hb8b9b432),
	.w8(32'h3922a12a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ebffad),
	.w1(32'h390db9c7),
	.w2(32'h38aa3d5e),
	.w3(32'hb9b72a34),
	.w4(32'h38ea605b),
	.w5(32'hb8c45501),
	.w6(32'h3898ae3b),
	.w7(32'hb8b0147c),
	.w8(32'h3749127c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cc18b),
	.w1(32'h3a601379),
	.w2(32'h3a3eae31),
	.w3(32'hba5af24f),
	.w4(32'h38ced05c),
	.w5(32'hb8f0103f),
	.w6(32'hb9bb895c),
	.w7(32'h38427b6a),
	.w8(32'h39cd8a57),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d37f5),
	.w1(32'hb95ce389),
	.w2(32'h3897bdb1),
	.w3(32'h3a156244),
	.w4(32'hb8c882a7),
	.w5(32'h38137ce3),
	.w6(32'hb9127e91),
	.w7(32'hb98dce5b),
	.w8(32'hb8a60fa0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4b19d),
	.w1(32'hb90331e3),
	.w2(32'hb7f7d441),
	.w3(32'hba0bc5a3),
	.w4(32'hb8895dc6),
	.w5(32'hb8694c21),
	.w6(32'hb89303ac),
	.w7(32'hb8fdc822),
	.w8(32'hb84d277b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82461e7),
	.w1(32'hb93a10be),
	.w2(32'hb91b0bd0),
	.w3(32'hb75580b0),
	.w4(32'hb8e207a0),
	.w5(32'hb94fe182),
	.w6(32'hb8a78308),
	.w7(32'hb9688762),
	.w8(32'hb9149414),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ca713a),
	.w1(32'h38a7b6f1),
	.w2(32'hb88ac3ee),
	.w3(32'hb915d150),
	.w4(32'h36859cd4),
	.w5(32'hb91bef8d),
	.w6(32'h39579613),
	.w7(32'h38d27f68),
	.w8(32'h390befef),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7986c94),
	.w1(32'hb9f9299a),
	.w2(32'hba65e729),
	.w3(32'hb9d5f67a),
	.w4(32'hba09f115),
	.w5(32'hba446087),
	.w6(32'hba7d74e6),
	.w7(32'hba72e84e),
	.w8(32'hb96c2b8c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7461bb),
	.w1(32'hb9ea523c),
	.w2(32'h390f6c59),
	.w3(32'hba191815),
	.w4(32'h390f5957),
	.w5(32'h3a9b8be4),
	.w6(32'h3815061c),
	.w7(32'h3968fdc7),
	.w8(32'h3a7ca5ea),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8c6d9),
	.w1(32'h39f09f2b),
	.w2(32'h39fe89ca),
	.w3(32'hba2ceffb),
	.w4(32'h37626e09),
	.w5(32'h38b502c1),
	.w6(32'hb904a03a),
	.w7(32'h382e490c),
	.w8(32'h3a0902e6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a97f3e),
	.w1(32'hb9d520cd),
	.w2(32'h385dd018),
	.w3(32'h38a12669),
	.w4(32'hb98ddae1),
	.w5(32'hb8a864f6),
	.w6(32'hb994fc67),
	.w7(32'hb87ada06),
	.w8(32'hb8cefbb2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c428a),
	.w1(32'h3a068b5c),
	.w2(32'h39b22b5d),
	.w3(32'hba7ce444),
	.w4(32'hb94c34c1),
	.w5(32'hb8b908c9),
	.w6(32'hb9fffc70),
	.w7(32'hb97f4208),
	.w8(32'h399c01fc),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8af6876),
	.w1(32'h34e5f552),
	.w2(32'hb9102c62),
	.w3(32'hba1fef87),
	.w4(32'hb9caac5c),
	.w5(32'hb9e8356f),
	.w6(32'hba02894b),
	.w7(32'hba208d74),
	.w8(32'hb9c5bdd6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb6bd4),
	.w1(32'h3a25cd29),
	.w2(32'h3a241888),
	.w3(32'hba162892),
	.w4(32'hb8634d22),
	.w5(32'hb9c1fef7),
	.w6(32'hba951d76),
	.w7(32'hb99d94ed),
	.w8(32'hb93621db),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3869317a),
	.w1(32'hb9009052),
	.w2(32'hb7bd9272),
	.w3(32'h36d13c07),
	.w4(32'hb8ae9be5),
	.w5(32'h376c68a2),
	.w6(32'hb940494f),
	.w7(32'hb90919db),
	.w8(32'h381b24cb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b62aa5),
	.w1(32'h38b73965),
	.w2(32'h391c1fed),
	.w3(32'h37d7fb54),
	.w4(32'h386dd1e5),
	.w5(32'hb8ee4a93),
	.w6(32'h3899d03f),
	.w7(32'h38f5bf93),
	.w8(32'h3847a32d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9185d0f),
	.w1(32'hb999a77b),
	.w2(32'hb8dd2edf),
	.w3(32'hb9475baf),
	.w4(32'hb90996a9),
	.w5(32'hb945ce3c),
	.w6(32'hb9f2ac9f),
	.w7(32'hb8b58d88),
	.w8(32'h3892ccca),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e0553),
	.w1(32'h3a356c19),
	.w2(32'h39a45a6a),
	.w3(32'hb9e56c1b),
	.w4(32'hb7c701b2),
	.w5(32'hb9b4f7cf),
	.w6(32'hba14e5cb),
	.w7(32'hb81f7779),
	.w8(32'hb9aaded9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39feaf8b),
	.w1(32'h39dc1c66),
	.w2(32'h3a16bc09),
	.w3(32'hb8f259ac),
	.w4(32'hb81725ef),
	.w5(32'h38cce6f1),
	.w6(32'hba3ddabc),
	.w7(32'hb99a0ba7),
	.w8(32'hb787f475),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389721b7),
	.w1(32'hb7c4d11e),
	.w2(32'h3953a9e8),
	.w3(32'hb7686999),
	.w4(32'h38d6a2dc),
	.w5(32'h39d9ed42),
	.w6(32'h396a70f0),
	.w7(32'h3959459a),
	.w8(32'h39a0cd8e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f705ff),
	.w1(32'hb8a5ae10),
	.w2(32'hb91703f8),
	.w3(32'h39fb83c7),
	.w4(32'hb8d1d3bb),
	.w5(32'hb932ee11),
	.w6(32'h37da6662),
	.w7(32'hb8e46d5d),
	.w8(32'h3824a861),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e9c533),
	.w1(32'hb9980131),
	.w2(32'hb97f9637),
	.w3(32'hb803b3c9),
	.w4(32'hb9639c6d),
	.w5(32'hb989b5fa),
	.w6(32'hb98da8e8),
	.w7(32'hb97a0e97),
	.w8(32'hb985e463),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9075b),
	.w1(32'hb812310a),
	.w2(32'hba0b8a8e),
	.w3(32'hba0ba448),
	.w4(32'hb8eb59c9),
	.w5(32'hba03f3e3),
	.w6(32'h398bdfc1),
	.w7(32'hb8f6ff60),
	.w8(32'hb86c4004),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c8838),
	.w1(32'h38560944),
	.w2(32'h3a864e31),
	.w3(32'hbadccefe),
	.w4(32'hba97fc82),
	.w5(32'hb9ca46f1),
	.w6(32'hbadfbff5),
	.w7(32'hba43fffe),
	.w8(32'h392f77bb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec8db4),
	.w1(32'h3a33c0ac),
	.w2(32'hb8afe7b7),
	.w3(32'hb9593e3b),
	.w4(32'h387c19bd),
	.w5(32'hb9e9cb70),
	.w6(32'h383a35d2),
	.w7(32'hb9d8fa10),
	.w8(32'hba262721),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba063cee),
	.w1(32'hb99c36cb),
	.w2(32'h36690360),
	.w3(32'hba16e3f5),
	.w4(32'h37a1e34f),
	.w5(32'h39988b6f),
	.w6(32'hb8f6e6b4),
	.w7(32'h3994cbd2),
	.w8(32'h3a1343db),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96cfbf7),
	.w1(32'h3922c89e),
	.w2(32'h39686e71),
	.w3(32'hb9dd41fd),
	.w4(32'h380fd326),
	.w5(32'h389f2bc4),
	.w6(32'h39a4d88a),
	.w7(32'h39f3becd),
	.w8(32'h3a6d72d9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3870a4ba),
	.w1(32'hb9290601),
	.w2(32'h3878d86c),
	.w3(32'hb8224f33),
	.w4(32'hb980563f),
	.w5(32'hb907402d),
	.w6(32'hb97071aa),
	.w7(32'hb91b6e4e),
	.w8(32'hb9b3033e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918f913),
	.w1(32'hb8ca2c84),
	.w2(32'hb9a06ee6),
	.w3(32'hb9c25975),
	.w4(32'h391ddaea),
	.w5(32'h39965841),
	.w6(32'h38d8fdb7),
	.w7(32'hb8cd70e8),
	.w8(32'hb9d1e598),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980d095),
	.w1(32'h398a9acb),
	.w2(32'h39c916f3),
	.w3(32'h398086f4),
	.w4(32'h38a81bf2),
	.w5(32'h39277cb7),
	.w6(32'h39bdee4d),
	.w7(32'h39b45474),
	.w8(32'h3959e443),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a5531),
	.w1(32'h37621f6e),
	.w2(32'h38a78ea0),
	.w3(32'hb8cf5d4b),
	.w4(32'hb708b9e4),
	.w5(32'h391ba3ce),
	.w6(32'hb950d8c0),
	.w7(32'h393e7a81),
	.w8(32'hb90b1c90),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d45fd),
	.w1(32'hba01b362),
	.w2(32'hb9db6de8),
	.w3(32'hb7d5faf9),
	.w4(32'hb9b69024),
	.w5(32'hb98d7c8c),
	.w6(32'hba069970),
	.w7(32'hb9e095c9),
	.w8(32'hb9c724c8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ac610),
	.w1(32'h399c06f2),
	.w2(32'h38760dcd),
	.w3(32'hba3f6df7),
	.w4(32'h3901195d),
	.w5(32'hb8c7cf8a),
	.w6(32'hb9fb8528),
	.w7(32'hba1165f0),
	.w8(32'hb8b0d6fa),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e5d5e6),
	.w1(32'h3a94bbe9),
	.w2(32'h37d701c6),
	.w3(32'hba02244b),
	.w4(32'hb893a7e1),
	.w5(32'hb94f583a),
	.w6(32'h39014a00),
	.w7(32'hb9c74d5b),
	.w8(32'hba0e6a39),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab0f52),
	.w1(32'hb8b1ab5f),
	.w2(32'hba410aa9),
	.w3(32'hb7090a8f),
	.w4(32'hb89b2f61),
	.w5(32'hb96c0d03),
	.w6(32'hb86f8a5f),
	.w7(32'hb9cbf55d),
	.w8(32'hb9bc280e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1df3d),
	.w1(32'h3a2f48a7),
	.w2(32'h393dd58a),
	.w3(32'h3836e68a),
	.w4(32'h3973ad7f),
	.w5(32'hb8fd172a),
	.w6(32'h38511421),
	.w7(32'hb9678d18),
	.w8(32'h386651fb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb6239),
	.w1(32'h3889f2bc),
	.w2(32'hb912dc16),
	.w3(32'h39a2f6c1),
	.w4(32'hb8fc153e),
	.w5(32'hb9d1b450),
	.w6(32'hb908396e),
	.w7(32'hb99e031f),
	.w8(32'hb9eb93a7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88dac6a),
	.w1(32'h390d4321),
	.w2(32'h38a2f670),
	.w3(32'hb8b61767),
	.w4(32'h38c4a218),
	.w5(32'h36a95d54),
	.w6(32'h39269160),
	.w7(32'h380b5dc4),
	.w8(32'h392533d4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ebe44c),
	.w1(32'h3865b7e9),
	.w2(32'hb8e02f97),
	.w3(32'h38e6529b),
	.w4(32'hb95983df),
	.w5(32'hb9b6888c),
	.w6(32'hb9930631),
	.w7(32'hb995b2d7),
	.w8(32'hb9204085),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f3f214),
	.w1(32'hb9a21b1b),
	.w2(32'hb8aac9c2),
	.w3(32'hb8efef0f),
	.w4(32'hb9ce16d6),
	.w5(32'hb9cbcc2f),
	.w6(32'hb99325af),
	.w7(32'hb91454c9),
	.w8(32'hb9b34e4b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9721c38),
	.w1(32'hb8d3dd29),
	.w2(32'hb93c565e),
	.w3(32'hb9f6362f),
	.w4(32'hb92526a3),
	.w5(32'hb95cfb1a),
	.w6(32'h38dd3cfb),
	.w7(32'hb8accad5),
	.w8(32'h38cf6e7b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86c5c27),
	.w1(32'h394c688d),
	.w2(32'h3908f556),
	.w3(32'hb89997ac),
	.w4(32'h391904a3),
	.w5(32'h3812d5e8),
	.w6(32'h394a97f0),
	.w7(32'h38a9d729),
	.w8(32'h39356f66),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d212c),
	.w1(32'hb9970121),
	.w2(32'h399c00c3),
	.w3(32'h392df2de),
	.w4(32'h3921dd17),
	.w5(32'h396c7a8b),
	.w6(32'hb8d44095),
	.w7(32'h3935bdd4),
	.w8(32'hb951c577),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9853cef),
	.w1(32'hb8128f41),
	.w2(32'hb95b640a),
	.w3(32'hb93cbf21),
	.w4(32'hb8e55b8a),
	.w5(32'hb92c7123),
	.w6(32'hb90b1d50),
	.w7(32'hb957f25d),
	.w8(32'h37a7edfe),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b476c2),
	.w1(32'h39a39ea4),
	.w2(32'hb8d7b768),
	.w3(32'hb95702c7),
	.w4(32'h3960b79f),
	.w5(32'h39537d15),
	.w6(32'hba5cbb21),
	.w7(32'hb9ec49e9),
	.w8(32'hba091905),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48ee89),
	.w1(32'h3a0a38c7),
	.w2(32'h399233cc),
	.w3(32'h3a6c07af),
	.w4(32'h3947cd06),
	.w5(32'hb7807bd6),
	.w6(32'hb9ba1c12),
	.w7(32'hb9376a2f),
	.w8(32'hb8b85d19),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c41c57),
	.w1(32'hb92bbab1),
	.w2(32'h3931dd16),
	.w3(32'hb9f300ab),
	.w4(32'hb9910bec),
	.w5(32'hb8a9112f),
	.w6(32'hba8b6a61),
	.w7(32'hba25e734),
	.w8(32'hba4cfa3c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96742ea),
	.w1(32'hb8977cc3),
	.w2(32'h3831e238),
	.w3(32'hb9f25c0e),
	.w4(32'hb87f371b),
	.w5(32'hb8eb3b5b),
	.w6(32'hb8b28069),
	.w7(32'h37f6fa7c),
	.w8(32'h35cc487f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c539e6),
	.w1(32'h3981022a),
	.w2(32'h3922ba02),
	.w3(32'hb8a89281),
	.w4(32'h39435490),
	.w5(32'h3817de9e),
	.w6(32'h398a7ffa),
	.w7(32'h38c5d1d0),
	.w8(32'h3980dcc1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39631f92),
	.w1(32'h38d51bb0),
	.w2(32'h380dfc76),
	.w3(32'h398222bc),
	.w4(32'h37c3d938),
	.w5(32'hb8c3b586),
	.w6(32'h38841cbd),
	.w7(32'hb79bfece),
	.w8(32'h37c7599d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73244be),
	.w1(32'h38a2a600),
	.w2(32'hb7988f67),
	.w3(32'hb8e4868d),
	.w4(32'hb71165c4),
	.w5(32'hb90b04b0),
	.w6(32'h386afb91),
	.w7(32'hb8b222e9),
	.w8(32'h37ea7a50),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f4038),
	.w1(32'h3a11cccb),
	.w2(32'hb9247f49),
	.w3(32'hb9b654cf),
	.w4(32'h393b37d6),
	.w5(32'h388300ce),
	.w6(32'hb9b55d87),
	.w7(32'hb80a0635),
	.w8(32'hb900db0e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c12665),
	.w1(32'hb9b8236c),
	.w2(32'hba1a05f2),
	.w3(32'h39fd0034),
	.w4(32'hb9b82966),
	.w5(32'hba2dfa48),
	.w6(32'hb9e18a56),
	.w7(32'hba0d5dc1),
	.w8(32'hba5a72ec),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93155b),
	.w1(32'h3866323b),
	.w2(32'hb8901c24),
	.w3(32'hba68f808),
	.w4(32'h38826254),
	.w5(32'hb70f201e),
	.w6(32'h3a017d87),
	.w7(32'h39262470),
	.w8(32'h39944100),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807a9bd),
	.w1(32'hb848af47),
	.w2(32'h36655a2f),
	.w3(32'h389f0445),
	.w4(32'h38d843c6),
	.w5(32'h38e44f8b),
	.w6(32'h37095e25),
	.w7(32'hb83041b2),
	.w8(32'h39bd0137),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39785d4f),
	.w1(32'hb8e863ba),
	.w2(32'hb8e5a423),
	.w3(32'h39b76829),
	.w4(32'hb902c133),
	.w5(32'hb9449d69),
	.w6(32'hb9253d08),
	.w7(32'hb9653206),
	.w8(32'hb8a64764),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97fa0ef),
	.w1(32'hb98b5c42),
	.w2(32'hba68652f),
	.w3(32'hb9a64720),
	.w4(32'h3763136d),
	.w5(32'hb97d2ba6),
	.w6(32'hb9a72cac),
	.w7(32'h38f283a0),
	.w8(32'hb9b0235c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56cfc9),
	.w1(32'h39726187),
	.w2(32'h393c53f5),
	.w3(32'h3820046c),
	.w4(32'h39801ad3),
	.w5(32'h38fafd64),
	.w6(32'h39cbf246),
	.w7(32'h388796ec),
	.w8(32'hb7b7a49e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f5ba42),
	.w1(32'hb8a6fe44),
	.w2(32'hb9e716ba),
	.w3(32'hb9465802),
	.w4(32'hb8d65ece),
	.w5(32'hb9cc54dc),
	.w6(32'hba1961ab),
	.w7(32'hb9d6be86),
	.w8(32'hb8da4584),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fd40a9),
	.w1(32'hb97dcc71),
	.w2(32'h37d00b14),
	.w3(32'h38e17d97),
	.w4(32'h377f02ee),
	.w5(32'hb72db14c),
	.w6(32'hb8d3cabc),
	.w7(32'h388e7f98),
	.w8(32'h389be374),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c33ee),
	.w1(32'hb90e52fa),
	.w2(32'hb938d079),
	.w3(32'hb8375e6b),
	.w4(32'h39a81a35),
	.w5(32'h3a2bd462),
	.w6(32'h37550f54),
	.w7(32'h38e92e0b),
	.w8(32'h398ef198),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule