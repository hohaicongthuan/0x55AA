module layer_8_featuremap_116(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e4004),
	.w1(32'h3c4b1c90),
	.w2(32'h3c1b18c7),
	.w3(32'hbbd299f6),
	.w4(32'h3cbe142a),
	.w5(32'hbbe2fff9),
	.w6(32'h3b288a6f),
	.w7(32'h3cbcb1c7),
	.w8(32'hbc841b34),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5c360),
	.w1(32'h3c9ac617),
	.w2(32'hbb7e16a1),
	.w3(32'h3becb1a6),
	.w4(32'hbbcd894d),
	.w5(32'hbc93c25c),
	.w6(32'h3ca11878),
	.w7(32'hb9074fd4),
	.w8(32'h3c10d019),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4fad8),
	.w1(32'hbc21e47f),
	.w2(32'hbaddc148),
	.w3(32'hba9006cb),
	.w4(32'hbc86f73f),
	.w5(32'hbac6d6b4),
	.w6(32'h3b99b45c),
	.w7(32'hbbb674dc),
	.w8(32'hbccdcd79),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87ba0a),
	.w1(32'h3cb6e235),
	.w2(32'h3c39116c),
	.w3(32'hbc7feca0),
	.w4(32'h3c15531c),
	.w5(32'hbc293002),
	.w6(32'h3c7d0859),
	.w7(32'h3c2bf64e),
	.w8(32'hbd157ff8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b74fa),
	.w1(32'h3cba8b96),
	.w2(32'hbadb7099),
	.w3(32'h3cac15ea),
	.w4(32'h3a3961c6),
	.w5(32'h3be80c3f),
	.w6(32'h3d01ee1b),
	.w7(32'hbc094e7f),
	.w8(32'hbbcb1997),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78c838),
	.w1(32'h3bdc2510),
	.w2(32'hb98ee738),
	.w3(32'hbb3e53e7),
	.w4(32'h3c4b05cb),
	.w5(32'hbbf08bed),
	.w6(32'hbbc3f816),
	.w7(32'h3c3d5f9f),
	.w8(32'hbc42a8ba),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d7b64e),
	.w1(32'hbb117131),
	.w2(32'h3c88ed90),
	.w3(32'hbb6e1915),
	.w4(32'h3c5916d5),
	.w5(32'h3a430889),
	.w6(32'hbc2cc847),
	.w7(32'h3c981e1c),
	.w8(32'hbc3aeae1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b7f7),
	.w1(32'h3c4c3851),
	.w2(32'hbc276ee3),
	.w3(32'h3cd61959),
	.w4(32'h3bfea272),
	.w5(32'h3c2bd5ab),
	.w6(32'h3c9df6a7),
	.w7(32'hbbee3548),
	.w8(32'h3bdace62),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15fbc2),
	.w1(32'hbc55bdb7),
	.w2(32'h3b94aa30),
	.w3(32'hbc1fe366),
	.w4(32'hbc1fdf3e),
	.w5(32'hbb558ef2),
	.w6(32'hbcb461d3),
	.w7(32'hbb7adaac),
	.w8(32'hbb2eeefd),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bc67e),
	.w1(32'hba83d2eb),
	.w2(32'hbb490ec6),
	.w3(32'h3a9274a2),
	.w4(32'hbc290fbd),
	.w5(32'h3c086bc3),
	.w6(32'h3c0f2459),
	.w7(32'hbbc480a1),
	.w8(32'hbcb411fa),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce4feec),
	.w1(32'h3c80609a),
	.w2(32'hbb91ec00),
	.w3(32'h3c9d2f04),
	.w4(32'hbc070451),
	.w5(32'h3c7668db),
	.w6(32'h3c8f9e58),
	.w7(32'hbbb482d1),
	.w8(32'h3ca676d9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb86205),
	.w1(32'hbbdb907e),
	.w2(32'h3b1f9d9f),
	.w3(32'hbb9271d8),
	.w4(32'h3b45aeb9),
	.w5(32'h3bce73ad),
	.w6(32'hbafc7649),
	.w7(32'h3c0321d1),
	.w8(32'h3cd7a198),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d005e65),
	.w1(32'hbb3e9f78),
	.w2(32'h3aee6ded),
	.w3(32'hbaf599d8),
	.w4(32'hb9d5900f),
	.w5(32'hb9838154),
	.w6(32'h3bafa15a),
	.w7(32'h3a94bc2c),
	.w8(32'h3bf34660),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9d4f5),
	.w1(32'h3ada4cff),
	.w2(32'hbba32740),
	.w3(32'hbad6ba9a),
	.w4(32'hbbab4f17),
	.w5(32'hbb94415b),
	.w6(32'h39aeaa5a),
	.w7(32'h398c111a),
	.w8(32'hba88d2ec),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe12304),
	.w1(32'hbb5d9fc9),
	.w2(32'hbbe5e918),
	.w3(32'hbc27cfd0),
	.w4(32'hbbc7e23f),
	.w5(32'hbb8ee603),
	.w6(32'hbac5c6ab),
	.w7(32'hbb84f713),
	.w8(32'hbb416bbe),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81eb28),
	.w1(32'hbbc13d43),
	.w2(32'h3c0036fe),
	.w3(32'hbc1fd2c6),
	.w4(32'hbb5679c8),
	.w5(32'h3be49e31),
	.w6(32'hbb8664fe),
	.w7(32'hbc155734),
	.w8(32'h3bcb24c6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b9a2f),
	.w1(32'h3c48c897),
	.w2(32'hba2bd79c),
	.w3(32'h3bbf3c03),
	.w4(32'h3b37ff57),
	.w5(32'hba965317),
	.w6(32'hbbdde509),
	.w7(32'hbc3c95d8),
	.w8(32'hbc9a0df5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89ea04),
	.w1(32'hbb5752ab),
	.w2(32'hba2c2f6e),
	.w3(32'hbb366e11),
	.w4(32'h3ca59efc),
	.w5(32'h3c23ae82),
	.w6(32'hbc0eae9b),
	.w7(32'h3bb0280b),
	.w8(32'h3cb1f34a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0d40f),
	.w1(32'h393ff8cc),
	.w2(32'h3c51d5b4),
	.w3(32'hbc462676),
	.w4(32'h3c1149e1),
	.w5(32'h3c57be5c),
	.w6(32'h3bfba64f),
	.w7(32'h3a503202),
	.w8(32'h3c43890d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70bcbc),
	.w1(32'h3b1c884c),
	.w2(32'h3aff5034),
	.w3(32'h3c8b695e),
	.w4(32'h3a4fcbee),
	.w5(32'h3c7c55f8),
	.w6(32'h3c1c0ac3),
	.w7(32'h3c0f88c1),
	.w8(32'h3b79a248),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb3170),
	.w1(32'hbadc239a),
	.w2(32'h3b777b06),
	.w3(32'hbba2cbca),
	.w4(32'h3c2cbc0d),
	.w5(32'hbb476117),
	.w6(32'h3c5a2df6),
	.w7(32'h3bc7a938),
	.w8(32'hbd03e601),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b947cae),
	.w1(32'hbbf4c788),
	.w2(32'h3bd59424),
	.w3(32'hbc0c44fa),
	.w4(32'hbb4c2ca1),
	.w5(32'hbc39b911),
	.w6(32'hbc5e8f1d),
	.w7(32'h3c6279e7),
	.w8(32'h3a761dc2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca49224),
	.w1(32'hbc0df71b),
	.w2(32'h3bbe391c),
	.w3(32'h3bae0e0e),
	.w4(32'hbb73d102),
	.w5(32'hbb9221dc),
	.w6(32'hbced0d6f),
	.w7(32'hbb0ee736),
	.w8(32'hbc4c5c3d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72bce3),
	.w1(32'h3c6085ea),
	.w2(32'hbb4f6e3b),
	.w3(32'h3ba3d1ed),
	.w4(32'hbb180d02),
	.w5(32'h3b036c8e),
	.w6(32'h3c2b48f4),
	.w7(32'h3ae35992),
	.w8(32'h3a8b91eb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae36e59),
	.w1(32'h39536d0e),
	.w2(32'h3bfe1bfd),
	.w3(32'hba2a6327),
	.w4(32'hbb33b58e),
	.w5(32'hbb27a365),
	.w6(32'hbb7e8637),
	.w7(32'h3b91d4dd),
	.w8(32'h3bacfb1c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fd7a0),
	.w1(32'hbbb8fac6),
	.w2(32'h3b7a702f),
	.w3(32'hbc8115d1),
	.w4(32'h3bc13231),
	.w5(32'h3b3ccfc8),
	.w6(32'hbc2a7306),
	.w7(32'h3c3f71c5),
	.w8(32'hbc70df7e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b26cd),
	.w1(32'hbb69835b),
	.w2(32'h3bda4a98),
	.w3(32'h3ae79c88),
	.w4(32'hbc3d6a5f),
	.w5(32'h3b9fd178),
	.w6(32'h3b2f940f),
	.w7(32'hbb7ef7c4),
	.w8(32'hbcaa5c66),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a3a38),
	.w1(32'h3b1e2e87),
	.w2(32'hbca0a730),
	.w3(32'hbbe3cb25),
	.w4(32'hbcd91f24),
	.w5(32'hbd140945),
	.w6(32'hbc808742),
	.w7(32'hbd01778c),
	.w8(32'hbd28a048),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb4234b),
	.w1(32'hbccd35d1),
	.w2(32'hbbd7a51d),
	.w3(32'hbcad96b0),
	.w4(32'h3c1192d0),
	.w5(32'h3c81c6f5),
	.w6(32'hbce84292),
	.w7(32'h3acc53de),
	.w8(32'h3c85c336),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf3243c),
	.w1(32'hbc230446),
	.w2(32'h3b1320fc),
	.w3(32'hbc02c4ac),
	.w4(32'h3b6fc4ef),
	.w5(32'hbc818c8e),
	.w6(32'hbbfce7e6),
	.w7(32'h3acc50c4),
	.w8(32'hbbbd4498),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77b86),
	.w1(32'hbc1a596e),
	.w2(32'hbb96251d),
	.w3(32'hbc7689fc),
	.w4(32'hbb9ba78e),
	.w5(32'hbb6a89bc),
	.w6(32'h3a306dd8),
	.w7(32'hbb91dfc8),
	.w8(32'hbb928979),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9449ea),
	.w1(32'hbb11fde5),
	.w2(32'hbc0b3b1c),
	.w3(32'hba684dcc),
	.w4(32'hbc8b5c2d),
	.w5(32'hbc34a112),
	.w6(32'hba263ee2),
	.w7(32'hbccb8294),
	.w8(32'h3c9b9c75),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2fa14),
	.w1(32'hbbbbe438),
	.w2(32'h3c058a57),
	.w3(32'hbc4347ac),
	.w4(32'h3bcc4681),
	.w5(32'hbc03acd8),
	.w6(32'hbcca711a),
	.w7(32'h3b066980),
	.w8(32'hbd0083db),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47fe96),
	.w1(32'h3b8353bf),
	.w2(32'h3bb6c22c),
	.w3(32'h3b6c156e),
	.w4(32'h3bf512da),
	.w5(32'h3c9427c1),
	.w6(32'hba9ecead),
	.w7(32'h3c01b822),
	.w8(32'hbb0b5957),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a7703),
	.w1(32'h3b510e59),
	.w2(32'h389e6f38),
	.w3(32'h3c104eaa),
	.w4(32'h3adbf54a),
	.w5(32'hbc161512),
	.w6(32'hbb17f96a),
	.w7(32'h3ba541b4),
	.w8(32'hbc12187e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cc3ab),
	.w1(32'h3b54d4f7),
	.w2(32'hbbc8ee8a),
	.w3(32'h3bfc70d7),
	.w4(32'hbb972422),
	.w5(32'hbca39749),
	.w6(32'h3c23bb50),
	.w7(32'hba152756),
	.w8(32'hbc8fa224),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70ee3f),
	.w1(32'hbc412b45),
	.w2(32'hbb99206c),
	.w3(32'hbbe4415f),
	.w4(32'hbcb605f9),
	.w5(32'hbcd975b3),
	.w6(32'hbbd3e657),
	.w7(32'hbc8e4830),
	.w8(32'hbd182ff2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b460383),
	.w1(32'hbcccd2ff),
	.w2(32'hbc55c06a),
	.w3(32'hbc9732d2),
	.w4(32'hbc351181),
	.w5(32'hbb825aa5),
	.w6(32'hbd1d620f),
	.w7(32'hbcb1c1ec),
	.w8(32'hbc0da4c1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34f3cd),
	.w1(32'hb9cef5d2),
	.w2(32'h3bee4774),
	.w3(32'hbabe9d5c),
	.w4(32'hbae293e8),
	.w5(32'hba1cf757),
	.w6(32'hbc01e7bd),
	.w7(32'hbb1322ae),
	.w8(32'h3c790f30),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeeead2),
	.w1(32'hbc0fcbea),
	.w2(32'h3bb5d4fd),
	.w3(32'hbc180ed6),
	.w4(32'hbba5dcf8),
	.w5(32'hbb876cb4),
	.w6(32'hbb1f80f7),
	.w7(32'hbb7c36d3),
	.w8(32'hbb44fcae),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c9d68),
	.w1(32'h3be9679e),
	.w2(32'hbba46033),
	.w3(32'hb9ca6e7c),
	.w4(32'hbbd6dd4d),
	.w5(32'h3ca58e90),
	.w6(32'hbb1fa507),
	.w7(32'hbb6b7e21),
	.w8(32'h3c633373),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc391),
	.w1(32'hb9935c5c),
	.w2(32'hbc1ee0dd),
	.w3(32'h3a8e400c),
	.w4(32'hbc6b8ac2),
	.w5(32'hbc0e5b49),
	.w6(32'hbc683ed0),
	.w7(32'hbc8b3bac),
	.w8(32'hbc2d55f9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2923d7),
	.w1(32'hbca5c629),
	.w2(32'h3c372933),
	.w3(32'hbc9a0424),
	.w4(32'h3c02b902),
	.w5(32'h3b3af8fa),
	.w6(32'hbcb408c3),
	.w7(32'h3c4c61ca),
	.w8(32'hbc8d0d57),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7879f6),
	.w1(32'h3bd2b0ca),
	.w2(32'h3a7d5f14),
	.w3(32'h3b23db5b),
	.w4(32'hba4c4e62),
	.w5(32'hba8152bc),
	.w6(32'hbb36802f),
	.w7(32'h38a710c9),
	.w8(32'h3b922786),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5db9a4),
	.w1(32'hba7b9e5f),
	.w2(32'h3ad0a77a),
	.w3(32'hbb1938ad),
	.w4(32'hbbacf9a6),
	.w5(32'h3bf6c656),
	.w6(32'hbaddf720),
	.w7(32'h3c16d13b),
	.w8(32'h3d17ead4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b3356),
	.w1(32'hbc41c94d),
	.w2(32'h3b7980b0),
	.w3(32'hbc2f1cd8),
	.w4(32'h3c1bce98),
	.w5(32'hbc303f19),
	.w6(32'hbba82aa6),
	.w7(32'hbb008604),
	.w8(32'hbc76ffcd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1153d),
	.w1(32'hba6ef037),
	.w2(32'hbc7bcfa9),
	.w3(32'hbb203d40),
	.w4(32'hbc350fa4),
	.w5(32'hbab71627),
	.w6(32'h3bd3afd3),
	.w7(32'hbbc3be64),
	.w8(32'h3cabbe9a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5ac59),
	.w1(32'hbc18806e),
	.w2(32'h3c1780a5),
	.w3(32'hbca93837),
	.w4(32'hbb432b70),
	.w5(32'h3c883a13),
	.w6(32'hbc0a60ba),
	.w7(32'h3bc6f7a2),
	.w8(32'h3c13b985),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8cac4),
	.w1(32'h3b30c11b),
	.w2(32'hbc4c69ec),
	.w3(32'h3af718e3),
	.w4(32'hba84d8ba),
	.w5(32'hbb0f358b),
	.w6(32'h3b1e23ab),
	.w7(32'hbaa009e0),
	.w8(32'h3d1fdfe1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a6562),
	.w1(32'hbc0ce86d),
	.w2(32'hbb8e2a57),
	.w3(32'hbc182343),
	.w4(32'hbc807397),
	.w5(32'h3c5e4f82),
	.w6(32'hbba044d5),
	.w7(32'hbb986098),
	.w8(32'h3d50c5c2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e3300),
	.w1(32'hbc7ac86a),
	.w2(32'h3bdf0aa5),
	.w3(32'hbce5a128),
	.w4(32'h3c5a2ab4),
	.w5(32'h3cc81af4),
	.w6(32'hbcd79a4b),
	.w7(32'h3ceb084b),
	.w8(32'h3a7a3bdf),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3580a1),
	.w1(32'h3bbcfae9),
	.w2(32'hbb637a12),
	.w3(32'h3bf43340),
	.w4(32'hbc544752),
	.w5(32'hbc50928a),
	.w6(32'h3c69e621),
	.w7(32'hb9e92f06),
	.w8(32'hbc8e0af7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b972189),
	.w1(32'hbc17267d),
	.w2(32'hbb3ec998),
	.w3(32'hbc683ed0),
	.w4(32'h3c045a7d),
	.w5(32'hbbdd9c0c),
	.w6(32'hbc693c64),
	.w7(32'hbad2a2fb),
	.w8(32'h3d0e0872),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba77c49),
	.w1(32'h3bfc13ec),
	.w2(32'hbac807bc),
	.w3(32'h3b4a8b7b),
	.w4(32'hbbcb1a21),
	.w5(32'hbb6bfd0f),
	.w6(32'h3c544570),
	.w7(32'hba87d4f2),
	.w8(32'h3be661af),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b002705),
	.w1(32'h3a627eea),
	.w2(32'h3c245fcb),
	.w3(32'hbb311376),
	.w4(32'h3bc0060e),
	.w5(32'h3c4dfdc4),
	.w6(32'h3a7311a6),
	.w7(32'hbad892be),
	.w8(32'hba26ad5c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c758533),
	.w1(32'h3b946819),
	.w2(32'h3c1b9601),
	.w3(32'h3b0dc385),
	.w4(32'h3b58b3fc),
	.w5(32'hbc10fa94),
	.w6(32'h3c11ab66),
	.w7(32'h3c246d90),
	.w8(32'hbbc379bc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68661a),
	.w1(32'h3a724e26),
	.w2(32'hbbabea56),
	.w3(32'h3bd1096c),
	.w4(32'hbc6aa820),
	.w5(32'h3a2cc77f),
	.w6(32'hbbe30d53),
	.w7(32'hbc3c26a2),
	.w8(32'h3a97df7e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4ab03),
	.w1(32'hbac41dea),
	.w2(32'h3c9fcc78),
	.w3(32'hbc118a7f),
	.w4(32'h3c7357d1),
	.w5(32'h3c272d44),
	.w6(32'hbbf52c74),
	.w7(32'h3c3ef588),
	.w8(32'hbca5cde2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b39b6),
	.w1(32'h3ba6fa61),
	.w2(32'hbab1148d),
	.w3(32'h3c221f17),
	.w4(32'hbb51b17e),
	.w5(32'hbae62ce8),
	.w6(32'h3c730d8d),
	.w7(32'hbad470c9),
	.w8(32'h3b89c131),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cdc08),
	.w1(32'h3afdabb5),
	.w2(32'h3c10a9df),
	.w3(32'hb9be8bda),
	.w4(32'h3bc37f51),
	.w5(32'hbc98baf2),
	.w6(32'h39ed2c85),
	.w7(32'h3c5e206a),
	.w8(32'hba1d7cb5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2708),
	.w1(32'hbb163f42),
	.w2(32'hba85804d),
	.w3(32'hbc11a68f),
	.w4(32'h3b89efb7),
	.w5(32'h3c27d918),
	.w6(32'h3b809597),
	.w7(32'h3ca83b39),
	.w8(32'hbbd6e06f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9c284),
	.w1(32'h3bb06a28),
	.w2(32'h3a208207),
	.w3(32'hbafaef40),
	.w4(32'hbb5d2f86),
	.w5(32'h3a49ed62),
	.w6(32'h3b3f7faf),
	.w7(32'hbb96816a),
	.w8(32'h3a3bc4ad),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf96b05),
	.w1(32'hbb0586f8),
	.w2(32'h3caa4963),
	.w3(32'hbb84d7c6),
	.w4(32'h3c8a23f7),
	.w5(32'h3cfb2a71),
	.w6(32'hbc01f7b3),
	.w7(32'h3c8a0545),
	.w8(32'h3d53dbbb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c892873),
	.w1(32'h3c0b7533),
	.w2(32'h3a8ec80b),
	.w3(32'h3b8fb42d),
	.w4(32'h3ae120d7),
	.w5(32'hbc8e824c),
	.w6(32'hbbc4ba1a),
	.w7(32'h3c75c7c3),
	.w8(32'h3cbd8cf2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc746a98),
	.w1(32'hbc819016),
	.w2(32'hbc23b302),
	.w3(32'hbb7c37e4),
	.w4(32'hbc957277),
	.w5(32'hbc215a2e),
	.w6(32'h38869ae6),
	.w7(32'hbc8c45a4),
	.w8(32'hbb17a8cd),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c648d4d),
	.w1(32'hbbe0bea8),
	.w2(32'h3a7cb40e),
	.w3(32'hbc433e4e),
	.w4(32'h3c11be85),
	.w5(32'h3cc2929e),
	.w6(32'hbc868080),
	.w7(32'hba4908c6),
	.w8(32'h3bb7c309),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c566027),
	.w1(32'h3b3b9e28),
	.w2(32'h3c865c82),
	.w3(32'hbb1082fb),
	.w4(32'h3c4df035),
	.w5(32'h3cb9530c),
	.w6(32'hbbdc6f18),
	.w7(32'h3bdbf625),
	.w8(32'h3bb096c1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb544277),
	.w1(32'h3c2289a6),
	.w2(32'hb9032ae2),
	.w3(32'h3c218089),
	.w4(32'hbba54248),
	.w5(32'hbc69e5b4),
	.w6(32'h3cf3d60e),
	.w7(32'hbc7c866b),
	.w8(32'hbc806696),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35b089),
	.w1(32'hbbae8272),
	.w2(32'hbb0e1582),
	.w3(32'hbc7c8334),
	.w4(32'hbc81913d),
	.w5(32'hbb3e7a62),
	.w6(32'hbc04d5b1),
	.w7(32'hbb9d75ed),
	.w8(32'h3cbee4eb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb092c),
	.w1(32'hbc935144),
	.w2(32'hbc2398f9),
	.w3(32'hbc22f446),
	.w4(32'h3c197b21),
	.w5(32'h3cacd80a),
	.w6(32'hbc8ca2df),
	.w7(32'h3c6c85e6),
	.w8(32'h3d0b1f3d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5562f3),
	.w1(32'hbb7b0422),
	.w2(32'hbc8dcc5f),
	.w3(32'hbc8d869d),
	.w4(32'hbc99a5a2),
	.w5(32'h3cb4a5f1),
	.w6(32'h3bb9608c),
	.w7(32'hbc025aec),
	.w8(32'h3ce3fcfe),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e8637),
	.w1(32'hbc9ff5e6),
	.w2(32'h3b9dfbf1),
	.w3(32'hbca5f356),
	.w4(32'h3b5b2326),
	.w5(32'h3c101a58),
	.w6(32'hbc764b8a),
	.w7(32'h3c8d542b),
	.w8(32'h3cc6419b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b046e),
	.w1(32'h3c8c4c3f),
	.w2(32'hbbd45df9),
	.w3(32'h3ca6366a),
	.w4(32'hbbb93ca0),
	.w5(32'hbbb5503a),
	.w6(32'hbb2dccb1),
	.w7(32'hbc54b6e0),
	.w8(32'hbaf271c3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45fd45),
	.w1(32'hba2f498f),
	.w2(32'hbac0ce53),
	.w3(32'hbbd74075),
	.w4(32'h3c0e54be),
	.w5(32'h3aef6b90),
	.w6(32'hbc5511f9),
	.w7(32'h3ba693af),
	.w8(32'hbae74791),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81980e),
	.w1(32'hbae4dbb9),
	.w2(32'hbc419e1f),
	.w3(32'hbc848dd4),
	.w4(32'hbc0e4aca),
	.w5(32'hbaa837cd),
	.w6(32'h3bb0b0fe),
	.w7(32'hbcbbd5a8),
	.w8(32'h3c3b4f88),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef2cbc),
	.w1(32'hbb77f830),
	.w2(32'h3b10554c),
	.w3(32'hbbf86422),
	.w4(32'h3c5afedb),
	.w5(32'hbb7d78f2),
	.w6(32'hbaf0875e),
	.w7(32'h3cde267d),
	.w8(32'h3c3272c9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9a2f),
	.w1(32'h3bb1c49f),
	.w2(32'h367015a6),
	.w3(32'h3ab2c557),
	.w4(32'h373359df),
	.w5(32'h36cac0f0),
	.w6(32'hbb9e68dd),
	.w7(32'hb6991bdc),
	.w8(32'h369a212f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08665a),
	.w1(32'hbafde814),
	.w2(32'hba63757e),
	.w3(32'hba13cccc),
	.w4(32'hb9afc3d6),
	.w5(32'h3a05f866),
	.w6(32'hb98c18db),
	.w7(32'hba6f79f5),
	.w8(32'hb9863cfb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f3587),
	.w1(32'hba037784),
	.w2(32'h39ddfbca),
	.w3(32'h38fcee2d),
	.w4(32'hba0269b6),
	.w5(32'h3920d530),
	.w6(32'hb8f85a1e),
	.w7(32'h39733ebe),
	.w8(32'h3a2e2e09),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57a5855),
	.w1(32'h3533d740),
	.w2(32'h373649bb),
	.w3(32'hb639227d),
	.w4(32'hb5fc5f2c),
	.w5(32'hb78d0c80),
	.w6(32'hb51ca586),
	.w7(32'hb78d78bf),
	.w8(32'hb6b13b33),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361ee97c),
	.w1(32'hb8046e97),
	.w2(32'h372bcd0c),
	.w3(32'hb8105345),
	.w4(32'hb81dd323),
	.w5(32'hb835f73e),
	.w6(32'h354f88ad),
	.w7(32'hb72c9770),
	.w8(32'hb7a98be5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05905d),
	.w1(32'hba672ee5),
	.w2(32'hb9411636),
	.w3(32'hba52d619),
	.w4(32'hbaa958b1),
	.w5(32'hba04f4ab),
	.w6(32'h3990c939),
	.w7(32'hb9aca0d7),
	.w8(32'h39ac515e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2d123),
	.w1(32'hba659543),
	.w2(32'hb776179a),
	.w3(32'hb907d4c9),
	.w4(32'h36f26899),
	.w5(32'h3a5c6140),
	.w6(32'hb8c87e11),
	.w7(32'hb9570fdf),
	.w8(32'h399f7c6d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b1763),
	.w1(32'h3bd0dbef),
	.w2(32'h3bc7eb49),
	.w3(32'h3ba33dcb),
	.w4(32'h3bde3ebb),
	.w5(32'h3baf5dda),
	.w6(32'h3b33107a),
	.w7(32'h3b6b6e71),
	.w8(32'h3bee778e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f3eea),
	.w1(32'hbb2dc67f),
	.w2(32'hba5f957f),
	.w3(32'hba2104ca),
	.w4(32'hba92c8c2),
	.w5(32'h39a14f7b),
	.w6(32'hba726675),
	.w7(32'hbae4c77c),
	.w8(32'h3a0f55f5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a9b14),
	.w1(32'hba29c66c),
	.w2(32'h39c51cc9),
	.w3(32'hba05add7),
	.w4(32'hba2addfd),
	.w5(32'h397c015d),
	.w6(32'h39414a28),
	.w7(32'hb9beb83b),
	.w8(32'h3a2f2b27),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69d33a9),
	.w1(32'h37cbb174),
	.w2(32'h37351845),
	.w3(32'h3864c177),
	.w4(32'hb65df244),
	.w5(32'hb68467de),
	.w6(32'h35928f88),
	.w7(32'h370e7dd5),
	.w8(32'h35d8f312),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37403fb2),
	.w1(32'hb6ae991d),
	.w2(32'hb7c65f7d),
	.w3(32'hb715b3ab),
	.w4(32'hb33b577e),
	.w5(32'h36b953ca),
	.w6(32'hb7c06db4),
	.w7(32'hb77af2fc),
	.w8(32'hb53eef1b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72f8775),
	.w1(32'hb6cc9b97),
	.w2(32'hb683a55c),
	.w3(32'hb52f2bfc),
	.w4(32'hb712067f),
	.w5(32'h378dd922),
	.w6(32'hb56862fe),
	.w7(32'h3746940a),
	.w8(32'h3782b1c2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb781cd0d),
	.w1(32'hb8012a78),
	.w2(32'hb859d38e),
	.w3(32'h3691b75d),
	.w4(32'hb8cfbb7e),
	.w5(32'hb62c80fd),
	.w6(32'hb689f6f8),
	.w7(32'h38885dc4),
	.w8(32'h322522b0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d6f83),
	.w1(32'h3a5fd46e),
	.w2(32'h3a325339),
	.w3(32'h3a2e1edd),
	.w4(32'h3a1494a5),
	.w5(32'h39b2e4c8),
	.w6(32'h3a3d7132),
	.w7(32'h3a66d94d),
	.w8(32'h3a34000a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881533b),
	.w1(32'h382ca8c6),
	.w2(32'h3823ff4b),
	.w3(32'h3863378f),
	.w4(32'h3730b75b),
	.w5(32'h382e2893),
	.w6(32'hb69b25a4),
	.w7(32'h38768a82),
	.w8(32'h385d1637),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4dab5),
	.w1(32'h38d50900),
	.w2(32'hb916a197),
	.w3(32'hb99eed6b),
	.w4(32'hb80aa9ee),
	.w5(32'h3914f2dd),
	.w6(32'h37731dba),
	.w7(32'h3857ab39),
	.w8(32'h3a08041f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d053d),
	.w1(32'hba000c94),
	.w2(32'hb7c7c282),
	.w3(32'hb9ae3a6e),
	.w4(32'hb95a7fb1),
	.w5(32'h391a5743),
	.w6(32'hb98b2510),
	.w7(32'hb98f2ce8),
	.w8(32'h39066020),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97d1c98),
	.w1(32'h3954ab7c),
	.w2(32'h39c49a91),
	.w3(32'hb8420151),
	.w4(32'h3820724c),
	.w5(32'h3963e8a4),
	.w6(32'hb7e30410),
	.w7(32'h399956c1),
	.w8(32'h39d5f14b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79a680),
	.w1(32'hba32265a),
	.w2(32'h3888ba43),
	.w3(32'hb96014b9),
	.w4(32'h389b5fd6),
	.w5(32'h395aa432),
	.w6(32'hb9a1fe97),
	.w7(32'hb9e61238),
	.w8(32'h39c4dda6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ace225),
	.w1(32'h390498ea),
	.w2(32'h3a27cd3c),
	.w3(32'h388017eb),
	.w4(32'h3935d702),
	.w5(32'h3a416063),
	.w6(32'hb8260911),
	.w7(32'hb85c85c6),
	.w8(32'h3a1478cb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb702ec00),
	.w1(32'h369a176d),
	.w2(32'h380eb739),
	.w3(32'h38277e85),
	.w4(32'hb7a9b03e),
	.w5(32'hb78bfb68),
	.w6(32'h3759ed7b),
	.w7(32'h35e5b9e0),
	.w8(32'hb73d472e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37826221),
	.w1(32'h3722c1b8),
	.w2(32'hb77ef994),
	.w3(32'hb751b19a),
	.w4(32'hb72ad11d),
	.w5(32'hb7758e07),
	.w6(32'hb827cc46),
	.w7(32'h343dea2d),
	.w8(32'h36f27d4d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d4b803),
	.w1(32'hb79a727a),
	.w2(32'hb809063e),
	.w3(32'hb7f7a647),
	.w4(32'hb71ff65a),
	.w5(32'hb7f4aeda),
	.w6(32'hb5952b09),
	.w7(32'hb7052775),
	.w8(32'hb725a9f6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33ef97f6),
	.w1(32'h37cfc99f),
	.w2(32'hb708476e),
	.w3(32'h375d7952),
	.w4(32'h36a848f5),
	.w5(32'hb68371e2),
	.w6(32'h37471ae5),
	.w7(32'hb6edb2ee),
	.w8(32'hb7aed406),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382bda35),
	.w1(32'h383cc403),
	.w2(32'h38c6ddee),
	.w3(32'h3906b9bb),
	.w4(32'h3889eb86),
	.w5(32'h388aa0cf),
	.w6(32'hb7c6bd1c),
	.w7(32'h37be6cc2),
	.w8(32'h38eeae94),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b157ab),
	.w1(32'hb6cecdfb),
	.w2(32'h37c58d76),
	.w3(32'hb7833cb0),
	.w4(32'h37f48e74),
	.w5(32'hb6c019bb),
	.w6(32'hb646f654),
	.w7(32'h354fc8d8),
	.w8(32'h37980476),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397558b4),
	.w1(32'h3947cc98),
	.w2(32'h37e4746c),
	.w3(32'hba287233),
	.w4(32'hb99e3071),
	.w5(32'h38d98cde),
	.w6(32'h39790e83),
	.w7(32'h393b003a),
	.w8(32'h3a2f277b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c4d7df),
	.w1(32'h3900598a),
	.w2(32'h37540ccb),
	.w3(32'h38a21281),
	.w4(32'h38d798af),
	.w5(32'hb83e7bda),
	.w6(32'h39280b98),
	.w7(32'h390d24f2),
	.w8(32'h383a5d99),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb28d6),
	.w1(32'hbb1b641a),
	.w2(32'hbab271ad),
	.w3(32'hb9c90996),
	.w4(32'hba92efb7),
	.w5(32'hb9cb712b),
	.w6(32'hba00d32d),
	.w7(32'hba8b9231),
	.w8(32'hb95bc7af),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379ce5f5),
	.w1(32'h37e247b3),
	.w2(32'h38804f0e),
	.w3(32'h37abd9d3),
	.w4(32'h38eea72d),
	.w5(32'h357ae471),
	.w6(32'hb8539e33),
	.w7(32'hb7e84235),
	.w8(32'h3822f6c5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cdd339),
	.w1(32'hb8f0d510),
	.w2(32'hb96dc191),
	.w3(32'hb9389b77),
	.w4(32'hb8e30bf9),
	.w5(32'hb9546bb9),
	.w6(32'h3884ada4),
	.w7(32'hb8c36fcc),
	.w8(32'hb8c5d3fe),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936b57e),
	.w1(32'h3934c0fe),
	.w2(32'h38c10672),
	.w3(32'h39166097),
	.w4(32'h39183530),
	.w5(32'h3840c768),
	.w6(32'h397e1f76),
	.w7(32'h39548003),
	.w8(32'h38f6bed2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38523f48),
	.w1(32'h36ff4d64),
	.w2(32'h3711df4f),
	.w3(32'h375ffe8a),
	.w4(32'h38da2ea8),
	.w5(32'hb754119d),
	.w6(32'h375e408b),
	.w7(32'h3841b74c),
	.w8(32'h38111be2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb811b427),
	.w1(32'h39309aa2),
	.w2(32'h39bc14c2),
	.w3(32'h3967ecf8),
	.w4(32'h39d995f1),
	.w5(32'h39c94f24),
	.w6(32'h37ba251c),
	.w7(32'h399dba58),
	.w8(32'h39ceff9f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3809933b),
	.w1(32'h397c2d16),
	.w2(32'h39924160),
	.w3(32'h3966a5d9),
	.w4(32'h39faa814),
	.w5(32'h3a06d1f6),
	.w6(32'hb7c68fc4),
	.w7(32'hb82073a6),
	.w8(32'h377af032),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d595d1),
	.w1(32'hb9a0beed),
	.w2(32'hb9b93404),
	.w3(32'hb9bbfa39),
	.w4(32'hb9c79ed2),
	.w5(32'hb9a938b7),
	.w6(32'hb931cb65),
	.w7(32'hb91c8d29),
	.w8(32'hb985e89c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885b4f6),
	.w1(32'h38cc8e77),
	.w2(32'h38060a8d),
	.w3(32'h38cc0ad8),
	.w4(32'h3839a304),
	.w5(32'h37e8d9d1),
	.w6(32'h382d68a5),
	.w7(32'h38035a63),
	.w8(32'h3801feb9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d50dc4),
	.w1(32'hb9d4d3e1),
	.w2(32'hb9d308dd),
	.w3(32'hb8effeda),
	.w4(32'hb970da9d),
	.w5(32'h38b5b6ba),
	.w6(32'hb8896adb),
	.w7(32'hb9b4a98c),
	.w8(32'h39131a48),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a19d85),
	.w1(32'h36a7b8f0),
	.w2(32'hb6b1f097),
	.w3(32'h387f41f1),
	.w4(32'hb78d3cb8),
	.w5(32'hb770c1ba),
	.w6(32'hb820b3db),
	.w7(32'hb7fc131c),
	.w8(32'hb798d9e9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0f400),
	.w1(32'h37cc28da),
	.w2(32'h3846afca),
	.w3(32'h391e6f69),
	.w4(32'h38441340),
	.w5(32'h3884f895),
	.w6(32'h37bcc271),
	.w7(32'hb8632788),
	.w8(32'h38564906),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e9b4b),
	.w1(32'hba2b5d5b),
	.w2(32'h376f7f08),
	.w3(32'hb8a05c5a),
	.w4(32'hb8edb920),
	.w5(32'h39d76253),
	.w6(32'hb8577f94),
	.w7(32'hb980f498),
	.w8(32'hb823eb1e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb1744f70),
	.w1(32'hb67fed54),
	.w2(32'hb7c3937f),
	.w3(32'hb6cc5022),
	.w4(32'hb43fb850),
	.w5(32'hb77726a6),
	.w6(32'hb634e5e3),
	.w7(32'hb78f96a3),
	.w8(32'hb3b79032),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91de81d),
	.w1(32'hb80d7807),
	.w2(32'h386b1035),
	.w3(32'h37148dd2),
	.w4(32'h37cf77f1),
	.w5(32'h3865ef8f),
	.w6(32'hb814ed56),
	.w7(32'h38034f5b),
	.w8(32'h388671d7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a298b37),
	.w1(32'h3a4ba963),
	.w2(32'h3a633708),
	.w3(32'hb7dc41be),
	.w4(32'h390f625b),
	.w5(32'h3995ed62),
	.w6(32'h39b4d51a),
	.w7(32'h3a90ef49),
	.w8(32'h3ab91268),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380df4da),
	.w1(32'h3895b682),
	.w2(32'hb8a9187b),
	.w3(32'h387c4302),
	.w4(32'h38bc5a93),
	.w5(32'hb726598e),
	.w6(32'hb5f0b04b),
	.w7(32'hb8468424),
	.w8(32'hb8a4e652),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3795a4a9),
	.w1(32'h381d4d44),
	.w2(32'h379439e6),
	.w3(32'hb5e35420),
	.w4(32'h38024d82),
	.w5(32'h3730c0c8),
	.w6(32'h3796ad2b),
	.w7(32'h37a79a8c),
	.w8(32'h3763db00),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e6f5ef),
	.w1(32'hb6c4d24b),
	.w2(32'hb7e324e0),
	.w3(32'hb717fbb2),
	.w4(32'hb86292ad),
	.w5(32'h3587cf9e),
	.w6(32'hb6da9642),
	.w7(32'h379cc170),
	.w8(32'hb887a799),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376b5a53),
	.w1(32'hb7e796b3),
	.w2(32'hb80ca194),
	.w3(32'hb7f16967),
	.w4(32'hb86ca957),
	.w5(32'hb7eaa576),
	.w6(32'h36ef9d34),
	.w7(32'hb7d773b9),
	.w8(32'hb8848103),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d09e7),
	.w1(32'hb9cd6d6e),
	.w2(32'hb9100dfe),
	.w3(32'hb9af84e5),
	.w4(32'hb8572aec),
	.w5(32'h3962a7c7),
	.w6(32'hb853bf66),
	.w7(32'h38a1d1e3),
	.w8(32'h398d2027),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952b4a5),
	.w1(32'hb88f5b1c),
	.w2(32'h399c19bc),
	.w3(32'hb83237ed),
	.w4(32'hb81a0424),
	.w5(32'h390029aa),
	.w6(32'hb900e954),
	.w7(32'h3949c7b9),
	.w8(32'h398fcb25),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba492c28),
	.w1(32'hba316f6d),
	.w2(32'hb9fc54f9),
	.w3(32'hb9dfb8b8),
	.w4(32'hb9861fc7),
	.w5(32'hb7af99b5),
	.w6(32'hb9078221),
	.w7(32'hb9acee39),
	.w8(32'h38782784),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule