module layer_8_featuremap_82(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacee723),
	.w1(32'hbb027ac6),
	.w2(32'hbacc42fe),
	.w3(32'h3ad070f8),
	.w4(32'hbb0bf9c9),
	.w5(32'hbba6335c),
	.w6(32'hbb304020),
	.w7(32'h3abf49f3),
	.w8(32'hbb23e825),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b45f0),
	.w1(32'h3ab0dabe),
	.w2(32'h3ad6054b),
	.w3(32'hb84f0463),
	.w4(32'h3ac8c5cd),
	.w5(32'hbae3e4ac),
	.w6(32'hbae583fc),
	.w7(32'h3a60e11d),
	.w8(32'hba804570),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa59497),
	.w1(32'h3adc192d),
	.w2(32'h3b084177),
	.w3(32'h3a8d0364),
	.w4(32'h3aa36e9e),
	.w5(32'hba768b0c),
	.w6(32'h3a546ca2),
	.w7(32'h3b1213d3),
	.w8(32'h3c5d19c1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90d12),
	.w1(32'h3c3fe6c2),
	.w2(32'h3c270bb4),
	.w3(32'hbc71d22e),
	.w4(32'h3bd87603),
	.w5(32'h3c081968),
	.w6(32'h3bd29baf),
	.w7(32'hbbcfdccd),
	.w8(32'hbaa76ea7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ec35),
	.w1(32'hbae5a487),
	.w2(32'h3a3ee925),
	.w3(32'hbb12f0d3),
	.w4(32'hba285117),
	.w5(32'hbb84e87f),
	.w6(32'hbb42a08e),
	.w7(32'hb9c1a0d5),
	.w8(32'hbcb09571),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabd3a1),
	.w1(32'h3bcf0257),
	.w2(32'h3cdee6e9),
	.w3(32'hbb5ee7ca),
	.w4(32'h3c73e947),
	.w5(32'h3c426762),
	.w6(32'hbc912bfc),
	.w7(32'hbaaf6bd5),
	.w8(32'hba981623),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae18d8a),
	.w1(32'hba6684e9),
	.w2(32'h3b1c691f),
	.w3(32'h3ad8f10b),
	.w4(32'h3a97c1b6),
	.w5(32'hbb9a6ff5),
	.w6(32'h3b0697d6),
	.w7(32'h3bd80996),
	.w8(32'hb9c6a6eb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5089f),
	.w1(32'hbb81865b),
	.w2(32'h38cf4f78),
	.w3(32'hbafb0022),
	.w4(32'h3a1054b7),
	.w5(32'hbb6095f7),
	.w6(32'hbb266310),
	.w7(32'hba06397c),
	.w8(32'hbad43a78),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbcebd),
	.w1(32'h3a48643a),
	.w2(32'h39900c2a),
	.w3(32'h3b1651b9),
	.w4(32'hb88fb9b8),
	.w5(32'hbbf4d6c9),
	.w6(32'h3acc1365),
	.w7(32'h3b8730fc),
	.w8(32'h3c7fc782),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce31dcb),
	.w1(32'hbc71de58),
	.w2(32'hbca4c245),
	.w3(32'hbc2355f7),
	.w4(32'h3ce877d9),
	.w5(32'h3c98470a),
	.w6(32'h3d1735f2),
	.w7(32'hbbfb4eb0),
	.w8(32'h3b87f48f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a84dc),
	.w1(32'h3aca22d1),
	.w2(32'h3a4e7750),
	.w3(32'h3a6508fa),
	.w4(32'h37da636c),
	.w5(32'hbbe2ab9a),
	.w6(32'h3b83a89d),
	.w7(32'h3acd0884),
	.w8(32'hbb493a28),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c89d),
	.w1(32'hb8eaa229),
	.w2(32'h3b431015),
	.w3(32'h39d792a2),
	.w4(32'h3b19af3a),
	.w5(32'hbb053374),
	.w6(32'hba786ed2),
	.w7(32'h3b6275c5),
	.w8(32'hba57e731),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf33847),
	.w1(32'h39ab376a),
	.w2(32'h3919cdc9),
	.w3(32'hba63d4a8),
	.w4(32'hba247662),
	.w5(32'hbbe12a9c),
	.w6(32'h3aef1c95),
	.w7(32'h3b50aaa9),
	.w8(32'hbcbf65c2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1d6fa),
	.w1(32'h3be542c2),
	.w2(32'h3cf5a4cd),
	.w3(32'hbb60d58f),
	.w4(32'h3c8031bb),
	.w5(32'h3c3d99af),
	.w6(32'hbca5ee94),
	.w7(32'hbb1829a9),
	.w8(32'hbc7c2003),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bca0f),
	.w1(32'hbab6c0ae),
	.w2(32'h3c9f08f7),
	.w3(32'hbb63a3d8),
	.w4(32'h3c40f13a),
	.w5(32'h3c4e96d8),
	.w6(32'hbc438557),
	.w7(32'h3ab62927),
	.w8(32'h38db88f7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396da3be),
	.w1(32'h3b7b937c),
	.w2(32'h3a294462),
	.w3(32'h3b33d316),
	.w4(32'hba84ed0e),
	.w5(32'hbaf752d8),
	.w6(32'hbb863dc6),
	.w7(32'hbaec74cf),
	.w8(32'h3b84c643),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca44595),
	.w1(32'h3b99809d),
	.w2(32'hbc989890),
	.w3(32'hbbbfe827),
	.w4(32'h3c143a35),
	.w5(32'h3c2db390),
	.w6(32'h3c378fce),
	.w7(32'hbbf07809),
	.w8(32'hba3be6f7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb863dc8),
	.w1(32'hba8955e2),
	.w2(32'hbb891c81),
	.w3(32'hbb2a5be7),
	.w4(32'hbb62ce71),
	.w5(32'hbbedd715),
	.w6(32'h3a119704),
	.w7(32'h39191a3a),
	.w8(32'hbacbbd52),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe873a3),
	.w1(32'hbb1d3116),
	.w2(32'hbc3c6dfc),
	.w3(32'hbb11d424),
	.w4(32'hbbd53cc2),
	.w5(32'hbc839da8),
	.w6(32'hbc035466),
	.w7(32'hbc167ca5),
	.w8(32'hbd48650f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd052247),
	.w1(32'h3b6ce8b9),
	.w2(32'hbd2118a8),
	.w3(32'hbd0e33ea),
	.w4(32'hbd56c881),
	.w5(32'hbcba5481),
	.w6(32'hbd3181da),
	.w7(32'hbd115d70),
	.w8(32'h3b1b9f3f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4866ea),
	.w1(32'hbbb8b7fc),
	.w2(32'hbb8b2982),
	.w3(32'h3b254ec2),
	.w4(32'hbb5bb758),
	.w5(32'hbb17c43d),
	.w6(32'hba8a3b56),
	.w7(32'h3a9a57c2),
	.w8(32'hbb320174),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78ca07),
	.w1(32'hb9b3b75d),
	.w2(32'h3b59a391),
	.w3(32'hbaf8d309),
	.w4(32'h3a9264a0),
	.w5(32'hbb135f02),
	.w6(32'hbac40ec1),
	.w7(32'h3b558451),
	.w8(32'h3cd2cf2c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0bdf5b),
	.w1(32'hbbd0dba8),
	.w2(32'hbce23277),
	.w3(32'h3bcf2ed6),
	.w4(32'hbcb38ac5),
	.w5(32'hbcce57a3),
	.w6(32'h3c3b5855),
	.w7(32'hbbc9daf1),
	.w8(32'h3b0ab478),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba127792),
	.w1(32'hbb4602d0),
	.w2(32'hbbee3080),
	.w3(32'hba804a7f),
	.w4(32'hbb4faa3d),
	.w5(32'hbc053b13),
	.w6(32'hbbeee4d8),
	.w7(32'hbc0cee7c),
	.w8(32'hbc014428),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb005e41),
	.w1(32'h3bac0d74),
	.w2(32'hbac4bafc),
	.w3(32'hbba6a281),
	.w4(32'hba999a04),
	.w5(32'h3a0c0652),
	.w6(32'hbbe32c5d),
	.w7(32'hbbc86db8),
	.w8(32'h3cc53b3a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02daf0),
	.w1(32'hbbc1fcb0),
	.w2(32'hbcd3ad21),
	.w3(32'h3bc21f2d),
	.w4(32'hbca7a898),
	.w5(32'hbcc0b817),
	.w6(32'h3c2f4ebe),
	.w7(32'hbbbc6268),
	.w8(32'h3ca8cae9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdfc380),
	.w1(32'hbba5314f),
	.w2(32'hbcb4cdfb),
	.w3(32'h3ba65033),
	.w4(32'hbc8f2745),
	.w5(32'hbca4b5c9),
	.w6(32'h3c15d277),
	.w7(32'hbba10408),
	.w8(32'h3a41910a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b552d1a),
	.w1(32'hbbdd7589),
	.w2(32'hbc0fbd19),
	.w3(32'h3b0cb31e),
	.w4(32'hbb8e70ec),
	.w5(32'hbba42c2b),
	.w6(32'hb98745ca),
	.w7(32'hb951231c),
	.w8(32'hbbd8d522),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c126c),
	.w1(32'h3ab44be1),
	.w2(32'hbac44209),
	.w3(32'h3c190775),
	.w4(32'hbc3423d0),
	.w5(32'hbc2069a6),
	.w6(32'hbb36f940),
	.w7(32'hbb8c8482),
	.w8(32'hbaf5084c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ed39f),
	.w1(32'h3aa542ee),
	.w2(32'h3b2054e7),
	.w3(32'h377d0019),
	.w4(32'h3b2aaa00),
	.w5(32'h3a66ef76),
	.w6(32'h39aa39df),
	.w7(32'h3acc1ded),
	.w8(32'hbb9c5593),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb12720),
	.w1(32'h3c5ce743),
	.w2(32'hbb8ef1ce),
	.w3(32'hbb509e41),
	.w4(32'hbb7eff72),
	.w5(32'hbbf405a6),
	.w6(32'h3aaf108a),
	.w7(32'h3bb20075),
	.w8(32'hbb6ba87a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0afa6),
	.w1(32'hbbdc8573),
	.w2(32'hbb883a58),
	.w3(32'h3bc1acdf),
	.w4(32'hbb0beb95),
	.w5(32'hba352334),
	.w6(32'h3ba7e0e7),
	.w7(32'h3c45614f),
	.w8(32'h3ad70678),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce6fb6a),
	.w1(32'hbc102ade),
	.w2(32'h3cde1bbd),
	.w3(32'hbc2a89c9),
	.w4(32'h3b5e6f3f),
	.w5(32'h3bc248f1),
	.w6(32'h3abceb57),
	.w7(32'h3babccd9),
	.w8(32'hbc4a4860),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f3c80),
	.w1(32'hba8bcfce),
	.w2(32'hbc6c89ac),
	.w3(32'hbbb2da48),
	.w4(32'hbc93bd3b),
	.w5(32'hbab4db97),
	.w6(32'hbb73055c),
	.w7(32'hbc49cf32),
	.w8(32'hbca83290),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c9632),
	.w1(32'h3bc9b7c0),
	.w2(32'h3cd7caf1),
	.w3(32'hbb45b4fa),
	.w4(32'h3c61c865),
	.w5(32'h3c2798f9),
	.w6(32'hbc917105),
	.w7(32'hbb02fa91),
	.w8(32'h395c725f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cb684),
	.w1(32'hbaf83e46),
	.w2(32'hbbef6b18),
	.w3(32'hba708273),
	.w4(32'hbbec31e3),
	.w5(32'hbc4ff12a),
	.w6(32'hbbd0070f),
	.w7(32'hbbce7d61),
	.w8(32'hbc078f5b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896ad8),
	.w1(32'hbb2014d6),
	.w2(32'hbbdd8299),
	.w3(32'hbb9c2d71),
	.w4(32'hbbcbab66),
	.w5(32'h3add8fda),
	.w6(32'hbb8fe8dc),
	.w7(32'hba24bdb2),
	.w8(32'hbaeccc7f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb515322),
	.w1(32'h3ad494f3),
	.w2(32'h3b48373b),
	.w3(32'h3aa379aa),
	.w4(32'h3b510be0),
	.w5(32'h3adc19ea),
	.w6(32'h3ab0f5d8),
	.w7(32'h3b3bee46),
	.w8(32'hbcde2772),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1e0cff),
	.w1(32'hbc2bd9ff),
	.w2(32'h3d16b343),
	.w3(32'hbc050d69),
	.w4(32'h3cbae346),
	.w5(32'h3cd8ed28),
	.w6(32'hbcdb45d2),
	.w7(32'h3ad91374),
	.w8(32'hbaafca54),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f8c54),
	.w1(32'hbb0f7ecb),
	.w2(32'hbb4603fd),
	.w3(32'h3b140494),
	.w4(32'hbb2e2f67),
	.w5(32'hbad0431d),
	.w6(32'hb98d940f),
	.w7(32'h3ad468a0),
	.w8(32'h3c22224c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52dbd8),
	.w1(32'hbb2232ef),
	.w2(32'hbc30203c),
	.w3(32'h3b1ad3db),
	.w4(32'hbc07a629),
	.w5(32'hbc192ea2),
	.w6(32'h3b9897fb),
	.w7(32'hbb0e48b6),
	.w8(32'h3a434883),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984f8f1),
	.w1(32'h3976f2a9),
	.w2(32'h3949a56e),
	.w3(32'h376d030d),
	.w4(32'h38a787ab),
	.w5(32'hb8451546),
	.w6(32'h3a04823c),
	.w7(32'h38a2a476),
	.w8(32'hbb24221a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10bbfa),
	.w1(32'hba60de8a),
	.w2(32'hbadbe4cd),
	.w3(32'hba8d4444),
	.w4(32'hba8a1470),
	.w5(32'hbb366f36),
	.w6(32'hbb0568b1),
	.w7(32'h3a395741),
	.w8(32'h3a286868),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39383ceb),
	.w1(32'hb90960be),
	.w2(32'hb811e3a6),
	.w3(32'hb8fcc32a),
	.w4(32'hb7e369a9),
	.w5(32'h38848b80),
	.w6(32'h39a3d67d),
	.w7(32'hb87bfe6c),
	.w8(32'h3a1e7893),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e984f4),
	.w1(32'h3a24aa94),
	.w2(32'h3a355d20),
	.w3(32'h38e02cbb),
	.w4(32'h3a006641),
	.w5(32'h3a12f940),
	.w6(32'h3a0a8cbd),
	.w7(32'h39da7ee6),
	.w8(32'hba4d69de),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd93d7),
	.w1(32'hbb1331b9),
	.w2(32'hbab648cb),
	.w3(32'hbade0413),
	.w4(32'hba97ccf0),
	.w5(32'hba8d9e7b),
	.w6(32'hba311df9),
	.w7(32'hba8fbabb),
	.w8(32'h3b248865),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06462e),
	.w1(32'hbb1a8c3a),
	.w2(32'hbac01a19),
	.w3(32'hb696f98e),
	.w4(32'hbb218d94),
	.w5(32'hbb1a83c1),
	.w6(32'h3b4dc1bb),
	.w7(32'h3aadee99),
	.w8(32'h3a930be4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc685),
	.w1(32'h39e0db55),
	.w2(32'h3a7a9fa5),
	.w3(32'h3a8e94a3),
	.w4(32'h39f8934e),
	.w5(32'h399b8cd4),
	.w6(32'h3a86a98c),
	.w7(32'h3a97705a),
	.w8(32'hba22e050),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c12f3),
	.w1(32'hba8bd14e),
	.w2(32'hba61ac29),
	.w3(32'hba4c8795),
	.w4(32'hba7cf4e3),
	.w5(32'hba234a94),
	.w6(32'hba53f57c),
	.w7(32'hba77e4a8),
	.w8(32'h3a358879),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39748a4c),
	.w1(32'h38eab2b7),
	.w2(32'h3a1afc3b),
	.w3(32'h3845d61b),
	.w4(32'h39771729),
	.w5(32'h39acb7ce),
	.w6(32'h3a26befe),
	.w7(32'h39e030fb),
	.w8(32'h39d8941c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ad78a),
	.w1(32'h38e9bc81),
	.w2(32'h39538d67),
	.w3(32'hb689d1e8),
	.w4(32'h38c7c92d),
	.w5(32'h39896124),
	.w6(32'h3968c67e),
	.w7(32'h3943e2f7),
	.w8(32'h3a88b516),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad2dbc),
	.w1(32'h38acbe59),
	.w2(32'h3987526a),
	.w3(32'h38bfdd4e),
	.w4(32'h392eec1c),
	.w5(32'h3a0239ef),
	.w6(32'h3a3047e2),
	.w7(32'h39c04a12),
	.w8(32'h3ab2f34d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32a426),
	.w1(32'h3b3890a9),
	.w2(32'hba32de8c),
	.w3(32'h3b292e8a),
	.w4(32'hb98adaaf),
	.w5(32'hba2ed93e),
	.w6(32'hba14e797),
	.w7(32'h3a872452),
	.w8(32'h390c3a48),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e22e9),
	.w1(32'hba55d8b7),
	.w2(32'hb9bbf94c),
	.w3(32'hb8a8998e),
	.w4(32'hb9a23283),
	.w5(32'h3932a557),
	.w6(32'hba040db6),
	.w7(32'hba79348a),
	.w8(32'hb9c81ef2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae768f),
	.w1(32'hbb760d57),
	.w2(32'hbabe3dc9),
	.w3(32'h39cac393),
	.w4(32'hbb12dba0),
	.w5(32'hbab87a87),
	.w6(32'hba1200b4),
	.w7(32'h3a87e685),
	.w8(32'hb9e50409),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3aeed),
	.w1(32'hbb095634),
	.w2(32'hbb025a81),
	.w3(32'hb89cdf04),
	.w4(32'hba918c82),
	.w5(32'hbaeca890),
	.w6(32'h395fe1c6),
	.w7(32'hb9957f21),
	.w8(32'h398fa417),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dd75c),
	.w1(32'h391f1fc8),
	.w2(32'h3b14c7c7),
	.w3(32'h3a845bea),
	.w4(32'h3b1175aa),
	.w5(32'h3aa66e12),
	.w6(32'h3a623de7),
	.w7(32'h3afa2e74),
	.w8(32'hbb366262),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3a023),
	.w1(32'hb8eccdc6),
	.w2(32'hbb1ad6e2),
	.w3(32'hba1ba78a),
	.w4(32'hbad99a34),
	.w5(32'hbb3ac83b),
	.w6(32'hbb2710e0),
	.w7(32'hb9188fa8),
	.w8(32'h38d0a852),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e855bc),
	.w1(32'h38be30f2),
	.w2(32'h39622257),
	.w3(32'h37c9373c),
	.w4(32'h39878da9),
	.w5(32'h39846e00),
	.w6(32'h3929ecb2),
	.w7(32'h391aad2a),
	.w8(32'h3a13a207),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a677f42),
	.w1(32'h3a5c32a3),
	.w2(32'h3980bb72),
	.w3(32'h3a326866),
	.w4(32'hb9388f2a),
	.w5(32'h37e0f238),
	.w6(32'h3a33d102),
	.w7(32'h39c58260),
	.w8(32'h388b244c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03fb15),
	.w1(32'hba834c5e),
	.w2(32'h3b2ab082),
	.w3(32'h3a53ceb1),
	.w4(32'h3b28c3eb),
	.w5(32'h392f09aa),
	.w6(32'h3a337f4d),
	.w7(32'h3a159689),
	.w8(32'hb9c54e3e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70d98c),
	.w1(32'hbb27193e),
	.w2(32'hbb263de3),
	.w3(32'hbaa17474),
	.w4(32'hbaef98cb),
	.w5(32'hbb0e5993),
	.w6(32'hba1796c4),
	.w7(32'hbaac674c),
	.w8(32'h3a8d0190),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27b25e),
	.w1(32'h39b4282a),
	.w2(32'h3a09ced1),
	.w3(32'h39bcd331),
	.w4(32'h3a4e0b6a),
	.w5(32'h3a74979c),
	.w6(32'h3a0554b5),
	.w7(32'h389dd0d7),
	.w8(32'hbaa0f417),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c8a7f),
	.w1(32'h3b73e897),
	.w2(32'hbacf0b8a),
	.w3(32'h3a60d31a),
	.w4(32'h3aa02d3e),
	.w5(32'h3ae3adc6),
	.w6(32'hbb2db976),
	.w7(32'h39610e71),
	.w8(32'h3a38421a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d39b03),
	.w1(32'h38f624ec),
	.w2(32'h39a1c7e5),
	.w3(32'hb9556f62),
	.w4(32'h38bdbdf5),
	.w5(32'h398a586b),
	.w6(32'h39aa5e0f),
	.w7(32'h3945f412),
	.w8(32'h39910c2d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940e6f8),
	.w1(32'h38f59cbd),
	.w2(32'h392c3477),
	.w3(32'hb78104f2),
	.w4(32'h38b22638),
	.w5(32'h393fc6ba),
	.w6(32'h39492e1d),
	.w7(32'h38cbb63f),
	.w8(32'h3a077600),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39849423),
	.w1(32'h3941cde0),
	.w2(32'h3976444d),
	.w3(32'h388d138e),
	.w4(32'h392e52ba),
	.w5(32'h39a91b67),
	.w6(32'h39ae97c9),
	.w7(32'h394c8943),
	.w8(32'hb9ca53c2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba971c2a),
	.w1(32'hbb15c029),
	.w2(32'hbaea5b82),
	.w3(32'h393af9e3),
	.w4(32'hbaba7f85),
	.w5(32'hba833446),
	.w6(32'h393c9de3),
	.w7(32'h39a06228),
	.w8(32'h3a0d96f7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6432c),
	.w1(32'h39b47dfe),
	.w2(32'h39fe1bb5),
	.w3(32'h37af4e83),
	.w4(32'h3994e3bc),
	.w5(32'h39b8847b),
	.w6(32'h39f9ec8f),
	.w7(32'h39bc8e5d),
	.w8(32'h3a5f07d7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90e8eb),
	.w1(32'h3aa68f11),
	.w2(32'h3ab2c48d),
	.w3(32'h3a71c127),
	.w4(32'h3ac20d3b),
	.w5(32'h3a93c79a),
	.w6(32'h3aa39724),
	.w7(32'h3ab4d105),
	.w8(32'h3a8027b4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5c267),
	.w1(32'h39fad8f6),
	.w2(32'h39a21d61),
	.w3(32'hb81d7028),
	.w4(32'h3960dda4),
	.w5(32'h39b81a1f),
	.w6(32'h3a1d8408),
	.w7(32'h38ff5190),
	.w8(32'h3a1ac8ce),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986d310),
	.w1(32'h397af5a1),
	.w2(32'h3a10e0f5),
	.w3(32'h38f1876c),
	.w4(32'h39682051),
	.w5(32'h39b16324),
	.w6(32'h3a250c32),
	.w7(32'h3a096de2),
	.w8(32'h3a89ce17),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2da501),
	.w1(32'h3a5a896c),
	.w2(32'h3a189dcc),
	.w3(32'h382b2113),
	.w4(32'h39aa7753),
	.w5(32'h3a0d5ea5),
	.w6(32'h3a53fe4b),
	.w7(32'h399356d6),
	.w8(32'hbb5fe9bd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b18ed),
	.w1(32'hbb2189dc),
	.w2(32'hbb2355e5),
	.w3(32'hbac78d37),
	.w4(32'hbb09a149),
	.w5(32'hbb25c4dc),
	.w6(32'hbb34f7b2),
	.w7(32'hbb1a71b0),
	.w8(32'h398db934),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bacfdb),
	.w1(32'hb91c3359),
	.w2(32'hb994b669),
	.w3(32'hb8c4d89c),
	.w4(32'hb7b67afd),
	.w5(32'hb8cd8756),
	.w6(32'h389679bb),
	.w7(32'h388a8142),
	.w8(32'h3a2d76fd),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940df38),
	.w1(32'h38995e8d),
	.w2(32'h39064b1a),
	.w3(32'hb7d82afd),
	.w4(32'h388224ec),
	.w5(32'h394b664d),
	.w6(32'h39df9d2e),
	.w7(32'h3905d6b9),
	.w8(32'h3a2145a8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399aa6d1),
	.w1(32'h393fd498),
	.w2(32'h380ee1aa),
	.w3(32'h38bfe1d9),
	.w4(32'h392a30f4),
	.w5(32'h390101fa),
	.w6(32'h39ece4a3),
	.w7(32'h38d1daab),
	.w8(32'h3a771e9c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa21060),
	.w1(32'h3abc112b),
	.w2(32'h3acde22b),
	.w3(32'h3a840bae),
	.w4(32'h3ad98408),
	.w5(32'h3aa853ed),
	.w6(32'h3ab1df95),
	.w7(32'h3ac72cc1),
	.w8(32'h3a524e8c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c10e8),
	.w1(32'h3a5d9741),
	.w2(32'h3a8b7b09),
	.w3(32'h3a19598d),
	.w4(32'h3a902b76),
	.w5(32'h3a63eaf8),
	.w6(32'h3a6d3481),
	.w7(32'h3a4d1876),
	.w8(32'h379a360b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa0a6c),
	.w1(32'hb9d6c2b2),
	.w2(32'hb9a9bb4b),
	.w3(32'hb9882c46),
	.w4(32'hb936f8eb),
	.w5(32'hb994060b),
	.w6(32'hb87e2cb8),
	.w7(32'hb8e98a7e),
	.w8(32'hba0d0241),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaecc7f),
	.w1(32'hbb01ca6e),
	.w2(32'hba9882f8),
	.w3(32'h39ff5e5b),
	.w4(32'hba889e55),
	.w5(32'hbaf10a15),
	.w6(32'hb9a8336b),
	.w7(32'h38063e3b),
	.w8(32'h394b613f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb960fd2e),
	.w1(32'hba4f9603),
	.w2(32'hba53ec7d),
	.w3(32'hba3f056e),
	.w4(32'hba150f20),
	.w5(32'hba1a1ef7),
	.w6(32'hb99130ac),
	.w7(32'hb9f5672f),
	.w8(32'h39226ced),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4f475),
	.w1(32'hba45e4f4),
	.w2(32'h3a1f0a20),
	.w3(32'hba18e1eb),
	.w4(32'hb995c7cc),
	.w5(32'h397890ae),
	.w6(32'h3a2bb134),
	.w7(32'h3a302381),
	.w8(32'hba7a8523),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e1d17),
	.w1(32'hbb886559),
	.w2(32'hbb4a3901),
	.w3(32'hba9f3cf5),
	.w4(32'hbb14ed49),
	.w5(32'hbaa274ca),
	.w6(32'hbac0956d),
	.w7(32'hbab9575c),
	.w8(32'hb9a99e50),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e5298),
	.w1(32'hba9282ed),
	.w2(32'hba30a5df),
	.w3(32'hb9cd3e7f),
	.w4(32'hba0b506e),
	.w5(32'hb8d90f55),
	.w6(32'hba5346ea),
	.w7(32'hba88c503),
	.w8(32'h3a55a3e1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3c4b1),
	.w1(32'h3a164e58),
	.w2(32'h3a2576a2),
	.w3(32'h396c421a),
	.w4(32'h39f9c7d9),
	.w5(32'h3a18df47),
	.w6(32'h3a19ccf8),
	.w7(32'h39a92680),
	.w8(32'hba5629ec),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba906983),
	.w1(32'hbab88f0e),
	.w2(32'hba950b60),
	.w3(32'hba86dfbb),
	.w4(32'hbaa78695),
	.w5(32'hba57730d),
	.w6(32'hba8b3371),
	.w7(32'hbaa3cf7d),
	.w8(32'h39b1d412),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9712aa7),
	.w1(32'hb982b577),
	.w2(32'h3a42a51d),
	.w3(32'hb9bcad93),
	.w4(32'hba12f5be),
	.w5(32'hb7a64d20),
	.w6(32'h398c853b),
	.w7(32'h3a5119ac),
	.w8(32'hb9bf7d8d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396145e3),
	.w1(32'h3a27aefa),
	.w2(32'h393de1e2),
	.w3(32'h39cbe7a7),
	.w4(32'hb94664c8),
	.w5(32'h35a8bcc8),
	.w6(32'h38eae8f7),
	.w7(32'h39e275a7),
	.w8(32'hba4ebd79),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87c715),
	.w1(32'hbaacc3a3),
	.w2(32'hba8b4844),
	.w3(32'hba7c8826),
	.w4(32'hba9d5a57),
	.w5(32'hba4b0215),
	.w6(32'hba8246b3),
	.w7(32'hba99beb6),
	.w8(32'hba326887),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69c51f),
	.w1(32'hba954f59),
	.w2(32'hba71dcfc),
	.w3(32'hba5a29b0),
	.w4(32'hba87e96e),
	.w5(32'hba2f3b2e),
	.w6(32'hba5fa516),
	.w7(32'hba82b313),
	.w8(32'hb9a0b9b8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19370b),
	.w1(32'hba73ae46),
	.w2(32'hba3597b9),
	.w3(32'hba3394fa),
	.w4(32'hba31726c),
	.w5(32'hb9b9232d),
	.w6(32'hba898a8e),
	.w7(32'hbab19b57),
	.w8(32'hb8d9000c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985586b),
	.w1(32'hba9b1f65),
	.w2(32'hb9a089b3),
	.w3(32'h398bff84),
	.w4(32'hb94f8ffa),
	.w5(32'hbb0262b8),
	.w6(32'hbaaef01d),
	.w7(32'h3a3da65c),
	.w8(32'h399f0408),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e03c6c),
	.w1(32'h382cdb34),
	.w2(32'h383e1e20),
	.w3(32'h3895c23f),
	.w4(32'h389fc3ff),
	.w5(32'h390dc862),
	.w6(32'h395eef79),
	.w7(32'h390544c3),
	.w8(32'h3a8e61b1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ea9d3),
	.w1(32'hbac5ebfb),
	.w2(32'hb7ec9331),
	.w3(32'h3ad7a1bf),
	.w4(32'h39f76af1),
	.w5(32'h3a1348da),
	.w6(32'h3927657c),
	.w7(32'h3ab60c3b),
	.w8(32'h3a12b428),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f71f0),
	.w1(32'hb980b8c2),
	.w2(32'hb88b6753),
	.w3(32'h398bc782),
	.w4(32'h3a0bac59),
	.w5(32'h3ab2c8b0),
	.w6(32'hba4e2845),
	.w7(32'hba952b9c),
	.w8(32'h3a9c3e38),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38997b07),
	.w1(32'hbaf5bdcc),
	.w2(32'hbab6c50c),
	.w3(32'h3a667731),
	.w4(32'hb97a4ef6),
	.w5(32'hbaf00895),
	.w6(32'h3ae87528),
	.w7(32'h3b098cb2),
	.w8(32'h3abcfda6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b259dea),
	.w1(32'h3a18a89a),
	.w2(32'hba43231b),
	.w3(32'h39d9aa87),
	.w4(32'hba8e1e33),
	.w5(32'hb9b70f93),
	.w6(32'h3b51ec31),
	.w7(32'h3b25113c),
	.w8(32'h3a58e153),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f0ed3),
	.w1(32'h3aa7cba4),
	.w2(32'h3ab53c6b),
	.w3(32'h3a6a94df),
	.w4(32'h3abf8b09),
	.w5(32'h3a92d8eb),
	.w6(32'h3a9ab5a7),
	.w7(32'h3aae4f7b),
	.w8(32'h3939c963),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961e22e),
	.w1(32'hb97b3f2a),
	.w2(32'h3a0794e6),
	.w3(32'hba2b4cc7),
	.w4(32'hb99a72dd),
	.w5(32'h389cb9bd),
	.w6(32'h3987802f),
	.w7(32'h3a035904),
	.w8(32'hb9fedf5d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92212b),
	.w1(32'hba8817b4),
	.w2(32'hba6c0593),
	.w3(32'hba1c0eeb),
	.w4(32'hbac52502),
	.w5(32'hba97bb2d),
	.w6(32'hba279ddf),
	.w7(32'hba09fc08),
	.w8(32'h39fbce9c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de0a90),
	.w1(32'h35a27e79),
	.w2(32'h39701c9d),
	.w3(32'hb897c590),
	.w4(32'h38ab44ee),
	.w5(32'h39a31f7e),
	.w6(32'h398f483a),
	.w7(32'h394055e7),
	.w8(32'h3a90eb74),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e89cb),
	.w1(32'h3a92aa64),
	.w2(32'h3aefd460),
	.w3(32'h3a6c0cc9),
	.w4(32'h3ae47803),
	.w5(32'h3aa7bdab),
	.w6(32'h3ab10f76),
	.w7(32'h3a98f6be),
	.w8(32'h3829f5a0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9842f42),
	.w1(32'hba13f41a),
	.w2(32'hb9a93e42),
	.w3(32'hb99620f4),
	.w4(32'hb9829333),
	.w5(32'h3816284b),
	.w6(32'hba1d1ac2),
	.w7(32'hba55d659),
	.w8(32'hb9adc158),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2ec70),
	.w1(32'hba0e32be),
	.w2(32'hb9ee4296),
	.w3(32'hb9d0d115),
	.w4(32'hba039af8),
	.w5(32'hb9ae1b90),
	.w6(32'hb9ddb79f),
	.w7(32'hba00a05c),
	.w8(32'hba676788),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbec0c5),
	.w1(32'h39fe3916),
	.w2(32'h380fecec),
	.w3(32'hba9f02b3),
	.w4(32'h3affac89),
	.w5(32'hbae75368),
	.w6(32'hbadb05ca),
	.w7(32'hbad757ad),
	.w8(32'hbbdb5fb2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4382d7),
	.w1(32'hbca5fcfb),
	.w2(32'h3cbc4b01),
	.w3(32'hbc4d7d23),
	.w4(32'hbd011ba3),
	.w5(32'h3aa458e3),
	.w6(32'hbca01b47),
	.w7(32'h3c4f07e8),
	.w8(32'h3aa64c23),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b966ef7),
	.w1(32'h3ab8b581),
	.w2(32'h3b7ce7ed),
	.w3(32'hb9e7a20f),
	.w4(32'h3b0a81cb),
	.w5(32'hba7dcd04),
	.w6(32'h3ba6aa0a),
	.w7(32'h3afe6ffa),
	.w8(32'hba3ecc1c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eadbca),
	.w1(32'hbb4e54c7),
	.w2(32'hba199b0d),
	.w3(32'h3aa3cb1a),
	.w4(32'h39dde0e5),
	.w5(32'hbaadb569),
	.w6(32'hbb0b447c),
	.w7(32'hbb675553),
	.w8(32'hbb08ba3d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf29ab),
	.w1(32'hbc0e7c0d),
	.w2(32'hbabb4b16),
	.w3(32'hba924a70),
	.w4(32'h3bdb543b),
	.w5(32'h3a69b498),
	.w6(32'hbb05e090),
	.w7(32'hbb6d74af),
	.w8(32'h3b6f2ba9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be45dcc),
	.w1(32'h392cda4d),
	.w2(32'hb9a1ad13),
	.w3(32'hbba480f0),
	.w4(32'hbbc1e47c),
	.w5(32'hb9a235de),
	.w6(32'h3c706296),
	.w7(32'hbbc419a2),
	.w8(32'h3c0256d9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4db71d),
	.w1(32'h3b04d0f3),
	.w2(32'h3b8c37d8),
	.w3(32'h3bb1cc6a),
	.w4(32'h3c2dba8b),
	.w5(32'h3c3f6bdf),
	.w6(32'h3b2e47c0),
	.w7(32'hba7b1386),
	.w8(32'h3c1b8314),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19c82c),
	.w1(32'h3a9dd726),
	.w2(32'h3ae97b7d),
	.w3(32'h3b4ff704),
	.w4(32'h391c0518),
	.w5(32'h3bef03dc),
	.w6(32'h3b471299),
	.w7(32'h3b3752d8),
	.w8(32'h3a411774),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad85291),
	.w1(32'hbbe4eec7),
	.w2(32'h3aa8ba68),
	.w3(32'h3ba2ad1b),
	.w4(32'h3b44aff6),
	.w5(32'h3ab860ff),
	.w6(32'hbaadf423),
	.w7(32'h3ada3ede),
	.w8(32'h3987a810),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabd76f),
	.w1(32'hbb7aea57),
	.w2(32'h3b40fdd7),
	.w3(32'h3a417a62),
	.w4(32'hb6c09516),
	.w5(32'h3a26728f),
	.w6(32'h393d1b0d),
	.w7(32'h3b1c2dc8),
	.w8(32'h3b1296bd),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba94d21),
	.w1(32'hbb8edd13),
	.w2(32'h3bb79b75),
	.w3(32'h398f51bc),
	.w4(32'hb980ba78),
	.w5(32'hb965dd41),
	.w6(32'h3b51fa46),
	.w7(32'h3bab9e66),
	.w8(32'hbbaf0558),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17713a),
	.w1(32'hbcd533f3),
	.w2(32'hbbb8f190),
	.w3(32'h3ca1de44),
	.w4(32'hbbc293c9),
	.w5(32'hb9b06b7e),
	.w6(32'hbcd9542d),
	.w7(32'h3ab18ecf),
	.w8(32'h3b1e9cf8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c62b8),
	.w1(32'hbbee7372),
	.w2(32'hbbbb8476),
	.w3(32'hbb076a61),
	.w4(32'hbbf12e4d),
	.w5(32'hbba63249),
	.w6(32'h3a7d2696),
	.w7(32'hba9badbc),
	.w8(32'h3b97cd07),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc4e6f),
	.w1(32'h3be477ae),
	.w2(32'hbb536cc7),
	.w3(32'h3bc478a1),
	.w4(32'h3c4a29ff),
	.w5(32'hbb3abb3a),
	.w6(32'hb9d55fa1),
	.w7(32'hbbe163d9),
	.w8(32'hbbf1f555),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c1bf1),
	.w1(32'hbbf4cdb5),
	.w2(32'hbd05c9fa),
	.w3(32'hbc6affd7),
	.w4(32'hbccf1e8d),
	.w5(32'hbca288e4),
	.w6(32'hbc86d0c6),
	.w7(32'hbc817ee0),
	.w8(32'hbc286cea),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fd6fe),
	.w1(32'h3c474710),
	.w2(32'h3c220e7f),
	.w3(32'h3bd9ad3d),
	.w4(32'h3c08c11d),
	.w5(32'hbc2b6c72),
	.w6(32'hbb60be1b),
	.w7(32'hba9635b3),
	.w8(32'hbad2e659),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc707fa1),
	.w1(32'h3c526411),
	.w2(32'hbbbffc31),
	.w3(32'hbca4e4bd),
	.w4(32'hbc62644e),
	.w5(32'hb896e8ee),
	.w6(32'hbc1e101f),
	.w7(32'hbace8d77),
	.w8(32'h3b90bcf5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc786a3),
	.w1(32'hbac03994),
	.w2(32'h3c0623bc),
	.w3(32'h3bad09dc),
	.w4(32'h3b007b30),
	.w5(32'h3bc55187),
	.w6(32'h3a8db62d),
	.w7(32'h3bce6d07),
	.w8(32'hbaa701b4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0042b9),
	.w1(32'h3bb1bce1),
	.w2(32'h3aa8aa7c),
	.w3(32'hbb69739c),
	.w4(32'hbb9e7de9),
	.w5(32'hbbb40b90),
	.w6(32'h39dc1f30),
	.w7(32'hbbd0d1c0),
	.w8(32'hbc7ac2fb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05af5e),
	.w1(32'hbc5f66c7),
	.w2(32'h3c823ca9),
	.w3(32'hbc420913),
	.w4(32'h3c4fc932),
	.w5(32'h3c152db7),
	.w6(32'hbd23e732),
	.w7(32'hbceeceb6),
	.w8(32'hbbc400e6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0055b),
	.w1(32'hbc04146a),
	.w2(32'h3aa3cec2),
	.w3(32'h39b2ed0d),
	.w4(32'hba567f90),
	.w5(32'hbac96e73),
	.w6(32'hbb6564a7),
	.w7(32'h3aa305cd),
	.w8(32'h3bfc7507),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd9ae),
	.w1(32'hbc010980),
	.w2(32'h3b5cee8b),
	.w3(32'h3c01ede8),
	.w4(32'h3b387fa6),
	.w5(32'h3b9befc2),
	.w6(32'h3935eb60),
	.w7(32'h3c0a9ef9),
	.w8(32'hbc98dd2a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd157531),
	.w1(32'hbc96fd5a),
	.w2(32'h3c516898),
	.w3(32'hba5cac02),
	.w4(32'hbc8e013a),
	.w5(32'hbbab2898),
	.w6(32'h3c486a3e),
	.w7(32'h3c2a52df),
	.w8(32'h39e62adb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule