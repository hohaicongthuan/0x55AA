module layer_8_featuremap_219(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b0ecb),
	.w1(32'hbbd75ec0),
	.w2(32'h3a9c5b22),
	.w3(32'hbc8e6ece),
	.w4(32'h3b691933),
	.w5(32'h3c36771a),
	.w6(32'hbaa8031d),
	.w7(32'h3bb1975b),
	.w8(32'h3c9d4a3f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c89e5),
	.w1(32'hbafa070e),
	.w2(32'h3afc8a10),
	.w3(32'hbc5b3ebe),
	.w4(32'hbabcc0e7),
	.w5(32'hbb1b291e),
	.w6(32'hbbe5b814),
	.w7(32'hbabd7a50),
	.w8(32'hbb139b4a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6188cf),
	.w1(32'hbbaeee3c),
	.w2(32'h3b0b3a0e),
	.w3(32'hbbc611bc),
	.w4(32'h3c3fbe91),
	.w5(32'h3c803729),
	.w6(32'hbb6fdcdd),
	.w7(32'hbbfc628b),
	.w8(32'hbc290e50),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88f582),
	.w1(32'hbb8caba4),
	.w2(32'hbbc749fe),
	.w3(32'h3c1136a2),
	.w4(32'hbb9e92c6),
	.w5(32'h3c908af5),
	.w6(32'h3c76736b),
	.w7(32'h3cbf731b),
	.w8(32'h3c635442),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc276aa3),
	.w1(32'hbb380f0b),
	.w2(32'hbbb27c5a),
	.w3(32'h3c4db0fa),
	.w4(32'hbb92e563),
	.w5(32'hbb2dfc4a),
	.w6(32'h3b500e58),
	.w7(32'h3b3c099f),
	.w8(32'hbabef779),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b47c),
	.w1(32'hbc347dec),
	.w2(32'hbca71ccb),
	.w3(32'h3b3f70b4),
	.w4(32'hbc831923),
	.w5(32'hbd121f33),
	.w6(32'hbca8baa6),
	.w7(32'hbcce8b6d),
	.w8(32'hbd022950),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc843b1f),
	.w1(32'hba5fbdbb),
	.w2(32'hbbed838c),
	.w3(32'hbc8e0cf7),
	.w4(32'hbb3c63a1),
	.w5(32'hb9966b24),
	.w6(32'h3b8e9e52),
	.w7(32'h3c00058f),
	.w8(32'h3b12ae27),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c0bc3),
	.w1(32'h3c183cd6),
	.w2(32'h3c1bdf9e),
	.w3(32'hbb9f1137),
	.w4(32'hbc689fad),
	.w5(32'hbc8a3743),
	.w6(32'h3c2098a0),
	.w7(32'h3cb8bbd3),
	.w8(32'h3c728974),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5e52c),
	.w1(32'hbc1cfee3),
	.w2(32'hbca74e87),
	.w3(32'hbc4dc3f8),
	.w4(32'hbbcd3e95),
	.w5(32'hbb45c245),
	.w6(32'h3c3250e8),
	.w7(32'h3c086c8a),
	.w8(32'h3b9fe664),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8f337),
	.w1(32'hbbe0938c),
	.w2(32'hbbed6f6e),
	.w3(32'hbb7a93be),
	.w4(32'hbb9777cd),
	.w5(32'hbb5749fb),
	.w6(32'hbb2dd00c),
	.w7(32'h3c116bf5),
	.w8(32'h3bdafc94),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd045af4),
	.w1(32'h3994807a),
	.w2(32'h3b8d8cf7),
	.w3(32'hbcaa24f4),
	.w4(32'hbbe3d75f),
	.w5(32'hbba654d9),
	.w6(32'hba181dec),
	.w7(32'h3c565ebe),
	.w8(32'h3caeed19),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc00248),
	.w1(32'hbc495c7a),
	.w2(32'h3bc8ffc9),
	.w3(32'hbc92ae9a),
	.w4(32'hbc2e491f),
	.w5(32'hbbc15da7),
	.w6(32'hbbd47b0f),
	.w7(32'h3be1ad7b),
	.w8(32'h3c25ea3d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c9cac),
	.w1(32'h3c80eb65),
	.w2(32'h3d015be8),
	.w3(32'hbca3a5da),
	.w4(32'hbbbf6d23),
	.w5(32'hbc323976),
	.w6(32'h3c549081),
	.w7(32'h3c973203),
	.w8(32'h3c4ed6ef),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74a561),
	.w1(32'hbb2990bb),
	.w2(32'hbc3f1387),
	.w3(32'hbc9d66d3),
	.w4(32'hbb0daf2b),
	.w5(32'hbac2918f),
	.w6(32'hbc8b61ed),
	.w7(32'hbcd3bfd7),
	.w8(32'hbc746a36),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc93d1d),
	.w1(32'hbbf9cc45),
	.w2(32'hbc895f6b),
	.w3(32'hbbed6aa6),
	.w4(32'hbbb95752),
	.w5(32'hb9ae3300),
	.w6(32'h3bc5096d),
	.w7(32'h3b8facc3),
	.w8(32'h3a06e941),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1185ca),
	.w1(32'hbb8dcf3d),
	.w2(32'hbba3c758),
	.w3(32'h3c05b1d5),
	.w4(32'hbaa34377),
	.w5(32'hbbd173e1),
	.w6(32'hb93b21b6),
	.w7(32'hbba1f461),
	.w8(32'h3a4dbf02),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e46ab),
	.w1(32'h3c1fd2b3),
	.w2(32'h3ba567e6),
	.w3(32'hbba9f12b),
	.w4(32'h39b530ed),
	.w5(32'h3c113fe7),
	.w6(32'hbc26ca34),
	.w7(32'hbb029ed0),
	.w8(32'hbae64ae5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb155cd8),
	.w1(32'h3a0e9063),
	.w2(32'h3c652689),
	.w3(32'hbc6ca696),
	.w4(32'h3b01267f),
	.w5(32'h3bb7c4c7),
	.w6(32'hbac54ea0),
	.w7(32'h3c3e1c82),
	.w8(32'h3c26c003),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfd7559),
	.w1(32'hbc5afdec),
	.w2(32'h3cd1a02a),
	.w3(32'hbd18c89a),
	.w4(32'h3bfa4686),
	.w5(32'h3d5834ac),
	.w6(32'hbcae154d),
	.w7(32'h3c95933c),
	.w8(32'h3d3d191d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17168c),
	.w1(32'hbc597443),
	.w2(32'hbc69499b),
	.w3(32'hba8656cd),
	.w4(32'hb9a48280),
	.w5(32'hbb063d96),
	.w6(32'hbb350a35),
	.w7(32'hbb9d0c36),
	.w8(32'hbb891f54),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1907eb),
	.w1(32'h3b9d54f4),
	.w2(32'hbca8c125),
	.w3(32'h3c81c2d4),
	.w4(32'h3a960a0f),
	.w5(32'hbca850b1),
	.w6(32'hbbe68f8c),
	.w7(32'hbc11662f),
	.w8(32'hbc506e06),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf4a0f),
	.w1(32'hbcb032a6),
	.w2(32'hbd12c336),
	.w3(32'hbbffe6cb),
	.w4(32'hbc9e069a),
	.w5(32'hbc41843f),
	.w6(32'hbbd33419),
	.w7(32'hbc8baefd),
	.w8(32'hbcfa525b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce73455),
	.w1(32'hbc987947),
	.w2(32'h3d24d635),
	.w3(32'hbc825b35),
	.w4(32'h3cd67e2c),
	.w5(32'h3d9d3da9),
	.w6(32'hbce7d781),
	.w7(32'h3bfe9355),
	.w8(32'h3cfb4183),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00d6df),
	.w1(32'hbc584b66),
	.w2(32'hbc75acdd),
	.w3(32'hbbae0549),
	.w4(32'hbc2fa0ec),
	.w5(32'hbc3abb7e),
	.w6(32'h3bef8b61),
	.w7(32'hbc8dbe85),
	.w8(32'hbca8d580),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ea49a),
	.w1(32'hbc8a97d6),
	.w2(32'h3bc3b67e),
	.w3(32'h3ab13e16),
	.w4(32'h377f8743),
	.w5(32'h3c3f7ec8),
	.w6(32'hbcafc9a3),
	.w7(32'hbcfd52b6),
	.w8(32'hbc6f6e30),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b829b6e),
	.w1(32'hbc34e3ee),
	.w2(32'h3a28bbd7),
	.w3(32'hbc5e3cab),
	.w4(32'hbc18ac69),
	.w5(32'hbb86f7d0),
	.w6(32'hbcda8217),
	.w7(32'hbc276598),
	.w8(32'h3c730757),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25c983),
	.w1(32'hbcd99051),
	.w2(32'hbd1c4aa5),
	.w3(32'hbbd03c48),
	.w4(32'hbc922627),
	.w5(32'hbc84706a),
	.w6(32'hbb9d0e7d),
	.w7(32'hbc8d504f),
	.w8(32'hbc8dcb29),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbde203d5),
	.w1(32'h3d7ecbb6),
	.w2(32'h3c544534),
	.w3(32'hbdfd4a20),
	.w4(32'h3cd2fcbf),
	.w5(32'hbb3c12d8),
	.w6(32'hbdd827b2),
	.w7(32'hbc929654),
	.w8(32'h3d5baed2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf0eca),
	.w1(32'hbac3a382),
	.w2(32'h3b8c28e2),
	.w3(32'hbc280753),
	.w4(32'hbc358b6c),
	.w5(32'hbc796892),
	.w6(32'hb886399a),
	.w7(32'h3ca6727e),
	.w8(32'h3c36904c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9292fa),
	.w1(32'hbb0ba534),
	.w2(32'hbbf1c2f8),
	.w3(32'hbc9e8bb7),
	.w4(32'h3b27c636),
	.w5(32'h3b233e0c),
	.w6(32'hbb1758ad),
	.w7(32'h3b01635d),
	.w8(32'h3bcd6079),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3244c2),
	.w1(32'h3c85bbaa),
	.w2(32'h3cc293bf),
	.w3(32'h3c485bcd),
	.w4(32'hbc90627a),
	.w5(32'hbd209845),
	.w6(32'h3bcde770),
	.w7(32'h3cb32144),
	.w8(32'h3c91c620),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e67d5),
	.w1(32'hba0f552c),
	.w2(32'h3c8b375d),
	.w3(32'hbd0434a4),
	.w4(32'hbb7a1159),
	.w5(32'hbb1f3ba2),
	.w6(32'hbc3ca5ca),
	.w7(32'hbc4f6477),
	.w8(32'h3aed8685),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbbfde6),
	.w1(32'hbbd6f611),
	.w2(32'hbc94be4d),
	.w3(32'hbad44e38),
	.w4(32'hbc215553),
	.w5(32'hbc3f05b7),
	.w6(32'hbc08a010),
	.w7(32'hbbf9f0ae),
	.w8(32'hbbaed030),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20a0d3),
	.w1(32'h3a1d9cf7),
	.w2(32'h3bdc21a6),
	.w3(32'hbc3b3a8e),
	.w4(32'h37898e77),
	.w5(32'hbab979f2),
	.w6(32'hbb846c1d),
	.w7(32'h3b4fbe8c),
	.w8(32'hbb82e95d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749c97),
	.w1(32'h3c169bde),
	.w2(32'h3bc638dc),
	.w3(32'h3b2c4c0e),
	.w4(32'hbc0cf63d),
	.w5(32'hbca4ce75),
	.w6(32'h3c9f4741),
	.w7(32'h3c1a14e7),
	.w8(32'h3b9b461c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e6da1),
	.w1(32'h3add6ce6),
	.w2(32'h3be4964c),
	.w3(32'hbd092f4b),
	.w4(32'hbb05d578),
	.w5(32'h3bd65e18),
	.w6(32'hbc79b07c),
	.w7(32'h3b886d14),
	.w8(32'h3bc9df6c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7a5d4),
	.w1(32'hbc037c3f),
	.w2(32'h399a9a2b),
	.w3(32'h3b6f56cb),
	.w4(32'hbb8ffae0),
	.w5(32'h3bbd19d4),
	.w6(32'hbbe6840a),
	.w7(32'hbb90f3fe),
	.w8(32'hbb5b4c06),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a13f7),
	.w1(32'hbbd898ab),
	.w2(32'hbc9a95d3),
	.w3(32'h3b7a0776),
	.w4(32'hbb742eae),
	.w5(32'hbb34c0da),
	.w6(32'h3b8697ae),
	.w7(32'h3bdd33eb),
	.w8(32'h3babf0b5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc301024),
	.w1(32'hbbe71d3e),
	.w2(32'hbbee1077),
	.w3(32'h3ba3b210),
	.w4(32'hba25b11c),
	.w5(32'h3b13773b),
	.w6(32'h3ba45e96),
	.w7(32'hbbf03ec0),
	.w8(32'hba71c493),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b535a52),
	.w1(32'h3bef3720),
	.w2(32'h3c14a085),
	.w3(32'h3b1f33ad),
	.w4(32'h3a71f51e),
	.w5(32'h3bda53e2),
	.w6(32'hba0fb3f9),
	.w7(32'h3ac11db0),
	.w8(32'h3b90a421),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0f222d),
	.w1(32'hbc80cefe),
	.w2(32'hba74d47b),
	.w3(32'hbd1b45f3),
	.w4(32'hbc5de303),
	.w5(32'hba2ce0fd),
	.w6(32'hbcfb9623),
	.w7(32'hbb56a988),
	.w8(32'hbc28bd62),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc080068),
	.w1(32'hbba0a997),
	.w2(32'h3bca8309),
	.w3(32'hbc3adca1),
	.w4(32'h3bb5316a),
	.w5(32'h3c05bb57),
	.w6(32'h3acdade1),
	.w7(32'hbc24d9b8),
	.w8(32'h3bb7e3c5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1942a),
	.w1(32'hbb4c170c),
	.w2(32'h3b0e3a7d),
	.w3(32'hbbac2a03),
	.w4(32'hbc2d05bb),
	.w5(32'hba3612a4),
	.w6(32'hbb75a41f),
	.w7(32'hba9909b9),
	.w8(32'hbb4a502f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc0697),
	.w1(32'hbc290928),
	.w2(32'hbbb5d7fe),
	.w3(32'hbc5a80f5),
	.w4(32'hbc294684),
	.w5(32'hbb3d387d),
	.w6(32'hbb83f363),
	.w7(32'h3c30eba3),
	.w8(32'h3c4880df),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a44a6),
	.w1(32'hbbcbe5ca),
	.w2(32'hbbb7b1e0),
	.w3(32'hbc942f2f),
	.w4(32'h3b821463),
	.w5(32'h3ca2f093),
	.w6(32'h3b006bfb),
	.w7(32'h3c9b5149),
	.w8(32'h3cceefae),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b509931),
	.w1(32'hbb1c5cad),
	.w2(32'h3bbf2f75),
	.w3(32'h3c882a25),
	.w4(32'h3b047171),
	.w5(32'h3c44ffcb),
	.w6(32'h3bd855a9),
	.w7(32'h3c3ae5e3),
	.w8(32'h3c811416),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f980a0),
	.w1(32'hbc28a9f3),
	.w2(32'hbab1f458),
	.w3(32'h3b43c597),
	.w4(32'hba24df0d),
	.w5(32'h3c420189),
	.w6(32'hbba344c5),
	.w7(32'hbafd0d17),
	.w8(32'hba858b06),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc56806),
	.w1(32'hbccfb74d),
	.w2(32'hbc1ca599),
	.w3(32'h3bc80bfb),
	.w4(32'hbc19af42),
	.w5(32'h3b0f8fa9),
	.w6(32'hba24d674),
	.w7(32'h3adb7739),
	.w8(32'h3b9094e9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42093),
	.w1(32'hbc918e37),
	.w2(32'hbcce250b),
	.w3(32'hbbb644a5),
	.w4(32'hbb822ec9),
	.w5(32'h3abee76b),
	.w6(32'h3bb74e74),
	.w7(32'hbc6431cb),
	.w8(32'hbcfe25a8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ac470),
	.w1(32'h3b209e10),
	.w2(32'h3c911c34),
	.w3(32'hbc141ff1),
	.w4(32'hbb8f5877),
	.w5(32'h3c15eadd),
	.w6(32'hbbccd1e0),
	.w7(32'h3c464555),
	.w8(32'h3bf02c15),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0314d),
	.w1(32'hbc128b24),
	.w2(32'hbc53f52e),
	.w3(32'hbbd4691d),
	.w4(32'hbb1369d4),
	.w5(32'hbc27986d),
	.w6(32'h3c1488f4),
	.w7(32'h3c4988cd),
	.w8(32'hbc808dec),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75d3f6),
	.w1(32'hbc972a96),
	.w2(32'h38c25ae5),
	.w3(32'hbd0e2cdb),
	.w4(32'h3b3e8ddf),
	.w5(32'h3ce608b6),
	.w6(32'hbd1af269),
	.w7(32'hbbec5a5e),
	.w8(32'h3c788992),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4a302),
	.w1(32'hbb54fec8),
	.w2(32'hbb11665a),
	.w3(32'h3a756cba),
	.w4(32'h3aada694),
	.w5(32'h3bcef788),
	.w6(32'h3bb3d7e0),
	.w7(32'h3c24c89d),
	.w8(32'h3c22e15c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08dea2),
	.w1(32'hbbd77738),
	.w2(32'h39d487b6),
	.w3(32'hbbc2205e),
	.w4(32'h3c39ab32),
	.w5(32'h3bc78905),
	.w6(32'h3b3aeb21),
	.w7(32'h3b4da60b),
	.w8(32'h3cc82afc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e5848),
	.w1(32'h3939db12),
	.w2(32'h3a69dcbe),
	.w3(32'hbbdb40e6),
	.w4(32'h3b29dd44),
	.w5(32'h3a7d57dd),
	.w6(32'h3b2da863),
	.w7(32'h3ab6d823),
	.w8(32'h3c36e902),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee5f6),
	.w1(32'hbcc2e8ff),
	.w2(32'hbbf43f68),
	.w3(32'hbca53714),
	.w4(32'h3b4e7c97),
	.w5(32'h3bbd5d1c),
	.w6(32'hbbb1367b),
	.w7(32'h3cf4ff1e),
	.w8(32'h3d1d79bc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b8097),
	.w1(32'hbba0780d),
	.w2(32'hbb41b4c1),
	.w3(32'hbc7be96f),
	.w4(32'hbc96603a),
	.w5(32'hbc57e65b),
	.w6(32'hbb93fdb5),
	.w7(32'hbc44c356),
	.w8(32'hbb1bac7f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca039d0),
	.w1(32'h3b1425f8),
	.w2(32'h3b7c724a),
	.w3(32'hbcb97103),
	.w4(32'hbc20546d),
	.w5(32'hbb89d618),
	.w6(32'hbbf9a4ce),
	.w7(32'h3c1d4cc1),
	.w8(32'h3c6386a7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f8296),
	.w1(32'hbc12bd79),
	.w2(32'hbb8f0323),
	.w3(32'hbc026003),
	.w4(32'hbbd91fe5),
	.w5(32'hba2efd75),
	.w6(32'hbbe436ac),
	.w7(32'h3913608c),
	.w8(32'h3c046b8b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c24a5),
	.w1(32'hbb9b3b2c),
	.w2(32'hbc8cf1b2),
	.w3(32'hbc0a7214),
	.w4(32'hbc35c9ad),
	.w5(32'h3aace493),
	.w6(32'hbbb3d4f4),
	.w7(32'hbc37d54f),
	.w8(32'hbc11a4fb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25cb45),
	.w1(32'hbcd18e1a),
	.w2(32'hbca7e7a4),
	.w3(32'h3c50f88b),
	.w4(32'hba52bb8c),
	.w5(32'h3c9ee4cb),
	.w6(32'hbc799ada),
	.w7(32'hbd0bd2ad),
	.w8(32'hbccfbec1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd9c74),
	.w1(32'hbcd7fc33),
	.w2(32'hbc94173f),
	.w3(32'h3c3085d6),
	.w4(32'h396231b9),
	.w5(32'h3cc9a1eb),
	.w6(32'hbb52bdb6),
	.w7(32'hbc3a1f1d),
	.w8(32'hbba03830),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b4198),
	.w1(32'h3a45a114),
	.w2(32'h3b5f74d8),
	.w3(32'h3bf73804),
	.w4(32'h3b86fcb5),
	.w5(32'hbc05d113),
	.w6(32'hbbecd0e0),
	.w7(32'h3c64ccc0),
	.w8(32'h3c84e904),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbf321),
	.w1(32'hbb49ea06),
	.w2(32'h39148cb8),
	.w3(32'hbcbd08b4),
	.w4(32'hbba89bf2),
	.w5(32'h3ade6c3f),
	.w6(32'hbc1bbcc6),
	.w7(32'hbb6e6187),
	.w8(32'hbb7c7a58),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4cd300),
	.w1(32'hbb84a676),
	.w2(32'h39a9b4e2),
	.w3(32'h39fc296c),
	.w4(32'hbbee6b5b),
	.w5(32'hbc09ebb2),
	.w6(32'hbbc9066a),
	.w7(32'hbb6aa1a4),
	.w8(32'hb9c7547d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c2225),
	.w1(32'h3a9be0c9),
	.w2(32'h3c1fcc78),
	.w3(32'hbca35cda),
	.w4(32'h3b115c73),
	.w5(32'h3c3e5b13),
	.w6(32'hbc0daa1c),
	.w7(32'h3c0b1d80),
	.w8(32'h3c19b869),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aab78),
	.w1(32'hbc943e61),
	.w2(32'hbcaf9ef4),
	.w3(32'hb98bbcf4),
	.w4(32'hbbbf0ae4),
	.w5(32'hbbbc92bd),
	.w6(32'hbb4e241a),
	.w7(32'hbbc7a84b),
	.w8(32'hba7ad67e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194a40),
	.w1(32'hbc3293f8),
	.w2(32'hbaf77086),
	.w3(32'h3b0a0078),
	.w4(32'h3b82f1f3),
	.w5(32'h3bbaed82),
	.w6(32'hba4aa9ba),
	.w7(32'hbb3b8aea),
	.w8(32'hbc01eb22),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25b97c),
	.w1(32'h3c05b340),
	.w2(32'h3c64b5ac),
	.w3(32'h3c0e7692),
	.w4(32'h3b865dbb),
	.w5(32'h3a0a3f4f),
	.w6(32'h3a8a65a3),
	.w7(32'h3bc797f6),
	.w8(32'h3c007b46),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39d378),
	.w1(32'hbb9d4f85),
	.w2(32'hbc9b82c8),
	.w3(32'hbcab86cf),
	.w4(32'hbc7864cf),
	.w5(32'h3caf5531),
	.w6(32'hbcb2804e),
	.w7(32'h3c164955),
	.w8(32'h3cbcff02),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc49ea1),
	.w1(32'hbb0f84ec),
	.w2(32'hbc47998b),
	.w3(32'h3d15e093),
	.w4(32'h3c3c881f),
	.w5(32'h3c3ff13a),
	.w6(32'h3be6552b),
	.w7(32'hb96f6734),
	.w8(32'hbbb751dd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0388a3),
	.w1(32'hbb66ef33),
	.w2(32'hbc404d64),
	.w3(32'h3be50d3d),
	.w4(32'hbb64157a),
	.w5(32'hbc0e1990),
	.w6(32'hbc83e339),
	.w7(32'hbc36548c),
	.w8(32'hbc81a57c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020d38),
	.w1(32'hbc99a1c1),
	.w2(32'hbc78337e),
	.w3(32'hbac4e064),
	.w4(32'hbc5056c3),
	.w5(32'h3b65b67b),
	.w6(32'hbc6455b3),
	.w7(32'hbc90d4e6),
	.w8(32'hbc39d159),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccee5c1),
	.w1(32'h3ca7f31a),
	.w2(32'h3b8321ec),
	.w3(32'hbc4e205d),
	.w4(32'h3c0cb0e1),
	.w5(32'hbc6cd51e),
	.w6(32'h3c558291),
	.w7(32'h3cb17531),
	.w8(32'h3c1bae8a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc521f36),
	.w1(32'hbcae3afa),
	.w2(32'hba16db2c),
	.w3(32'hbc913cc4),
	.w4(32'h39fb9501),
	.w5(32'h3c5669c9),
	.w6(32'hbccdc7d8),
	.w7(32'hbceaab66),
	.w8(32'hbc4aaa0a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee59e2),
	.w1(32'hbbf23074),
	.w2(32'hbbc64979),
	.w3(32'h3c437f13),
	.w4(32'hbbb8194e),
	.w5(32'h3c18e4d5),
	.w6(32'hbb203019),
	.w7(32'h3b37922d),
	.w8(32'hbb4d739d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf66476),
	.w1(32'h3c1413ae),
	.w2(32'h3bfd29fe),
	.w3(32'h3b896f46),
	.w4(32'hbb54f8bf),
	.w5(32'hbc1f1832),
	.w6(32'h3bc90786),
	.w7(32'h3b603e09),
	.w8(32'h3a3c6f83),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9751ec),
	.w1(32'hbb47f3bd),
	.w2(32'h3bef4cb0),
	.w3(32'hbced809f),
	.w4(32'hbb2a7344),
	.w5(32'h3b7490df),
	.w6(32'hbb2f5052),
	.w7(32'h3cac924e),
	.w8(32'h3c96c024),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc597c16),
	.w1(32'h3c3d7c7f),
	.w2(32'h3c957a4e),
	.w3(32'hbc2e5928),
	.w4(32'h3b194418),
	.w5(32'h3b86b4e3),
	.w6(32'h3c06a228),
	.w7(32'h3c863c52),
	.w8(32'h3c7fbf4f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c5eea),
	.w1(32'h3a841847),
	.w2(32'hbb468db4),
	.w3(32'hbc359f23),
	.w4(32'hbc1bc706),
	.w5(32'hbc188810),
	.w6(32'h3b8c81ec),
	.w7(32'h3b9346f2),
	.w8(32'hbbe48143),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7bdab),
	.w1(32'hbc5676c8),
	.w2(32'hbc564edf),
	.w3(32'hbc8e1d95),
	.w4(32'hba92a49c),
	.w5(32'h3be31921),
	.w6(32'hbb0d0aa7),
	.w7(32'hbc07f13f),
	.w8(32'hbb9ed6d9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27cacd),
	.w1(32'h3c3cb3f2),
	.w2(32'h3b460504),
	.w3(32'h3ba50eb3),
	.w4(32'hba459dab),
	.w5(32'hbc091354),
	.w6(32'hbc445ed4),
	.w7(32'hba15bff3),
	.w8(32'h3b32916d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31cc6e),
	.w1(32'hbcbaccce),
	.w2(32'hbc42406c),
	.w3(32'hbc6db3f9),
	.w4(32'hbb8f7e28),
	.w5(32'h3c66417e),
	.w6(32'hbb3d2636),
	.w7(32'hbc01960f),
	.w8(32'hbbe34fbb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd03f1f),
	.w1(32'hbc863ad8),
	.w2(32'hbd0ec353),
	.w3(32'hbcc4bb54),
	.w4(32'hbca15dc6),
	.w5(32'hbc7b8847),
	.w6(32'h3c39c287),
	.w7(32'h3ccd613b),
	.w8(32'hbc8a5fab),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17ec06),
	.w1(32'hbc9f0f54),
	.w2(32'hbc4a20e4),
	.w3(32'hbccf99ee),
	.w4(32'hbc219166),
	.w5(32'h3ccfa8cd),
	.w6(32'hbcb05cb6),
	.w7(32'h3c43d5f0),
	.w8(32'h3c96c4b1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ec7a0),
	.w1(32'h3c98be56),
	.w2(32'h3c7a3133),
	.w3(32'hbbd434b7),
	.w4(32'hbb04e342),
	.w5(32'hbc5b919f),
	.w6(32'h3bd17401),
	.w7(32'h3c9a2662),
	.w8(32'h3c7afcfc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c135f3e),
	.w1(32'h3c0b51c4),
	.w2(32'h3b189ca5),
	.w3(32'hbc8f6f84),
	.w4(32'h3af8acb7),
	.w5(32'hbc405c5a),
	.w6(32'h3c5ae402),
	.w7(32'h3c81314d),
	.w8(32'h3c183cb8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b410c),
	.w1(32'hbbf72bab),
	.w2(32'h3c6d6d3a),
	.w3(32'hbc8ac539),
	.w4(32'h3bc38fbf),
	.w5(32'h3c6f0c00),
	.w6(32'hbc670d00),
	.w7(32'hbcb7829b),
	.w8(32'hbc075f45),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb72996),
	.w1(32'h3aef6dfd),
	.w2(32'hbb19ec1a),
	.w3(32'hbb7ae48a),
	.w4(32'hbc30c1e6),
	.w5(32'hbc9ab66a),
	.w6(32'h3b3d6b64),
	.w7(32'h3c33a961),
	.w8(32'h3bee12eb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a8f7f),
	.w1(32'hbc033fb9),
	.w2(32'hbb9c1840),
	.w3(32'hbcba0965),
	.w4(32'hbc20445c),
	.w5(32'h3c4714df),
	.w6(32'h3bc0bcdc),
	.w7(32'h3b277f24),
	.w8(32'hb95380e6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf80ee),
	.w1(32'hba2d96ee),
	.w2(32'hbafeee6c),
	.w3(32'hba4f3bec),
	.w4(32'hbba1ed70),
	.w5(32'h3c04d44c),
	.w6(32'hbaeb309f),
	.w7(32'hbc109014),
	.w8(32'hbbff9178),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7152ad),
	.w1(32'h3a9b45c0),
	.w2(32'h3c0812c2),
	.w3(32'h3b1cef83),
	.w4(32'h3b6408f9),
	.w5(32'h3b0b3bf2),
	.w6(32'h3b0b342d),
	.w7(32'h3b882250),
	.w8(32'hb9d3ff87),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7b5ad),
	.w1(32'h3bd1a0c8),
	.w2(32'hb9cc35a4),
	.w3(32'hbb375ef7),
	.w4(32'hbad00528),
	.w5(32'hbbf0c559),
	.w6(32'hbc1b3a89),
	.w7(32'hbbdcfe3b),
	.w8(32'hbb699011),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7568c9),
	.w1(32'hbb7173c6),
	.w2(32'h3baab1cb),
	.w3(32'hbc0f844d),
	.w4(32'h3b19f29f),
	.w5(32'h3b887be0),
	.w6(32'h39d1594a),
	.w7(32'h3bce653f),
	.w8(32'h3bf1f275),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4aeba),
	.w1(32'h3c163a67),
	.w2(32'hb968a92d),
	.w3(32'hbb0299d7),
	.w4(32'hbc02a123),
	.w5(32'hbcc6a4a5),
	.w6(32'h3c7c73db),
	.w7(32'h3cb4fca8),
	.w8(32'h3c617d5f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0619cf),
	.w1(32'h3b981e3a),
	.w2(32'h3aeece54),
	.w3(32'hbc9a270d),
	.w4(32'hbbf63e74),
	.w5(32'hbc4ea7b0),
	.w6(32'h3c4f5b67),
	.w7(32'h3cb1cc47),
	.w8(32'h3c981550),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc929a62),
	.w1(32'hbc4da719),
	.w2(32'hbc0d8ba8),
	.w3(32'hbcdf07e6),
	.w4(32'hbb53393c),
	.w5(32'h3c0c40fd),
	.w6(32'hbc060637),
	.w7(32'hbba81fad),
	.w8(32'hba6a40f7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cfb10),
	.w1(32'h3ba331f3),
	.w2(32'h3a607e01),
	.w3(32'hbc0c2d3e),
	.w4(32'h3bcc4a57),
	.w5(32'hba8d167e),
	.w6(32'h3b9abda3),
	.w7(32'h3b4c0f99),
	.w8(32'hbb9abc51),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a672282),
	.w1(32'hbb807069),
	.w2(32'h3b2e991a),
	.w3(32'h3bd2130e),
	.w4(32'h3ba49f99),
	.w5(32'h3b8e12b6),
	.w6(32'h3b0d2d88),
	.w7(32'h3b024fe5),
	.w8(32'h3be59a3f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c053fd8),
	.w1(32'h3ba3b104),
	.w2(32'h3c5d530a),
	.w3(32'h3c150ca0),
	.w4(32'h3c277530),
	.w5(32'h3c5fee5b),
	.w6(32'hbc186a7a),
	.w7(32'hbb9c0bf9),
	.w8(32'hbb6556f7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5c9e4),
	.w1(32'hbba84c87),
	.w2(32'hbbaf4e2b),
	.w3(32'h3b1d65a4),
	.w4(32'h38786f8a),
	.w5(32'hbb80f8c7),
	.w6(32'h3b36d1c3),
	.w7(32'hb74fdea0),
	.w8(32'h3b314ad7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc070bce),
	.w1(32'hbb8a6ea3),
	.w2(32'hbc034136),
	.w3(32'h3b06a3f7),
	.w4(32'hbc4a14d3),
	.w5(32'hbc7c183e),
	.w6(32'h3a520402),
	.w7(32'h3b11821e),
	.w8(32'h3c372b6c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cfea9),
	.w1(32'h3b1613e0),
	.w2(32'h3b61228e),
	.w3(32'hbaf86d5c),
	.w4(32'hbaa17b3b),
	.w5(32'hbab0f39d),
	.w6(32'hb9fb8e77),
	.w7(32'hbbbda11d),
	.w8(32'h3b9d285d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfe68d),
	.w1(32'hbc3a6608),
	.w2(32'hbc9dcf8b),
	.w3(32'h3a889e1e),
	.w4(32'h3baf335e),
	.w5(32'h3c29414f),
	.w6(32'hbc25d684),
	.w7(32'hbc97b072),
	.w8(32'hbca6088c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6e531),
	.w1(32'h3b0a1b2e),
	.w2(32'h3c189643),
	.w3(32'h3cb528b1),
	.w4(32'hb98d56f6),
	.w5(32'h3c006377),
	.w6(32'h3b0b2df3),
	.w7(32'hbbc353ac),
	.w8(32'hbbe73844),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfa3e2),
	.w1(32'hbbe712f4),
	.w2(32'hbb91b43d),
	.w3(32'h3b552424),
	.w4(32'hbbc4d6a2),
	.w5(32'h3a40ec2b),
	.w6(32'hbc2f3230),
	.w7(32'h3b80a8fe),
	.w8(32'h3c526bb4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1aa5da),
	.w1(32'hba9ceace),
	.w2(32'h3c1c850a),
	.w3(32'hbb7e7adb),
	.w4(32'hbbae65db),
	.w5(32'hbc4e4350),
	.w6(32'h39367e40),
	.w7(32'h3c8d6d85),
	.w8(32'h3bedd3da),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20d1e4),
	.w1(32'hbc796399),
	.w2(32'hbb805bf5),
	.w3(32'hbc006719),
	.w4(32'hbbd3544f),
	.w5(32'h3c510a26),
	.w6(32'hbc08f6d4),
	.w7(32'hbb89c133),
	.w8(32'hbb8781fb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c478382),
	.w1(32'h3bf9c485),
	.w2(32'h3b9cc256),
	.w3(32'h3c905453),
	.w4(32'hbb1c8acb),
	.w5(32'hbc18a3c3),
	.w6(32'h3b8c5e32),
	.w7(32'h3c1d0a94),
	.w8(32'h3c0361e8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eb44f),
	.w1(32'h3a06dc2b),
	.w2(32'h3bfb9104),
	.w3(32'hbc64efed),
	.w4(32'h3a84981d),
	.w5(32'h3b80f504),
	.w6(32'hbbd13877),
	.w7(32'h39612894),
	.w8(32'h3b8c4c2f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93dc0e3),
	.w1(32'h3c06d5be),
	.w2(32'hbbc84600),
	.w3(32'hbbebb133),
	.w4(32'h3c6d9049),
	.w5(32'h3ae91c27),
	.w6(32'hbb371665),
	.w7(32'hbbdf3825),
	.w8(32'hbbf91cb6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb127d19),
	.w1(32'hb9933139),
	.w2(32'hbb0af10e),
	.w3(32'h3c0d23f8),
	.w4(32'hba34a265),
	.w5(32'hbbaa8372),
	.w6(32'hb95ddbcd),
	.w7(32'h3b777e9d),
	.w8(32'hbacc30b0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c073a9b),
	.w1(32'h3bdfd13c),
	.w2(32'h3c038011),
	.w3(32'h3b0554ed),
	.w4(32'hbbd17bc4),
	.w5(32'hb8b38b3d),
	.w6(32'h3b8ceb6a),
	.w7(32'h3ba06d99),
	.w8(32'hb9bb2ec4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b9b40),
	.w1(32'hbb84fd82),
	.w2(32'h3cf977c8),
	.w3(32'hbab7c655),
	.w4(32'h3c4d541b),
	.w5(32'h3cc2d82a),
	.w6(32'hbc43e585),
	.w7(32'hbc05d768),
	.w8(32'h3bac7a38),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17d4b6),
	.w1(32'h3b779fc5),
	.w2(32'hba880501),
	.w3(32'h3c204297),
	.w4(32'hbc2d42e3),
	.w5(32'hbc8c5661),
	.w6(32'h3bfbbc88),
	.w7(32'h3bfda39d),
	.w8(32'h3be02aeb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20fd38),
	.w1(32'hba71985b),
	.w2(32'h3b2eb56a),
	.w3(32'hbca2e465),
	.w4(32'hba85e4e9),
	.w5(32'hbb27be8f),
	.w6(32'hbb63a72a),
	.w7(32'hb8eb4df8),
	.w8(32'h3a3b657c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b677861),
	.w1(32'hba6a8752),
	.w2(32'h3b695018),
	.w3(32'hbbc2a346),
	.w4(32'h3c9715bd),
	.w5(32'h3d04c056),
	.w6(32'hbc61cbb7),
	.w7(32'hbc6f4729),
	.w8(32'hbc97b169),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a6218),
	.w1(32'hbb61fbf4),
	.w2(32'h3ae6df1a),
	.w3(32'h3d101502),
	.w4(32'hbb1aef64),
	.w5(32'h3b66b1ee),
	.w6(32'hbb9269c9),
	.w7(32'h3b6898cf),
	.w8(32'h3b5ab1ef),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5331a9),
	.w1(32'hbc1e77b1),
	.w2(32'hbbb75fea),
	.w3(32'hbaee7253),
	.w4(32'hbc26c5e0),
	.w5(32'hbc6b5347),
	.w6(32'hbbdc51c5),
	.w7(32'hbc58879a),
	.w8(32'hbb85f002),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a5b83),
	.w1(32'hbc642cba),
	.w2(32'hbb47f305),
	.w3(32'hbbb56c60),
	.w4(32'h3b7ebf3e),
	.w5(32'h3c3bad44),
	.w6(32'hbc57d9e7),
	.w7(32'hbc8dad19),
	.w8(32'hbb6532f4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cd69a),
	.w1(32'h3bda8af8),
	.w2(32'h3bc786e1),
	.w3(32'h3c4b931e),
	.w4(32'h3b4c967a),
	.w5(32'h3c0a2064),
	.w6(32'h3c1a8fce),
	.w7(32'h3c03e2b6),
	.w8(32'h3c21c362),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c07fc),
	.w1(32'hbc2e74e9),
	.w2(32'hba8fef10),
	.w3(32'hbc9b511b),
	.w4(32'hbbde0d39),
	.w5(32'h3c4020c1),
	.w6(32'hbc10a83d),
	.w7(32'hbc0e9a95),
	.w8(32'hbb5132bd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4fa83),
	.w1(32'hbb14c038),
	.w2(32'h3b1974ae),
	.w3(32'h3b8d9b08),
	.w4(32'hbb137710),
	.w5(32'hbb2169f8),
	.w6(32'hbb8c5186),
	.w7(32'hbb17816e),
	.w8(32'h38901013),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29589c),
	.w1(32'h3aa11141),
	.w2(32'h3b6e116b),
	.w3(32'hbb978e44),
	.w4(32'hbb474820),
	.w5(32'h39748b2e),
	.w6(32'hba35b4b5),
	.w7(32'hbb1dbf29),
	.w8(32'hbb1d66d3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558682),
	.w1(32'h39412c30),
	.w2(32'h3c202a26),
	.w3(32'hbbd19325),
	.w4(32'h3c6aba52),
	.w5(32'h3cf91eec),
	.w6(32'h3a8677ad),
	.w7(32'h3b8431ec),
	.w8(32'h3b9f7d9e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c166762),
	.w1(32'hbb940f1c),
	.w2(32'hbc5648d6),
	.w3(32'h3cbca6e7),
	.w4(32'hbc9a63a6),
	.w5(32'hbc474a4e),
	.w6(32'h3b85f110),
	.w7(32'hbbc7c583),
	.w8(32'h3a5e5d00),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d499e),
	.w1(32'hbabb89d6),
	.w2(32'h3b8b13b1),
	.w3(32'hbb97f4f8),
	.w4(32'h3b01ffda),
	.w5(32'h3bbea85d),
	.w6(32'hb872d543),
	.w7(32'h3a86ab24),
	.w8(32'h3ae1c2f1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ea7e3),
	.w1(32'hbc016c1a),
	.w2(32'hbba9de7f),
	.w3(32'hbbad85e5),
	.w4(32'hbbef4773),
	.w5(32'hbbc9286b),
	.w6(32'hbb01ad43),
	.w7(32'hbbd8b686),
	.w8(32'h3c2c8d78),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule