module layer_8_featuremap_190(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d0916),
	.w1(32'hbc15f797),
	.w2(32'hbc423576),
	.w3(32'h3bd454ad),
	.w4(32'h3b276c0f),
	.w5(32'h3b0e7607),
	.w6(32'hbbd6e08c),
	.w7(32'hbb2aa4e7),
	.w8(32'h3b09e674),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba15111),
	.w1(32'h3aa63241),
	.w2(32'h3b697e6d),
	.w3(32'h3be5c304),
	.w4(32'hba90a61f),
	.w5(32'hbade6367),
	.w6(32'h3a13de4f),
	.w7(32'h3a1bc51c),
	.w8(32'h3b3a1799),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5890d),
	.w1(32'hbb500642),
	.w2(32'h3b16c31b),
	.w3(32'h39e6e85d),
	.w4(32'h3c8fb872),
	.w5(32'h3c54c646),
	.w6(32'h3bd112fb),
	.w7(32'h3886fc97),
	.w8(32'hbbf7ca75),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca03924),
	.w1(32'hb8a278f8),
	.w2(32'hbb35b5c3),
	.w3(32'h3c2bbf2c),
	.w4(32'h3c10ef81),
	.w5(32'h3c82b17f),
	.w6(32'h3b8d4fcd),
	.w7(32'h3c4a44b5),
	.w8(32'h3b27b701),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89fafc),
	.w1(32'hbbcf2379),
	.w2(32'hbba331bb),
	.w3(32'h3cdf5f39),
	.w4(32'hbac7a619),
	.w5(32'hba29a2b8),
	.w6(32'h3a738ee1),
	.w7(32'hbaaa36e4),
	.w8(32'hbaebbdc2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82844b),
	.w1(32'hbb654900),
	.w2(32'hbc7aa6e7),
	.w3(32'hbb0e2e55),
	.w4(32'hbc967aa8),
	.w5(32'hbc428e3e),
	.w6(32'hbbb6cb6a),
	.w7(32'hbb41bfa8),
	.w8(32'h3af2783c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e05ff),
	.w1(32'hbaa6b91b),
	.w2(32'hbb3f31dd),
	.w3(32'hb9c83e7a),
	.w4(32'h3a592667),
	.w5(32'hba8680b9),
	.w6(32'h3b3c711d),
	.w7(32'h3a093ae1),
	.w8(32'hba8d4190),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fd0b9),
	.w1(32'hbc7b4214),
	.w2(32'hbd112935),
	.w3(32'hbad533ab),
	.w4(32'h398075bc),
	.w5(32'h3d1f5320),
	.w6(32'h3c7f2886),
	.w7(32'h3ca10d38),
	.w8(32'h3a696a8b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ff161),
	.w1(32'hbbe0794a),
	.w2(32'hbb7701fd),
	.w3(32'h3d50ff7c),
	.w4(32'h3b2e6f32),
	.w5(32'h3a93c611),
	.w6(32'hbb6c3cbe),
	.w7(32'hbbf3e442),
	.w8(32'hbbbf4ae8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b963c),
	.w1(32'hbc1e89f4),
	.w2(32'hb9ed63b5),
	.w3(32'hbaf78380),
	.w4(32'hba9b0a30),
	.w5(32'hbc8c1e64),
	.w6(32'hbc2a9807),
	.w7(32'hbc014cfe),
	.w8(32'hba35f488),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1dbc7),
	.w1(32'hbb97e71b),
	.w2(32'h390062ac),
	.w3(32'hbc8ca326),
	.w4(32'h37d0e0d9),
	.w5(32'h3bec3b99),
	.w6(32'hbb410b88),
	.w7(32'hbb9d1822),
	.w8(32'hbc03faf8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb22bd),
	.w1(32'hbadb2971),
	.w2(32'hba00fbec),
	.w3(32'h3c07862e),
	.w4(32'hbb6eeda4),
	.w5(32'hba1c14c5),
	.w6(32'hba8c4727),
	.w7(32'hbbec75c6),
	.w8(32'hbb715f41),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba848298),
	.w1(32'h3ba0d0d6),
	.w2(32'hb9dc127b),
	.w3(32'h3b8dbafd),
	.w4(32'hbb601bc6),
	.w5(32'hbc09a1de),
	.w6(32'h3b4e5a65),
	.w7(32'h3b663b99),
	.w8(32'h3b824d32),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12a28d),
	.w1(32'hbb468199),
	.w2(32'hbc3dd67f),
	.w3(32'h3b4a82d4),
	.w4(32'hbc595aca),
	.w5(32'hbcd7dec4),
	.w6(32'h3ae27e68),
	.w7(32'hbb2d25ef),
	.w8(32'h3c140b36),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d9315),
	.w1(32'h3836ad0d),
	.w2(32'hbacebb16),
	.w3(32'hbd018f92),
	.w4(32'h3b02c31a),
	.w5(32'hba3c2d40),
	.w6(32'hbb15c146),
	.w7(32'hbadd0cae),
	.w8(32'hbb46f9bf),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f88ff),
	.w1(32'hbc3c6546),
	.w2(32'hbb1cfe03),
	.w3(32'hbb3f1a6c),
	.w4(32'h3c51d6b3),
	.w5(32'hbb10fe3c),
	.w6(32'hbb88ebbe),
	.w7(32'hbc77ea82),
	.w8(32'hbc46a49f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc022440),
	.w1(32'h3c1c7c5b),
	.w2(32'h3c03b002),
	.w3(32'hbb3c6dd0),
	.w4(32'hbc35ddb0),
	.w5(32'hbc5cee27),
	.w6(32'hbaf127e3),
	.w7(32'h3b36f65f),
	.w8(32'h3c44b8c9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02b2d5),
	.w1(32'h3bf3cd4e),
	.w2(32'h3bc4affb),
	.w3(32'h3a70cf7c),
	.w4(32'hbb384369),
	.w5(32'hbbe8f0dc),
	.w6(32'hbc25f7a2),
	.w7(32'hbc2ef1de),
	.w8(32'hbbb4047e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22839b),
	.w1(32'h3c2e22d1),
	.w2(32'h3b0dbe64),
	.w3(32'h3b7c46fd),
	.w4(32'hbc7f138b),
	.w5(32'hbcaf0b2f),
	.w6(32'hbadae085),
	.w7(32'h38f7d253),
	.w8(32'h3bf0ad6f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21b923),
	.w1(32'h3ba4814d),
	.w2(32'h3a84c12e),
	.w3(32'hbc418283),
	.w4(32'h3b1ffa93),
	.w5(32'h394db2ef),
	.w6(32'h3b0c3926),
	.w7(32'h3a92a12c),
	.w8(32'hb9a4260f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02d176),
	.w1(32'hbbc88a45),
	.w2(32'hbb3153fc),
	.w3(32'h3a2a832f),
	.w4(32'h3c04c0fc),
	.w5(32'h3b2c7680),
	.w6(32'hbb10e9c5),
	.w7(32'hbbb7f1d5),
	.w8(32'hbbe90347),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b7e1a),
	.w1(32'hbbdb1749),
	.w2(32'hbca0fdde),
	.w3(32'hbb738c28),
	.w4(32'hbbb1d4ca),
	.w5(32'hbc6658cb),
	.w6(32'h3b04d723),
	.w7(32'h3ad76df4),
	.w8(32'hbba6e4d4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83724b),
	.w1(32'hbbd42d3d),
	.w2(32'hba0e9ef7),
	.w3(32'hbc5918f4),
	.w4(32'hbc33b949),
	.w5(32'hbcd06a1f),
	.w6(32'hbbc7eb0d),
	.w7(32'hbc680ff2),
	.w8(32'hbb2fa75b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf13973),
	.w1(32'hbb8407fd),
	.w2(32'hbc611267),
	.w3(32'hbcbd7cb5),
	.w4(32'hbc734f21),
	.w5(32'hbc585221),
	.w6(32'h3bcad809),
	.w7(32'h3c13e357),
	.w8(32'hba0c9acf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4339da),
	.w1(32'h3a142056),
	.w2(32'h3bfe1981),
	.w3(32'hbaf4ff26),
	.w4(32'h3c1bb1d0),
	.w5(32'h3bfbdca3),
	.w6(32'hbba8046b),
	.w7(32'hbb8666bd),
	.w8(32'hbae324d3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5fa018),
	.w1(32'hbb1cea43),
	.w2(32'hba799b38),
	.w3(32'hbc056b2e),
	.w4(32'h3b97a6eb),
	.w5(32'hba414792),
	.w6(32'hba997799),
	.w7(32'hbb81721f),
	.w8(32'hbb9fa26f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c286b50),
	.w1(32'hbb849bac),
	.w2(32'hbc236bf2),
	.w3(32'hbbaa40db),
	.w4(32'h38431dd4),
	.w5(32'h3d24a60f),
	.w6(32'hbb24be22),
	.w7(32'hbafb088a),
	.w8(32'hbb7cd597),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6aa9e6),
	.w1(32'h3c66a56d),
	.w2(32'h3b816fe8),
	.w3(32'h3d585246),
	.w4(32'hbc0d86c3),
	.w5(32'hbc3695eb),
	.w6(32'hbb4ed2a0),
	.w7(32'h3b9c0ba9),
	.w8(32'h3c380b84),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ed984),
	.w1(32'h3bb247c9),
	.w2(32'hbb631411),
	.w3(32'hba2e9cae),
	.w4(32'h3b9b7d64),
	.w5(32'hbb62c596),
	.w6(32'hbb0ce16e),
	.w7(32'hbb6bb5c1),
	.w8(32'hb947ea81),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0746b),
	.w1(32'hbb8f3645),
	.w2(32'hbb57283b),
	.w3(32'hbaacfe7a),
	.w4(32'hbb4e779f),
	.w5(32'h3a9d59b1),
	.w6(32'hbb249b94),
	.w7(32'hbab72d81),
	.w8(32'hbabca545),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3958afd5),
	.w1(32'hbbc4425e),
	.w2(32'hbc17d135),
	.w3(32'h39ff1581),
	.w4(32'h3ae830bc),
	.w5(32'h3b7d449f),
	.w6(32'h3b7da083),
	.w7(32'h3b763ac8),
	.w8(32'h3b57eb82),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1498ac),
	.w1(32'h3bbb8819),
	.w2(32'h3bdfab51),
	.w3(32'h3b072144),
	.w4(32'hbc22fa33),
	.w5(32'hbc6df2c3),
	.w6(32'hbc6444bd),
	.w7(32'hbc079173),
	.w8(32'h3b8ea31b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9f682),
	.w1(32'hbb104321),
	.w2(32'hbbd3bc7b),
	.w3(32'hbb8176c4),
	.w4(32'hbc4141fc),
	.w5(32'hbca99e53),
	.w6(32'hbc55ae40),
	.w7(32'hbbd13122),
	.w8(32'hbad804c0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a5cba),
	.w1(32'h3c35e128),
	.w2(32'h3bd851fc),
	.w3(32'hbc4cf6dd),
	.w4(32'h3b724da1),
	.w5(32'hbb5b18f1),
	.w6(32'h3a8eca85),
	.w7(32'h3bdfbc90),
	.w8(32'h3c11be81),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab72b4),
	.w1(32'hbb7c30a5),
	.w2(32'hbbf1c880),
	.w3(32'hbba19958),
	.w4(32'h3b4534e0),
	.w5(32'h3bf24b91),
	.w6(32'h3b9989dd),
	.w7(32'hbacb91b6),
	.w8(32'hbb13ec1c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96904f),
	.w1(32'hbc231e11),
	.w2(32'hbbff5e7a),
	.w3(32'h3c02c476),
	.w4(32'h3c15f078),
	.w5(32'h3d321977),
	.w6(32'h3ad46e1e),
	.w7(32'h3b4465e5),
	.w8(32'hbae46ef6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4c55f),
	.w1(32'hb9ee0266),
	.w2(32'h3a8b565c),
	.w3(32'h3cfeb4a4),
	.w4(32'hbb10a1f4),
	.w5(32'hbae924d2),
	.w6(32'hba2c6866),
	.w7(32'h3896e1e5),
	.w8(32'h3b334bc3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a267f9d),
	.w1(32'h39e57b0d),
	.w2(32'h3b18e147),
	.w3(32'hbb3b8d3b),
	.w4(32'h3af888c2),
	.w5(32'h3a0acfd9),
	.w6(32'h3b5c55e7),
	.w7(32'h3b9b7912),
	.w8(32'h3b0e8d86),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78db37),
	.w1(32'h3c69c490),
	.w2(32'h3c2b50f9),
	.w3(32'hb9a48ca1),
	.w4(32'h3a378c84),
	.w5(32'hbb63580b),
	.w6(32'h3be5a94f),
	.w7(32'h3c373b58),
	.w8(32'h3bf678f3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50b218),
	.w1(32'hbbbe2c00),
	.w2(32'hbc75365a),
	.w3(32'h3c16ad9e),
	.w4(32'hbbafb0e3),
	.w5(32'hbbecb59e),
	.w6(32'h3b6dc2fa),
	.w7(32'h3bbf94f9),
	.w8(32'hbadd5c95),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc003ea2),
	.w1(32'hbb170707),
	.w2(32'hbb0ac945),
	.w3(32'hbc48bea7),
	.w4(32'hbb88e430),
	.w5(32'hbaf3088d),
	.w6(32'hbb2532d4),
	.w7(32'hbb1962eb),
	.w8(32'hbae33013),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba882226),
	.w1(32'h3af2941a),
	.w2(32'h3a99dce8),
	.w3(32'hb56ddd18),
	.w4(32'hbbe89a6c),
	.w5(32'hbbe260c0),
	.w6(32'h3a6c083c),
	.w7(32'h39f5dfa9),
	.w8(32'hb9af9650),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d62a2),
	.w1(32'h3bf0eea4),
	.w2(32'h3bc9ec0f),
	.w3(32'h3bb3b2bd),
	.w4(32'hbbdc151a),
	.w5(32'hbb8bdb38),
	.w6(32'hbae2bd9e),
	.w7(32'h3a06573e),
	.w8(32'h3b7a42a5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cce32d),
	.w1(32'h3ac9963f),
	.w2(32'hb858ee2a),
	.w3(32'hb70605e8),
	.w4(32'hbc0cc3e1),
	.w5(32'hbc516411),
	.w6(32'hbc479c67),
	.w7(32'hbc1e4bfb),
	.w8(32'hbc1f8037),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d7cfb),
	.w1(32'hbc5b3c1f),
	.w2(32'hbbf7ff2c),
	.w3(32'hba90c1c7),
	.w4(32'h3c465c61),
	.w5(32'h3c64f75f),
	.w6(32'h3bf9c8e0),
	.w7(32'hbbd9fd7c),
	.w8(32'hbaf56e0e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9e692),
	.w1(32'h3b903f22),
	.w2(32'hbb0a21ea),
	.w3(32'hbbb70649),
	.w4(32'h3a1933a6),
	.w5(32'hbb67d078),
	.w6(32'hba42400b),
	.w7(32'hbb3c62c6),
	.w8(32'hbb10ded1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72b7b4),
	.w1(32'h39d079be),
	.w2(32'hba4fa068),
	.w3(32'hbb5f06c5),
	.w4(32'hbc08e4d6),
	.w5(32'hbc31191b),
	.w6(32'h3bbe2877),
	.w7(32'h3a7b9e2e),
	.w8(32'h3b22e7f3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c6101),
	.w1(32'hbc8069cb),
	.w2(32'h3b9d3063),
	.w3(32'hbc1aa1f2),
	.w4(32'h3cc3043c),
	.w5(32'h3d077d40),
	.w6(32'hbbce605a),
	.w7(32'hbb0dd0ec),
	.w8(32'hbc610e2d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8c7eb),
	.w1(32'hbc87a476),
	.w2(32'h3a083f8f),
	.w3(32'h3c758190),
	.w4(32'h3d121912),
	.w5(32'h3d2ad7d5),
	.w6(32'hba946e16),
	.w7(32'hb8f572c5),
	.w8(32'hbbdea216),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb91941),
	.w1(32'h3ba488fd),
	.w2(32'h3bb1fd85),
	.w3(32'h3c6cb95e),
	.w4(32'hbc117b01),
	.w5(32'hbc33a845),
	.w6(32'h3ab40244),
	.w7(32'hbb126de9),
	.w8(32'h3a6741af),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17df5c),
	.w1(32'h3bf8f419),
	.w2(32'h3b8466b5),
	.w3(32'hba6aaba3),
	.w4(32'hba5b6c9c),
	.w5(32'hb92276d2),
	.w6(32'hb961b81f),
	.w7(32'hbaf21bc1),
	.w8(32'h3ae8d421),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc552c7),
	.w1(32'h3b840a00),
	.w2(32'h3a90ea8a),
	.w3(32'h3a683e1d),
	.w4(32'hbbebff42),
	.w5(32'hbc17aea1),
	.w6(32'hbb08014e),
	.w7(32'hbba158c4),
	.w8(32'hb9954de8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29df86),
	.w1(32'hba4c0933),
	.w2(32'h3b7a3b58),
	.w3(32'h3b6bce79),
	.w4(32'hbb7861b2),
	.w5(32'hbb24642f),
	.w6(32'hbad8dd8c),
	.w7(32'h3aaa77d5),
	.w8(32'h3b19a7b2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b8399),
	.w1(32'h3b89f7a6),
	.w2(32'hbb40ffeb),
	.w3(32'hb9ee6b07),
	.w4(32'hbbe5bafa),
	.w5(32'hbbcc9617),
	.w6(32'h3b23b9f1),
	.w7(32'h3b5a02bd),
	.w8(32'h3b0a370f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40a6bb),
	.w1(32'h3c44cfb2),
	.w2(32'h39d78ccd),
	.w3(32'hbc058519),
	.w4(32'hba20c257),
	.w5(32'hbc2f96d7),
	.w6(32'hb9ea4743),
	.w7(32'h3ba7ead9),
	.w8(32'h3c0e9d22),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc001fb5),
	.w1(32'hbc2a34d0),
	.w2(32'hbbe45ea4),
	.w3(32'h3b870a64),
	.w4(32'hbc0ff66a),
	.w5(32'hbc000ea5),
	.w6(32'hbc2adacb),
	.w7(32'hbc734537),
	.w8(32'hbc24180c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51aeaa),
	.w1(32'hbc300ad2),
	.w2(32'hbc973a43),
	.w3(32'hbb420070),
	.w4(32'h3a91d127),
	.w5(32'h3ab51c5f),
	.w6(32'h3b52e528),
	.w7(32'hbb018b7f),
	.w8(32'hbbafbd45),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d30d6),
	.w1(32'h3a6c2452),
	.w2(32'hb9dc0628),
	.w3(32'hbadb4a4f),
	.w4(32'hb999eb0d),
	.w5(32'hb87a1ba5),
	.w6(32'hbb3fe7de),
	.w7(32'hb993a550),
	.w8(32'h3ad733bd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb322aa8),
	.w1(32'h3a5112a8),
	.w2(32'hb8e3c263),
	.w3(32'hba879531),
	.w4(32'h3a6041d2),
	.w5(32'hbb295864),
	.w6(32'hb9c48aed),
	.w7(32'hbaa6642f),
	.w8(32'hba37d04f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf54f22),
	.w1(32'h3bf7dd4d),
	.w2(32'hbc0a1dd6),
	.w3(32'hbadd8068),
	.w4(32'hbb800608),
	.w5(32'hbbfc31de),
	.w6(32'h3c3fe156),
	.w7(32'h3c446a47),
	.w8(32'hbbf35a9f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b257d93),
	.w1(32'h3b9e9f38),
	.w2(32'h3bcd11f0),
	.w3(32'hbbe0832a),
	.w4(32'h3be5c5d7),
	.w5(32'h3a2b8a17),
	.w6(32'hbb9b546c),
	.w7(32'hbbc8dec2),
	.w8(32'hbb3e45f4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf42794),
	.w1(32'h3ab99ba2),
	.w2(32'h3b856c20),
	.w3(32'h3baaea16),
	.w4(32'h3b635fdf),
	.w5(32'hbb89e916),
	.w6(32'h3c4286bb),
	.w7(32'h3ba68cc8),
	.w8(32'h3bb02aca),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8b5ea),
	.w1(32'h3b8ab9ae),
	.w2(32'h3ba6ee75),
	.w3(32'hbc01e451),
	.w4(32'h3a10ecd4),
	.w5(32'h3b812bd1),
	.w6(32'hba94f6f8),
	.w7(32'hbb47b2fb),
	.w8(32'h3b20c87f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b39dd5),
	.w1(32'hbaeb22d6),
	.w2(32'hbb1d8ba3),
	.w3(32'h3c10f547),
	.w4(32'hbb3e3194),
	.w5(32'h3b2b4b97),
	.w6(32'h38bab5c1),
	.w7(32'hbab66f6e),
	.w8(32'hbb1b2ecb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d431b),
	.w1(32'h3bddea31),
	.w2(32'h3b8fa3cd),
	.w3(32'h3a8258c6),
	.w4(32'hb9cef94e),
	.w5(32'h3aa6f196),
	.w6(32'hba31cc54),
	.w7(32'h3affcc3b),
	.w8(32'h3ab3f303),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2d24e),
	.w1(32'hbc4c2eb3),
	.w2(32'hbc33c775),
	.w3(32'h3b82f759),
	.w4(32'hbc928c37),
	.w5(32'hbc414fda),
	.w6(32'hba10e84d),
	.w7(32'hbb99657c),
	.w8(32'hbb3d4da4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04f98f),
	.w1(32'h3abe8104),
	.w2(32'h3ca449e2),
	.w3(32'hbc0316d7),
	.w4(32'h3c6169ae),
	.w5(32'hbbfaf731),
	.w6(32'hbc6b8146),
	.w7(32'hbca338f1),
	.w8(32'hbbffb4a6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceeee61),
	.w1(32'h3a30c7b9),
	.w2(32'hbb0083e6),
	.w3(32'hbcdc892a),
	.w4(32'hb8c1b889),
	.w5(32'hbc3a2695),
	.w6(32'hbb04ccb9),
	.w7(32'hbb12ef79),
	.w8(32'hbb49620a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9209f),
	.w1(32'h3ccaef48),
	.w2(32'h3c5c2809),
	.w3(32'hb8a69315),
	.w4(32'h3beff8d6),
	.w5(32'hb90203cb),
	.w6(32'h3bd35cf8),
	.w7(32'h3c3732e2),
	.w8(32'h3c56cdda),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c308690),
	.w1(32'h3976341b),
	.w2(32'h3bbc0e1a),
	.w3(32'h398f7a43),
	.w4(32'h3c02eec4),
	.w5(32'h3c589eb6),
	.w6(32'h3b1680dc),
	.w7(32'h3ba7abcf),
	.w8(32'hbb9bf52d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c857795),
	.w1(32'h3b7dd0f0),
	.w2(32'h3b98f23d),
	.w3(32'h3c31da14),
	.w4(32'hbb3265de),
	.w5(32'hbac91c3e),
	.w6(32'h3a0ccb7e),
	.w7(32'hbb629856),
	.w8(32'hbb3c3f1f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b333b),
	.w1(32'hbc0be497),
	.w2(32'hbb902277),
	.w3(32'h39e493ad),
	.w4(32'hb9b7dc85),
	.w5(32'hbbf5dd5e),
	.w6(32'h3a5a898c),
	.w7(32'hbbde81db),
	.w8(32'hbc679d53),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95e748),
	.w1(32'hbc63015b),
	.w2(32'hbc819cb4),
	.w3(32'hbc2a29fc),
	.w4(32'h3cb4919a),
	.w5(32'h3cbb4a20),
	.w6(32'h388a806b),
	.w7(32'h3b4e3224),
	.w8(32'hbba6efcd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23b8b2),
	.w1(32'hbb995d65),
	.w2(32'hbc18ccd9),
	.w3(32'hbb50caea),
	.w4(32'hbad74556),
	.w5(32'h3b89325d),
	.w6(32'h3be6d45e),
	.w7(32'h3bf45e72),
	.w8(32'hbbd0eaa5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc211e14),
	.w1(32'hba8b154f),
	.w2(32'hbaa4181a),
	.w3(32'h3ac1a438),
	.w4(32'h3c2e3247),
	.w5(32'h3b219e5e),
	.w6(32'hbb6183cc),
	.w7(32'h3b5d0b92),
	.w8(32'hba9236ca),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9b617),
	.w1(32'h3a5dbe2a),
	.w2(32'hbc445acd),
	.w3(32'hbb889cd2),
	.w4(32'hbc26124a),
	.w5(32'hbb9b8412),
	.w6(32'h3add18cc),
	.w7(32'h3a744850),
	.w8(32'hbaef86c3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bf4a3),
	.w1(32'h3a90ca4d),
	.w2(32'hbb6249dd),
	.w3(32'h3ad3edf8),
	.w4(32'h3b08ab3b),
	.w5(32'h3b37c3b9),
	.w6(32'h3b176a29),
	.w7(32'h3b4ce9ba),
	.w8(32'hbb6ab7bf),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb180854),
	.w1(32'hbb2b5e77),
	.w2(32'hbbf58dbc),
	.w3(32'h3bd3a62b),
	.w4(32'hbaece1ad),
	.w5(32'hbb8b9c7a),
	.w6(32'hb9ec9326),
	.w7(32'hba882242),
	.w8(32'hba3522a7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc78a24),
	.w1(32'hbb92e5da),
	.w2(32'hbc139291),
	.w3(32'h3a2c631d),
	.w4(32'hbc1ff9ff),
	.w5(32'hbb8b1b28),
	.w6(32'h3b57a2db),
	.w7(32'h3b7090f9),
	.w8(32'h3b5ef3af),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21073c),
	.w1(32'hbb9d64fc),
	.w2(32'hbc5bdafc),
	.w3(32'hbb781e24),
	.w4(32'hbc48b809),
	.w5(32'hbc4aa689),
	.w6(32'hbc7e7b28),
	.w7(32'hbc76254c),
	.w8(32'hbb30790b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37cff4),
	.w1(32'hbb9fed41),
	.w2(32'hbbf03152),
	.w3(32'hbad9594a),
	.w4(32'h3c19bb3f),
	.w5(32'h398da991),
	.w6(32'hbbe60c1c),
	.w7(32'hbacbb766),
	.w8(32'hbb8514f1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdbb54),
	.w1(32'h3c640992),
	.w2(32'h3c0ec1c5),
	.w3(32'hbbb0f36b),
	.w4(32'h3b53c76d),
	.w5(32'hbb99bb0f),
	.w6(32'h3bbfda6d),
	.w7(32'h3bed14ee),
	.w8(32'h3c7f41ec),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00226c),
	.w1(32'h3c2d6a4f),
	.w2(32'h3bbb51a7),
	.w3(32'hbb41da84),
	.w4(32'hbbef7c71),
	.w5(32'hbc1a7e4b),
	.w6(32'h3a8d9aba),
	.w7(32'hba1a7df1),
	.w8(32'h3b3c8ccd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a627d5c),
	.w1(32'h3b0a29ad),
	.w2(32'hbc08137d),
	.w3(32'hbc1fa740),
	.w4(32'hbbef627d),
	.w5(32'h3b75cde5),
	.w6(32'h3bacc735),
	.w7(32'h3b286636),
	.w8(32'hba720a61),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c934c),
	.w1(32'h37463b62),
	.w2(32'hbbd74463),
	.w3(32'h3b679c9c),
	.w4(32'hbc236f1b),
	.w5(32'hbc6eccb0),
	.w6(32'hbc3bc121),
	.w7(32'h39a9f8ff),
	.w8(32'h3b4efe62),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4a04),
	.w1(32'h3a84bd34),
	.w2(32'hbc0ec803),
	.w3(32'hbc4e4d73),
	.w4(32'h3b676bd4),
	.w5(32'h3ca98d25),
	.w6(32'h3aefc18a),
	.w7(32'h3c67e5de),
	.w8(32'h3c277693),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9308cd),
	.w1(32'hbb38d2ab),
	.w2(32'h3b21242c),
	.w3(32'h3d11985b),
	.w4(32'h3b016245),
	.w5(32'h3b812665),
	.w6(32'hb90e7e38),
	.w7(32'hbb164a5a),
	.w8(32'h38e050a6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab34106),
	.w1(32'h3b15d782),
	.w2(32'h393eab09),
	.w3(32'hbb30572b),
	.w4(32'hbc0bfbaf),
	.w5(32'hbb64b366),
	.w6(32'hbb081af8),
	.w7(32'hbb100337),
	.w8(32'hbaae2ed8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99317a5),
	.w1(32'hbbe33990),
	.w2(32'hbbd9679f),
	.w3(32'h3bb44d91),
	.w4(32'h3bb9df96),
	.w5(32'h3c0a1458),
	.w6(32'h39a58c5c),
	.w7(32'h39a2e4f0),
	.w8(32'hb90669ad),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17ff3d),
	.w1(32'h3a09843a),
	.w2(32'h3c5dc646),
	.w3(32'h3b96c591),
	.w4(32'h3ccc6251),
	.w5(32'h3d0fcf07),
	.w6(32'h3bd67529),
	.w7(32'hbb80941f),
	.w8(32'hbc4f0269),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd7c16b),
	.w1(32'hbc18bfee),
	.w2(32'hba6c205c),
	.w3(32'h3ca9bcd6),
	.w4(32'h3c9bf30e),
	.w5(32'h3c51a96f),
	.w6(32'h3bb56efd),
	.w7(32'hbbdfbbf7),
	.w8(32'hbb58651c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b846249),
	.w1(32'h3b3dd696),
	.w2(32'h3c231b22),
	.w3(32'h3b64c950),
	.w4(32'h3c18b21c),
	.w5(32'hbb0af643),
	.w6(32'h3b1b4215),
	.w7(32'h3aece8fd),
	.w8(32'h3c00a7b1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be68e49),
	.w1(32'h3aa67730),
	.w2(32'h3a136929),
	.w3(32'hbbb61941),
	.w4(32'hbb251c60),
	.w5(32'hbb2f4347),
	.w6(32'h3a722df4),
	.w7(32'hba383385),
	.w8(32'hba62f02f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6fc43),
	.w1(32'h3b284ace),
	.w2(32'h3892bf65),
	.w3(32'hbb7b83c4),
	.w4(32'hba17f42f),
	.w5(32'hbb3de7ea),
	.w6(32'h3b5b54be),
	.w7(32'h39380f01),
	.w8(32'h3a93e3d7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b4e32),
	.w1(32'h3ac31251),
	.w2(32'h3aabea3e),
	.w3(32'hbaccd420),
	.w4(32'h3c41e57a),
	.w5(32'h3bbca9f4),
	.w6(32'hbaf1725e),
	.w7(32'h3c114a6b),
	.w8(32'hb9b86915),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030857),
	.w1(32'h3a91269a),
	.w2(32'hbb74abfb),
	.w3(32'h3c19126c),
	.w4(32'hba99d2af),
	.w5(32'hbb58f642),
	.w6(32'h3aa788e9),
	.w7(32'hb8aec943),
	.w8(32'h3935091d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba979001),
	.w1(32'hb994ade3),
	.w2(32'hba68cb36),
	.w3(32'h3b43015a),
	.w4(32'hbb15a564),
	.w5(32'hbb60b226),
	.w6(32'h3afa087f),
	.w7(32'hb98fb769),
	.w8(32'hbb232314),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac59b31),
	.w1(32'h3c124b4d),
	.w2(32'h3bd73ee4),
	.w3(32'h3b176394),
	.w4(32'h3a9728ea),
	.w5(32'hbb38fba8),
	.w6(32'h3adbbcc3),
	.w7(32'h3bc68fd1),
	.w8(32'h3b9df3ee),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085fc9),
	.w1(32'h3c1e5e59),
	.w2(32'h3ba4fcc5),
	.w3(32'h3c1c45f0),
	.w4(32'h3b31bce3),
	.w5(32'h3a886d80),
	.w6(32'h3b5f4a61),
	.w7(32'h3bdedfb4),
	.w8(32'h3c05255e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2b6d0),
	.w1(32'h3bd3de3a),
	.w2(32'h3c735cec),
	.w3(32'h3c846a34),
	.w4(32'hbc7fb7a3),
	.w5(32'hbcf79859),
	.w6(32'hbc2d95fa),
	.w7(32'hba9db034),
	.w8(32'h3a9b5a29),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e4544),
	.w1(32'h3a4618fd),
	.w2(32'hba7d8734),
	.w3(32'hbc4900a6),
	.w4(32'hbc20f899),
	.w5(32'hbb851e7d),
	.w6(32'h39d38458),
	.w7(32'h3b834c57),
	.w8(32'hbbec0fec),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af03a0f),
	.w1(32'h3c432b08),
	.w2(32'h3b56c5c1),
	.w3(32'hbba0f6e5),
	.w4(32'hbbca9dae),
	.w5(32'hbc1f0916),
	.w6(32'h39d9e68d),
	.w7(32'hbba63e2a),
	.w8(32'h3c39f6f2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc154395),
	.w1(32'h3bf364fc),
	.w2(32'h3b413e03),
	.w3(32'hbad2cfe2),
	.w4(32'hbb8bec02),
	.w5(32'hbcc2b272),
	.w6(32'h3be5f295),
	.w7(32'h3c22c4e9),
	.w8(32'h3c11e613),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d72c7),
	.w1(32'h3a5702ce),
	.w2(32'h3d04443a),
	.w3(32'hbca9ac9e),
	.w4(32'h3c96dfbb),
	.w5(32'h3b1610ca),
	.w6(32'hba250745),
	.w7(32'hbc8fd6cf),
	.w8(32'hbc72ed60),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c8d4c),
	.w1(32'h3cb70ffd),
	.w2(32'h3c68eaf8),
	.w3(32'hbc899c1b),
	.w4(32'h3ad1f423),
	.w5(32'h3c229298),
	.w6(32'h3bed3dac),
	.w7(32'h3b77b7e0),
	.w8(32'h3c0e9cc0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c044015),
	.w1(32'h3a6e545a),
	.w2(32'hba30b1cb),
	.w3(32'h3cb29ac2),
	.w4(32'hbade9785),
	.w5(32'hbbe23e70),
	.w6(32'hbba513b0),
	.w7(32'hbb9b13cb),
	.w8(32'hbab979fe),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad900c5),
	.w1(32'hbc90f56e),
	.w2(32'hbc45cae2),
	.w3(32'hbbac7740),
	.w4(32'h3c35fc87),
	.w5(32'h3c5556b0),
	.w6(32'h3aa8f6b6),
	.w7(32'hba7be4d3),
	.w8(32'hbc08a3bc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af13552),
	.w1(32'hbbce1eba),
	.w2(32'hbbbd8c31),
	.w3(32'h3bb6aab5),
	.w4(32'hbc36cb52),
	.w5(32'hbc6ed895),
	.w6(32'hbbd767d4),
	.w7(32'hbba77569),
	.w8(32'h3aa2a329),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28e798),
	.w1(32'hbbb6c411),
	.w2(32'hbb9d0966),
	.w3(32'hbc4dab79),
	.w4(32'h3b50d7a3),
	.w5(32'h3bd798ab),
	.w6(32'hba84e4b3),
	.w7(32'hbbae47ec),
	.w8(32'hbadeef43),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fac757),
	.w1(32'hbb0df919),
	.w2(32'hba5edc75),
	.w3(32'h3c14ebb4),
	.w4(32'hbb612e79),
	.w5(32'hbb19532e),
	.w6(32'hbae47f28),
	.w7(32'hbaa90106),
	.w8(32'hb8a6b788),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94b164),
	.w1(32'h3bfdb085),
	.w2(32'h3c0a008a),
	.w3(32'hbad03a44),
	.w4(32'hbbb22711),
	.w5(32'hbc8c1be5),
	.w6(32'h3b3e7a9a),
	.w7(32'h3c09bcaf),
	.w8(32'h3c0ee78c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c170c82),
	.w1(32'h3b1f5ff3),
	.w2(32'hbb0af7b5),
	.w3(32'hbca29a62),
	.w4(32'hb90daf57),
	.w5(32'h3a8be251),
	.w6(32'h3afaf4ff),
	.w7(32'h3a2722ca),
	.w8(32'h399399eb),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04635a),
	.w1(32'h3b7580cf),
	.w2(32'hbb35a310),
	.w3(32'h3ac789e7),
	.w4(32'hbb688c68),
	.w5(32'hbc338a1f),
	.w6(32'h3b52db87),
	.w7(32'h3bdaea81),
	.w8(32'h3c0d4e53),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2f07c),
	.w1(32'h3c6149c7),
	.w2(32'h3cea923c),
	.w3(32'hbac26761),
	.w4(32'hbc0d0553),
	.w5(32'hbcf7f16d),
	.w6(32'hbc2b4e79),
	.w7(32'hbbafb1c5),
	.w8(32'h3bf302f7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c940679),
	.w1(32'hbbc1c41e),
	.w2(32'hbbced879),
	.w3(32'hbcd91daa),
	.w4(32'h3afbc972),
	.w5(32'h3c157079),
	.w6(32'h3b88366a),
	.w7(32'hbac176d6),
	.w8(32'h3891dd92),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc089434),
	.w1(32'h3a2da36b),
	.w2(32'h3aad28a5),
	.w3(32'h3b9361fb),
	.w4(32'hbba7b8b6),
	.w5(32'hbb5bbc9e),
	.w6(32'hbb2e849f),
	.w7(32'hb9db1cd8),
	.w8(32'h3a23204a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb841ec5b),
	.w1(32'hbb39dc89),
	.w2(32'h3aa14836),
	.w3(32'hb90f97cb),
	.w4(32'hbb25dbf3),
	.w5(32'hbbabf72a),
	.w6(32'hb9d5584b),
	.w7(32'hbb63937a),
	.w8(32'h3992a76f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba098ec),
	.w1(32'h3b1ba0d5),
	.w2(32'hbaa38676),
	.w3(32'hbbc6388a),
	.w4(32'hbadf9c5b),
	.w5(32'hbbc4ec11),
	.w6(32'hb9b4f12e),
	.w7(32'h3b776641),
	.w8(32'h3b9fd0ee),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c640a),
	.w1(32'hbbec7105),
	.w2(32'hbc4555d2),
	.w3(32'hb984b1f4),
	.w4(32'hbc189177),
	.w5(32'hbc82cbaa),
	.w6(32'hbb4ceffa),
	.w7(32'hbb07e275),
	.w8(32'h39cd517e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46aa7a),
	.w1(32'hbb08afb8),
	.w2(32'hbb3a7d76),
	.w3(32'hbc999a1a),
	.w4(32'h3b5cb694),
	.w5(32'hbba41dcf),
	.w6(32'hbbd723de),
	.w7(32'hbb24cdd2),
	.w8(32'hbb9c2383),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20e240),
	.w1(32'h3c4e2f82),
	.w2(32'h3c3e3a55),
	.w3(32'hbc06a51a),
	.w4(32'h3b4974f8),
	.w5(32'hbbb39649),
	.w6(32'hbbaf2265),
	.w7(32'hbba375a7),
	.w8(32'h3b648004),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92f48f),
	.w1(32'hbb7445db),
	.w2(32'hbb9f8581),
	.w3(32'h3b90a85b),
	.w4(32'hbb4fa992),
	.w5(32'hbc02de4f),
	.w6(32'h3b041ae3),
	.w7(32'hbb8f99ff),
	.w8(32'hbbd672bb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f5c0f),
	.w1(32'h3b177b77),
	.w2(32'h3a8f8320),
	.w3(32'hbb17d7e9),
	.w4(32'h3ad8b9c1),
	.w5(32'h3aaa9556),
	.w6(32'h3afbb951),
	.w7(32'h3af613a9),
	.w8(32'h3a06659b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913782c),
	.w1(32'hbad71bb2),
	.w2(32'hbbce7c2d),
	.w3(32'h3ac159d3),
	.w4(32'h3b1035ea),
	.w5(32'hbae1700d),
	.w6(32'h3badc80a),
	.w7(32'hb9d6f8ea),
	.w8(32'h3b3865f7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc371c),
	.w1(32'h3cd62df8),
	.w2(32'h3c87772d),
	.w3(32'h3afca93b),
	.w4(32'hbc27e1cf),
	.w5(32'hbb0e01ff),
	.w6(32'h3be3b19a),
	.w7(32'h3c5f4b8b),
	.w8(32'h3c8e8109),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb1640),
	.w1(32'hbc58746e),
	.w2(32'hbbedf599),
	.w3(32'h3c08aff8),
	.w4(32'h3c993698),
	.w5(32'h3caa2176),
	.w6(32'hbb20e2b3),
	.w7(32'hbb5fe2e6),
	.w8(32'hbc5bab63),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca71c45),
	.w1(32'h3ad75ea1),
	.w2(32'h3bb248db),
	.w3(32'hbc1e9cdb),
	.w4(32'h3b05b174),
	.w5(32'h3b98e62a),
	.w6(32'h3ae376f3),
	.w7(32'h3b5ea395),
	.w8(32'h3ab69c16),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7543aa),
	.w1(32'h3b64e012),
	.w2(32'hbc3c9b5a),
	.w3(32'h3a50136a),
	.w4(32'h3bb5628c),
	.w5(32'hbc562b3b),
	.w6(32'h3ba7a97a),
	.w7(32'hbc1635c9),
	.w8(32'h3bcdaa77),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule