module layer_8_featuremap_65(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43f249),
	.w1(32'hba11a868),
	.w2(32'hb8dd9cf5),
	.w3(32'hba1ee514),
	.w4(32'hb9ec2ccd),
	.w5(32'hb8acf8ee),
	.w6(32'hb921d9c7),
	.w7(32'hb99deca7),
	.w8(32'hb97e3301),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9544067),
	.w1(32'hb97d8f0a),
	.w2(32'hb9af5f1b),
	.w3(32'hb9a07d75),
	.w4(32'hb9aa6a1c),
	.w5(32'hb9c0de9f),
	.w6(32'hb883815d),
	.w7(32'hb9a55d0c),
	.w8(32'hb983f5b0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f47a3),
	.w1(32'hb95479e6),
	.w2(32'hb90c25b7),
	.w3(32'hb904c7c5),
	.w4(32'hb912bac4),
	.w5(32'hb90f4955),
	.w6(32'hb81b89b2),
	.w7(32'hb973d5c9),
	.w8(32'h3a112d9b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3be84a),
	.w1(32'h3b781c00),
	.w2(32'h3a9f8bfb),
	.w3(32'h3acfa964),
	.w4(32'h3b13485e),
	.w5(32'h3b22d436),
	.w6(32'hba789c91),
	.w7(32'hbae62daa),
	.w8(32'h39531a21),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d1f9b),
	.w1(32'hb92bf376),
	.w2(32'h39be2c8d),
	.w3(32'h38ccfcbf),
	.w4(32'hb8e90c02),
	.w5(32'h394173be),
	.w6(32'hb93014fa),
	.w7(32'h38f0d012),
	.w8(32'hbac72983),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b63bd8),
	.w1(32'hb9c0883a),
	.w2(32'hb998606a),
	.w3(32'hb8e38b67),
	.w4(32'h39b37e08),
	.w5(32'h3a7421c7),
	.w6(32'hb806d5aa),
	.w7(32'hbacab5b9),
	.w8(32'hb9a12c85),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9274255),
	.w1(32'hba108a0d),
	.w2(32'hb9aec763),
	.w3(32'hb9651286),
	.w4(32'hba1b0ab2),
	.w5(32'hb9fd9e67),
	.w6(32'hb8f480e3),
	.w7(32'hb9337b0b),
	.w8(32'h39b0cf89),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391854ec),
	.w1(32'hb947b936),
	.w2(32'h39fea322),
	.w3(32'h392e0997),
	.w4(32'h397748c7),
	.w5(32'h39ad924d),
	.w6(32'hb98e4942),
	.w7(32'h39ae8436),
	.w8(32'hb7f03c81),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a3c6d5),
	.w1(32'hb9b7d10a),
	.w2(32'hb930a6a9),
	.w3(32'hb899f010),
	.w4(32'hba234f17),
	.w5(32'hba0764e1),
	.w6(32'h392b7eac),
	.w7(32'h38154263),
	.w8(32'h3a8e4dc6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7080b),
	.w1(32'h3b27ae4b),
	.w2(32'h3a91e5e0),
	.w3(32'hba2f4c90),
	.w4(32'hb811c126),
	.w5(32'hbae5547c),
	.w6(32'h396c1a16),
	.w7(32'h3836ded5),
	.w8(32'h3a5f078d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fc5ad),
	.w1(32'h3a286550),
	.w2(32'h3a3729c0),
	.w3(32'h3a39fc11),
	.w4(32'h3a420b58),
	.w5(32'h3a44af64),
	.w6(32'h39e1d03e),
	.w7(32'h394d26cf),
	.w8(32'hb9b21059),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942a3cc),
	.w1(32'hb9b5c6d2),
	.w2(32'hb92832dc),
	.w3(32'hb951a4b3),
	.w4(32'hb980eb9c),
	.w5(32'hb92b0d10),
	.w6(32'hb9344b78),
	.w7(32'hb9a4a91f),
	.w8(32'hb80f1114),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c01902),
	.w1(32'h39600f07),
	.w2(32'h391625d5),
	.w3(32'h39480e51),
	.w4(32'h38d3a813),
	.w5(32'hb6de6ebd),
	.w6(32'h393a377e),
	.w7(32'h396fa7fb),
	.w8(32'hbad4f5e3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3b116),
	.w1(32'hb9e20b6c),
	.w2(32'hb96c0f93),
	.w3(32'hb90717d0),
	.w4(32'h39cd5d2f),
	.w5(32'h3a9b0c9d),
	.w6(32'h38ab8826),
	.w7(32'hbad06786),
	.w8(32'hbaadbb48),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdba18),
	.w1(32'hb83ae23f),
	.w2(32'hb9992a85),
	.w3(32'hb98fda58),
	.w4(32'hb82930f7),
	.w5(32'h3a2663e5),
	.w6(32'hb9ceef16),
	.w7(32'hba8d7877),
	.w8(32'h3978dbd3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab7fed),
	.w1(32'h3905bb19),
	.w2(32'h3a0af5d4),
	.w3(32'hb9c1e5c5),
	.w4(32'h383fd44b),
	.w5(32'hb8b2468c),
	.w6(32'h39ae32e2),
	.w7(32'h38b03bec),
	.w8(32'h3afe3811),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ae90b),
	.w1(32'h39378041),
	.w2(32'hbb8d7d1c),
	.w3(32'h3baf4dd2),
	.w4(32'h3bcfa296),
	.w5(32'h3b074744),
	.w6(32'h3b1ceb89),
	.w7(32'h3a98e872),
	.w8(32'hb98f2212),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904a37d),
	.w1(32'h3a1326b7),
	.w2(32'h39608584),
	.w3(32'h38df1f8b),
	.w4(32'hb96887fb),
	.w5(32'h390693ae),
	.w6(32'hb928e6a4),
	.w7(32'h38e530dd),
	.w8(32'h39c4d75f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10e0d1),
	.w1(32'h3aa02011),
	.w2(32'h3acd2c11),
	.w3(32'h3a0f5963),
	.w4(32'h3aad6726),
	.w5(32'h3a189506),
	.w6(32'h39428bba),
	.w7(32'h3a783bb4),
	.w8(32'h3b8bf6d1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac07564),
	.w1(32'hbb80da40),
	.w2(32'hbb5cc4d6),
	.w3(32'h39a0ad21),
	.w4(32'h39b74eed),
	.w5(32'h38f2e187),
	.w6(32'h3b05286a),
	.w7(32'hbb2f8732),
	.w8(32'h3a5dd1ea),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b8dc0),
	.w1(32'h38bd0ac0),
	.w2(32'h39ddf8be),
	.w3(32'h3a0d6d84),
	.w4(32'h391ae68a),
	.w5(32'h3a1c6adc),
	.w6(32'h39f67d06),
	.w7(32'h3a9967e1),
	.w8(32'hba3014f2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed06ee),
	.w1(32'hba64f709),
	.w2(32'hb94d6329),
	.w3(32'hb9b5ce86),
	.w4(32'hb9db0e1f),
	.w5(32'hb96189ca),
	.w6(32'hba6f0614),
	.w7(32'hba0e2775),
	.w8(32'h3abea74c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0c4a),
	.w1(32'hb98728c6),
	.w2(32'h3a206fe5),
	.w3(32'hba58cf7c),
	.w4(32'hb9a15b6e),
	.w5(32'hb881fcde),
	.w6(32'h399af85a),
	.w7(32'h3b2ead46),
	.w8(32'hba1030d4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2922c),
	.w1(32'hba4e98c8),
	.w2(32'h3a55705e),
	.w3(32'hba770e85),
	.w4(32'hb947cf91),
	.w5(32'h3a7ce2d7),
	.w6(32'hb9d4e820),
	.w7(32'h390419bd),
	.w8(32'h3b266a16),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d9b6c),
	.w1(32'hbb23c695),
	.w2(32'hbae1a296),
	.w3(32'hbaf5b2da),
	.w4(32'hbb911245),
	.w5(32'hbb32abc2),
	.w6(32'h3aafa83e),
	.w7(32'h39df2982),
	.w8(32'h3abb4e01),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d59fdc),
	.w1(32'hb95fdbf9),
	.w2(32'h3a17a16e),
	.w3(32'hba320e92),
	.w4(32'hb9aa0b6b),
	.w5(32'hb924b0a2),
	.w6(32'h39e1d276),
	.w7(32'h3b2651f7),
	.w8(32'h3a9b7756),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9408a9c),
	.w1(32'hb8ec2579),
	.w2(32'h3a0840f5),
	.w3(32'hb9e0a51a),
	.w4(32'hb9626492),
	.w5(32'hb8f06f4b),
	.w6(32'h3a0cfffb),
	.w7(32'h3b150603),
	.w8(32'h3a4e8220),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba707da2),
	.w1(32'hbad3a505),
	.w2(32'hba6856d7),
	.w3(32'hba2b4132),
	.w4(32'hba7fbc08),
	.w5(32'hba013619),
	.w6(32'hb9dd1199),
	.w7(32'h391e7256),
	.w8(32'hbb1f8b61),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54ab6a),
	.w1(32'hbb71e0e2),
	.w2(32'h3a92d962),
	.w3(32'hbb53f0e2),
	.w4(32'hb9d11949),
	.w5(32'h39075408),
	.w6(32'hbaf7b9b7),
	.w7(32'hbb2f94b7),
	.w8(32'hb98bb963),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a26560),
	.w1(32'h372e0362),
	.w2(32'hb900f228),
	.w3(32'hb856bf72),
	.w4(32'h3805484b),
	.w5(32'hb8b37c54),
	.w6(32'hb81c27f0),
	.w7(32'hb991bab3),
	.w8(32'hb9945624),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a8f2a),
	.w1(32'h3a33043b),
	.w2(32'hbb4127c4),
	.w3(32'hba76a2ef),
	.w4(32'h39b7c922),
	.w5(32'h39b02411),
	.w6(32'hb9234233),
	.w7(32'hbb14625a),
	.w8(32'h3b073576),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b4496),
	.w1(32'hba76034a),
	.w2(32'hba479b04),
	.w3(32'hb9d8cc9b),
	.w4(32'hbb171342),
	.w5(32'hbabac638),
	.w6(32'h3ac0a4ca),
	.w7(32'h3ae0987d),
	.w8(32'hbb009cf5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb068448),
	.w1(32'hba78eb6a),
	.w2(32'hbb6648e4),
	.w3(32'hba148bab),
	.w4(32'hbabf8def),
	.w5(32'hba9b0af6),
	.w6(32'hbb0dbff6),
	.w7(32'hbb76381b),
	.w8(32'h3aeccf9a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb217aa),
	.w1(32'h3bb89fff),
	.w2(32'h3b2531fc),
	.w3(32'h3b018bed),
	.w4(32'h3b4a1b66),
	.w5(32'h39dc3d93),
	.w6(32'h3b3ee244),
	.w7(32'h3a9c2598),
	.w8(32'hbab7b712),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba0daf),
	.w1(32'hb9bf3aa4),
	.w2(32'hb9692c1e),
	.w3(32'hb8cc54a6),
	.w4(32'h39cb87ad),
	.w5(32'h3a859017),
	.w6(32'h38ae0bcd),
	.w7(32'hbab1db89),
	.w8(32'hb9c3b8dc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2057b4),
	.w1(32'hb93f770d),
	.w2(32'h3a0f4c94),
	.w3(32'hb9a467ae),
	.w4(32'hb8fb3237),
	.w5(32'h39d8339e),
	.w6(32'hb8c7c0eb),
	.w7(32'h3903790d),
	.w8(32'h3b25d927),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6263fa),
	.w1(32'hbb05b4e3),
	.w2(32'hb997a24d),
	.w3(32'hba3cfab7),
	.w4(32'hbaa44177),
	.w5(32'hba529cf1),
	.w6(32'hb8dc3c73),
	.w7(32'h3a71ed9d),
	.w8(32'hba01546f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0baac4),
	.w1(32'hb9ea0151),
	.w2(32'hb9b4fc40),
	.w3(32'hb992a5f0),
	.w4(32'hb9556d53),
	.w5(32'hb922381a),
	.w6(32'hb99f76f4),
	.w7(32'hba0eda9e),
	.w8(32'hbb30abf9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60d316),
	.w1(32'h3810f9da),
	.w2(32'hb9dcab77),
	.w3(32'hba64b233),
	.w4(32'hba178a0f),
	.w5(32'h3acfee47),
	.w6(32'hba95c96a),
	.w7(32'hbb03937e),
	.w8(32'h3a7fdf02),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dc222),
	.w1(32'hbad3e734),
	.w2(32'hba08a676),
	.w3(32'hba764c4f),
	.w4(32'hbb05d5d2),
	.w5(32'hba6fe73c),
	.w6(32'h388d931f),
	.w7(32'h3a2f85f2),
	.w8(32'h3a1b7529),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96943b8),
	.w1(32'hb8a88017),
	.w2(32'h39092771),
	.w3(32'hb9a636b3),
	.w4(32'hb9127aa6),
	.w5(32'hb956bea8),
	.w6(32'h374bebac),
	.w7(32'h3a812a14),
	.w8(32'hbb8b71d4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ff8e5),
	.w1(32'hbb83530c),
	.w2(32'hbb33d92b),
	.w3(32'hbb00acdb),
	.w4(32'hbb85c8c8),
	.w5(32'hb9d2175a),
	.w6(32'hbb582c45),
	.w7(32'hbb7ddfc5),
	.w8(32'hbbc8b466),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfb590),
	.w1(32'hbaaa5bc5),
	.w2(32'h3b554f99),
	.w3(32'h3c52cbe2),
	.w4(32'h3b73d44b),
	.w5(32'hbbe0e825),
	.w6(32'hbc18343b),
	.w7(32'h3b4bca0f),
	.w8(32'h3aa3a658),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e2a4b),
	.w1(32'hbaea6d8c),
	.w2(32'h3a8b9e83),
	.w3(32'hbbe97d9c),
	.w4(32'hbc29d463),
	.w5(32'hbb3056ba),
	.w6(32'h3b81efad),
	.w7(32'h3b33a5b4),
	.w8(32'hb7574ffa),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3891a),
	.w1(32'hbb0bc735),
	.w2(32'hbabbcc3e),
	.w3(32'hbb6840af),
	.w4(32'hbbe1a5cd),
	.w5(32'hbb2ae2cc),
	.w6(32'h3ac43031),
	.w7(32'hba07d64c),
	.w8(32'hbb4b618e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abca2b0),
	.w1(32'hbb7ce723),
	.w2(32'hbb907750),
	.w3(32'h3bec4c3b),
	.w4(32'h3b808962),
	.w5(32'h3b6acc05),
	.w6(32'hbc3a6297),
	.w7(32'hbbec6a6e),
	.w8(32'h3c0a89b8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcac20a),
	.w1(32'hbb4b2e4c),
	.w2(32'h3bbcb58c),
	.w3(32'h3bb4daf4),
	.w4(32'h3c63c116),
	.w5(32'h3c2f42bf),
	.w6(32'hbc4ebcf6),
	.w7(32'hbc7e5784),
	.w8(32'hbb8e75cd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1283fa),
	.w1(32'h3a74134e),
	.w2(32'hbbc9fe3a),
	.w3(32'h3a17524f),
	.w4(32'hbb5ef196),
	.w5(32'h3a29054e),
	.w6(32'hbbff4c51),
	.w7(32'hbc12eab2),
	.w8(32'hbc36dff3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db70bf),
	.w1(32'hbaa2b10a),
	.w2(32'hbc8129cb),
	.w3(32'h3cca8114),
	.w4(32'h3d00dff5),
	.w5(32'h3c1d6b2f),
	.w6(32'hbc8901d6),
	.w7(32'hbc9ab1b1),
	.w8(32'hba985d16),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8784bc),
	.w1(32'hbab2ead5),
	.w2(32'hba53e923),
	.w3(32'hbadcb3ed),
	.w4(32'hbb8421b7),
	.w5(32'h399903b8),
	.w6(32'hb8d58de5),
	.w7(32'hbaeee289),
	.w8(32'h3a4ee742),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad79822),
	.w1(32'hb9f51a54),
	.w2(32'h393a3bd1),
	.w3(32'hbb9234b4),
	.w4(32'hbbbb8372),
	.w5(32'hbb44a841),
	.w6(32'h3b16ad5d),
	.w7(32'h3a8894bd),
	.w8(32'h3a7c63b9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb998fe2),
	.w1(32'hbad1280b),
	.w2(32'h3a684aa8),
	.w3(32'hbc2af073),
	.w4(32'hbc509ba4),
	.w5(32'hbbb74748),
	.w6(32'h3bb5dac8),
	.w7(32'h3b5c961c),
	.w8(32'h39c394ca),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31510d),
	.w1(32'h3b8c76b7),
	.w2(32'h3c8089b4),
	.w3(32'hbb76a996),
	.w4(32'h3b45eb36),
	.w5(32'h3c2e5448),
	.w6(32'hbbeb3756),
	.w7(32'h3bd133f6),
	.w8(32'hbc53ebb0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a50f3),
	.w1(32'h3a295d7e),
	.w2(32'hbc024ad0),
	.w3(32'h3c8a51bb),
	.w4(32'h3cbb76bb),
	.w5(32'h3c0f2d60),
	.w6(32'hbc8b2a11),
	.w7(32'hbc8b4ecb),
	.w8(32'hbba3a5d6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd79abe),
	.w1(32'h3b97d738),
	.w2(32'h3c4a2da8),
	.w3(32'h3c2129cc),
	.w4(32'hba838063),
	.w5(32'hbb6012fd),
	.w6(32'hbbdf61ac),
	.w7(32'h3c1d7bc5),
	.w8(32'h3c39952a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47325a),
	.w1(32'h3c75a996),
	.w2(32'h3c25801c),
	.w3(32'h3bb47641),
	.w4(32'h3c17319d),
	.w5(32'h3bd84fbd),
	.w6(32'h3c8b26e6),
	.w7(32'h3c201e5f),
	.w8(32'hba70fcee),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aae362),
	.w1(32'hbae3aee8),
	.w2(32'hbb115bb1),
	.w3(32'hbc1a51a3),
	.w4(32'hbc1f9d3c),
	.w5(32'h3b70eb4e),
	.w6(32'hba55e6e2),
	.w7(32'hbb763ec6),
	.w8(32'hbc26bd8a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e534fb),
	.w1(32'hbc351011),
	.w2(32'h3b150ee3),
	.w3(32'h3b14ae5a),
	.w4(32'hbc3d864b),
	.w5(32'hbc0babbd),
	.w6(32'hbc4a0c4b),
	.w7(32'hbba35b27),
	.w8(32'h3c008bf4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b69c4),
	.w1(32'hbb1fe2b1),
	.w2(32'hbc1a2685),
	.w3(32'hbbc523eb),
	.w4(32'hbb9d3764),
	.w5(32'hbbd9e319),
	.w6(32'h3c82c567),
	.w7(32'h3c0158ce),
	.w8(32'h39c0b268),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c07c5),
	.w1(32'hba8ffeda),
	.w2(32'h3ac18803),
	.w3(32'h3c0e66af),
	.w4(32'h3c650e7a),
	.w5(32'h3c4000ea),
	.w6(32'hbc4c1f01),
	.w7(32'hbada2773),
	.w8(32'h3c13e034),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab985f),
	.w1(32'h3ab2fd9c),
	.w2(32'hbc4dbd7d),
	.w3(32'h3c03b5b9),
	.w4(32'h3a6a6a32),
	.w5(32'h3c5885c1),
	.w6(32'h3b5eefff),
	.w7(32'hbc3895ab),
	.w8(32'hbbb9418d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f5681),
	.w1(32'h3851245f),
	.w2(32'hbacfab42),
	.w3(32'hb9d6704d),
	.w4(32'h3b10b5a9),
	.w5(32'h3c04c77d),
	.w6(32'hbc407666),
	.w7(32'hbc0a15ea),
	.w8(32'hba2ad8bf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b0cdf),
	.w1(32'h3b18fed0),
	.w2(32'h3b64ae1d),
	.w3(32'hbc1e8a88),
	.w4(32'hbc0b31be),
	.w5(32'hbb73d6fa),
	.w6(32'h3bc45911),
	.w7(32'h3b7b2fc9),
	.w8(32'hbbbdc8d6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73154e),
	.w1(32'hbc2d3979),
	.w2(32'hbbbca45f),
	.w3(32'hbc1fc681),
	.w4(32'hbcad3728),
	.w5(32'hbcf08144),
	.w6(32'hbc1aae51),
	.w7(32'hbb8f05b5),
	.w8(32'hb6e5eeb9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bda56),
	.w1(32'hbb2d58d6),
	.w2(32'hbadfffa2),
	.w3(32'hbb8ae228),
	.w4(32'hbbfdf13f),
	.w5(32'hbb2a55e4),
	.w6(32'hb98ca50a),
	.w7(32'hba422efe),
	.w8(32'h3ab4b6c2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa209aa),
	.w1(32'hba0a1425),
	.w2(32'h3a7568c9),
	.w3(32'hbb47fc74),
	.w4(32'hbb95e34e),
	.w5(32'hba7f5d63),
	.w6(32'h3b4dad34),
	.w7(32'h3b070a4f),
	.w8(32'h3883c8c3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa9628),
	.w1(32'hba58ba02),
	.w2(32'hb93b4b6e),
	.w3(32'hbb410c00),
	.w4(32'hbb797963),
	.w5(32'hbae05ba6),
	.w6(32'h3a6e9ee7),
	.w7(32'h399ffa2b),
	.w8(32'hbbf22c73),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1102c8),
	.w1(32'hbb942b8f),
	.w2(32'hbc12a4f5),
	.w3(32'h3a0e58c2),
	.w4(32'h3b974055),
	.w5(32'h3c0a7045),
	.w6(32'hbc1e3af8),
	.w7(32'hbc4a834c),
	.w8(32'hb9cf62d8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988eb3d),
	.w1(32'hba9074d2),
	.w2(32'hb89ac16e),
	.w3(32'hba8fe813),
	.w4(32'hbb8487d8),
	.w5(32'hb992d165),
	.w6(32'h398cdbf1),
	.w7(32'hba958a5c),
	.w8(32'h3cd5ddba),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f5bf9),
	.w1(32'hbadbb0d7),
	.w2(32'h3b1e0dbe),
	.w3(32'hbd10220c),
	.w4(32'hbd22622e),
	.w5(32'hbca4a3b3),
	.w6(32'h3d36aabf),
	.w7(32'h3d07fe32),
	.w8(32'hbb312278),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4336b9),
	.w1(32'hbb4e5820),
	.w2(32'hbaf837b9),
	.w3(32'hbb3e96c6),
	.w4(32'hbba9d6f1),
	.w5(32'hbaeb06c8),
	.w6(32'hbab83b3f),
	.w7(32'hbb044205),
	.w8(32'hba9f89ca),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381d1d02),
	.w1(32'hbb0ca85d),
	.w2(32'hbaf404ff),
	.w3(32'h38c66224),
	.w4(32'hbb60eecb),
	.w5(32'hba1e313d),
	.w6(32'hbb007830),
	.w7(32'hbb3e823c),
	.w8(32'hba38cd48),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5406e),
	.w1(32'hbaffac03),
	.w2(32'hb8abf074),
	.w3(32'hbb08f15d),
	.w4(32'hbba3fff5),
	.w5(32'hba95243f),
	.w6(32'h39a19323),
	.w7(32'hb9b6fceb),
	.w8(32'hbb872ed5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d946e),
	.w1(32'hbc3ff518),
	.w2(32'hbba17929),
	.w3(32'h3bad40d6),
	.w4(32'h3c724f06),
	.w5(32'h3c80e66b),
	.w6(32'hbc138cfe),
	.w7(32'hbc0a45b1),
	.w8(32'hbb6a381b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad24ae0),
	.w1(32'hbbae7980),
	.w2(32'hbb9a3d82),
	.w3(32'h3a7f379e),
	.w4(32'hbb82fd70),
	.w5(32'hbb058e43),
	.w6(32'hbbb1c4ef),
	.w7(32'hbbcf98bf),
	.w8(32'hba5eca9d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb278b58),
	.w1(32'hbac8c84c),
	.w2(32'h38dbf335),
	.w3(32'hbba7017e),
	.w4(32'hbbd9dd99),
	.w5(32'hbb1be585),
	.w6(32'h3a7ffdc5),
	.w7(32'h39e1a69b),
	.w8(32'hbb66ddbc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ec00e),
	.w1(32'hbb7aa6ab),
	.w2(32'hbb4f0f49),
	.w3(32'hbaf924bb),
	.w4(32'hbb8bd2fc),
	.w5(32'hbaa06f05),
	.w6(32'hbb6f84ca),
	.w7(32'hbb769886),
	.w8(32'h3cf63c5e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85a3f6),
	.w1(32'hbb0baf76),
	.w2(32'h3a3016ff),
	.w3(32'hbd201aeb),
	.w4(32'hbd32d12a),
	.w5(32'hbcbd18ae),
	.w6(32'h3d54af8a),
	.w7(32'h3d1ab521),
	.w8(32'h3c4c4f7d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0ccb8),
	.w1(32'h392b2b2b),
	.w2(32'h3b65d381),
	.w3(32'hbca8c157),
	.w4(32'hbcc3e0a1),
	.w5(32'hbc360d1d),
	.w6(32'h3cceae65),
	.w7(32'h3c913d90),
	.w8(32'h3b8b0b0d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fea255),
	.w1(32'hba98d907),
	.w2(32'h3ac9849d),
	.w3(32'hba7a1d0e),
	.w4(32'hbb83196e),
	.w5(32'h3b77d526),
	.w6(32'h3b030ea3),
	.w7(32'h3ae8ecde),
	.w8(32'h3ac79c7b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6456c),
	.w1(32'hbc801af0),
	.w2(32'hbca564b5),
	.w3(32'hbc6592de),
	.w4(32'hbc2bf9af),
	.w5(32'hbbd9688b),
	.w6(32'hba46d01e),
	.w7(32'hbbb1a6ce),
	.w8(32'hbac00230),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b1b0d),
	.w1(32'hbb0276a8),
	.w2(32'hbabf63c4),
	.w3(32'hba818e50),
	.w4(32'hbb3f2642),
	.w5(32'hba277fe0),
	.w6(32'hbb48bd4c),
	.w7(32'hbb32cc18),
	.w8(32'h3a89c18a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d319e),
	.w1(32'hb9fbbc95),
	.w2(32'hbad85243),
	.w3(32'h3b83b801),
	.w4(32'h3a4947c8),
	.w5(32'h3bc6e3f8),
	.w6(32'hbbb359a3),
	.w7(32'hbb934f55),
	.w8(32'h3a1ce8fb),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920e18),
	.w1(32'h3b2d80f7),
	.w2(32'h3be85ec2),
	.w3(32'hbc8abdac),
	.w4(32'hbbb22ed5),
	.w5(32'hba970062),
	.w6(32'hbc06ac62),
	.w7(32'h3af861e4),
	.w8(32'hbc373bb2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb149da),
	.w1(32'hb9eb9627),
	.w2(32'hbc0c1315),
	.w3(32'h3c9c5364),
	.w4(32'h3c94f726),
	.w5(32'h3bce0dee),
	.w6(32'hbca70110),
	.w7(32'hbcb17e76),
	.w8(32'hb9162c9a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f1737),
	.w1(32'hba5569c7),
	.w2(32'h38a8e53d),
	.w3(32'hbb5f5060),
	.w4(32'hbbcf5328),
	.w5(32'hbaf9fe9d),
	.w6(32'h3b52c014),
	.w7(32'h3aa8b09c),
	.w8(32'hbc723bd4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c97db),
	.w1(32'hbadbc6e6),
	.w2(32'hbcab7b9e),
	.w3(32'h3d0624d7),
	.w4(32'h3d2a9a13),
	.w5(32'h3c4ffdb7),
	.w6(32'hbcb4380e),
	.w7(32'hbccc53e2),
	.w8(32'hbb17f348),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05e898),
	.w1(32'hba691dfb),
	.w2(32'hbb9c71e9),
	.w3(32'hba56a42a),
	.w4(32'hbb9a6885),
	.w5(32'hbb293541),
	.w6(32'hbad51d9c),
	.w7(32'hbb990221),
	.w8(32'hbaaa077b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba95581),
	.w1(32'hbae9f109),
	.w2(32'hbb70842d),
	.w3(32'h3be3eb72),
	.w4(32'h3c4ed2a8),
	.w5(32'h3c04dcbf),
	.w6(32'hbc2b2037),
	.w7(32'hbc0074df),
	.w8(32'hbc624040),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f31afb),
	.w1(32'hbad4f64b),
	.w2(32'hbca08b92),
	.w3(32'h3cfa53bd),
	.w4(32'h3d1f54fa),
	.w5(32'h3c424a8e),
	.w6(32'hbca9947b),
	.w7(32'hbcbfd9bf),
	.w8(32'hbc4243df),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec36c0),
	.w1(32'hbab03cfd),
	.w2(32'hbc88d816),
	.w3(32'h3cd66d4b),
	.w4(32'h3d087bc7),
	.w5(32'h3c26d405),
	.w6(32'hbc912719),
	.w7(32'hbca3def2),
	.w8(32'hbc20d446),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc30c53),
	.w1(32'h3afecbaf),
	.w2(32'hbbc534d2),
	.w3(32'h3ca04dfb),
	.w4(32'h3cb5f7a7),
	.w5(32'h3c118e05),
	.w6(32'hbc6f1b9f),
	.w7(32'hbc7cf147),
	.w8(32'h3b2e72e3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d75d0),
	.w1(32'h3b627c82),
	.w2(32'h3c196f2e),
	.w3(32'hbbf91af7),
	.w4(32'hbbfb947a),
	.w5(32'h3c8ea5b8),
	.w6(32'hbbe7f7fc),
	.w7(32'hbc2e6e67),
	.w8(32'h3a132cb5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98ecaf),
	.w1(32'hb980580a),
	.w2(32'h3a2c9204),
	.w3(32'hbb6a3873),
	.w4(32'hbb8cdc49),
	.w5(32'hbaebec45),
	.w6(32'h3aec30d8),
	.w7(32'h3aa3ff2b),
	.w8(32'hbc5bdcfb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae2a3),
	.w1(32'hbbab8a81),
	.w2(32'hbb63d424),
	.w3(32'hbc58dfcc),
	.w4(32'hbc570c5a),
	.w5(32'hbc508e94),
	.w6(32'hbc427eab),
	.w7(32'hbc3a0c74),
	.w8(32'hbca0402f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedfa65),
	.w1(32'hbb63f94a),
	.w2(32'hbc880914),
	.w3(32'h3cd78c95),
	.w4(32'h3cd5f375),
	.w5(32'h3bc02a98),
	.w6(32'hbd06fd3f),
	.w7(32'hbd094327),
	.w8(32'hbce26fb3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a15a7),
	.w1(32'hbc3bbfe2),
	.w2(32'hbc4e7f25),
	.w3(32'hbbc95692),
	.w4(32'hbb8c3a02),
	.w5(32'h3ad3f520),
	.w6(32'hbce9f6d7),
	.w7(32'hbcdd88b3),
	.w8(32'hba76b2f0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84aed8),
	.w1(32'h3b60e790),
	.w2(32'h3be30da5),
	.w3(32'hbbb16d43),
	.w4(32'hbb0f1f33),
	.w5(32'hbc09fe08),
	.w6(32'hb9f26c83),
	.w7(32'h3b545d3f),
	.w8(32'h3cd7ccda),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66f532),
	.w1(32'hbae7760c),
	.w2(32'h3a45c9c9),
	.w3(32'hbd0c1294),
	.w4(32'hbd1cde15),
	.w5(32'hbca55392),
	.w6(32'h3d3b0984),
	.w7(32'h3d084435),
	.w8(32'hb8420416),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdf06d),
	.w1(32'hbab92b38),
	.w2(32'hba9a09bf),
	.w3(32'hba87efec),
	.w4(32'hbb9d3525),
	.w5(32'hb92262a7),
	.w6(32'hb98ffb08),
	.w7(32'hbaceea60),
	.w8(32'hbbdb537d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b085d76),
	.w1(32'hbb998d39),
	.w2(32'hbbdced3d),
	.w3(32'h3c4f9044),
	.w4(32'h3c936b9f),
	.w5(32'h3c407b50),
	.w6(32'hbca95c57),
	.w7(32'hbc512c54),
	.w8(32'h3a31910d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd3ede),
	.w1(32'hba14fbf5),
	.w2(32'hb905ebef),
	.w3(32'hbb89fd7d),
	.w4(32'hbbb593d0),
	.w5(32'hbb4ce800),
	.w6(32'h3ae9c87f),
	.w7(32'h39c3f352),
	.w8(32'h3c90b798),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d1e17),
	.w1(32'hba0190d6),
	.w2(32'h3bc6313b),
	.w3(32'hbd0c24ea),
	.w4(32'hbd2916f7),
	.w5(32'hbc8e8d6d),
	.w6(32'h3d226434),
	.w7(32'h3cd53123),
	.w8(32'hbc1daf41),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f359),
	.w1(32'hba4d43f1),
	.w2(32'hbbfdd2fd),
	.w3(32'h3caf0163),
	.w4(32'h3cba86a1),
	.w5(32'h3c27382b),
	.w6(32'hbc8b01e6),
	.w7(32'hbc90d015),
	.w8(32'hbbc89279),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a262eee),
	.w1(32'hba0ec82c),
	.w2(32'hbbf70581),
	.w3(32'h3c526bd5),
	.w4(32'h3c8478d6),
	.w5(32'h3baa85b1),
	.w6(32'hbc18e285),
	.w7(32'hbc23b955),
	.w8(32'hbb78ff50),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b495724),
	.w1(32'h3b0c5662),
	.w2(32'h3a922732),
	.w3(32'h3b63f826),
	.w4(32'h3c386cfa),
	.w5(32'h3bc4f64b),
	.w6(32'hbc325769),
	.w7(32'hbc00e715),
	.w8(32'h3c2462dc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f80c2),
	.w1(32'hbbd57460),
	.w2(32'hbb386dc6),
	.w3(32'hbb6e4515),
	.w4(32'h3ba80ba5),
	.w5(32'h3c7b86d3),
	.w6(32'hbc8a188a),
	.w7(32'hbcc0e30b),
	.w8(32'hbc1a6695),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0696bc),
	.w1(32'hbba7468a),
	.w2(32'hbbcbe076),
	.w3(32'h3c230722),
	.w4(32'h3c8a403a),
	.w5(32'h3bb987c4),
	.w6(32'hbc9f1fa6),
	.w7(32'hbc43cdb3),
	.w8(32'hbc916d14),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ff2f8),
	.w1(32'h3ba091db),
	.w2(32'h3b90e4ac),
	.w3(32'h3ca700d4),
	.w4(32'h3d04c29f),
	.w5(32'h3cb64ac3),
	.w6(32'hbcba9540),
	.w7(32'hbc8411c6),
	.w8(32'hbc2272ed),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77ef29),
	.w1(32'h3b970791),
	.w2(32'hbbc076d9),
	.w3(32'h3bd0f040),
	.w4(32'h3c8493c7),
	.w5(32'h3bd115cf),
	.w6(32'hbc83117e),
	.w7(32'hbca121be),
	.w8(32'h3b12e4aa),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c242687),
	.w1(32'h3bd1e6b4),
	.w2(32'hbc3ec97d),
	.w3(32'h3bc0c2dc),
	.w4(32'h3ba3c92f),
	.w5(32'h3b1c3138),
	.w6(32'hb7f43906),
	.w7(32'hbc28367f),
	.w8(32'hbbf49355),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f6394),
	.w1(32'h3a829a73),
	.w2(32'hbab99d0d),
	.w3(32'h3b155afb),
	.w4(32'h3c450174),
	.w5(32'h3b4a3cf9),
	.w6(32'hbbbb676e),
	.w7(32'hbc282831),
	.w8(32'h3cea5c93),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc263afe),
	.w1(32'hbb65a2b1),
	.w2(32'hbc216747),
	.w3(32'hbcfe2c41),
	.w4(32'hbd39f798),
	.w5(32'hbd0884bb),
	.w6(32'h3d425ebd),
	.w7(32'h3cebfe88),
	.w8(32'hbc91d75b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb23aa),
	.w1(32'h395f19af),
	.w2(32'hbb4faed1),
	.w3(32'h3c7b5af5),
	.w4(32'h3ce115fa),
	.w5(32'h3c7f1565),
	.w6(32'hbcd45a59),
	.w7(32'hbcb10300),
	.w8(32'hbc27b517),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3580ab),
	.w1(32'hbb3144e8),
	.w2(32'hbaf0ffa2),
	.w3(32'h3beafa9d),
	.w4(32'h3c33165b),
	.w5(32'h3bd3e89c),
	.w6(32'hbc7f40ac),
	.w7(32'hbc316b63),
	.w8(32'hbc8d297f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0e48f),
	.w1(32'hbbe2bc1e),
	.w2(32'hbbbfb571),
	.w3(32'h3c69ac5a),
	.w4(32'h3cbe8969),
	.w5(32'h3c3e486c),
	.w6(32'hbd022556),
	.w7(32'hbcb7f45d),
	.w8(32'hbca4c257),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd61eb8),
	.w1(32'h3c075b5f),
	.w2(32'h3bdafa96),
	.w3(32'h3c8ef1c6),
	.w4(32'h3c86a9f5),
	.w5(32'hbb09cd10),
	.w6(32'hbc88d455),
	.w7(32'hb97d8e9c),
	.w8(32'h3ab97b1c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22461a),
	.w1(32'h3c747ea0),
	.w2(32'h3c0a9a53),
	.w3(32'h3c446bdf),
	.w4(32'h3bce9cbc),
	.w5(32'h3c2d2b09),
	.w6(32'h3c08a9df),
	.w7(32'hba09d7b1),
	.w8(32'h3b59b53f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba646ffa),
	.w1(32'h3c0a92ac),
	.w2(32'h3a31e8d5),
	.w3(32'hbbaf5f21),
	.w4(32'h3b879693),
	.w5(32'h3c7d0e60),
	.w6(32'hbbfd3a9a),
	.w7(32'hbc8b6454),
	.w8(32'h3affb25d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc281490),
	.w1(32'h3bc2ed09),
	.w2(32'hbc409346),
	.w3(32'hba8ad109),
	.w4(32'h3c3bbf8b),
	.w5(32'hbc5f3cdc),
	.w6(32'h3b94d26f),
	.w7(32'h3af4e052),
	.w8(32'hbbab9a92),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bc623),
	.w1(32'h3b870594),
	.w2(32'hbbdcba06),
	.w3(32'h3bc85c4d),
	.w4(32'h3ba6d793),
	.w5(32'hbc18c7e3),
	.w6(32'hbbec752b),
	.w7(32'hbbba0a22),
	.w8(32'hbb999aac),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11bb48),
	.w1(32'h3b62d719),
	.w2(32'h3c08ef8f),
	.w3(32'hbbf2ac23),
	.w4(32'h3c0a853c),
	.w5(32'h3c22be81),
	.w6(32'hbb5a6f8d),
	.w7(32'hbb577988),
	.w8(32'h3b4f8379),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb1c04),
	.w1(32'hba864d3e),
	.w2(32'hbc1b3c59),
	.w3(32'h3be4ac6f),
	.w4(32'h3c837bc3),
	.w5(32'h3b7c2bd0),
	.w6(32'h3bd677c3),
	.w7(32'hb9756da6),
	.w8(32'hbc4e9676),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e64c6),
	.w1(32'h3a8b1c19),
	.w2(32'h3c327fe5),
	.w3(32'h3cbb9d80),
	.w4(32'h3ce7a5ab),
	.w5(32'h3ce0addc),
	.w6(32'hbcae498e),
	.w7(32'hbc0dd443),
	.w8(32'h3aa43c6c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d0448),
	.w1(32'hb9c71659),
	.w2(32'hbb84e2d0),
	.w3(32'hbb272e61),
	.w4(32'hbbfb64f7),
	.w5(32'h3ab4532f),
	.w6(32'hbb2920d2),
	.w7(32'hbba09981),
	.w8(32'h3b63a8f9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04b4ca),
	.w1(32'hbb7447db),
	.w2(32'hbc6acee2),
	.w3(32'hbb2ec900),
	.w4(32'hba06862b),
	.w5(32'hbc05947f),
	.w6(32'h3aa1043c),
	.w7(32'hbbe8ea98),
	.w8(32'hbc2a883a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86d743),
	.w1(32'h3c81fb02),
	.w2(32'h3c7064b0),
	.w3(32'h3d0eedb2),
	.w4(32'h3d2b0489),
	.w5(32'h3d0ec1a4),
	.w6(32'hbc61112c),
	.w7(32'hbbffa130),
	.w8(32'hbc82b9bb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86ab90),
	.w1(32'hbcee3f24),
	.w2(32'hbc87c5e1),
	.w3(32'h3c139b81),
	.w4(32'h3c423112),
	.w5(32'h399b1138),
	.w6(32'hbc94eff2),
	.w7(32'hbc7e8afd),
	.w8(32'hbc2f58c5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule