module layer_10_featuremap_92(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa76ec),
	.w1(32'h3a656f7f),
	.w2(32'h39acce72),
	.w3(32'hba85eb05),
	.w4(32'h3a8df070),
	.w5(32'hbb61580a),
	.w6(32'hba0e9d97),
	.w7(32'hba0cc282),
	.w8(32'hbb857ab6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34804a),
	.w1(32'hbba3f6c8),
	.w2(32'h3ae787c6),
	.w3(32'h3bb6d708),
	.w4(32'h3b5a3020),
	.w5(32'hbbca87e3),
	.w6(32'h3b01b4bb),
	.w7(32'h39b6775e),
	.w8(32'hbc082c9c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67971f8),
	.w1(32'hbb4a8075),
	.w2(32'h3aecf7b6),
	.w3(32'hbb17ee96),
	.w4(32'hbb0be36b),
	.w5(32'hbb958502),
	.w6(32'hba8558c9),
	.w7(32'h3ae663fd),
	.w8(32'h3baa8157),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc3600),
	.w1(32'h3b34e90c),
	.w2(32'hbb2835ac),
	.w3(32'h3b546537),
	.w4(32'hbb6b94a3),
	.w5(32'hbaa96712),
	.w6(32'hba0ca803),
	.w7(32'h3b478efb),
	.w8(32'h3bdb4748),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5af5f),
	.w1(32'hbae6e4a0),
	.w2(32'h3b381cfb),
	.w3(32'h3b3c2cad),
	.w4(32'h3af54fe3),
	.w5(32'hb982d8b2),
	.w6(32'h3bb53f81),
	.w7(32'h3b88e3af),
	.w8(32'h3c7c20b9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567533),
	.w1(32'hbb05ed59),
	.w2(32'h3a0aa5e6),
	.w3(32'h3ad7b93c),
	.w4(32'h3c080494),
	.w5(32'hbc3452b3),
	.w6(32'hbb4b76ec),
	.w7(32'h3abaf440),
	.w8(32'h3aa99b85),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9ebae),
	.w1(32'h3b3fb34f),
	.w2(32'h3bd5565d),
	.w3(32'hbb58b718),
	.w4(32'hbc1e4b6d),
	.w5(32'h3d3c754e),
	.w6(32'h3ba719ea),
	.w7(32'hbb3f15be),
	.w8(32'hbbf1ab95),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5078d),
	.w1(32'hba9d154c),
	.w2(32'hbb5b6426),
	.w3(32'h39fe9c7f),
	.w4(32'h3973b120),
	.w5(32'hb9d56bb2),
	.w6(32'h3b90fae7),
	.w7(32'hbbe5ed6b),
	.w8(32'hbb7277e2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ab9c5),
	.w1(32'h3c6879e3),
	.w2(32'h3b24c8e7),
	.w3(32'hba357585),
	.w4(32'hbae8c482),
	.w5(32'hba5b8e3e),
	.w6(32'hbb32464c),
	.w7(32'h3a4b7f74),
	.w8(32'h36eea140),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe46136),
	.w1(32'hb9823c24),
	.w2(32'h3ad9f380),
	.w3(32'hbb3dec48),
	.w4(32'hbbefcfb9),
	.w5(32'hba261f21),
	.w6(32'hbb47ecf4),
	.w7(32'hbc82d45e),
	.w8(32'h3a364068),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b38a1),
	.w1(32'hbab4028f),
	.w2(32'h3954b2d7),
	.w3(32'hbb3964b9),
	.w4(32'hbc78354f),
	.w5(32'hbb9a2737),
	.w6(32'hbac8ffe5),
	.w7(32'hb9515e2e),
	.w8(32'hba7ba487),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb481b58),
	.w1(32'hba8f1b29),
	.w2(32'h3a482cc6),
	.w3(32'hbbd819b3),
	.w4(32'hbbb91076),
	.w5(32'h3b016e46),
	.w6(32'hbac1f57a),
	.w7(32'h3ad32c5f),
	.w8(32'hbab3fed2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb613854),
	.w1(32'hbb010e53),
	.w2(32'h3be44b1d),
	.w3(32'hbb91df05),
	.w4(32'h38b72d80),
	.w5(32'hbaf05d2e),
	.w6(32'hb9a5a141),
	.w7(32'hbb7799f6),
	.w8(32'hba3ac4af),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38dd92),
	.w1(32'hbbbca4b6),
	.w2(32'hbb2dff49),
	.w3(32'hba8b2dbf),
	.w4(32'h3c048e19),
	.w5(32'h3aa11327),
	.w6(32'h3ad36282),
	.w7(32'hbc0f205b),
	.w8(32'hbb5cbf5b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf77971),
	.w1(32'hbb819507),
	.w2(32'hbb918ede),
	.w3(32'h3a1152d5),
	.w4(32'hba2f07de),
	.w5(32'h3b06a130),
	.w6(32'h3b8262f7),
	.w7(32'h3afaa958),
	.w8(32'h3b905482),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b377993),
	.w1(32'hbb35f758),
	.w2(32'h3c111cc0),
	.w3(32'h3d18365a),
	.w4(32'hba123ea7),
	.w5(32'h38d0875d),
	.w6(32'h39141c0d),
	.w7(32'h3a702f38),
	.w8(32'h3c130a55),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c6787),
	.w1(32'h3c1601ea),
	.w2(32'hba9ba908),
	.w3(32'hba8a3ef8),
	.w4(32'hb81bc608),
	.w5(32'hbc82a429),
	.w6(32'h3bb57992),
	.w7(32'h3af389ce),
	.w8(32'hbb8d3acf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb661e),
	.w1(32'h3aad3302),
	.w2(32'h3ba1bc91),
	.w3(32'hba71f0e5),
	.w4(32'h3ad6109d),
	.w5(32'h3a9a378b),
	.w6(32'h3b22226f),
	.w7(32'h3c5f922c),
	.w8(32'hbad45312),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac79a45),
	.w1(32'h3c45a31a),
	.w2(32'h3b8d41eb),
	.w3(32'hbab4188d),
	.w4(32'hba018810),
	.w5(32'hbb4c9535),
	.w6(32'hbb979f6d),
	.w7(32'h3b87a901),
	.w8(32'hbaba3c8a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed4ca0),
	.w1(32'h3942732d),
	.w2(32'hbb924141),
	.w3(32'hba74ba2d),
	.w4(32'hbb824250),
	.w5(32'hba041fe8),
	.w6(32'hbb6ee254),
	.w7(32'h3a69a9bc),
	.w8(32'hbbabb8d5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afca907),
	.w1(32'hbb430a1e),
	.w2(32'hbc6cbd84),
	.w3(32'hbb097237),
	.w4(32'hbaf807fc),
	.w5(32'hbb51c6ce),
	.w6(32'h3ca16c84),
	.w7(32'h3abe65f1),
	.w8(32'hbadd6141),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45b672),
	.w1(32'hbab08f40),
	.w2(32'hbb974ae1),
	.w3(32'h3a43d40d),
	.w4(32'h3a8da76c),
	.w5(32'hba8efc12),
	.w6(32'h3b5059d2),
	.w7(32'hb92418c6),
	.w8(32'hb8f559ff),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ca898),
	.w1(32'hba8c2b81),
	.w2(32'h3b27290a),
	.w3(32'hbaaed074),
	.w4(32'hba8b782e),
	.w5(32'hbc874800),
	.w6(32'hbb8961d6),
	.w7(32'h3977c1a9),
	.w8(32'hbc00d84a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39849304),
	.w1(32'h3b2653de),
	.w2(32'hbac7b593),
	.w3(32'hbb3582dd),
	.w4(32'h3994be37),
	.w5(32'hbb408e6a),
	.w6(32'h3acd1981),
	.w7(32'h3a814361),
	.w8(32'hbab8280f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b5ecd),
	.w1(32'hbbad4743),
	.w2(32'h3850dbbe),
	.w3(32'hbb4fe875),
	.w4(32'hbbb74ccf),
	.w5(32'h3a7415c6),
	.w6(32'h387406f6),
	.w7(32'hbab92d06),
	.w8(32'hbc2ef189),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa56c32),
	.w1(32'h3bda9332),
	.w2(32'hbbc7dedc),
	.w3(32'hbb41b8ff),
	.w4(32'h3b95f1b4),
	.w5(32'hba84e93b),
	.w6(32'hbc2f9704),
	.w7(32'hb9690d35),
	.w8(32'h3b3476eb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ad07f),
	.w1(32'h3b0e3614),
	.w2(32'hb9c8c227),
	.w3(32'hbad82da0),
	.w4(32'hbba48310),
	.w5(32'h3b208941),
	.w6(32'hba367fec),
	.w7(32'hbb4f5eeb),
	.w8(32'h3a2f33d7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3a7c4),
	.w1(32'hbbafa4ac),
	.w2(32'h3b2f7e22),
	.w3(32'h3b4008a5),
	.w4(32'hbba48005),
	.w5(32'h3ce52606),
	.w6(32'h3b47d1f0),
	.w7(32'hbc08a0b6),
	.w8(32'hba5b0a01),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b325f5c),
	.w1(32'h3b2efae7),
	.w2(32'hbca09b7d),
	.w3(32'hbb9979d9),
	.w4(32'h39afaa6f),
	.w5(32'h3a3f4daf),
	.w6(32'hb97dd07c),
	.w7(32'hb98312ce),
	.w8(32'h3b200b6b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04b9e0),
	.w1(32'hb9464ec6),
	.w2(32'hbb3ec9b3),
	.w3(32'h3ac68122),
	.w4(32'hbca5c3d6),
	.w5(32'hb9663ed3),
	.w6(32'h3a7b11fa),
	.w7(32'h3a01bd93),
	.w8(32'hbaa88cbe),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0556a1),
	.w1(32'h3ad8cd0d),
	.w2(32'h3ae5e960),
	.w3(32'h3b084b4e),
	.w4(32'h3b8c2b64),
	.w5(32'h3af58fcc),
	.w6(32'h3ab3b33e),
	.w7(32'h3a85545d),
	.w8(32'hbb0d79bd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bdff4),
	.w1(32'hbaa84ec5),
	.w2(32'h38a72f39),
	.w3(32'h3b887537),
	.w4(32'hb82c02f8),
	.w5(32'hbb1d4c1b),
	.w6(32'h3aaa1fe1),
	.w7(32'hbaac6a6b),
	.w8(32'h3b12f13f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b297b70),
	.w1(32'hbb55de56),
	.w2(32'h3af366c9),
	.w3(32'h3a132880),
	.w4(32'h3b44759b),
	.w5(32'h3af9fb9b),
	.w6(32'hba0e4ce8),
	.w7(32'h3ad2671d),
	.w8(32'hba4c7dbd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80fc23),
	.w1(32'h3b1c78c2),
	.w2(32'hbbf2a125),
	.w3(32'h3b52e4ba),
	.w4(32'h3b0d553e),
	.w5(32'hbb0ac2bf),
	.w6(32'hb738c86e),
	.w7(32'h3af11d59),
	.w8(32'hba0e24c0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa0420),
	.w1(32'h3ac1e365),
	.w2(32'hb76eb7cf),
	.w3(32'h3b7a3800),
	.w4(32'h3a5b62e9),
	.w5(32'hba0ad610),
	.w6(32'h3b72abb8),
	.w7(32'h3b2510ef),
	.w8(32'hbba9101b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a238),
	.w1(32'h3ba9a28a),
	.w2(32'h3ad5beb3),
	.w3(32'h3a485a66),
	.w4(32'hbb07731c),
	.w5(32'h3b71cf96),
	.w6(32'h3c880eaf),
	.w7(32'hbb399715),
	.w8(32'hbb2a5cfe),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91155cd),
	.w1(32'h3b387f5b),
	.w2(32'hbb30bdd2),
	.w3(32'hbc03657e),
	.w4(32'hbc33d9a3),
	.w5(32'h3cb63724),
	.w6(32'h3aceb97f),
	.w7(32'h3b42f689),
	.w8(32'hbacffc41),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0570e7),
	.w1(32'h3a67ac75),
	.w2(32'hba9a58ab),
	.w3(32'hb90b5fc2),
	.w4(32'hbbace801),
	.w5(32'hba8b8975),
	.w6(32'hbae3d5a3),
	.w7(32'hb9f9cff5),
	.w8(32'h3addc848),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1227eb),
	.w1(32'h388f49e8),
	.w2(32'hbb0d71aa),
	.w3(32'h3b08948e),
	.w4(32'h3b6e8e4d),
	.w5(32'h39013c01),
	.w6(32'hba1b4cbe),
	.w7(32'h3adf5f57),
	.w8(32'h3a578ee8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8aead7),
	.w1(32'h39de9286),
	.w2(32'hbacde2f6),
	.w3(32'h3b219046),
	.w4(32'hbc85ebdc),
	.w5(32'hb8be0aee),
	.w6(32'hbcdcbd82),
	.w7(32'h3a2ead52),
	.w8(32'hba7ac900),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb617bf35),
	.w1(32'h3acaab06),
	.w2(32'hba9bff12),
	.w3(32'hbb2dc65d),
	.w4(32'h3b143b34),
	.w5(32'hb7ac3c0e),
	.w6(32'hb88e5c55),
	.w7(32'hba343a7a),
	.w8(32'hb9b9d6c7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fa561),
	.w1(32'h3a3fe6b9),
	.w2(32'h3b43d33e),
	.w3(32'hbac4bafe),
	.w4(32'h3d198cac),
	.w5(32'hbb949c1b),
	.w6(32'h3b4bf02b),
	.w7(32'hbb3a0d22),
	.w8(32'hbb206b14),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87fbbc),
	.w1(32'hb8b089d2),
	.w2(32'hb9769bdf),
	.w3(32'h3a01efb2),
	.w4(32'hbadeab0b),
	.w5(32'hbad7dd42),
	.w6(32'h393d15a2),
	.w7(32'hbb4b9fd3),
	.w8(32'h3b287722),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9b8c8),
	.w1(32'h3a81e71a),
	.w2(32'h3b492d35),
	.w3(32'h3a5af60b),
	.w4(32'hba8e4871),
	.w5(32'h3a1a000e),
	.w6(32'h3b7c540f),
	.w7(32'h3c22fe02),
	.w8(32'hb99a0a27),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38506af3),
	.w1(32'h3ccd91f4),
	.w2(32'h3ae77598),
	.w3(32'h3a841529),
	.w4(32'h3a39a336),
	.w5(32'h3cf9604d),
	.w6(32'hba1c0210),
	.w7(32'hbb386eb3),
	.w8(32'hba3ff0c5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8568f),
	.w1(32'h39a7411a),
	.w2(32'hbad2d9a7),
	.w3(32'h3aeb42d3),
	.w4(32'hbb025ee8),
	.w5(32'hbccb2dec),
	.w6(32'hbc8ed0b2),
	.w7(32'hb9debf02),
	.w8(32'hbb68df71),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e95f7),
	.w1(32'h3a396559),
	.w2(32'hba14d304),
	.w3(32'hbc7abcd4),
	.w4(32'h3b81d836),
	.w5(32'hbc463a52),
	.w6(32'h3818dd9c),
	.w7(32'h3a3bb0de),
	.w8(32'hb99e5c22),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdab1ca),
	.w1(32'hb9e26df4),
	.w2(32'h3a3869d5),
	.w3(32'hbae413f9),
	.w4(32'hbc4a5d1e),
	.w5(32'h3ac19b9a),
	.w6(32'h39fb7efb),
	.w7(32'h3ace3dfa),
	.w8(32'hba4bf99d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab2464),
	.w1(32'hba8f7c78),
	.w2(32'h3a91dae2),
	.w3(32'hb9e390ca),
	.w4(32'hbb2a5ebd),
	.w5(32'h3b05cf39),
	.w6(32'hb9e0f7be),
	.w7(32'h3a1836de),
	.w8(32'h3a24a68d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad76385),
	.w1(32'hba79142f),
	.w2(32'hba21a8da),
	.w3(32'hba9abebb),
	.w4(32'h3b9e465c),
	.w5(32'h39d12985),
	.w6(32'hba7978f2),
	.w7(32'h3924f62d),
	.w8(32'hb9fe2955),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f9150),
	.w1(32'h3af6afd5),
	.w2(32'hba928a08),
	.w3(32'h3b465117),
	.w4(32'h3a870468),
	.w5(32'h3936f945),
	.w6(32'hba3e7869),
	.w7(32'h3b07c9c3),
	.w8(32'h39294fa6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ae13f),
	.w1(32'h385051b8),
	.w2(32'h3b1767cb),
	.w3(32'hbb1a2342),
	.w4(32'hbaabf47e),
	.w5(32'hbac1a64f),
	.w6(32'hbc85d614),
	.w7(32'h3afbf8e1),
	.w8(32'hba706132),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7fccb),
	.w1(32'hbb08d30f),
	.w2(32'hb91bd16a),
	.w3(32'hbaa17f22),
	.w4(32'h3939852a),
	.w5(32'hb992bdc6),
	.w6(32'hb8f650aa),
	.w7(32'hba3f75c4),
	.w8(32'hbaaa9e3d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12dd36),
	.w1(32'h39a6bfd6),
	.w2(32'hba397f3d),
	.w3(32'hb99ebe77),
	.w4(32'h3ad5c5c1),
	.w5(32'hba5318fd),
	.w6(32'hb9f78176),
	.w7(32'h3b634840),
	.w8(32'hbb985c33),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0296c2),
	.w1(32'h3b2efb57),
	.w2(32'h3b09c600),
	.w3(32'h3a5a2ccc),
	.w4(32'hba24f4be),
	.w5(32'h3b10583e),
	.w6(32'h39e62923),
	.w7(32'h3b046da3),
	.w8(32'h3b13c9f8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdf1a3),
	.w1(32'hbc81d778),
	.w2(32'h3b9da6f1),
	.w3(32'hbc62f54c),
	.w4(32'h3c0370fe),
	.w5(32'hbc2d20eb),
	.w6(32'h398364ba),
	.w7(32'hbc0b7902),
	.w8(32'hba104059),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfbb764),
	.w1(32'h399e2f8f),
	.w2(32'h3ab8d7a6),
	.w3(32'h3c400d3e),
	.w4(32'hbaac64c3),
	.w5(32'hbbd0350a),
	.w6(32'h39199445),
	.w7(32'hbb798e87),
	.w8(32'hbbba351b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ad92e),
	.w1(32'h39b6e089),
	.w2(32'h3c0930ee),
	.w3(32'h3b13126f),
	.w4(32'hbaf73cf2),
	.w5(32'h3b043a49),
	.w6(32'h3c3c733e),
	.w7(32'h3c29e401),
	.w8(32'h3c4454f4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2eaff),
	.w1(32'h3b8e0f00),
	.w2(32'hba9c6bec),
	.w3(32'h3aff1602),
	.w4(32'h3bd10c54),
	.w5(32'h395e9b29),
	.w6(32'hbc010478),
	.w7(32'hba0901e8),
	.w8(32'h3c079718),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac1f3a),
	.w1(32'h3adcf0c1),
	.w2(32'h3c1257e7),
	.w3(32'h3d9091b1),
	.w4(32'hbb7405a7),
	.w5(32'hbbc411da),
	.w6(32'hbb267b4e),
	.w7(32'hbbc5cfe9),
	.w8(32'hb9f180c4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd206c32),
	.w1(32'hbc0ca3af),
	.w2(32'hbb233973),
	.w3(32'hbbffd90e),
	.w4(32'h3b6d94bf),
	.w5(32'h39c82e92),
	.w6(32'hbb8b9abf),
	.w7(32'hbbebe9b6),
	.w8(32'h3beefe6c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb86ea),
	.w1(32'h3a06533f),
	.w2(32'h3a9e081a),
	.w3(32'hba137516),
	.w4(32'h38b77225),
	.w5(32'hbc84e146),
	.w6(32'h3bf07328),
	.w7(32'hbba7c4d3),
	.w8(32'h3be95438),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dca5d),
	.w1(32'hbad9e835),
	.w2(32'h3be9f3e4),
	.w3(32'hbb6d92eb),
	.w4(32'hbb312141),
	.w5(32'h3bb52217),
	.w6(32'hbb26d392),
	.w7(32'h3b4e1f1c),
	.w8(32'hbb8c887d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ab16e),
	.w1(32'hba9100c3),
	.w2(32'h3b736e61),
	.w3(32'hba498898),
	.w4(32'hbc080e34),
	.w5(32'hbafdb2d0),
	.w6(32'hbc0a329e),
	.w7(32'h3be4a222),
	.w8(32'h3c25be9b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e3bce),
	.w1(32'hbb4d5ae3),
	.w2(32'h3b3771c6),
	.w3(32'hbca3f25b),
	.w4(32'h3bd557f7),
	.w5(32'hbbfdc3e8),
	.w6(32'hbb7d0cc7),
	.w7(32'hbb9026ff),
	.w8(32'hb96f237d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfbcd3),
	.w1(32'hbc7a59ac),
	.w2(32'hbbd245b8),
	.w3(32'h3a93b4df),
	.w4(32'hbb2abff0),
	.w5(32'h37a967fa),
	.w6(32'hbbb7063c),
	.w7(32'hbc232ae3),
	.w8(32'hbd752af6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a3843),
	.w1(32'h39aafffd),
	.w2(32'h3a9cb78c),
	.w3(32'h3acae974),
	.w4(32'hbc147f36),
	.w5(32'hbc32f20b),
	.w6(32'h3b12c1d7),
	.w7(32'h3a83f7e1),
	.w8(32'h3b8b3fd1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd07a88),
	.w1(32'hbba6f350),
	.w2(32'hbb309a58),
	.w3(32'h3a82dbe7),
	.w4(32'hb9e55f10),
	.w5(32'hbb09930e),
	.w6(32'hbaeeefb6),
	.w7(32'hbc04c383),
	.w8(32'hb9df0b94),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a7912),
	.w1(32'hbd42e89c),
	.w2(32'h3a1403cb),
	.w3(32'hbbc70fdd),
	.w4(32'h39e9204c),
	.w5(32'hbb76d29b),
	.w6(32'h3b0ddbe5),
	.w7(32'hbd94d350),
	.w8(32'hbc59e849),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78cdbc),
	.w1(32'hbb817b25),
	.w2(32'h3b829169),
	.w3(32'h3c8b1d2d),
	.w4(32'hbc0566d4),
	.w5(32'hbc0f3839),
	.w6(32'hbbf395d0),
	.w7(32'h3a13bb81),
	.w8(32'h3b135435),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf50fc9),
	.w1(32'h3d38e790),
	.w2(32'h3ac3f249),
	.w3(32'h3a85b834),
	.w4(32'h39e01fa7),
	.w5(32'hbbaadc24),
	.w6(32'hbcaa554c),
	.w7(32'hbbd4745f),
	.w8(32'hbcf4947d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba889100),
	.w1(32'hbc39b7c7),
	.w2(32'h3b8dbbf5),
	.w3(32'hbac17bc4),
	.w4(32'hbc17871b),
	.w5(32'hb8be401e),
	.w6(32'h3a52e2ed),
	.w7(32'hbaa5d0fb),
	.w8(32'hbb44449d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb692558),
	.w1(32'h3a01cc9d),
	.w2(32'hbbfc3ed7),
	.w3(32'h3b5b2796),
	.w4(32'h39d16596),
	.w5(32'h3c4acd6f),
	.w6(32'hbc005e9c),
	.w7(32'hbae25387),
	.w8(32'hbac96762),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a863630),
	.w1(32'hb8cbfaee),
	.w2(32'hbabe7d64),
	.w3(32'h3b77a83e),
	.w4(32'hbba18041),
	.w5(32'hbc191403),
	.w6(32'hb93c4a20),
	.w7(32'hbaf9eb58),
	.w8(32'hbc20b206),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac79a68),
	.w1(32'hbb8931f6),
	.w2(32'hb826aa64),
	.w3(32'h3ae5f304),
	.w4(32'hbc910e70),
	.w5(32'hbbcfb25b),
	.w6(32'h3ac4f11a),
	.w7(32'hbbab1260),
	.w8(32'hbb898616),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae03fef),
	.w1(32'hb9133257),
	.w2(32'hbd1fcb6d),
	.w3(32'hba81b375),
	.w4(32'hbbddcf7a),
	.w5(32'hbb2580cf),
	.w6(32'hbc3c1fb5),
	.w7(32'hbb49632a),
	.w8(32'hbae3e530),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc048e0d),
	.w1(32'hbc02db0f),
	.w2(32'hbbdfbddc),
	.w3(32'hbbb8051a),
	.w4(32'hbbcc4dc5),
	.w5(32'hbb7739b0),
	.w6(32'hbcde9291),
	.w7(32'hbc3ca8e0),
	.w8(32'hbb842772),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2f6a7),
	.w1(32'hbc33077f),
	.w2(32'hba901c09),
	.w3(32'hbb3f0d3f),
	.w4(32'hbc920ca9),
	.w5(32'hbc1f1a77),
	.w6(32'hbbb7630e),
	.w7(32'hbb97ce22),
	.w8(32'hbc83479d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7c60c),
	.w1(32'hbb962b27),
	.w2(32'h3b06dc44),
	.w3(32'hbba82fb5),
	.w4(32'hb84d5513),
	.w5(32'h3b5484de),
	.w6(32'hbb13da3b),
	.w7(32'h3b881029),
	.w8(32'hbc29926e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd210ef),
	.w1(32'hba06933e),
	.w2(32'h3c4dde46),
	.w3(32'hbb20c153),
	.w4(32'hbb959b20),
	.w5(32'hbce60755),
	.w6(32'h388fa47e),
	.w7(32'h3c3def1a),
	.w8(32'h3b9a1eb1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7cfda),
	.w1(32'h3c034db5),
	.w2(32'hbbd96aad),
	.w3(32'h3c2f9837),
	.w4(32'hbcd07c7e),
	.w5(32'h3bac704c),
	.w6(32'hbb12b5e9),
	.w7(32'h3c0c66cb),
	.w8(32'h3b1f54ee),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b478),
	.w1(32'hbd1e353f),
	.w2(32'h3b89a011),
	.w3(32'h3bcb3390),
	.w4(32'hba9842da),
	.w5(32'h3c27a9e2),
	.w6(32'h3bad7103),
	.w7(32'hbb9ed7c3),
	.w8(32'hbc765753),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8b1da),
	.w1(32'hbae20e7d),
	.w2(32'h3b5747a2),
	.w3(32'h3aa77958),
	.w4(32'hbb68e2c9),
	.w5(32'hbbc66cc3),
	.w6(32'h3b807f09),
	.w7(32'h3bcb8f88),
	.w8(32'hbbccad9e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2eca7),
	.w1(32'hbab0eb13),
	.w2(32'h3c0daeb5),
	.w3(32'h3995f95c),
	.w4(32'hbbd1f769),
	.w5(32'hbbb63655),
	.w6(32'hb9c0d7f2),
	.w7(32'h3ba79e90),
	.w8(32'hbab23e7f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a6b4e),
	.w1(32'hba625ae0),
	.w2(32'hbb8c1ab7),
	.w3(32'h3acdef54),
	.w4(32'hbd3cf55e),
	.w5(32'hbb834ee3),
	.w6(32'hbbe3f3b3),
	.w7(32'hbb6585f7),
	.w8(32'h3a2834ce),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab91e8),
	.w1(32'hbb0779b2),
	.w2(32'h3adcc26e),
	.w3(32'hbb46a560),
	.w4(32'hbb3b3091),
	.w5(32'h3b45ed99),
	.w6(32'h3b946e5b),
	.w7(32'h3c3c51d7),
	.w8(32'h3ba1b2b0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf35230),
	.w1(32'h3c92f467),
	.w2(32'hbc504aa1),
	.w3(32'h3bb70c29),
	.w4(32'h3c0737c1),
	.w5(32'hbb558ba0),
	.w6(32'h3b72accf),
	.w7(32'hbaceb308),
	.w8(32'hbbad44d0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fdd1c),
	.w1(32'hbbfa2b45),
	.w2(32'hbbe34d73),
	.w3(32'hbb238bc1),
	.w4(32'h3b904e3c),
	.w5(32'hbbbc5b9e),
	.w6(32'h3ac78def),
	.w7(32'hbbedb967),
	.w8(32'h3b013c40),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add9bfd),
	.w1(32'h3bef1ba5),
	.w2(32'h3b4bd213),
	.w3(32'hbb70830d),
	.w4(32'h3be8ec08),
	.w5(32'hbb1d0eb5),
	.w6(32'hbb4847a6),
	.w7(32'hbb606d69),
	.w8(32'hba352f8d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a819f),
	.w1(32'hb9846ec5),
	.w2(32'h3bebc678),
	.w3(32'hbb23fd69),
	.w4(32'hbc116a0d),
	.w5(32'hbad484dd),
	.w6(32'hbafab409),
	.w7(32'hb88deded),
	.w8(32'h3c096b4a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c501f),
	.w1(32'hbadaa0ce),
	.w2(32'hb915b871),
	.w3(32'h3adfe9eb),
	.w4(32'h3ac0acc9),
	.w5(32'h3b8d9587),
	.w6(32'hbd07b499),
	.w7(32'h3c7d9008),
	.w8(32'hbb51c258),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cbc3a),
	.w1(32'hb976b5d6),
	.w2(32'h3bc4cd56),
	.w3(32'hbbe7c094),
	.w4(32'h3b0f9a1d),
	.w5(32'h3a379616),
	.w6(32'h3a145ae6),
	.w7(32'hba94fe8e),
	.w8(32'hbbacd43f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b313ffe),
	.w1(32'h386f8b75),
	.w2(32'h3bc7331b),
	.w3(32'h3dc843be),
	.w4(32'h3b18ec3f),
	.w5(32'hbb2a958c),
	.w6(32'hbc0952d6),
	.w7(32'hbb30497f),
	.w8(32'hbb38f832),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c111b54),
	.w1(32'hbb8f41e9),
	.w2(32'h3cefdfaf),
	.w3(32'h381838a7),
	.w4(32'h3b8bf819),
	.w5(32'hbb7c5670),
	.w6(32'hbb07393b),
	.w7(32'hbc0dfd9c),
	.w8(32'hbb5bf631),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5cdbf),
	.w1(32'hbcaf8eff),
	.w2(32'h3a2497d5),
	.w3(32'hbb25eb52),
	.w4(32'h3b97331b),
	.w5(32'hbb23ff79),
	.w6(32'h3a77269d),
	.w7(32'hbaf6b885),
	.w8(32'hbd1151fb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ba437),
	.w1(32'hbb89726c),
	.w2(32'hbb4949de),
	.w3(32'hb8f31ae7),
	.w4(32'h38c98a95),
	.w5(32'hbd08c01c),
	.w6(32'h3ba47923),
	.w7(32'h3bb3267e),
	.w8(32'h3ac130ca),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5135c),
	.w1(32'h3bba427e),
	.w2(32'hbaa2708f),
	.w3(32'h3b6f79fe),
	.w4(32'hba10f97b),
	.w5(32'hbc5f0a6f),
	.w6(32'h3b28a82f),
	.w7(32'h3bd10b67),
	.w8(32'h37dec3a6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d8754),
	.w1(32'hbba87229),
	.w2(32'hbb23bddd),
	.w3(32'hb986ba4e),
	.w4(32'h3b62d3ef),
	.w5(32'h3b27ded4),
	.w6(32'hbb9eabcc),
	.w7(32'hbba45fc5),
	.w8(32'hbb595e43),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7f9f1),
	.w1(32'h3c8b769f),
	.w2(32'hbc4ab57e),
	.w3(32'h3aa476e8),
	.w4(32'hbbe261bd),
	.w5(32'h3c0ca9ab),
	.w6(32'h3af1d460),
	.w7(32'hbbbeefe7),
	.w8(32'hbc829f22),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ba4b7),
	.w1(32'hbb34a0ef),
	.w2(32'h3a52fdfd),
	.w3(32'hbb410440),
	.w4(32'hbbd8be81),
	.w5(32'hba6c6875),
	.w6(32'hbae5548c),
	.w7(32'hbb56b50f),
	.w8(32'hbbe4ca86),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c100b52),
	.w1(32'h3a8f0293),
	.w2(32'hbbb98c02),
	.w3(32'h3b96a44b),
	.w4(32'h3db17bba),
	.w5(32'hba910a12),
	.w6(32'h3c7efb72),
	.w7(32'h3ba677b1),
	.w8(32'hbb0831fd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fca80),
	.w1(32'h3aa61f2a),
	.w2(32'h3ce4fa60),
	.w3(32'hba2db597),
	.w4(32'h3bb545dd),
	.w5(32'hb9dc8d4b),
	.w6(32'h3c510749),
	.w7(32'h3a85094d),
	.w8(32'hb9232e74),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacb254),
	.w1(32'hbbc39be1),
	.w2(32'h3adc5e2c),
	.w3(32'hbd2f3623),
	.w4(32'hbb36ad5c),
	.w5(32'h3b9fe9f3),
	.w6(32'hbb3a1494),
	.w7(32'h3b375e54),
	.w8(32'hbc9cafb1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accefa3),
	.w1(32'h3c87b1f9),
	.w2(32'h3cda4a59),
	.w3(32'h3afdfb28),
	.w4(32'h3b5f2125),
	.w5(32'hb98049db),
	.w6(32'h39084e8f),
	.w7(32'hbbd81cca),
	.w8(32'h3ac935bf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e6819),
	.w1(32'h3c88e73f),
	.w2(32'h3b0e9d27),
	.w3(32'hbb023770),
	.w4(32'hbbbabdd8),
	.w5(32'hba936ed7),
	.w6(32'h3ad366ef),
	.w7(32'h3b823052),
	.w8(32'hba9b68a3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff530d),
	.w1(32'hbb96e01b),
	.w2(32'hbb8b4ae3),
	.w3(32'hbb59935f),
	.w4(32'hbc23e0d3),
	.w5(32'h3a138953),
	.w6(32'hbc44c900),
	.w7(32'h3d557c59),
	.w8(32'h3bc990bc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48571f),
	.w1(32'hbbfd4d16),
	.w2(32'h3bac708c),
	.w3(32'hbb067515),
	.w4(32'h39524b65),
	.w5(32'h3b930131),
	.w6(32'hbb897963),
	.w7(32'h3b24fc3c),
	.w8(32'hba02e60b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad3e35),
	.w1(32'h3aaaf894),
	.w2(32'h396fd1e1),
	.w3(32'hba517726),
	.w4(32'h3b69d90b),
	.w5(32'hbb93bd9f),
	.w6(32'h3bd4d1fd),
	.w7(32'hbb030506),
	.w8(32'hbbc92c7a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf4dd12),
	.w1(32'hbb64b71e),
	.w2(32'h3a0fd908),
	.w3(32'hbc079553),
	.w4(32'h3b447705),
	.w5(32'hbbca4789),
	.w6(32'hbbadaa43),
	.w7(32'h39f0519e),
	.w8(32'hbb8cb6fc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b91f4),
	.w1(32'hbb385842),
	.w2(32'hbac6cf3e),
	.w3(32'h3a6ec1ae),
	.w4(32'h3b95c8d1),
	.w5(32'h3b107fd8),
	.w6(32'hbbd1c2ae),
	.w7(32'hbc06ecde),
	.w8(32'hbafc7f43),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a3341),
	.w1(32'h3bc64e79),
	.w2(32'hbbb41acc),
	.w3(32'h3ba31313),
	.w4(32'hbb5b9c4d),
	.w5(32'h3c7c5c29),
	.w6(32'hbb885a94),
	.w7(32'hbd01d20e),
	.w8(32'h3b8dda4a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78b823),
	.w1(32'hba9d8145),
	.w2(32'h39ae7f36),
	.w3(32'hbb936853),
	.w4(32'hbb782701),
	.w5(32'hb8b03443),
	.w6(32'hba93265b),
	.w7(32'h3beb18b7),
	.w8(32'h3b8e37da),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc014a19),
	.w1(32'h3a873637),
	.w2(32'hbadf04c7),
	.w3(32'h3b410427),
	.w4(32'h3aa65bf4),
	.w5(32'h3b900743),
	.w6(32'hbaa89439),
	.w7(32'hba4c0e1b),
	.w8(32'hbbb73c84),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ad71d),
	.w1(32'h3aab9d6f),
	.w2(32'h3af437a5),
	.w3(32'h3c8d847f),
	.w4(32'hbb1456b8),
	.w5(32'hba557794),
	.w6(32'hbabf5cdd),
	.w7(32'hbb901e6b),
	.w8(32'h380450fc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb224b06),
	.w1(32'hbb9aae5b),
	.w2(32'h39dcbb4a),
	.w3(32'hbbcab165),
	.w4(32'h3aeab68a),
	.w5(32'hbc2411f6),
	.w6(32'h39e46839),
	.w7(32'hba8c1bbe),
	.w8(32'hba04a7ea),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ca3d5),
	.w1(32'hb8c9bbbd),
	.w2(32'h3abddeb7),
	.w3(32'hbb6d73da),
	.w4(32'h3a8f0ea9),
	.w5(32'hbb696512),
	.w6(32'h3af82766),
	.w7(32'h3b048e2d),
	.w8(32'hbb3368cf),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bb8df),
	.w1(32'h3a7a6218),
	.w2(32'h3b96ccba),
	.w3(32'h3b389b15),
	.w4(32'hb9e84e91),
	.w5(32'hb971c00d),
	.w6(32'h3c912e09),
	.w7(32'h3b38e54c),
	.w8(32'h3ba34feb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0efb4),
	.w1(32'hbb2c98f8),
	.w2(32'h3a81cb47),
	.w3(32'h3bec057e),
	.w4(32'hbb22d17e),
	.w5(32'hba52090f),
	.w6(32'hbb5cd8f3),
	.w7(32'hbbd6d131),
	.w8(32'h3b687fb3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba298c1d),
	.w1(32'h3b283418),
	.w2(32'h3b70d46b),
	.w3(32'hbb183a54),
	.w4(32'hbb2f2303),
	.w5(32'hbb8192f9),
	.w6(32'hb93ce84e),
	.w7(32'h3a05b65a),
	.w8(32'h35edb344),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c6733),
	.w1(32'hbb49f9c3),
	.w2(32'hba288896),
	.w3(32'h3b164b3e),
	.w4(32'h3840da86),
	.w5(32'h39e2cf61),
	.w6(32'h3a89dcf8),
	.w7(32'hbabf6b9a),
	.w8(32'hba0281e9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0dfb7),
	.w1(32'hbb6faa2c),
	.w2(32'h39fb9315),
	.w3(32'hbad2558e),
	.w4(32'hbae78fe5),
	.w5(32'h3b740af6),
	.w6(32'hbc02bf57),
	.w7(32'h3ce5c6da),
	.w8(32'h3b97fca8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22be1a),
	.w1(32'h3b90ef16),
	.w2(32'hba339fa8),
	.w3(32'h3b14463b),
	.w4(32'hbbc81187),
	.w5(32'hbb8a3646),
	.w6(32'hbae13588),
	.w7(32'h3a856c4c),
	.w8(32'h3b08c06e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacc99c),
	.w1(32'h3ae46268),
	.w2(32'hba9601e1),
	.w3(32'h3c8d96ec),
	.w4(32'hbb14db6f),
	.w5(32'hbadf64a0),
	.w6(32'hb86c4089),
	.w7(32'h3acaf8bb),
	.w8(32'hbb3b90de),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc56adf),
	.w1(32'hbc6b05eb),
	.w2(32'h3b7e556a),
	.w3(32'h37d9cdbc),
	.w4(32'h3a7113f7),
	.w5(32'hbb68b392),
	.w6(32'hbb883613),
	.w7(32'h3a024643),
	.w8(32'h3b300f89),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dad72),
	.w1(32'hbb01e5f0),
	.w2(32'hbb44ee3a),
	.w3(32'hba6afc13),
	.w4(32'hb8e3d77b),
	.w5(32'hbb6dec7a),
	.w6(32'hbbae8083),
	.w7(32'hbb44b0b9),
	.w8(32'hba89e228),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56c121),
	.w1(32'h34cea334),
	.w2(32'hbb09c061),
	.w3(32'hbb124222),
	.w4(32'h3b4a4449),
	.w5(32'h3a75b202),
	.w6(32'hbbce5280),
	.w7(32'h37e48a48),
	.w8(32'h3bbaffa2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a8a1b),
	.w1(32'hbb1629c5),
	.w2(32'h38ef4ec6),
	.w3(32'hba99ad92),
	.w4(32'h3b0a1c09),
	.w5(32'h3d015906),
	.w6(32'h3b1068aa),
	.w7(32'h3b2faac1),
	.w8(32'hbb0cb36b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafd00e),
	.w1(32'h3bba1d74),
	.w2(32'h3b527526),
	.w3(32'hbbbff91f),
	.w4(32'hbb60cfe1),
	.w5(32'h3c0de643),
	.w6(32'hbc9b19c7),
	.w7(32'hba15ff68),
	.w8(32'h39c5056d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb625a91),
	.w1(32'h3a27c40b),
	.w2(32'h3a406e54),
	.w3(32'hb9cf71e1),
	.w4(32'hbb02070b),
	.w5(32'h3abebd91),
	.w6(32'hbac319bd),
	.w7(32'h3aaec3c6),
	.w8(32'h3c59e082),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ffa91),
	.w1(32'hbb0740dc),
	.w2(32'h3ccd367f),
	.w3(32'hbb06d805),
	.w4(32'hb96c07e8),
	.w5(32'h3a4c042d),
	.w6(32'h3a74c008),
	.w7(32'h3b7890af),
	.w8(32'hba839f68),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb911c),
	.w1(32'hb989cfd7),
	.w2(32'hbafddacf),
	.w3(32'h3ca7f05e),
	.w4(32'h3a83f397),
	.w5(32'hbb3c5d3c),
	.w6(32'hb98d9a0a),
	.w7(32'hbc3882d9),
	.w8(32'hba29327f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb112533),
	.w1(32'h3a95885a),
	.w2(32'h39e5ff20),
	.w3(32'hbbc92ed7),
	.w4(32'h3a60ed46),
	.w5(32'h3caa6ec4),
	.w6(32'hba4152d3),
	.w7(32'h397f3342),
	.w8(32'hbab4ee47),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba172f0d),
	.w1(32'h3bb17b6b),
	.w2(32'h3a0ecb4c),
	.w3(32'h3b45cd5f),
	.w4(32'h3b2a637d),
	.w5(32'h3b059df9),
	.w6(32'h3bad0226),
	.w7(32'hbbae8d2f),
	.w8(32'hba9950f1),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada4064),
	.w1(32'h3b0ff3bc),
	.w2(32'hbac388a9),
	.w3(32'hb9962d26),
	.w4(32'hbb3e1597),
	.w5(32'hbb2cb8fb),
	.w6(32'hbbb20a5e),
	.w7(32'hb97347e2),
	.w8(32'hb989ee5a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a941d0a),
	.w1(32'hbae2bf57),
	.w2(32'hbadcf968),
	.w3(32'hbb713bd3),
	.w4(32'hbbf6eb81),
	.w5(32'h3bc8e618),
	.w6(32'h3b03704e),
	.w7(32'h3b0b33c4),
	.w8(32'h3a269721),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb055ce6),
	.w1(32'hb9d25b49),
	.w2(32'h3b02c07f),
	.w3(32'h3b699bb2),
	.w4(32'h398ffabc),
	.w5(32'hbb7214d3),
	.w6(32'h3b05d6cf),
	.w7(32'hba74bc20),
	.w8(32'h3bdb774f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb159d53),
	.w1(32'hbb094079),
	.w2(32'h3a492c31),
	.w3(32'hba1cd9c0),
	.w4(32'hbb93020d),
	.w5(32'h3a968881),
	.w6(32'hba3b5148),
	.w7(32'hbc8b0f3c),
	.w8(32'hbb14b111),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ac6d7),
	.w1(32'h3a2f6380),
	.w2(32'h3a3d88d4),
	.w3(32'hbb1ccb11),
	.w4(32'h39fee356),
	.w5(32'h3a2532dc),
	.w6(32'hbacaeb8f),
	.w7(32'hbb099a5f),
	.w8(32'hbbb1235a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc63072),
	.w1(32'hbab4e40e),
	.w2(32'hbbd44388),
	.w3(32'hba9489b0),
	.w4(32'h3c32b061),
	.w5(32'hbb85290c),
	.w6(32'hbb12c156),
	.w7(32'hb9a56afc),
	.w8(32'hbb9db405),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe7fc2),
	.w1(32'h3b5d77bb),
	.w2(32'h3b4b07fc),
	.w3(32'h3b946ef7),
	.w4(32'hbb42fb04),
	.w5(32'h3ad50f47),
	.w6(32'h3b9290c5),
	.w7(32'hbbc363c2),
	.w8(32'hbb4bfe73),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e6d4e),
	.w1(32'hba39c87e),
	.w2(32'hbf19f260),
	.w3(32'h3ae41a54),
	.w4(32'hbf028551),
	.w5(32'hbf01fbad),
	.w6(32'h3b0c7fa3),
	.w7(32'hbe701ea3),
	.w8(32'hbf36c1cb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeeb6423),
	.w1(32'hbfbf6dbe),
	.w2(32'hbe96a8ef),
	.w3(32'hbf0718e5),
	.w4(32'hbfc7f03b),
	.w5(32'hbf035d34),
	.w6(32'hbf290dc4),
	.w7(32'h3f04f976),
	.w8(32'hbf0f950d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf0f6def),
	.w1(32'hbf1a192f),
	.w2(32'hbf131c39),
	.w3(32'hbeeb6959),
	.w4(32'h3e149779),
	.w5(32'hbf026288),
	.w6(32'hbe8ee2a1),
	.w7(32'hbeecaedb),
	.w8(32'hbedff42e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf147f22),
	.w1(32'hbebdc47f),
	.w2(32'hbe881f8b),
	.w3(32'hbf0683d0),
	.w4(32'hbf042d5e),
	.w5(32'hbf347828),
	.w6(32'h3f901a01),
	.w7(32'hbf0f2d17),
	.w8(32'hbecc16c3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1eec5e),
	.w1(32'hbf055f4d),
	.w2(32'hbf333402),
	.w3(32'hbedb85cf),
	.w4(32'h3e101577),
	.w5(32'hbf310db7),
	.w6(32'hbeafaff9),
	.w7(32'hbe9ab31b),
	.w8(32'hbf05ff38),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf00bbcb),
	.w1(32'hbf07cd52),
	.w2(32'hbe5258c3),
	.w3(32'hbf159cb3),
	.w4(32'hbf06fb99),
	.w5(32'hbf3b5bcb),
	.w6(32'hbf0dc81d),
	.w7(32'hbf15abcf),
	.w8(32'hbf06cc4c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf0b1e96),
	.w1(32'hbead3793),
	.w2(32'hbf06708d),
	.w3(32'hbf1e81f4),
	.w4(32'hbf5077ec),
	.w5(32'hbf102a53),
	.w6(32'hbefa1a23),
	.w7(32'hbf04db0d),
	.w8(32'hbedb81a2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf13d9c5),
	.w1(32'hbee425ab),
	.w2(32'hbf14c0fd),
	.w3(32'hbcb2a31a),
	.w4(32'hbf0c4b04),
	.w5(32'hbebd765b),
	.w6(32'hbece51e5),
	.w7(32'hbef01f39),
	.w8(32'hbf148a13),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf223291),
	.w1(32'hbf01d494),
	.w2(32'hbeb11bdc),
	.w3(32'hbf72c2fa),
	.w4(32'hbef3c349),
	.w5(32'hbf143dda),
	.w6(32'hbefc7ec9),
	.w7(32'hbf052659),
	.w8(32'hbf0eb771),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf05d008),
	.w1(32'hbf32ccbc),
	.w2(32'hbf0bc25b),
	.w3(32'hbeb13705),
	.w4(32'hbd09ad92),
	.w5(32'hbd948c34),
	.w6(32'hbeec5750),
	.w7(32'hbf07fbe1),
	.w8(32'hbeb3196f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbee23839),
	.w1(32'hbee290b8),
	.w2(32'hbec9c758),
	.w3(32'hbe9f3bf5),
	.w4(32'hbf059e7f),
	.w5(32'hbee26c01),
	.w6(32'h3f001d5e),
	.w7(32'h3f387281),
	.w8(32'hbf577917),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf0b715a),
	.w1(32'hbf3af9e7),
	.w2(32'hbf0e525e),
	.w3(32'hbe77101c),
	.w4(32'hbefffbc6),
	.w5(32'hbf1f5260),
	.w6(32'h3e5661d0),
	.w7(32'hbf032a77),
	.w8(32'hbeb76a08),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf17899c),
	.w1(32'hbe002757),
	.w2(32'hbf01a8a8),
	.w3(32'hbedd79ad),
	.w4(32'hbec25b58),
	.w5(32'hbefe571a),
	.w6(32'hbf219ae5),
	.w7(32'hbec31e01),
	.w8(32'hbede65ca),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f639a64),
	.w1(32'hbf07bf1a),
	.w2(32'hbdac1cfd),
	.w3(32'hbf05af80),
	.w4(32'hbecd341b),
	.w5(32'hbf0dd2e9),
	.w6(32'hbd95a5df),
	.w7(32'hbee263dd),
	.w8(32'h3d67ff4c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbecb3cb8),
	.w1(32'hbed0e397),
	.w2(32'hbf054fe2),
	.w3(32'hbf585c26),
	.w4(32'hbd05863d),
	.w5(32'hbf020c06),
	.w6(32'hbf48daea),
	.w7(32'hbed48253),
	.w8(32'hbf7e3529),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeede05c),
	.w1(32'hbf00125a),
	.w2(32'hbca67b21),
	.w3(32'hbf7c2cda),
	.w4(32'hbed3c0c6),
	.w5(32'hbfd54531),
	.w6(32'h3f540b05),
	.w7(32'hbdace2b2),
	.w8(32'hbf5c8f85),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf162fa5),
	.w1(32'hbf0173e9),
	.w2(32'hbeff27ce),
	.w3(32'hbf2bd5a5),
	.w4(32'hbf1f6858),
	.w5(32'hbf0512f8),
	.w6(32'hbe885d5f),
	.w7(32'hbf0c367d),
	.w8(32'hbf0a4616),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbed9e9dd),
	.w1(32'hbee032ed),
	.w2(32'hbee85055),
	.w3(32'hbf1b6f2e),
	.w4(32'hbf08db3e),
	.w5(32'hbf0ed28a),
	.w6(32'hbefef282),
	.w7(32'hbe9dc46c),
	.w8(32'hbeb6b814),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1ea02a),
	.w1(32'hbf1130cb),
	.w2(32'hbf0d6af0),
	.w3(32'h3f097777),
	.w4(32'hbf0ee65d),
	.w5(32'hbef845c3),
	.w6(32'hbecf0cfc),
	.w7(32'hbf5f9427),
	.w8(32'hbee6716c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf453b84),
	.w1(32'hbf0c4bba),
	.w2(32'hbee6c725),
	.w3(32'hbe65e502),
	.w4(32'hbf3a3fd5),
	.w5(32'hbdf7918b),
	.w6(32'hbebaf31f),
	.w7(32'hbe672876),
	.w8(32'hbe3c3573),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbefb00db),
	.w1(32'hbf01759d),
	.w2(32'hbf083a7c),
	.w3(32'hbf030354),
	.w4(32'hbec91b96),
	.w5(32'hbf334a79),
	.w6(32'hbefe27b2),
	.w7(32'hbe9cff6f),
	.w8(32'hbf0b7e28),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeee5bf5),
	.w1(32'hbe04ff16),
	.w2(32'h3dbc0864),
	.w3(32'hbf0bedbc),
	.w4(32'hbf16386c),
	.w5(32'hbee13f0e),
	.w6(32'h3f186eb6),
	.w7(32'hbf1a39a9),
	.w8(32'hbf00286a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf009d27),
	.w1(32'hbeef06d3),
	.w2(32'hbee72506),
	.w3(32'hbf00544b),
	.w4(32'hbf775dcf),
	.w5(32'hbf082929),
	.w6(32'hbea97a2d),
	.w7(32'hbe2b9b37),
	.w8(32'hbeb8dace),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeba96c4),
	.w1(32'hbf0e2615),
	.w2(32'hbf0e8de0),
	.w3(32'hbf6f49b1),
	.w4(32'hbedd2f4e),
	.w5(32'hbefb658c),
	.w6(32'hbe1404a1),
	.w7(32'hbf2318fa),
	.w8(32'hbef16d07),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf3202a1),
	.w1(32'hbf0c1356),
	.w2(32'hbf03cf46),
	.w3(32'hbeb0a4f9),
	.w4(32'hbf116df1),
	.w5(32'hbf014e52),
	.w6(32'hbf0ce41d),
	.w7(32'hbe9c92e9),
	.w8(32'h3eeac74e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7ab3d9),
	.w1(32'hbf4a3f0e),
	.w2(32'hbf212ba1),
	.w3(32'hbf417a82),
	.w4(32'hbecd6912),
	.w5(32'hbec9354b),
	.w6(32'hbedd1ce0),
	.w7(32'hbf281722),
	.w8(32'hbed4c17e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf3861df),
	.w1(32'hbf54ad5b),
	.w2(32'hbeadfa13),
	.w3(32'hbf0b15b9),
	.w4(32'hbeba083b),
	.w5(32'hbf00f9d7),
	.w6(32'hbf09448e),
	.w7(32'hbf088c9f),
	.w8(32'hbf3dc1a9),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbedfa1cb),
	.w1(32'hbef5cb9b),
	.w2(32'hbf36a228),
	.w3(32'hbe9f6849),
	.w4(32'hbf7b3699),
	.w5(32'hbef6fd2f),
	.w6(32'h3dce298c),
	.w7(32'hbf109cdb),
	.w8(32'hbf2034c0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec5525a),
	.w1(32'hbeb76990),
	.w2(32'hbeea22cf),
	.w3(32'hbed4a475),
	.w4(32'hbed12bfa),
	.w5(32'hbf197af7),
	.w6(32'hbf15e285),
	.w7(32'hbea220cb),
	.w8(32'h3c279260),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e46248a),
	.w1(32'h3eb6aa46),
	.w2(32'hb8daf3a1),
	.w3(32'hb64ce45c),
	.w4(32'hb7f4f37f),
	.w5(32'h3fbbd00c),
	.w6(32'h3ec447ba),
	.w7(32'h3ea504f3),
	.w8(32'h3f63a9b0),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fa7c3d2),
	.w1(32'hb98f5612),
	.w2(32'h3e8546dd),
	.w3(32'h3d2ab357),
	.w4(32'h39c83049),
	.w5(32'h3ce3d63e),
	.w6(32'h396c4af4),
	.w7(32'h391d23f5),
	.w8(32'h3faeb930),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87fd2ec),
	.w1(32'h3c6dc016),
	.w2(32'h3f997478),
	.w3(32'hb96037e5),
	.w4(32'hba0dba11),
	.w5(32'h3ce9e401),
	.w6(32'h3cce7ce0),
	.w7(32'h3dc3d3b1),
	.w8(32'h3d887481),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1d915a),
	.w1(32'h3f50fb72),
	.w2(32'h3a494e1b),
	.w3(32'h38ecbf5a),
	.w4(32'h3c046b4b),
	.w5(32'h3dd63f63),
	.w6(32'h3e9fe897),
	.w7(32'hb962031d),
	.w8(32'h3f158b7b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfae13),
	.w1(32'h3eec9443),
	.w2(32'h3c06e00c),
	.w3(32'h3ec01b7d),
	.w4(32'hba3c08d9),
	.w5(32'hba7bae12),
	.w6(32'h3df5e509),
	.w7(32'h3cb840ba),
	.w8(32'h3dacd10f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bdc66),
	.w1(32'hb9c6f036),
	.w2(32'h3d47b33e),
	.w3(32'h3e114045),
	.w4(32'h3d146ee7),
	.w5(32'h3ea2ef94),
	.w6(32'h3f055622),
	.w7(32'hba022b22),
	.w8(32'h3f195c66),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6405e5a),
	.w1(32'h36484d43),
	.w2(32'h3c83a812),
	.w3(32'h3d97a317),
	.w4(32'hb480a146),
	.w5(32'h3e5a2ca6),
	.w6(32'h3763ce0a),
	.w7(32'h3f1fbce2),
	.w8(32'h38135f9d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f5cb8af),
	.w1(32'hb9df826a),
	.w2(32'h3da58f39),
	.w3(32'hb7c86238),
	.w4(32'h3f0fff3d),
	.w5(32'h3d922cd3),
	.w6(32'h39d0ba6a),
	.w7(32'h3f30ef48),
	.w8(32'h3d7c89e3),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75361ad),
	.w1(32'h3e952ec9),
	.w2(32'hb7a84681),
	.w3(32'h3f238b4e),
	.w4(32'h3fcc2090),
	.w5(32'h3e60fc43),
	.w6(32'h37da193c),
	.w7(32'h3f1fa24c),
	.w8(32'h3c4e3803),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd4f0db),
	.w1(32'hb906ff6f),
	.w2(32'h3f559bbb),
	.w3(32'hb997a594),
	.w4(32'hb9902dfa),
	.w5(32'hb94e5fad),
	.w6(32'h3e312619),
	.w7(32'h3d55f912),
	.w8(32'hb88ac576),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3eeffe9e),
	.w1(32'h3e8ee382),
	.w2(32'h3eed1c5c),
	.w3(32'hb7427c03),
	.w4(32'h383e93a2),
	.w5(32'h3ee97918),
	.w6(32'h3e5a740c),
	.w7(32'h3e869a20),
	.w8(32'hb9197515),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962b982),
	.w1(32'hb921cb84),
	.w2(32'h3d002c2d),
	.w3(32'h393546eb),
	.w4(32'h3ee0a830),
	.w5(32'hba589ab4),
	.w6(32'h3f247b84),
	.w7(32'hb9121274),
	.w8(32'h3d252ff1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6c2639),
	.w1(32'h3bff3275),
	.w2(32'h3ec4aed8),
	.w3(32'hb79943de),
	.w4(32'h3f8e2c2a),
	.w5(32'h3d72f8d4),
	.w6(32'h3d4d2274),
	.w7(32'h36f099e7),
	.w8(32'hb687887d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb549c3e5),
	.w1(32'h3ed5489a),
	.w2(32'h3eed79bb),
	.w3(32'h3f11dec9),
	.w4(32'h3e86c70b),
	.w5(32'h3645706b),
	.w6(32'h35d32515),
	.w7(32'h3e84cac6),
	.w8(32'h372b36f6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ec5cffa),
	.w1(32'h3e88eaba),
	.w2(32'h3fad2e91),
	.w3(32'h3969400d),
	.w4(32'h388993be),
	.w5(32'h3c95edd5),
	.w6(32'hb8e8cf2d),
	.w7(32'h3f2ae413),
	.w8(32'h3f0ad479),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ec6ef33),
	.w1(32'h3ef680e8),
	.w2(32'h3f3ece08),
	.w3(32'h3f396529),
	.w4(32'h3f163665),
	.w5(32'hba0ba707),
	.w6(32'h3fa74504),
	.w7(32'h3bd873a6),
	.w8(32'hb91ed991),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2c8199),
	.w1(32'hb9477c08),
	.w2(32'h3c3f0157),
	.w3(32'h3d1ca8a6),
	.w4(32'hb9d9440a),
	.w5(32'h3f4979f1),
	.w6(32'h3a7a0436),
	.w7(32'h3a84fe35),
	.w8(32'h391850e5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e2ed0f5),
	.w1(32'h3d8eec4f),
	.w2(32'hb45e75fd),
	.w3(32'h3d73f1b7),
	.w4(32'h3b74c598),
	.w5(32'h3c63b30c),
	.w6(32'h3e4f0b42),
	.w7(32'h3faa2d98),
	.w8(32'h3d0268e0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f51969f),
	.w1(32'h3d7c862a),
	.w2(32'h3ef15b62),
	.w3(32'hba6c6b00),
	.w4(32'h3f30f98a),
	.w5(32'h3cab3fd8),
	.w6(32'hbabf5f31),
	.w7(32'h3d27e6f7),
	.w8(32'h3ea04b65),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fbd0433),
	.w1(32'h3f0443f9),
	.w2(32'h3d3351a8),
	.w3(32'h3c01a602),
	.w4(32'hba66cb8b),
	.w5(32'hba882da9),
	.w6(32'h3f162eb0),
	.w7(32'h3a24368b),
	.w8(32'h3a3e8124),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ea6fbbd),
	.w1(32'h381c7083),
	.w2(32'h3f80d744),
	.w3(32'hba6b017c),
	.w4(32'h3ea45cee),
	.w5(32'h398afe27),
	.w6(32'h3e5b3044),
	.w7(32'h3a24d1e9),
	.w8(32'h3d5913f3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbadc07),
	.w1(32'h3ea41731),
	.w2(32'h387623a6),
	.w3(32'h3f4ceadf),
	.w4(32'h3d80158d),
	.w5(32'h35d151c4),
	.w6(32'h36f2445d),
	.w7(32'h3b5a0c96),
	.w8(32'h3f08ce3c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370e1fed),
	.w1(32'h3f05dc45),
	.w2(32'h3e489009),
	.w3(32'h35c263b0),
	.w4(32'h3e752d12),
	.w5(32'h3d1e2b96),
	.w6(32'h3741551d),
	.w7(32'h3f26f71b),
	.w8(32'h3f72c1fb),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d945a5b),
	.w1(32'hb4e3610d),
	.w2(32'h3de4bc67),
	.w3(32'h3b6d374b),
	.w4(32'h3e7b5122),
	.w5(32'h36b92555),
	.w6(32'h3679237b),
	.w7(32'h3e063d60),
	.w8(32'h3be8d93e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabed083),
	.w1(32'h3f41e015),
	.w2(32'h3f3d0a51),
	.w3(32'h3e5e54a4),
	.w4(32'h3ebf282d),
	.w5(32'h3e6e13f0),
	.w6(32'h3d312dcc),
	.w7(32'h3ddc3721),
	.w8(32'h3e40d335),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e2312d1),
	.w1(32'hb98cc646),
	.w2(32'h3c4131ee),
	.w3(32'h3d6bf970),
	.w4(32'h3e245735),
	.w5(32'h3e200869),
	.w6(32'h3f572ff4),
	.w7(32'h3cefec97),
	.w8(32'h3db6148f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d57fb1c),
	.w1(32'h3f067518),
	.w2(32'h3ea40231),
	.w3(32'h3a4f13a2),
	.w4(32'h3cce3e3b),
	.w5(32'hb9d2a5b6),
	.w6(32'h3e9e7a5b),
	.w7(32'h3f330dd0),
	.w8(32'h3e3caa9b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf425b7),
	.w1(32'h3d779c81),
	.w2(32'h3db9d2b3),
	.w3(32'hb8d7a5ba),
	.w4(32'hb93a03e0),
	.w5(32'h3e469f5d),
	.w6(32'hb9871626),
	.w7(32'h3db345e7),
	.w8(32'hb99e76da),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f6899e2),
	.w1(32'h3cd64a10),
	.w2(32'hbdd9705e),
	.w3(32'hba8a1cd4),
	.w4(32'hbd039a2e),
	.w5(32'h3dfa6ba6),
	.w6(32'h3ddea665),
	.w7(32'hb8740213),
	.w8(32'h394e9972),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e382613),
	.w1(32'h3ce3bd7a),
	.w2(32'h38359d9e),
	.w3(32'hba46dfae),
	.w4(32'h3edfc160),
	.w5(32'h38ca89e6),
	.w6(32'hbefc459a),
	.w7(32'h3c122018),
	.w8(32'hb916f6ab),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c72ace),
	.w1(32'hbd544b21),
	.w2(32'h3caf3c86),
	.w3(32'h3d7a8717),
	.w4(32'hb80a5252),
	.w5(32'h3c690829),
	.w6(32'h3d04aea2),
	.w7(32'hb811a6e7),
	.w8(32'hba71ad4e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf45e2),
	.w1(32'h389a04a3),
	.w2(32'h3e0b7743),
	.w3(32'h3cc3e2f9),
	.w4(32'h3cf331c2),
	.w5(32'h3d720aac),
	.w6(32'h3c6b1ea2),
	.w7(32'hb8a806c7),
	.w8(32'h3c6cff70),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386eecec),
	.w1(32'h3d8238cf),
	.w2(32'h3b9ae001),
	.w3(32'h34776fc2),
	.w4(32'h3be05cf0),
	.w5(32'h3b9724b9),
	.w6(32'h3d196111),
	.w7(32'hbe19e718),
	.w8(32'hb91586e2),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2897e6),
	.w1(32'hba1754d3),
	.w2(32'hbd9545a8),
	.w3(32'hbc4e52d7),
	.w4(32'h3997a52b),
	.w5(32'h390ebb8b),
	.w6(32'hb9ed72c2),
	.w7(32'hbcacdefc),
	.w8(32'hbafcd4ca),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d213b),
	.w1(32'h3d3af3c3),
	.w2(32'h391e9f94),
	.w3(32'h3c0c6a34),
	.w4(32'h39a0f348),
	.w5(32'hb922d365),
	.w6(32'h3d847758),
	.w7(32'h3b604977),
	.w8(32'hb68df45e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4bc892),
	.w1(32'h3a237982),
	.w2(32'hb9cf45e2),
	.w3(32'h3c5d3fb0),
	.w4(32'h3d1c3b38),
	.w5(32'hb95dcc58),
	.w6(32'hbbce2f2f),
	.w7(32'hb9905dc3),
	.w8(32'hbec2ab03),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d068580),
	.w1(32'h3d318616),
	.w2(32'hba368d61),
	.w3(32'hbcc8c24c),
	.w4(32'hba06f960),
	.w5(32'hbc91917b),
	.w6(32'hbca98d2f),
	.w7(32'hbd7e9b21),
	.w8(32'h3da9725b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe3be0e1),
	.w1(32'h3c99c863),
	.w2(32'h3caca92a),
	.w3(32'h3a4f141d),
	.w4(32'h3c92bd75),
	.w5(32'hb9e02378),
	.w6(32'hb96cbb16),
	.w7(32'hb954bcbd),
	.w8(32'hb9bb6b6a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e62d7),
	.w1(32'hb98937c9),
	.w2(32'h3ccaad63),
	.w3(32'hbd30fb11),
	.w4(32'h3eabc19f),
	.w5(32'h3df0f05b),
	.w6(32'hb9a51d48),
	.w7(32'hb781a86c),
	.w8(32'hb87ec395),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdcf7127),
	.w1(32'hb999a79d),
	.w2(32'hbe91092c),
	.w3(32'h3dd9d7b8),
	.w4(32'h385d4ed5),
	.w5(32'h391a63c5),
	.w6(32'hbc5ee048),
	.w7(32'hb9865a7b),
	.w8(32'h3c9737d0),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1bc81),
	.w1(32'hbd2afb87),
	.w2(32'h3b5df02b),
	.w3(32'h3c696b4e),
	.w4(32'hb9a594fb),
	.w5(32'h3c21dbbe),
	.w6(32'h3853f958),
	.w7(32'hb9d51b78),
	.w8(32'hbcf01cd1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39045cb1),
	.w1(32'hb7c6bfe4),
	.w2(32'h3867285a),
	.w3(32'h3d267c09),
	.w4(32'h38958dfe),
	.w5(32'hbd2bfbfe),
	.w6(32'h3cc40843),
	.w7(32'hbdeb7329),
	.w8(32'hbc57faff),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd96de07),
	.w1(32'hb9a1bc5c),
	.w2(32'h399ae76f),
	.w3(32'hbd76fe29),
	.w4(32'hbbef4283),
	.w5(32'h3bb5f718),
	.w6(32'hbb2fcb5f),
	.w7(32'hbb032c62),
	.w8(32'hbab55966),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3df1b978),
	.w1(32'hbe8215bf),
	.w2(32'hbdf04867),
	.w3(32'h3e048549),
	.w4(32'hbc84b862),
	.w5(32'h3d9887ba),
	.w6(32'h3d0239dd),
	.w7(32'h3ce971b6),
	.w8(32'h3bc62f86),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c499975),
	.w1(32'hba204622),
	.w2(32'hba6b2a91),
	.w3(32'hbd859d7e),
	.w4(32'h39d33e96),
	.w5(32'hba169f53),
	.w6(32'hb9961034),
	.w7(32'h3d129ec3),
	.w8(32'h3925b5c5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee9045),
	.w1(32'hba796f27),
	.w2(32'h3d195f06),
	.w3(32'h3baecd5c),
	.w4(32'hbda715b8),
	.w5(32'h3d0e71d4),
	.w6(32'hbe832e81),
	.w7(32'h3b86a026),
	.w8(32'h3bf69128),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e66f751),
	.w1(32'h3d046812),
	.w2(32'h37a1eca4),
	.w3(32'hb8313db5),
	.w4(32'hbe83aea1),
	.w5(32'h3d18bd1b),
	.w6(32'h3b745009),
	.w7(32'h38a32e89),
	.w8(32'hbea1d80d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1397a2),
	.w1(32'hbd7e4539),
	.w2(32'hbd2a1903),
	.w3(32'h3d84c388),
	.w4(32'h3c929258),
	.w5(32'h3e05b804),
	.w6(32'h3bd6a113),
	.w7(32'h3a9c4100),
	.w8(32'hb98b189e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba97da2),
	.w1(32'hbac89d66),
	.w2(32'h3e0d05bb),
	.w3(32'h3c256e41),
	.w4(32'hbe091bbc),
	.w5(32'h3b38a20a),
	.w6(32'hbad7e1e7),
	.w7(32'hba77df10),
	.w8(32'h3bad4da1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb4b87),
	.w1(32'h3d17cbde),
	.w2(32'hb89359a6),
	.w3(32'h3dbb4d7d),
	.w4(32'h3c39d8eb),
	.w5(32'hbb88d68d),
	.w6(32'hbadfe41e),
	.w7(32'hbd47d570),
	.w8(32'h3cc7a316),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c240ce0),
	.w1(32'h3e31a4cb),
	.w2(32'hba27dfb0),
	.w3(32'hbac310c9),
	.w4(32'hba83a631),
	.w5(32'hbd83c059),
	.w6(32'hba878dfd),
	.w7(32'h3884014d),
	.w8(32'hbd086e3e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c898f28),
	.w1(32'hbd9bcaa6),
	.w2(32'hba84170a),
	.w3(32'hbd8bb9e7),
	.w4(32'h3b9d698e),
	.w5(32'hb9264b9b),
	.w6(32'h3c1d9774),
	.w7(32'h3b434813),
	.w8(32'h3b56f23e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd085c2f),
	.w1(32'h3c142e63),
	.w2(32'h3d59d1cc),
	.w3(32'h3d036bcb),
	.w4(32'h3a2892cb),
	.w5(32'hb9fb8791),
	.w6(32'h3a22a6ed),
	.w7(32'hbcc4ec20),
	.w8(32'hbed6dfdf),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dbd9da9),
	.w1(32'hbd76170e),
	.w2(32'hbe1322e9),
	.w3(32'h3df9ca82),
	.w4(32'h3dc5a5d8),
	.w5(32'hb80ad51d),
	.w6(32'hbc9255ca),
	.w7(32'h3d54f605),
	.w8(32'hbcff7cad),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c923b12),
	.w1(32'h3c0b17ee),
	.w2(32'hbdab8d03),
	.w3(32'h3b43ec9b),
	.w4(32'h3ab07e32),
	.w5(32'hbe505705),
	.w6(32'h3d825317),
	.w7(32'hb6b647d5),
	.w8(32'h3d02e5bd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbea0792b),
	.w1(32'h3d9c548a),
	.w2(32'hba2bc735),
	.w3(32'hbf54de2d),
	.w4(32'h3c8b04e0),
	.w5(32'hbd1b93d0),
	.w6(32'hb99b2493),
	.w7(32'h3a66aa9f),
	.w8(32'h3903278f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdac2f0),
	.w1(32'hb7a51176),
	.w2(32'h3d1aef90),
	.w3(32'h3d24f98c),
	.w4(32'h3e035964),
	.w5(32'h3987e015),
	.w6(32'hbc96f0ac),
	.w7(32'h380924d7),
	.w8(32'h3c18715d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f94a43),
	.w1(32'h3a08d334),
	.w2(32'h3e850cf8),
	.w3(32'h3ca92427),
	.w4(32'h3c3bd4a0),
	.w5(32'h3d34eaa8),
	.w6(32'h3c829006),
	.w7(32'h39816635),
	.w8(32'h3e476777),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3176a8),
	.w1(32'hb8f4be84),
	.w2(32'h39eccd8d),
	.w3(32'hb9884603),
	.w4(32'h3a568f12),
	.w5(32'h3e77948a),
	.w6(32'hba1a2047),
	.w7(32'h3c11c3cf),
	.w8(32'hba874dce),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de9a41),
	.w1(32'hb99e20f0),
	.w2(32'h3a801028),
	.w3(32'h3909549f),
	.w4(32'h3b55009f),
	.w5(32'h3a50a08f),
	.w6(32'hb7b22430),
	.w7(32'h3e25193f),
	.w8(32'h3a2e80d3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34c0c294),
	.w1(32'h39ae4188),
	.w2(32'h3b6c3366),
	.w3(32'h3bb3f1dc),
	.w4(32'hb62d64b2),
	.w5(32'h3d8f2eb2),
	.w6(32'h3d9d66aa),
	.w7(32'hb5c85020),
	.w8(32'h3994bc08),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c622a0e),
	.w1(32'hbac73625),
	.w2(32'hba0f1930),
	.w3(32'h3b3dafb4),
	.w4(32'h3a0c7759),
	.w5(32'h3b5806bb),
	.w6(32'h3cd6ef14),
	.w7(32'hb5f70fc8),
	.w8(32'hba5f0ea8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86d9b9),
	.w1(32'h3a226568),
	.w2(32'h3c581066),
	.w3(32'h3c9fb54e),
	.w4(32'h392cf023),
	.w5(32'h3c9e4703),
	.w6(32'hb9ecb9b1),
	.w7(32'h3a891cae),
	.w8(32'h393d0600),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29564b),
	.w1(32'h3715e36b),
	.w2(32'h3c383f05),
	.w3(32'h342b00c2),
	.w4(32'h3daed730),
	.w5(32'h3648789d),
	.w6(32'hb4ff147c),
	.w7(32'h39fd8824),
	.w8(32'h3d8a158f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba885fa1),
	.w1(32'h3d22d613),
	.w2(32'h3b064f3c),
	.w3(32'hba9d3cb3),
	.w4(32'h3c77d55c),
	.w5(32'h3af4df8a),
	.w6(32'hba814ef8),
	.w7(32'h3b08bae7),
	.w8(32'h39058be8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0a1f5),
	.w1(32'h3e671dae),
	.w2(32'h3bf6b3cd),
	.w3(32'h349157cd),
	.w4(32'h3e3a516d),
	.w5(32'h3a25d099),
	.w6(32'h3c19a05b),
	.w7(32'hb3f736d3),
	.w8(32'h3a7ca48f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc5088),
	.w1(32'hb8b28b17),
	.w2(32'h36d118b3),
	.w3(32'h3d25f85d),
	.w4(32'h3a20a6f0),
	.w5(32'hb848ec7e),
	.w6(32'hb84ddb2c),
	.w7(32'h3e7e0fad),
	.w8(32'h3e181b73),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35578325),
	.w1(32'h33f0ff69),
	.w2(32'h3c302533),
	.w3(32'h3beae005),
	.w4(32'h3cb507e5),
	.w5(32'hb79e4012),
	.w6(32'h3ca119e7),
	.w7(32'h3d110f52),
	.w8(32'h374721bc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e29423),
	.w1(32'h3c65bf11),
	.w2(32'hb6e9647f),
	.w3(32'h3e08fccc),
	.w4(32'hb6278ba3),
	.w5(32'h3aa86404),
	.w6(32'hb6636a3a),
	.w7(32'h3ab72129),
	.w8(32'h3aa3b81d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb1b42),
	.w1(32'h3e05a545),
	.w2(32'h3a90d50c),
	.w3(32'h3b156516),
	.w4(32'h36eb6ae4),
	.w5(32'hb7d5d9af),
	.w6(32'h39c305bd),
	.w7(32'h3e3e7721),
	.w8(32'hb8e59004),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d186e49),
	.w1(32'h3c0ad6a6),
	.w2(32'h3a9ae7c1),
	.w3(32'hba73862b),
	.w4(32'h3bce0421),
	.w5(32'hb9c3dd92),
	.w6(32'h3d16220f),
	.w7(32'h3ce3c209),
	.w8(32'h3ca81d63),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba516142),
	.w1(32'hb9cd2167),
	.w2(32'h39f87c97),
	.w3(32'hba4990a1),
	.w4(32'h3c93fae8),
	.w5(32'h3cf143c6),
	.w6(32'h3bd2c81c),
	.w7(32'h3e087989),
	.w8(32'h3d0ac4dd),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d06a42b),
	.w1(32'h3cc95a9b),
	.w2(32'h3a132dfd),
	.w3(32'h3e6cf132),
	.w4(32'h37f6a62d),
	.w5(32'h398682dd),
	.w6(32'h3bfcd840),
	.w7(32'h3d992706),
	.w8(32'h3aff9bad),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81570c),
	.w1(32'h35031b16),
	.w2(32'h3e2cb393),
	.w3(32'h365a5077),
	.w4(32'h36603582),
	.w5(32'hb69d9a8c),
	.w6(32'h36823183),
	.w7(32'h39932c12),
	.w8(32'h3c428711),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcc38b),
	.w1(32'h39a5ee63),
	.w2(32'h3979180a),
	.w3(32'h3c02622e),
	.w4(32'h3e6629a0),
	.w5(32'h3a9a0d8a),
	.w6(32'h3b73cda5),
	.w7(32'hb802c27b),
	.w8(32'h3e389f19),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35549930),
	.w1(32'h3e14fe6d),
	.w2(32'h39f16cca),
	.w3(32'hb59882a2),
	.w4(32'h3b0b6d88),
	.w5(32'h3c1b0fce),
	.w6(32'h3b3a97c9),
	.w7(32'h3cbfaa76),
	.w8(32'h3e36720d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913eecc),
	.w1(32'h354da32e),
	.w2(32'h35f93387),
	.w3(32'h3d641384),
	.w4(32'hb4f0dd48),
	.w5(32'h3534afb1),
	.w6(32'h3ddacb57),
	.w7(32'h3b077e30),
	.w8(32'h3da24cca),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85b1dfd),
	.w1(32'h3c6cf631),
	.w2(32'hb9840b13),
	.w3(32'h3bffe606),
	.w4(32'h37e79d33),
	.w5(32'h39b9e56f),
	.w6(32'h38aca0e8),
	.w7(32'h3e185277),
	.w8(32'h39595c7f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ddd2e00),
	.w1(32'h3afcc325),
	.w2(32'h3641a974),
	.w3(32'hb6906997),
	.w4(32'h389b8eff),
	.w5(32'h3d903fab),
	.w6(32'h3c66689d),
	.w7(32'h3593eff3),
	.w8(32'h363dec06),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364d603a),
	.w1(32'h3cd1f7a8),
	.w2(32'h3b0e1489),
	.w3(32'h36a9f5d6),
	.w4(32'h3c6d3ab6),
	.w5(32'h3d73d576),
	.w6(32'h3d2a06e1),
	.w7(32'h3d190d16),
	.w8(32'h3a3011ce),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc5c4f),
	.w1(32'h3bec822f),
	.w2(32'hb95b97bb),
	.w3(32'h39cd45c4),
	.w4(32'h3c0054e4),
	.w5(32'h38a13bff),
	.w6(32'h3929f40d),
	.w7(32'h3b37d69e),
	.w8(32'h392d6c8d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31f62f),
	.w1(32'h3d872cbd),
	.w2(32'h3bed6965),
	.w3(32'h3a5e2b8f),
	.w4(32'h3b21f3ab),
	.w5(32'h3c0eaa78),
	.w6(32'h3db290f7),
	.w7(32'h3d3437b1),
	.w8(32'h3b520337),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cf0d7),
	.w1(32'h3bd97bb2),
	.w2(32'h3b8d5123),
	.w3(32'h3d8eabed),
	.w4(32'h3aba3079),
	.w5(32'h3b9be04e),
	.w6(32'hb9841339),
	.w7(32'h398fcebb),
	.w8(32'h3a8006b4),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382650a7),
	.w1(32'h3a2a726a),
	.w2(32'h3836a67f),
	.w3(32'h3bda176d),
	.w4(32'h3d5d072d),
	.w5(32'h3bff7e1b),
	.w6(32'h3c4510c6),
	.w7(32'h3d50aba4),
	.w8(32'h3933187b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39857562),
	.w1(32'h3a8aad2f),
	.w2(32'h3c455f4a),
	.w3(32'h3a598961),
	.w4(32'h3b7cbf99),
	.w5(32'hb9a8dd5e),
	.w6(32'h3b40a370),
	.w7(32'h3b0d139b),
	.w8(32'h3dedf038),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374cbf6b),
	.w1(32'hb8ad082f),
	.w2(32'hb5ea750a),
	.w3(32'h3b2ff09b),
	.w4(32'h391675e2),
	.w5(32'hb632e42a),
	.w6(32'hb84211bb),
	.w7(32'h38103a04),
	.w8(32'h397d381a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba921be4),
	.w1(32'hb8f6ccce),
	.w2(32'hb9745750),
	.w3(32'hb98fda9d),
	.w4(32'h39932ae6),
	.w5(32'h3982daf2),
	.w6(32'hba917ad1),
	.w7(32'hbab335e4),
	.w8(32'hba59f4a0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule