module layer_8_featuremap_53(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b796c8d),
	.w1(32'hbb8baacd),
	.w2(32'h3b0bcf15),
	.w3(32'h3b840ab0),
	.w4(32'hbb6ea5c5),
	.w5(32'hbb3a3a07),
	.w6(32'hbaea265e),
	.w7(32'h3b01633e),
	.w8(32'h3a0eb4b1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ee5cf),
	.w1(32'h3a856e31),
	.w2(32'h3b814ae4),
	.w3(32'hb9c9c9b8),
	.w4(32'h3b95c0f8),
	.w5(32'hba123ba0),
	.w6(32'hbc14eed1),
	.w7(32'h3a339b02),
	.w8(32'hbb7af9e4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ef760),
	.w1(32'h3ac70989),
	.w2(32'h3bebc0e2),
	.w3(32'hbb6855ed),
	.w4(32'hba9b0fc8),
	.w5(32'hba671d4f),
	.w6(32'hbc3fd2f2),
	.w7(32'hbbab3b7f),
	.w8(32'h3c265d19),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d129f),
	.w1(32'h3c005ba6),
	.w2(32'hbb4bcc59),
	.w3(32'hbb7312c5),
	.w4(32'hba96546f),
	.w5(32'hbbe6d6c2),
	.w6(32'h3b278112),
	.w7(32'h3b49e739),
	.w8(32'hba841ea9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1144d8),
	.w1(32'hbaae8c69),
	.w2(32'hb9ff85fe),
	.w3(32'hbc56f975),
	.w4(32'hbc1d0244),
	.w5(32'hbc376de5),
	.w6(32'h3b22724e),
	.w7(32'h3c15fb1a),
	.w8(32'hbd3c6d6f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3864088b),
	.w1(32'h3c14ecaf),
	.w2(32'hbc297bbc),
	.w3(32'h3cf4ee0b),
	.w4(32'h3d883cfc),
	.w5(32'h3cb3fc50),
	.w6(32'hbd7a8d6d),
	.w7(32'hbd11b0d4),
	.w8(32'hbc0d4718),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0a4af),
	.w1(32'hbabc4fc2),
	.w2(32'hbaa8594d),
	.w3(32'hbb878b3b),
	.w4(32'hbb079786),
	.w5(32'hbbc932ea),
	.w6(32'hbb19382b),
	.w7(32'h3b0a48d7),
	.w8(32'h3bb30f21),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63d5fb),
	.w1(32'hbc01ef18),
	.w2(32'h3aff1312),
	.w3(32'hbcc92c51),
	.w4(32'hbcf0df5c),
	.w5(32'hbc809f2c),
	.w6(32'hbbfdffb6),
	.w7(32'hbb97c60e),
	.w8(32'hbc1fb5c5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb081bc6),
	.w1(32'hbb4750b5),
	.w2(32'hb99e0095),
	.w3(32'hbbccfe26),
	.w4(32'hbb9c988f),
	.w5(32'hbc0b8cb7),
	.w6(32'hbc24a97e),
	.w7(32'h3acd615b),
	.w8(32'hbc80cedd),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca84156),
	.w1(32'hbc5d46f9),
	.w2(32'hbc013a76),
	.w3(32'h3bb5ce5b),
	.w4(32'hbb6f9c56),
	.w5(32'hbca0bbad),
	.w6(32'h3c3d0cc9),
	.w7(32'h3b8a81fb),
	.w8(32'h3bb160c7),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39112277),
	.w1(32'hbbe23bf4),
	.w2(32'hbb7008d7),
	.w3(32'hbc6c1e8e),
	.w4(32'hbce7d1b0),
	.w5(32'hbc96d0f9),
	.w6(32'h3b160501),
	.w7(32'h395920f9),
	.w8(32'hbc3038a8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92f016),
	.w1(32'hbc32d694),
	.w2(32'hbc23034c),
	.w3(32'hba9d9e9d),
	.w4(32'hbb89fa49),
	.w5(32'hbc4c7156),
	.w6(32'hba1b775b),
	.w7(32'h3b72381a),
	.w8(32'hba82da07),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd36e86),
	.w1(32'hbbd7ceb7),
	.w2(32'hbbbe3135),
	.w3(32'hbbfcb928),
	.w4(32'hbac76171),
	.w5(32'hbb8fb4da),
	.w6(32'hbbf8cbe9),
	.w7(32'hba109ee7),
	.w8(32'hbd617a4e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a0709),
	.w1(32'h3a2b2cf3),
	.w2(32'hbbc0f667),
	.w3(32'h3d1535db),
	.w4(32'h3d918bdc),
	.w5(32'h3d035c40),
	.w6(32'hbd8ccafe),
	.w7(32'hbd19d738),
	.w8(32'hbc9647a5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5afa14),
	.w1(32'hbb35e696),
	.w2(32'hbb7c7dbe),
	.w3(32'h3c73e782),
	.w4(32'h3cff9f55),
	.w5(32'h3c2ae40b),
	.w6(32'hbd1e89d9),
	.w7(32'hbc912530),
	.w8(32'hbb7d2a2e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb572ab0),
	.w1(32'hba4cf399),
	.w2(32'h38ca6894),
	.w3(32'hbad25c2c),
	.w4(32'h3b6c2d9d),
	.w5(32'h394e1662),
	.w6(32'hbbf74bea),
	.w7(32'h3a0668e3),
	.w8(32'hbb69672b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13bb6d),
	.w1(32'h3ad87928),
	.w2(32'hbcba5ea7),
	.w3(32'h3c45ca95),
	.w4(32'h3b27a7be),
	.w5(32'hbb53d83d),
	.w6(32'hbb7a5d51),
	.w7(32'hbc30fe15),
	.w8(32'hbb819226),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4780db),
	.w1(32'hbc7c3cf1),
	.w2(32'hbbecaf65),
	.w3(32'hbc2b3acc),
	.w4(32'hbc859795),
	.w5(32'hbc33db32),
	.w6(32'hbabdc30d),
	.w7(32'h39950248),
	.w8(32'h3c37b097),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc922557),
	.w1(32'hbd3ec660),
	.w2(32'hbb674567),
	.w3(32'hbd031138),
	.w4(32'hbda0ac2c),
	.w5(32'hbcd85cd3),
	.w6(32'h3ce1945a),
	.w7(32'h3ca6f1b1),
	.w8(32'hbc7a2181),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfe9f1),
	.w1(32'hbc2fa53d),
	.w2(32'h3b066208),
	.w3(32'h3c2e3d42),
	.w4(32'h3acc11ed),
	.w5(32'h3a5ea9dd),
	.w6(32'h3a66d3e2),
	.w7(32'h3c7e6389),
	.w8(32'h3d0161df),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15545f),
	.w1(32'hbb13b58c),
	.w2(32'hbbb1dd3f),
	.w3(32'hbc93829c),
	.w4(32'hbcf6502c),
	.w5(32'hbce7dbf1),
	.w6(32'h3d56930f),
	.w7(32'h3d1aa50f),
	.w8(32'hbb646538),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f41ca),
	.w1(32'h3c77705f),
	.w2(32'h3c7d01b2),
	.w3(32'hbc188628),
	.w4(32'h3a25ae4a),
	.w5(32'hba8a6cf0),
	.w6(32'h3929790f),
	.w7(32'h3c03b345),
	.w8(32'h3cb9613c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d04a61f),
	.w1(32'h3b730fa0),
	.w2(32'h3c6f7f88),
	.w3(32'h3cc631ae),
	.w4(32'hbd155a99),
	.w5(32'hbb8a7353),
	.w6(32'h3dbc48c0),
	.w7(32'h3cda690e),
	.w8(32'h3c3ce172),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2474d9),
	.w1(32'h3b96e683),
	.w2(32'h3b7211b2),
	.w3(32'h3bb2d03d),
	.w4(32'h3b889776),
	.w5(32'hba517108),
	.w6(32'hbb4777c7),
	.w7(32'h3be09d8a),
	.w8(32'h3c207105),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcb917),
	.w1(32'h3b9f9055),
	.w2(32'hbafec9ae),
	.w3(32'hbc27707f),
	.w4(32'hbd096f89),
	.w5(32'hbca77618),
	.w6(32'h3cd4fc66),
	.w7(32'h3be38205),
	.w8(32'h3c8a67cd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6809f5),
	.w1(32'hbc1ebdca),
	.w2(32'hbbedbca1),
	.w3(32'hbbf99ee2),
	.w4(32'hbd2c18d8),
	.w5(32'hbcac2614),
	.w6(32'h3d87e908),
	.w7(32'h3c861253),
	.w8(32'h3b368770),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd82166),
	.w1(32'h39a83686),
	.w2(32'hba9b8c89),
	.w3(32'hbc27d3e0),
	.w4(32'hbc95b1b0),
	.w5(32'hbb3d5633),
	.w6(32'h3d316765),
	.w7(32'h3c777a88),
	.w8(32'h3ce7d25a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd93c63e),
	.w1(32'hbd89b128),
	.w2(32'hbd825e74),
	.w3(32'hbd42de95),
	.w4(32'hbdeba263),
	.w5(32'hbdc0eba6),
	.w6(32'h3d85c349),
	.w7(32'h3c01a88e),
	.w8(32'hbdbbbfea),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd6a2a),
	.w1(32'hbc9b237f),
	.w2(32'h3c00139f),
	.w3(32'h3c9e01a1),
	.w4(32'hbc557fed),
	.w5(32'hbccd8062),
	.w6(32'hbc3bcb28),
	.w7(32'h3ca01e65),
	.w8(32'hbb3101f7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a606464),
	.w1(32'h3afc69cd),
	.w2(32'h3a2978b4),
	.w3(32'h39b360cc),
	.w4(32'h3b556a76),
	.w5(32'hb9e64e41),
	.w6(32'hbbcc1559),
	.w7(32'hbb18a592),
	.w8(32'hbcaf434f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5ab6bc),
	.w1(32'hbd3a17e6),
	.w2(32'hbd61a26d),
	.w3(32'hbc3186b5),
	.w4(32'h3a8ab3fc),
	.w5(32'hbc5374d9),
	.w6(32'hbc5a77fa),
	.w7(32'hbcacdba1),
	.w8(32'h3d0c13ab),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befb2ac),
	.w1(32'h3c3a7f7b),
	.w2(32'hbbcbb493),
	.w3(32'hbd15f9d0),
	.w4(32'hbd6cfe3b),
	.w5(32'hbd20b561),
	.w6(32'h3d82c78c),
	.w7(32'h3cfa84d4),
	.w8(32'hbac33076),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfc43f5),
	.w1(32'hbcd4db33),
	.w2(32'hbd1ebde4),
	.w3(32'hbc2500b0),
	.w4(32'hbc9a3a1c),
	.w5(32'hbcbd3c4e),
	.w6(32'h3b323112),
	.w7(32'hbb9f1e91),
	.w8(32'hbbdef3d3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05cf3f),
	.w1(32'hbb717369),
	.w2(32'hb982c49b),
	.w3(32'hbc23bd23),
	.w4(32'h3bbb3b04),
	.w5(32'hbb629266),
	.w6(32'h39a4e43c),
	.w7(32'h3a1e7ec9),
	.w8(32'hbd3711c3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e42bf),
	.w1(32'h3bd7b8f0),
	.w2(32'hbb543f32),
	.w3(32'h3d35c711),
	.w4(32'h3d9fd83e),
	.w5(32'h3d1b2c9e),
	.w6(32'hbd637cff),
	.w7(32'hbcc68ad0),
	.w8(32'h3c694f2f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1434a5),
	.w1(32'hbc93e4af),
	.w2(32'hbc2b3e02),
	.w3(32'hbc60c9f9),
	.w4(32'hbc9f457f),
	.w5(32'hbcafb38f),
	.w6(32'hbba7ac61),
	.w7(32'h3b8c3c89),
	.w8(32'h3c4699f9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba559e2),
	.w1(32'hbb39a4b4),
	.w2(32'hbc5e2bd7),
	.w3(32'hbcf7765f),
	.w4(32'hbd3ae62b),
	.w5(32'hbcb771a5),
	.w6(32'h3cd224d6),
	.w7(32'h3b72f606),
	.w8(32'hba459fdc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85fe54),
	.w1(32'h3b9936c8),
	.w2(32'h3b979c02),
	.w3(32'h3a20b490),
	.w4(32'h3b5fa62f),
	.w5(32'h3b222fab),
	.w6(32'hbbbf0bc6),
	.w7(32'h3a5b45ac),
	.w8(32'hbcf548d7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6abd2),
	.w1(32'hbbdf038e),
	.w2(32'hbc0143dd),
	.w3(32'h3c8b3efe),
	.w4(32'h3d459c1d),
	.w5(32'h3c3425e1),
	.w6(32'hbd84de12),
	.w7(32'hbcd22758),
	.w8(32'h3ce997ce),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2b7a5),
	.w1(32'hbb544115),
	.w2(32'hb881d183),
	.w3(32'hbceb040f),
	.w4(32'hbd332363),
	.w5(32'hbca0da1b),
	.w6(32'h3d1c67c1),
	.w7(32'h3c99297a),
	.w8(32'h3c11b1e9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee76af),
	.w1(32'hbbfa2838),
	.w2(32'hbc8254ea),
	.w3(32'hbc540e9a),
	.w4(32'hbcb72ec0),
	.w5(32'hbca9159a),
	.w6(32'h3cc96688),
	.w7(32'h3c4a6e85),
	.w8(32'hbc15d736),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9c4f8),
	.w1(32'hbc4e71dd),
	.w2(32'hba9d81e8),
	.w3(32'hbbda39e4),
	.w4(32'hbc149b15),
	.w5(32'h3ae6e423),
	.w6(32'hbbd04ff4),
	.w7(32'hbb535cb4),
	.w8(32'hbbb75c92),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1af56a),
	.w1(32'hbbf9c288),
	.w2(32'hbbeadf1d),
	.w3(32'h3b70b6cf),
	.w4(32'hbc17f28c),
	.w5(32'hbbbc4bc1),
	.w6(32'hbc2ce304),
	.w7(32'h3bf4a079),
	.w8(32'h3aa75294),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b34fb),
	.w1(32'hbc32c9ce),
	.w2(32'hbb86e737),
	.w3(32'hba83a3df),
	.w4(32'hbc159f32),
	.w5(32'hbb35a5b3),
	.w6(32'hba998453),
	.w7(32'hbad8a22d),
	.w8(32'hba0fa5f2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92be47),
	.w1(32'hbc8d4729),
	.w2(32'hbbc05993),
	.w3(32'hbbe54650),
	.w4(32'hbccb95f7),
	.w5(32'hbc418beb),
	.w6(32'h3bf03e80),
	.w7(32'hbb64f8db),
	.w8(32'hbc3ddd7f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc08bea),
	.w1(32'hbca83670),
	.w2(32'hbb81cdc4),
	.w3(32'hbc8645f1),
	.w4(32'hbca5c85e),
	.w5(32'hbb349bd5),
	.w6(32'hbc1b665d),
	.w7(32'hbb7ff300),
	.w8(32'hbbb55f35),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc808f23),
	.w1(32'hbc6683fc),
	.w2(32'h3c393366),
	.w3(32'h3bbe438a),
	.w4(32'h3bc552a1),
	.w5(32'h3a9b6dd2),
	.w6(32'hbc51a151),
	.w7(32'h3a8bacca),
	.w8(32'hbc24b155),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08b72a),
	.w1(32'hbba27e62),
	.w2(32'hbc2f1d46),
	.w3(32'h3b0c9025),
	.w4(32'hbca5068e),
	.w5(32'hbc42ef71),
	.w6(32'h3c66d29a),
	.w7(32'h3a1337c9),
	.w8(32'hbca47f29),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d35bf),
	.w1(32'hbbc6526d),
	.w2(32'hbc308d85),
	.w3(32'hbca106da),
	.w4(32'hbc8118d2),
	.w5(32'hbc985093),
	.w6(32'hbc72d0c8),
	.w7(32'hbc69c144),
	.w8(32'hbb9455e5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95d23f),
	.w1(32'hbc2815ca),
	.w2(32'hbbca46f4),
	.w3(32'hbc2f622a),
	.w4(32'hbc7a3fc8),
	.w5(32'hbc065beb),
	.w6(32'h3b49c829),
	.w7(32'h3ab1a634),
	.w8(32'hba98b2a0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c651f9a),
	.w1(32'h3c5c12fb),
	.w2(32'h3be32457),
	.w3(32'h3c1dcda3),
	.w4(32'h3c6a58df),
	.w5(32'h3c1c6d16),
	.w6(32'h3c5a4226),
	.w7(32'h3c8adb97),
	.w8(32'h3c659a22),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc5ba9),
	.w1(32'h3c0f1572),
	.w2(32'h3c698340),
	.w3(32'hbba49f36),
	.w4(32'hbd0da05f),
	.w5(32'hbb15f582),
	.w6(32'h3c87d8ab),
	.w7(32'hbc8e2bdd),
	.w8(32'hbca5558b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc534511),
	.w1(32'hbc95dbfe),
	.w2(32'h3cb088c6),
	.w3(32'hbc453864),
	.w4(32'hbd11c9eb),
	.w5(32'hbc5e05a8),
	.w6(32'hbc2c05b1),
	.w7(32'h3c24711d),
	.w8(32'hbb95c1f9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3c959),
	.w1(32'hbcd935b2),
	.w2(32'hbc927d3d),
	.w3(32'hbc36feea),
	.w4(32'hbc7a6eee),
	.w5(32'hbc622e37),
	.w6(32'hbc57b10d),
	.w7(32'hbbdba269),
	.w8(32'hbc358f85),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49345d),
	.w1(32'hbb2e2676),
	.w2(32'h3c18e6f9),
	.w3(32'hbbb1bf2e),
	.w4(32'hbc86dd29),
	.w5(32'h38ddf7b1),
	.w6(32'hbc319afd),
	.w7(32'h3bb67f5f),
	.w8(32'hbab3b583),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfb15ee),
	.w1(32'hbd5fc352),
	.w2(32'hbc912c05),
	.w3(32'h3c3a9771),
	.w4(32'hbcaefb47),
	.w5(32'hbc8c046d),
	.w6(32'hbb45b479),
	.w7(32'hba9fd803),
	.w8(32'hbbdec180),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a995664),
	.w1(32'hbc40a0e8),
	.w2(32'h3a9f704d),
	.w3(32'h398cda52),
	.w4(32'h3a963e39),
	.w5(32'h3bead7d5),
	.w6(32'h3c6cac72),
	.w7(32'hba938612),
	.w8(32'hbb9ce581),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5ecb9),
	.w1(32'hbada4284),
	.w2(32'h3c2ee71d),
	.w3(32'hbc9003ad),
	.w4(32'hbd0b9b99),
	.w5(32'hbc1c9635),
	.w6(32'hbc6924dd),
	.w7(32'h3b1a0ba6),
	.w8(32'hbca02438),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3840fa),
	.w1(32'h3aac2722),
	.w2(32'hbc0f94a2),
	.w3(32'hbbfa9b3e),
	.w4(32'hbc5d41af),
	.w5(32'hbc995841),
	.w6(32'hba56e820),
	.w7(32'hbc992f44),
	.w8(32'hbc3e3c87),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc193933),
	.w1(32'hbcbe34f7),
	.w2(32'hbbe37c14),
	.w3(32'h395d1ecf),
	.w4(32'hbbf44c7c),
	.w5(32'hbbd2af9d),
	.w6(32'hbc731cb3),
	.w7(32'hb9fc4a17),
	.w8(32'h3a538899),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e08a0),
	.w1(32'hbc39e1b5),
	.w2(32'h3b833ffa),
	.w3(32'hb9491e6f),
	.w4(32'hbc172cfc),
	.w5(32'h3c37e40c),
	.w6(32'h3c4441c3),
	.w7(32'h3c3c28d0),
	.w8(32'hbc60e70b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bdd2c),
	.w1(32'hbc434c45),
	.w2(32'hbbcfd838),
	.w3(32'hbc2ce8f9),
	.w4(32'hbc73ad19),
	.w5(32'hbb9c6d34),
	.w6(32'hbc132f80),
	.w7(32'hbc17c6ed),
	.w8(32'h3b797954),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b652d),
	.w1(32'hbc85f67e),
	.w2(32'hbc8a864f),
	.w3(32'hbc28dc45),
	.w4(32'hbca6065b),
	.w5(32'hbca5ea61),
	.w6(32'h3c3e64c8),
	.w7(32'h3b7a153e),
	.w8(32'hbcb556af),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11da7d),
	.w1(32'hbc07296b),
	.w2(32'hbc2b4c0b),
	.w3(32'h3c4256f0),
	.w4(32'h3a333db0),
	.w5(32'hbbdf9ac3),
	.w6(32'hbc54c4b9),
	.w7(32'hbac8dd7a),
	.w8(32'hbb649d83),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab626db),
	.w1(32'hbb9c3414),
	.w2(32'hba6dd54b),
	.w3(32'hba68926b),
	.w4(32'hbb6c5a97),
	.w5(32'hb9798926),
	.w6(32'hbb16cb5e),
	.w7(32'hba829177),
	.w8(32'h3a7ba428),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21177b),
	.w1(32'hbbbb84a4),
	.w2(32'h3ae17a73),
	.w3(32'hba948839),
	.w4(32'hbbbd2b2f),
	.w5(32'hbb0e71b1),
	.w6(32'h3b6c3eaa),
	.w7(32'h3b5d2901),
	.w8(32'h39d0bd18),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cd172),
	.w1(32'h3ac8985d),
	.w2(32'hbb430698),
	.w3(32'h3b693963),
	.w4(32'h3a4083cf),
	.w5(32'hbb4fc61f),
	.w6(32'h3b14c6d4),
	.w7(32'hba3f43f6),
	.w8(32'hbc9ddb57),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac2c30),
	.w1(32'hbc20a94c),
	.w2(32'hbbfe6e8b),
	.w3(32'h3b226280),
	.w4(32'hbbdc825d),
	.w5(32'hbb2b1e0a),
	.w6(32'hb805320d),
	.w7(32'h3c023eb4),
	.w8(32'h3b15e02c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57e6f3),
	.w1(32'hbb9a40c7),
	.w2(32'hbaf0f336),
	.w3(32'hbb1577a2),
	.w4(32'hbb546b9a),
	.w5(32'hba968775),
	.w6(32'h396a014f),
	.w7(32'h3a6024fd),
	.w8(32'hba96a111),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d110e67),
	.w1(32'h3c51c31e),
	.w2(32'hbb5178f5),
	.w3(32'h3b03e128),
	.w4(32'hbcb5f365),
	.w5(32'hbce2fa09),
	.w6(32'h3c1d3402),
	.w7(32'hbc92b922),
	.w8(32'hbbc68fa9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3e004),
	.w1(32'hbb5f2d96),
	.w2(32'h3b067ec6),
	.w3(32'h3b17ceef),
	.w4(32'h3a839949),
	.w5(32'h3bc564b0),
	.w6(32'h3ace1e98),
	.w7(32'h3b733f82),
	.w8(32'hb9adfa21),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b087fae),
	.w1(32'hbab4dfeb),
	.w2(32'hbb5b7943),
	.w3(32'hbaabc38c),
	.w4(32'hbc07cd24),
	.w5(32'hbc1dbcfa),
	.w6(32'h3b7102fb),
	.w7(32'hba7b8a33),
	.w8(32'h3b86104c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84a480),
	.w1(32'hb993e6f1),
	.w2(32'h3be1dc6c),
	.w3(32'h3bd8ef42),
	.w4(32'h3ba40174),
	.w5(32'h3c332526),
	.w6(32'h3bc9fde6),
	.w7(32'h3c06a4a5),
	.w8(32'hbcb0fe0e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6de19),
	.w1(32'hbd0e0602),
	.w2(32'hbc9919c4),
	.w3(32'h3b0dac83),
	.w4(32'hbc479cc9),
	.w5(32'hbc44946e),
	.w6(32'hbc89b393),
	.w7(32'h3c84a8f4),
	.w8(32'h3c2bf4af),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24ef78),
	.w1(32'h3c2d1f03),
	.w2(32'h3c3ce4e8),
	.w3(32'h3c3be770),
	.w4(32'h3c2eb8c0),
	.w5(32'h3c4c1001),
	.w6(32'h3c4f65fb),
	.w7(32'h3c462dbe),
	.w8(32'h3aa4e6d8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c4a04),
	.w1(32'h3a04932b),
	.w2(32'h3b6ed9c0),
	.w3(32'h3c066875),
	.w4(32'h3b4f8359),
	.w5(32'h3bc13435),
	.w6(32'h3c4a429d),
	.w7(32'h3c00cc2c),
	.w8(32'h3ba34ddb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39685912),
	.w1(32'h39c7827e),
	.w2(32'h3b7361e9),
	.w3(32'h3b483092),
	.w4(32'h3b2174ed),
	.w5(32'h3bc687b9),
	.w6(32'h3b1a279a),
	.w7(32'h3b590553),
	.w8(32'hbbad368d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72158d),
	.w1(32'h3be20839),
	.w2(32'hbbd4cf97),
	.w3(32'hbba2f7e4),
	.w4(32'hbc61f4cc),
	.w5(32'hbc9c8d33),
	.w6(32'h3c5d950e),
	.w7(32'hbc5bd74d),
	.w8(32'hbbaa1789),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe6307),
	.w1(32'hbbb239b7),
	.w2(32'h3a5858cd),
	.w3(32'h3a7d3c63),
	.w4(32'hba1e915e),
	.w5(32'h3b1821c4),
	.w6(32'h3be75662),
	.w7(32'hbb46da77),
	.w8(32'hbb826dd5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc91e08),
	.w1(32'hbc4a42dd),
	.w2(32'hbbf96536),
	.w3(32'hbad9c47c),
	.w4(32'hbb974980),
	.w5(32'hbb034833),
	.w6(32'hbbfec334),
	.w7(32'hbaa15ace),
	.w8(32'hbb53fa8c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9df79f),
	.w1(32'hbc8a7bc6),
	.w2(32'hbb9f17dc),
	.w3(32'hb8a1bfe5),
	.w4(32'hbc64cf33),
	.w5(32'h3b6eca11),
	.w6(32'h3ba2bea8),
	.w7(32'h3c6b6b74),
	.w8(32'h3ac51924),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9a5c0),
	.w1(32'h3a0c9b67),
	.w2(32'h3b16f065),
	.w3(32'h3b823fea),
	.w4(32'hbabcdf58),
	.w5(32'hba033f5f),
	.w6(32'hbb203fa3),
	.w7(32'hbbf9cd10),
	.w8(32'hbc2ce5bd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee7c28),
	.w1(32'hbc39351a),
	.w2(32'hbbdb6933),
	.w3(32'hbbda6fe3),
	.w4(32'hbcc59c94),
	.w5(32'hbc7037be),
	.w6(32'h3c47a791),
	.w7(32'h3b11191a),
	.w8(32'h397f990c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd6525f),
	.w1(32'hbd685610),
	.w2(32'hbcc8ab73),
	.w3(32'hbd19ebf8),
	.w4(32'hbc62e684),
	.w5(32'hbc1786e0),
	.w6(32'hbcb9ab6e),
	.w7(32'hbc58c35e),
	.w8(32'hbc304b11),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6886f0),
	.w1(32'hbc8d618b),
	.w2(32'hbbac8937),
	.w3(32'hbc1c6f55),
	.w4(32'hbd0e2341),
	.w5(32'hbca0f600),
	.w6(32'h3c70c006),
	.w7(32'h3bc1719e),
	.w8(32'h3aa1d72b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcff657),
	.w1(32'hba4c85f9),
	.w2(32'hbb3e8805),
	.w3(32'h3bc30ba6),
	.w4(32'hbc4084f8),
	.w5(32'hbc1f86b6),
	.w6(32'h3c81e2e6),
	.w7(32'hbbec8bb7),
	.w8(32'hbd378cee),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bf13d),
	.w1(32'hbbc4e7e1),
	.w2(32'hbc4f406f),
	.w3(32'hbcc59060),
	.w4(32'hbc9e7bb1),
	.w5(32'hbcaf6ba6),
	.w6(32'hbc90db45),
	.w7(32'hbc944018),
	.w8(32'hbb251f8c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8672b),
	.w1(32'hbbcfe31e),
	.w2(32'hbbbc48db),
	.w3(32'hbbbb7e15),
	.w4(32'hbbe13457),
	.w5(32'hbb806463),
	.w6(32'hb93a7e87),
	.w7(32'hbb25ea39),
	.w8(32'h3c069b35),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd91289),
	.w1(32'hbcdc4abf),
	.w2(32'hbc5f8f46),
	.w3(32'h3b1f262f),
	.w4(32'hbc4c9384),
	.w5(32'hbbe60ac3),
	.w6(32'h39c156da),
	.w7(32'h3c1f9782),
	.w8(32'hbcdd1cd4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ad963),
	.w1(32'hbbf2ad74),
	.w2(32'hbc92120e),
	.w3(32'hbc9b2b14),
	.w4(32'hbcac8383),
	.w5(32'hbce2cb99),
	.w6(32'hbc42c38d),
	.w7(32'hbc94d967),
	.w8(32'hbce94b62),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89f72c),
	.w1(32'hbc32dd16),
	.w2(32'hbc78e71a),
	.w3(32'hbca06b8f),
	.w4(32'hbcac78b1),
	.w5(32'hbcc5504a),
	.w6(32'hbc718deb),
	.w7(32'hbca373d6),
	.w8(32'hbb558bf0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4ecf4),
	.w1(32'hbb1f7424),
	.w2(32'h3af36434),
	.w3(32'h3b603d96),
	.w4(32'h3b203aee),
	.w5(32'h3b6dce80),
	.w6(32'hb9ce1b6b),
	.w7(32'h3c07c5a5),
	.w8(32'h3b53e823),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5869a),
	.w1(32'hba8b7669),
	.w2(32'hbc141a65),
	.w3(32'h3b8380a2),
	.w4(32'hbb71c3f4),
	.w5(32'hbbed9882),
	.w6(32'hbc690df2),
	.w7(32'hbc0bcd99),
	.w8(32'h3b25be78),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa633d5),
	.w1(32'hbb84049c),
	.w2(32'hbb29cc58),
	.w3(32'hb9dae60e),
	.w4(32'hbbcc955e),
	.w5(32'hbbb661a0),
	.w6(32'h3b230009),
	.w7(32'hbaa84ac1),
	.w8(32'hbae414f2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d29e8),
	.w1(32'hbc878d23),
	.w2(32'h3b66edab),
	.w3(32'h3b917f29),
	.w4(32'hbc046eb7),
	.w5(32'hbbad4daa),
	.w6(32'h3c5de68e),
	.w7(32'h3c52a45f),
	.w8(32'hbc14b708),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91fe3a),
	.w1(32'hbd13b8a7),
	.w2(32'hbd0f9be0),
	.w3(32'hbbe14cc6),
	.w4(32'hbccca5fa),
	.w5(32'hbcecdac6),
	.w6(32'hbc2e0832),
	.w7(32'hbc29f196),
	.w8(32'hbc8b9c8d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c915b0c),
	.w1(32'h3b255b19),
	.w2(32'h3c31647e),
	.w3(32'h3aa8a5d4),
	.w4(32'hbc6d283d),
	.w5(32'h3b2c65f7),
	.w6(32'h3bb7d7fe),
	.w7(32'h3b67141f),
	.w8(32'h3a868299),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74de23),
	.w1(32'hbcaf77b7),
	.w2(32'h3c38063d),
	.w3(32'h3c264122),
	.w4(32'h3cc0cbd8),
	.w5(32'h3c644753),
	.w6(32'hbc3b8d26),
	.w7(32'h3bb0137c),
	.w8(32'hbb9643b3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d6055),
	.w1(32'h3c7981f2),
	.w2(32'h3aae8219),
	.w3(32'h3a9031dc),
	.w4(32'h3c16c804),
	.w5(32'hba2c34ba),
	.w6(32'h3bfb6666),
	.w7(32'hbc1a35bd),
	.w8(32'h3a371ecd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcac69c),
	.w1(32'hbc059248),
	.w2(32'hbb08587b),
	.w3(32'hbb2fd5f4),
	.w4(32'hbb7ae04d),
	.w5(32'h3a8711b0),
	.w6(32'hb9abb4fc),
	.w7(32'hb9e95729),
	.w8(32'hbb002189),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8de630),
	.w1(32'hbca4e943),
	.w2(32'hbaffe8fd),
	.w3(32'hbae58fa3),
	.w4(32'hbb8a9480),
	.w5(32'h3b51ebdc),
	.w6(32'hbbff73e4),
	.w7(32'h3c219d76),
	.w8(32'h3a3d1355),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6b06d),
	.w1(32'hba8be9a7),
	.w2(32'hba431e0e),
	.w3(32'h3b5ea56c),
	.w4(32'h3b83b06b),
	.w5(32'h3b816d84),
	.w6(32'hba94f783),
	.w7(32'hbb440a1c),
	.w8(32'h3b2d2b3a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca9ef97),
	.w1(32'h3c97dd65),
	.w2(32'h3c1809d3),
	.w3(32'h3c26193f),
	.w4(32'h3c87b12a),
	.w5(32'h3c3a3444),
	.w6(32'h3cabf706),
	.w7(32'h3c0ee29f),
	.w8(32'h3b2b0447),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5da40),
	.w1(32'hbc08b8e6),
	.w2(32'h3b85966b),
	.w3(32'hbbe2125c),
	.w4(32'hbb842dbd),
	.w5(32'h3c1b2aba),
	.w6(32'hbc38b80a),
	.w7(32'hba495056),
	.w8(32'hbc2d9ccb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd2a43),
	.w1(32'h39b9b7fe),
	.w2(32'hbb09f603),
	.w3(32'hbbab0874),
	.w4(32'hbacc125b),
	.w5(32'hbb5c6cf1),
	.w6(32'hbbf2cb20),
	.w7(32'hbbacd2d7),
	.w8(32'hb8537d55),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a10f8),
	.w1(32'h3b8abed3),
	.w2(32'h3c0b36b7),
	.w3(32'h3ac30f60),
	.w4(32'hbc77f89c),
	.w5(32'hbbaea024),
	.w6(32'h3c06362b),
	.w7(32'hbb580fb9),
	.w8(32'hbba349cc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bbc2f),
	.w1(32'h3b3ca833),
	.w2(32'h3babfcf2),
	.w3(32'h3bb89620),
	.w4(32'hba13f425),
	.w5(32'h3b7a18ac),
	.w6(32'h3bceb572),
	.w7(32'h3b8899fe),
	.w8(32'hbab59fc7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf10e3),
	.w1(32'h3c022ff1),
	.w2(32'h3ba25807),
	.w3(32'h3b9d9269),
	.w4(32'h3bbdd90e),
	.w5(32'h3b560397),
	.w6(32'h3b2e3dfc),
	.w7(32'h3997f82a),
	.w8(32'hbb0c58a8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2276e7),
	.w1(32'h3ac28f38),
	.w2(32'hbb195470),
	.w3(32'hba1c84c6),
	.w4(32'h3b88efb7),
	.w5(32'hb875cf66),
	.w6(32'hbb821f07),
	.w7(32'hbb57a328),
	.w8(32'hbbd3dbe9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65d713),
	.w1(32'h3a67f684),
	.w2(32'h3b612ff8),
	.w3(32'hbb6042b4),
	.w4(32'hbb45d137),
	.w5(32'hba5f9633),
	.w6(32'h3a5a7fd3),
	.w7(32'hbb02a7e1),
	.w8(32'hbab409d1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152238),
	.w1(32'h3bb4bedc),
	.w2(32'h3b870691),
	.w3(32'h3c01fb1e),
	.w4(32'h3c2ddc3e),
	.w5(32'h38c5b490),
	.w6(32'h3b8783a9),
	.w7(32'h3c1b2dfb),
	.w8(32'h3b6219be),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8fae7),
	.w1(32'h39a301f5),
	.w2(32'hbb3f6463),
	.w3(32'hbb8e2c32),
	.w4(32'h3a810d43),
	.w5(32'hb93bd564),
	.w6(32'hbb36464a),
	.w7(32'hbb75b95d),
	.w8(32'hbb4e1bf9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a1be8),
	.w1(32'h3b30d66e),
	.w2(32'h3bf363f4),
	.w3(32'h3b306d53),
	.w4(32'h3bcd5c20),
	.w5(32'h3c1dc74e),
	.w6(32'hbbbd442c),
	.w7(32'hbad486b0),
	.w8(32'hb95c9ca5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5f8f4),
	.w1(32'h3b03896e),
	.w2(32'h39740066),
	.w3(32'hbaf615ba),
	.w4(32'h3a32bfc5),
	.w5(32'hbaa8614c),
	.w6(32'h3a4f12a4),
	.w7(32'hba68b5e9),
	.w8(32'hbac3aaf4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e8b84),
	.w1(32'hb9116683),
	.w2(32'hbb0c4db0),
	.w3(32'hbaacdc05),
	.w4(32'hbaa26a1a),
	.w5(32'hbb2c7daa),
	.w6(32'hb9540de3),
	.w7(32'hbb5b769a),
	.w8(32'hbbbc3dd2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec4635),
	.w1(32'h38d7f179),
	.w2(32'hbafcab65),
	.w3(32'h3aa5f2ab),
	.w4(32'h3b0f4138),
	.w5(32'hbaa93a85),
	.w6(32'h3b676693),
	.w7(32'h3843df79),
	.w8(32'h3956d0ee),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8ba95),
	.w1(32'hba657c9b),
	.w2(32'hbba55a0c),
	.w3(32'h3b229fa5),
	.w4(32'hba2f1381),
	.w5(32'hbb3b8327),
	.w6(32'hbb033bbe),
	.w7(32'hbb9b578e),
	.w8(32'hbba1293a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63416e),
	.w1(32'hbc12a521),
	.w2(32'hbc220b72),
	.w3(32'hbc0d166e),
	.w4(32'hbc7ae241),
	.w5(32'hbc5e23ed),
	.w6(32'hbb87de5d),
	.w7(32'hbbd6a92f),
	.w8(32'hbbe94f08),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26c64f),
	.w1(32'h3b7fad20),
	.w2(32'h3b461716),
	.w3(32'hba0175fc),
	.w4(32'h3b398834),
	.w5(32'h3a4c6452),
	.w6(32'h3b587399),
	.w7(32'h3bac61b5),
	.w8(32'h3b0eb80c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b502111),
	.w1(32'h3a7324a9),
	.w2(32'h3b3b5dde),
	.w3(32'h3b956b66),
	.w4(32'h3b29e06c),
	.w5(32'h3b2b0a4c),
	.w6(32'h3b1d78ab),
	.w7(32'h3b3efc1f),
	.w8(32'h39b2e2e6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc0801),
	.w1(32'hbb8725d1),
	.w2(32'hbb8ad10b),
	.w3(32'h3bef32f1),
	.w4(32'h3a412467),
	.w5(32'hbb766407),
	.w6(32'h398e28b7),
	.w7(32'hbbf14a46),
	.w8(32'hbc109d01),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d618),
	.w1(32'hba7a406a),
	.w2(32'h3a3ddefd),
	.w3(32'hba368cfe),
	.w4(32'h3b40cb59),
	.w5(32'h3c106f9f),
	.w6(32'h3b8f581d),
	.w7(32'h3b8975dc),
	.w8(32'h3b8bbf14),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb175b0e),
	.w1(32'hbb58c4db),
	.w2(32'hbb1d7d9f),
	.w3(32'h3a40dbf1),
	.w4(32'h3a755953),
	.w5(32'h3b66eb89),
	.w6(32'hbb136098),
	.w7(32'h3992a9d7),
	.w8(32'hbb15a775),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39850283),
	.w1(32'h3b42f5b4),
	.w2(32'hba7569b9),
	.w3(32'h3b811444),
	.w4(32'h3bc4fd7e),
	.w5(32'h3a99cd50),
	.w6(32'h398da85c),
	.w7(32'h3a353d84),
	.w8(32'hbb79359f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fbb80),
	.w1(32'h3b1aa28c),
	.w2(32'h3b94f704),
	.w3(32'h3ac7d6ba),
	.w4(32'h3b99ee6b),
	.w5(32'h3b8b3b28),
	.w6(32'h3a71fac5),
	.w7(32'h3b72cfe4),
	.w8(32'hbac1abdc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2991b0),
	.w1(32'hba60ff47),
	.w2(32'hbbb17117),
	.w3(32'hbb8253f8),
	.w4(32'hbb96e109),
	.w5(32'hbc0a2138),
	.w6(32'hbba72681),
	.w7(32'hbbbf5ed6),
	.w8(32'hbb8f4180),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf4cc2),
	.w1(32'h3aa55900),
	.w2(32'h3b94d147),
	.w3(32'h3b980f24),
	.w4(32'h3bafb133),
	.w5(32'h3bbec692),
	.w6(32'h3bbb037f),
	.w7(32'h3be2b13b),
	.w8(32'h3b865658),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c8b86),
	.w1(32'hbb97ed81),
	.w2(32'hbc00bb1a),
	.w3(32'h3a2c966d),
	.w4(32'hbbcae278),
	.w5(32'hbba659e7),
	.w6(32'h39480e22),
	.w7(32'hbbea3b62),
	.w8(32'hbb84b805),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule