module layer_8_featuremap_63(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886db75),
	.w1(32'hb845109d),
	.w2(32'h39ab6d1a),
	.w3(32'hb99f3ebf),
	.w4(32'hb759c6e5),
	.w5(32'h395c80b5),
	.w6(32'h3828880c),
	.w7(32'hb86ec466),
	.w8(32'h391307f7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d00f74),
	.w1(32'h390aed3a),
	.w2(32'h393b716f),
	.w3(32'hb8b2d41c),
	.w4(32'h381be35c),
	.w5(32'h39394a8f),
	.w6(32'h38d5e19a),
	.w7(32'h3802b651),
	.w8(32'h39cf3676),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6851e),
	.w1(32'h38f76bbe),
	.w2(32'h38edf204),
	.w3(32'hb90e303b),
	.w4(32'hb8f281c5),
	.w5(32'h386b18c8),
	.w6(32'h39362cf6),
	.w7(32'h38b53008),
	.w8(32'hba3c73da),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac116d1),
	.w1(32'hbb093f30),
	.w2(32'hbb0b5010),
	.w3(32'h3a8310ce),
	.w4(32'hb98c68cc),
	.w5(32'hba98d3b6),
	.w6(32'h3957338f),
	.w7(32'h38efcd73),
	.w8(32'h39fda859),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00245d),
	.w1(32'h39c0d99c),
	.w2(32'h39c3781d),
	.w3(32'h398bd823),
	.w4(32'h39a6ab3b),
	.w5(32'h39b28149),
	.w6(32'h39b5f4c9),
	.w7(32'h399dd0ca),
	.w8(32'h39cf706e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8edaf1),
	.w1(32'h3a910217),
	.w2(32'h3a92bd08),
	.w3(32'h3a5f6430),
	.w4(32'h3a83cad6),
	.w5(32'h3a0f62d8),
	.w6(32'h3a3a21a5),
	.w7(32'h3a63d48b),
	.w8(32'h3a3a5230),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a141ebc),
	.w1(32'h3a18bc1b),
	.w2(32'h39a5251b),
	.w3(32'hb83e65ee),
	.w4(32'h397b11b2),
	.w5(32'h39a31e62),
	.w6(32'h39c449e0),
	.w7(32'hb791057d),
	.w8(32'h3a0b9f0d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a013027),
	.w1(32'h39da0579),
	.w2(32'h3a15a8de),
	.w3(32'h39bcb10b),
	.w4(32'h39e2e8e6),
	.w5(32'h39e24305),
	.w6(32'h39f3130f),
	.w7(32'h3a193304),
	.w8(32'h3a6599da),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a367cb1),
	.w1(32'h3a4bb133),
	.w2(32'h39f8de84),
	.w3(32'h38ea3318),
	.w4(32'h398f2841),
	.w5(32'h39e5dac4),
	.w6(32'h3a09ec00),
	.w7(32'h3850b9a2),
	.w8(32'hbb788014),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d1adc),
	.w1(32'hba4e8288),
	.w2(32'hbb266a83),
	.w3(32'h39a0e658),
	.w4(32'hba9c1c91),
	.w5(32'hba8e20a4),
	.w6(32'hbb5cfb1d),
	.w7(32'hba5dfcb5),
	.w8(32'h3998e4fb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e5c39c),
	.w1(32'hb9353134),
	.w2(32'hb972c612),
	.w3(32'hb996616b),
	.w4(32'hb9877723),
	.w5(32'hb9c50ef1),
	.w6(32'hb8ea1169),
	.w7(32'h37d2cf5a),
	.w8(32'h3a0446b9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee1c9f),
	.w1(32'h36f78070),
	.w2(32'h3844cfef),
	.w3(32'hb95c034f),
	.w4(32'hb91cd6ad),
	.w5(32'h37b8a0e8),
	.w6(32'h38fbe5a2),
	.w7(32'hb9051698),
	.w8(32'h3a04fc60),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b932a),
	.w1(32'h38d4c50c),
	.w2(32'h3851db2b),
	.w3(32'hb86128b6),
	.w4(32'h3746890f),
	.w5(32'hb816a22a),
	.w6(32'h39aa719f),
	.w7(32'h38cf935e),
	.w8(32'h39e6187a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93ba04),
	.w1(32'h3a9e4bf6),
	.w2(32'h3aa91b13),
	.w3(32'h3a7bd6d5),
	.w4(32'h3a9ad599),
	.w5(32'h3a3b7d47),
	.w6(32'h3a58f6cc),
	.w7(32'h3a84345a),
	.w8(32'h392eea1b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f1f93),
	.w1(32'h3a0c2a04),
	.w2(32'h3a161e7f),
	.w3(32'h3a00f145),
	.w4(32'h3a309a10),
	.w5(32'h39b66b97),
	.w6(32'h398b2363),
	.w7(32'h39c707cc),
	.w8(32'hb84714cc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75f719b),
	.w1(32'hb97dad69),
	.w2(32'hb93746b8),
	.w3(32'hb92293f9),
	.w4(32'h37a6e832),
	.w5(32'h38c78e5b),
	.w6(32'hb89981c6),
	.w7(32'h389b6052),
	.w8(32'h3a6c4004),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba348d88),
	.w1(32'hbae1e558),
	.w2(32'hbb1c359e),
	.w3(32'h39fa9c81),
	.w4(32'hba9d2eab),
	.w5(32'hbb27032b),
	.w6(32'h3aaa7067),
	.w7(32'h3a7514fe),
	.w8(32'h38f706af),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2e39d),
	.w1(32'hba457e6d),
	.w2(32'hba33ddba),
	.w3(32'hba66eadd),
	.w4(32'hba3eb5e8),
	.w5(32'hba2877fe),
	.w6(32'hb9b6eb79),
	.w7(32'hb9f32191),
	.w8(32'hb9410b2f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21d9ea),
	.w1(32'hba458828),
	.w2(32'h3a0d4267),
	.w3(32'hba4d5cdb),
	.w4(32'hb9c6091b),
	.w5(32'h37e82027),
	.w6(32'hb9c9cd24),
	.w7(32'h39b828b3),
	.w8(32'h39877576),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba561e1c),
	.w1(32'hbb60ca1e),
	.w2(32'hbb2176b9),
	.w3(32'hbb1ea176),
	.w4(32'hbb4d9256),
	.w5(32'hba83071e),
	.w6(32'hba972a87),
	.w7(32'hbac655b1),
	.w8(32'hba91032f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad3a7f),
	.w1(32'hbb064e0e),
	.w2(32'hba9ae210),
	.w3(32'hbaae5252),
	.w4(32'hbae6d8c0),
	.w5(32'hba7ef197),
	.w6(32'hbaff274a),
	.w7(32'hbac4165d),
	.w8(32'h3a404758),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41ef5b),
	.w1(32'h39facd09),
	.w2(32'h39da7ad9),
	.w3(32'h3a016df8),
	.w4(32'h3a144963),
	.w5(32'h39d5b48e),
	.w6(32'h39d304f8),
	.w7(32'h398df5c1),
	.w8(32'hb9f32956),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e63be),
	.w1(32'hba905bbb),
	.w2(32'hb9b20136),
	.w3(32'hba9901ec),
	.w4(32'hba88dd4a),
	.w5(32'hb9b0e158),
	.w6(32'hba544ad9),
	.w7(32'hba4de8df),
	.w8(32'h39af63a3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8093793),
	.w1(32'hba0ff28c),
	.w2(32'h39d2d91a),
	.w3(32'hb9c31acc),
	.w4(32'hba37e45a),
	.w5(32'hb8821115),
	.w6(32'hb94d1625),
	.w7(32'h399f7f83),
	.w8(32'hbabee59c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8757ae),
	.w1(32'hba117216),
	.w2(32'hba64e611),
	.w3(32'hba15aeed),
	.w4(32'hbab85615),
	.w5(32'hba81867e),
	.w6(32'hba876746),
	.w7(32'hb9ee3d6d),
	.w8(32'hba020b19),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba602e8f),
	.w1(32'hba7bcd90),
	.w2(32'hb9d9c581),
	.w3(32'hba876658),
	.w4(32'hba86ea14),
	.w5(32'hb9d398a7),
	.w6(32'hba45d890),
	.w7(32'hba442ff2),
	.w8(32'hb9adc1e7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43d20a),
	.w1(32'hba73821e),
	.w2(32'hba03b119),
	.w3(32'hba67ffa2),
	.w4(32'hba825e94),
	.w5(32'hb9f1de28),
	.w6(32'hba2bdec6),
	.w7(32'hba367474),
	.w8(32'hba987a21),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb078637),
	.w1(32'hba9ac438),
	.w2(32'h36969511),
	.w3(32'hbaef58ec),
	.w4(32'hba63abb2),
	.w5(32'h38d3b1e6),
	.w6(32'hbb190597),
	.w7(32'hbac41406),
	.w8(32'h39ed0b48),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5aa14d),
	.w1(32'hba4c9e5f),
	.w2(32'h3a9d37f7),
	.w3(32'hb92bd06a),
	.w4(32'h374dce9e),
	.w5(32'h39f82574),
	.w6(32'h38cc8171),
	.w7(32'h3b22514e),
	.w8(32'h398c342a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68b52ee),
	.w1(32'hb8b0598d),
	.w2(32'hb824c8ca),
	.w3(32'hb87e08af),
	.w4(32'hb8efb275),
	.w5(32'hb8903393),
	.w6(32'h38741d92),
	.w7(32'h374afc6a),
	.w8(32'h3b47be1f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3777ae),
	.w1(32'hbb0c0f50),
	.w2(32'hba5d9f5e),
	.w3(32'h3ab856c5),
	.w4(32'h39bf851f),
	.w5(32'hba8d6adf),
	.w6(32'h3b146aec),
	.w7(32'h3b39cdeb),
	.w8(32'hbadac650),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3a714),
	.w1(32'hbb0d7c39),
	.w2(32'hbaac4c43),
	.w3(32'hbb0889ea),
	.w4(32'hbb19bc3f),
	.w5(32'hba2a05da),
	.w6(32'hbb4d7840),
	.w7(32'hbb1534de),
	.w8(32'h3b04ba38),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad17f2),
	.w1(32'hbab1c96f),
	.w2(32'hbb1cd045),
	.w3(32'h3a13d2a5),
	.w4(32'hba84a9b8),
	.w5(32'hbb57d1b5),
	.w6(32'h3b14a48d),
	.w7(32'h3aa90099),
	.w8(32'h398e6e45),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e0feb),
	.w1(32'hb9dfd061),
	.w2(32'hbae89ddf),
	.w3(32'hb9840995),
	.w4(32'hbae2a577),
	.w5(32'hba4199aa),
	.w6(32'h3b2a5df1),
	.w7(32'h3b019d64),
	.w8(32'h39bcd744),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8558e5),
	.w1(32'h3a8b163e),
	.w2(32'h3a936b3d),
	.w3(32'h3a668382),
	.w4(32'h3a87cac8),
	.w5(32'h3a26a675),
	.w6(32'h3a4804bb),
	.w7(32'h3a72799f),
	.w8(32'hb78c359d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9537625),
	.w1(32'hb9e68f9d),
	.w2(32'h3985a9f2),
	.w3(32'hba4d95ad),
	.w4(32'hb9c09f95),
	.w5(32'h381ea5d9),
	.w6(32'hb9664dab),
	.w7(32'h37d70bf3),
	.w8(32'hbaae8fab),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaede475),
	.w1(32'hbb052259),
	.w2(32'hbabaf24f),
	.w3(32'hbac2ef3e),
	.w4(32'hbb20ae7c),
	.w5(32'hbacef5de),
	.w6(32'hba9d602e),
	.w7(32'hba9aa97f),
	.w8(32'h39356ac8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937cf5a),
	.w1(32'hb9710d1c),
	.w2(32'hb81cf3f3),
	.w3(32'hb9c141bc),
	.w4(32'hb9c9eaff),
	.w5(32'hb8cfcf9b),
	.w6(32'hb8680c97),
	.w7(32'hb8e257d1),
	.w8(32'hb93a9106),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e2ef2),
	.w1(32'h3a106243),
	.w2(32'h3a4903f0),
	.w3(32'h3a3cd3b8),
	.w4(32'h3a8b1c7e),
	.w5(32'h39731670),
	.w6(32'h38899592),
	.w7(32'h39a96805),
	.w8(32'hba750b9f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba847125),
	.w1(32'hba89baeb),
	.w2(32'hba3ce2b3),
	.w3(32'hba98942a),
	.w4(32'hba94ade8),
	.w5(32'hba0e9d51),
	.w6(32'hbab37d6a),
	.w7(32'hba939c85),
	.w8(32'hb95356a1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10ed9e),
	.w1(32'hba37d5e4),
	.w2(32'hb9ca48f8),
	.w3(32'hba3e3d71),
	.w4(32'hba39b55a),
	.w5(32'hb9c0e19e),
	.w6(32'hba173815),
	.w7(32'hba2551db),
	.w8(32'hba46d2f2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb0587),
	.w1(32'hba20c934),
	.w2(32'h3839ce60),
	.w3(32'h3a11f658),
	.w4(32'h3a8b6bfd),
	.w5(32'hb9ae8f9f),
	.w6(32'hb9a7b2fb),
	.w7(32'hb99e6a86),
	.w8(32'hbb66558e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7740cd),
	.w1(32'h3c020cb8),
	.w2(32'h3896c820),
	.w3(32'hbb8a8ce4),
	.w4(32'h3b6c3c23),
	.w5(32'hba9e3d43),
	.w6(32'h3b32a724),
	.w7(32'hbba77a70),
	.w8(32'hb518e88c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba980ff1),
	.w1(32'h37c67adb),
	.w2(32'hb96f5544),
	.w3(32'h3a2fa400),
	.w4(32'h390a2c90),
	.w5(32'hba803bbd),
	.w6(32'hba93020c),
	.w7(32'hbac85f11),
	.w8(32'hb9e30284),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfcd80),
	.w1(32'hb9b33cb2),
	.w2(32'hba7117a0),
	.w3(32'h378d55cf),
	.w4(32'hb7c59a3c),
	.w5(32'hbadaa85c),
	.w6(32'hba135cc2),
	.w7(32'hbaab5fec),
	.w8(32'hbad94251),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a6230),
	.w1(32'h3af8b7f4),
	.w2(32'h3a413192),
	.w3(32'hb9f7db39),
	.w4(32'h3a98dd76),
	.w5(32'h3af35eb3),
	.w6(32'hb9cb68f5),
	.w7(32'hba9b610d),
	.w8(32'hbc326fc8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e825e),
	.w1(32'h3bca6471),
	.w2(32'h3b55b778),
	.w3(32'h3aa72c12),
	.w4(32'hbb8418d9),
	.w5(32'hbae3f062),
	.w6(32'hbb26d447),
	.w7(32'hba329f4b),
	.w8(32'hbadd7995),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67b125),
	.w1(32'h39a5d680),
	.w2(32'h3b535338),
	.w3(32'hba49a535),
	.w4(32'h3ad569b6),
	.w5(32'h3a82b106),
	.w6(32'hbaf65221),
	.w7(32'h3b1958f3),
	.w8(32'hb9fd8243),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04c94c),
	.w1(32'h391d214b),
	.w2(32'h3acfa332),
	.w3(32'hba17a691),
	.w4(32'h39c3355a),
	.w5(32'h3b49644a),
	.w6(32'hba43c765),
	.w7(32'h3b151822),
	.w8(32'hba2df9df),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11b4d9),
	.w1(32'hb7f553da),
	.w2(32'hb9305c9f),
	.w3(32'hba07a840),
	.w4(32'h394b0240),
	.w5(32'hb9cdcf32),
	.w6(32'hb99a2d89),
	.w7(32'hba5a1853),
	.w8(32'h39b6adde),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0657b),
	.w1(32'h392b5f65),
	.w2(32'hb9f42c1c),
	.w3(32'h3a5f5e9a),
	.w4(32'h3a067b3a),
	.w5(32'hb9e7472b),
	.w6(32'h39225839),
	.w7(32'hba1eccad),
	.w8(32'h3a2d2427),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab09e9),
	.w1(32'h39a9e097),
	.w2(32'hba32fd66),
	.w3(32'h3ab86c0a),
	.w4(32'h3a74d8a1),
	.w5(32'hba9dce7a),
	.w6(32'hba077fb8),
	.w7(32'hbaf8c7d8),
	.w8(32'h3bb6958c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a535e15),
	.w1(32'hbba61e69),
	.w2(32'hba9d6426),
	.w3(32'h3b77eb9b),
	.w4(32'hbba41b67),
	.w5(32'hbb5cbf62),
	.w6(32'hbb2da813),
	.w7(32'hbb86f1aa),
	.w8(32'hb935f7d0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e11615),
	.w1(32'h3a08c4b2),
	.w2(32'h3a251af8),
	.w3(32'hba91cc8c),
	.w4(32'h3a74e45e),
	.w5(32'h3b018cee),
	.w6(32'h3a9cf7a9),
	.w7(32'h3ac4f980),
	.w8(32'hbbed562c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cd9623),
	.w1(32'h3bdde248),
	.w2(32'h3c1b8aeb),
	.w3(32'hba16590d),
	.w4(32'h3af71da6),
	.w5(32'h3bbedb06),
	.w6(32'h3b5875cc),
	.w7(32'h3bd01b4a),
	.w8(32'hbb0ed530),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb018941),
	.w1(32'hbb2c5c6d),
	.w2(32'h3a991df7),
	.w3(32'hbae39974),
	.w4(32'h3ae0c2ff),
	.w5(32'h3a4b8bfa),
	.w6(32'hbb0ad71b),
	.w7(32'hbb51d17f),
	.w8(32'h3b03124b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63a191),
	.w1(32'hbb8bea43),
	.w2(32'hba8a45a0),
	.w3(32'hbadc425e),
	.w4(32'hbb6bfcdb),
	.w5(32'h3abfdb48),
	.w6(32'h3a8b0af1),
	.w7(32'hbb056e1f),
	.w8(32'hba7ddb94),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab746d8),
	.w1(32'h3b0b729d),
	.w2(32'h3b2ee0fe),
	.w3(32'hbbb94fbe),
	.w4(32'hb96000e2),
	.w5(32'h3b9bda4f),
	.w6(32'hbba83f65),
	.w7(32'hba24cbcc),
	.w8(32'h3a2b2c2c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a130aa1),
	.w1(32'h39f94268),
	.w2(32'h3ada3d70),
	.w3(32'h3a09ab84),
	.w4(32'hb92f4032),
	.w5(32'h39f056f7),
	.w6(32'hb9c393fd),
	.w7(32'h3a841618),
	.w8(32'h39dd16a7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2675ab),
	.w1(32'hba9a149e),
	.w2(32'hbb32bcf1),
	.w3(32'hbab7e832),
	.w4(32'hbb4bfcdb),
	.w5(32'hbb8dd153),
	.w6(32'hbb392f91),
	.w7(32'hbb0f180e),
	.w8(32'hbb6046a6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c4c2),
	.w1(32'h3c259136),
	.w2(32'h3ab6d22c),
	.w3(32'h3b6372c9),
	.w4(32'h3a977559),
	.w5(32'hbbe83d46),
	.w6(32'hbbb30943),
	.w7(32'h39f42a99),
	.w8(32'hbb32fe5a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2d1ba),
	.w1(32'h3a6cee8f),
	.w2(32'h3a0cd1da),
	.w3(32'hbaef7626),
	.w4(32'h3904601c),
	.w5(32'hba39eb6c),
	.w6(32'h3a2666cd),
	.w7(32'hba6dee84),
	.w8(32'hb795ed8e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93793c),
	.w1(32'h3a202999),
	.w2(32'h3a89ca58),
	.w3(32'hb9cff106),
	.w4(32'h3a3a7bc4),
	.w5(32'h39469405),
	.w6(32'h3abc73ec),
	.w7(32'h3a523c45),
	.w8(32'h39c52ab3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bc89a),
	.w1(32'h3b9e49c5),
	.w2(32'hbad15709),
	.w3(32'hbb8cdf9a),
	.w4(32'hbbbca12a),
	.w5(32'hbb988741),
	.w6(32'hbaa07291),
	.w7(32'hbbd68a38),
	.w8(32'h399abe81),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3344e7),
	.w1(32'hb91ba2cc),
	.w2(32'hba91c3ae),
	.w3(32'h3a5cd888),
	.w4(32'hb8efbc0e),
	.w5(32'hbaae8b6d),
	.w6(32'hb990ad84),
	.w7(32'hba55895d),
	.w8(32'hb888f72b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2152fd),
	.w1(32'hb9901752),
	.w2(32'hb9f8a425),
	.w3(32'h399bd75b),
	.w4(32'hb96b73fb),
	.w5(32'hba59a8c5),
	.w6(32'hba176931),
	.w7(32'hba5a318c),
	.w8(32'h3997677c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9842d75),
	.w1(32'hb990aed8),
	.w2(32'hb9e269b7),
	.w3(32'h3a4e8b6d),
	.w4(32'h3968dce8),
	.w5(32'hba293d2d),
	.w6(32'hb902c745),
	.w7(32'hba1c72f7),
	.w8(32'hba371a5b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99d8b1),
	.w1(32'h3ab03b86),
	.w2(32'h3b09c8d8),
	.w3(32'hbb02ec91),
	.w4(32'hba38d38b),
	.w5(32'h39c21310),
	.w6(32'hbaca2f36),
	.w7(32'hba1f8ca8),
	.w8(32'hba526ae4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf032fa),
	.w1(32'hb93e9fef),
	.w2(32'hba1f8a38),
	.w3(32'hba0199ca),
	.w4(32'h394dbe14),
	.w5(32'hba00c652),
	.w6(32'hb9cfd477),
	.w7(32'hba5b0ec2),
	.w8(32'h3aafb31b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3a792),
	.w1(32'h39d9a71c),
	.w2(32'h3aacfd95),
	.w3(32'h3aad066b),
	.w4(32'hb9ed8dc9),
	.w5(32'hbaee510c),
	.w6(32'h39707694),
	.w7(32'hba3b71ff),
	.w8(32'hb9ef4356),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91fbd6),
	.w1(32'hba055af4),
	.w2(32'hb9f8035f),
	.w3(32'h3a1ead00),
	.w4(32'h3a37f8e4),
	.w5(32'hba54092b),
	.w6(32'hba11f793),
	.w7(32'hba033859),
	.w8(32'hba4e8bce),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f5737),
	.w1(32'hb981d401),
	.w2(32'hb9c5c0e5),
	.w3(32'hb9d6c6da),
	.w4(32'h3a107511),
	.w5(32'hb9285c5c),
	.w6(32'hba3f480d),
	.w7(32'hba6e2132),
	.w8(32'hb8972067),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20651c),
	.w1(32'hba89ad1d),
	.w2(32'hbaa7df30),
	.w3(32'h3a9a03d2),
	.w4(32'h398cd763),
	.w5(32'hbac59c48),
	.w6(32'hba79edf9),
	.w7(32'hba87cf50),
	.w8(32'hbaa61805),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b0d3),
	.w1(32'hbbb01f30),
	.w2(32'hba3cf1b3),
	.w3(32'hbbb21f5a),
	.w4(32'h3a605806),
	.w5(32'hbaccf016),
	.w6(32'h3a855fbf),
	.w7(32'hbab40df8),
	.w8(32'h3a06113f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba852533),
	.w1(32'hba05c135),
	.w2(32'hbb1570e3),
	.w3(32'h3aa82787),
	.w4(32'h3abd342a),
	.w5(32'hbb07e6bd),
	.w6(32'hba61a0f2),
	.w7(32'hbaf9836b),
	.w8(32'hb9d8fbd9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba770421),
	.w1(32'h38f2dbaa),
	.w2(32'h389fbb29),
	.w3(32'h39e1a0de),
	.w4(32'h3a0e7be3),
	.w5(32'hba0ab614),
	.w6(32'hba22499f),
	.w7(32'hba805e65),
	.w8(32'hb8cc71af),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b9ae4),
	.w1(32'hb92fffaa),
	.w2(32'hba3ccaeb),
	.w3(32'h3a493c62),
	.w4(32'h3a627548),
	.w5(32'hba872b9d),
	.w6(32'hba078403),
	.w7(32'hba86446a),
	.w8(32'h3acaa153),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfb1e5),
	.w1(32'h3a41a7c9),
	.w2(32'h3aef9f33),
	.w3(32'h3acfdef3),
	.w4(32'hba09f4ea),
	.w5(32'hbaf46333),
	.w6(32'h398c6eae),
	.w7(32'hb9d7fa46),
	.w8(32'h39dfd14c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad51641),
	.w1(32'h3a21b405),
	.w2(32'h3adb1204),
	.w3(32'h39814f40),
	.w4(32'h398c678c),
	.w5(32'h376b6762),
	.w6(32'h3a89c09c),
	.w7(32'h3a575c9d),
	.w8(32'h3ab3fb6f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39395891),
	.w1(32'hba4de08a),
	.w2(32'hba23c6da),
	.w3(32'h3a79a806),
	.w4(32'hb9f4f835),
	.w5(32'hbaec7ae6),
	.w6(32'hba8987d0),
	.w7(32'hba5e961f),
	.w8(32'hbaf82db0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b9d65),
	.w1(32'hbad426b6),
	.w2(32'hbb9905ce),
	.w3(32'hbaefa70e),
	.w4(32'hbaede024),
	.w5(32'hbb7b82ed),
	.w6(32'hbb678be2),
	.w7(32'hbb0ef3f3),
	.w8(32'hb9bc5327),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d984b2),
	.w1(32'h38d6d64c),
	.w2(32'hb9c6133e),
	.w3(32'h3a4bad22),
	.w4(32'h39adfed8),
	.w5(32'hba9e5073),
	.w6(32'h3966177f),
	.w7(32'hba9a96fa),
	.w8(32'h3a3ce3c5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0d6cd),
	.w1(32'hb99920c3),
	.w2(32'hba04ed9f),
	.w3(32'h3ab0d697),
	.w4(32'h38f3a336),
	.w5(32'hbac7d3eb),
	.w6(32'hbaca8e28),
	.w7(32'hbb217e3c),
	.w8(32'h3b48abed),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac41690),
	.w1(32'hbbeedb30),
	.w2(32'hba9c2685),
	.w3(32'h3aa3569e),
	.w4(32'h3a16da61),
	.w5(32'hbbf7d5d7),
	.w6(32'hbbab0a6f),
	.w7(32'hbc15a7de),
	.w8(32'h38d86d56),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97aa3e),
	.w1(32'h392a6720),
	.w2(32'h3a7269aa),
	.w3(32'h3903aa2f),
	.w4(32'h3a8655a3),
	.w5(32'h3aabfe22),
	.w6(32'h39f5df0f),
	.w7(32'h3a2b637e),
	.w8(32'hba80ef7a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e2876),
	.w1(32'hb99b183a),
	.w2(32'hba3ef279),
	.w3(32'hba354644),
	.w4(32'h3929ffe8),
	.w5(32'hba9b2289),
	.w6(32'hb942b38f),
	.w7(32'hba51fe06),
	.w8(32'hba5d4b2c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30ca09),
	.w1(32'h3925312a),
	.w2(32'h3b050d9c),
	.w3(32'hba40ab4f),
	.w4(32'h39effc6d),
	.w5(32'h3b83da78),
	.w6(32'hba7c0091),
	.w7(32'h3b441a33),
	.w8(32'h3a474b27),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba085adb),
	.w1(32'h3abba590),
	.w2(32'hb9e40de0),
	.w3(32'h3a86f56d),
	.w4(32'h3a03f321),
	.w5(32'hbac3f7e1),
	.w6(32'h3a3d2c89),
	.w7(32'hb9e71bc4),
	.w8(32'hba89ff4d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6beda9),
	.w1(32'hbab0f793),
	.w2(32'hbb315f7f),
	.w3(32'hbb7fc5c9),
	.w4(32'hbb3327f6),
	.w5(32'hbbaa779e),
	.w6(32'hbb230a09),
	.w7(32'hbba1556f),
	.w8(32'hba3e7f51),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b262715),
	.w1(32'h39290fab),
	.w2(32'h3afb238b),
	.w3(32'hba31d1e5),
	.w4(32'h39f59ecf),
	.w5(32'h3b797a06),
	.w6(32'hba6b8ba5),
	.w7(32'h3b3812c4),
	.w8(32'hba1b7d1e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10f6a0),
	.w1(32'h391ee999),
	.w2(32'h3ad9812d),
	.w3(32'hba18f173),
	.w4(32'h39c29cfd),
	.w5(32'h3b54c46f),
	.w6(32'hba445dcd),
	.w7(32'h3b1c12f3),
	.w8(32'hbacb4699),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16bca7),
	.w1(32'h3984fa87),
	.w2(32'h3852cfc0),
	.w3(32'hbb0579fa),
	.w4(32'h39503b98),
	.w5(32'h3a56600f),
	.w6(32'h39423fb9),
	.w7(32'h3a445789),
	.w8(32'h3c278140),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c026bc9),
	.w1(32'hbba62574),
	.w2(32'h3baea9ba),
	.w3(32'h3b9b9ad3),
	.w4(32'hbb97f66d),
	.w5(32'h3b8a494e),
	.w6(32'hbb384d47),
	.w7(32'h3b890199),
	.w8(32'h39378113),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbbdaf),
	.w1(32'h3904b612),
	.w2(32'hb96a8426),
	.w3(32'h3a04cb92),
	.w4(32'h39b77c0f),
	.w5(32'hb9bd9a5b),
	.w6(32'h36d62fa1),
	.w7(32'hba0cb105),
	.w8(32'hbae2cc5c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964c467),
	.w1(32'hba711268),
	.w2(32'hbb1d4010),
	.w3(32'hbb4de761),
	.w4(32'h3a22b163),
	.w5(32'h3a1ff7a6),
	.w6(32'hbb1cff0a),
	.w7(32'hbc08efcb),
	.w8(32'hb8a1e690),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fb614),
	.w1(32'hb9df3909),
	.w2(32'hba9f6a6e),
	.w3(32'hba4d80cb),
	.w4(32'h3a6be305),
	.w5(32'hba180edd),
	.w6(32'h3ad7a0c6),
	.w7(32'h3987ed1b),
	.w8(32'hbb1158f1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1123c),
	.w1(32'hba160109),
	.w2(32'h3983da87),
	.w3(32'hbb34e68f),
	.w4(32'h39e6362d),
	.w5(32'h3b295de9),
	.w6(32'hbb4b837e),
	.w7(32'hbb569756),
	.w8(32'hba4eadf1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c24021),
	.w1(32'hb831c01a),
	.w2(32'h3aa5012a),
	.w3(32'hbb8c3be4),
	.w4(32'hbb7147f7),
	.w5(32'hbb5f1075),
	.w6(32'hba219819),
	.w7(32'hbb2b5148),
	.w8(32'h3ab17a96),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba978c88),
	.w1(32'h3a2bd929),
	.w2(32'h3ac1de4a),
	.w3(32'h3abe80cc),
	.w4(32'hba099126),
	.w5(32'hbae28784),
	.w6(32'h39b5e77b),
	.w7(32'hb9a24f91),
	.w8(32'hb75a5430),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36336b),
	.w1(32'h39d0f26c),
	.w2(32'hb90e52a2),
	.w3(32'h3a54a4b3),
	.w4(32'hb993024f),
	.w5(32'hba8fc9c0),
	.w6(32'hb9936f5c),
	.w7(32'hba8bf537),
	.w8(32'hbaef0fc4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe5d3a),
	.w1(32'h3abd8d36),
	.w2(32'hbb082d13),
	.w3(32'hbad022ca),
	.w4(32'hbaa1f720),
	.w5(32'hbad55160),
	.w6(32'hbb01164a),
	.w7(32'hb94aa020),
	.w8(32'h39e3000a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4e0f1),
	.w1(32'hb740dc1a),
	.w2(32'hb9dad8a7),
	.w3(32'h3a94a567),
	.w4(32'h3a260028),
	.w5(32'hba11a5a1),
	.w6(32'h3893ed55),
	.w7(32'hba391518),
	.w8(32'h39c25db7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e6054),
	.w1(32'h3a272618),
	.w2(32'h3b5e5a39),
	.w3(32'hb9b92854),
	.w4(32'h3a13c145),
	.w5(32'h3a81bda8),
	.w6(32'h3b0484c6),
	.w7(32'h3b19eccd),
	.w8(32'hbaff5d9d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba809f9c),
	.w1(32'hba0afbea),
	.w2(32'hba0cb88c),
	.w3(32'hbb2f05e3),
	.w4(32'hba4740ad),
	.w5(32'hba2f44ff),
	.w6(32'hba3801cb),
	.w7(32'hba207456),
	.w8(32'hb9a39f50),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a861158),
	.w1(32'h38079087),
	.w2(32'h3a31ae5c),
	.w3(32'hb99d58ba),
	.w4(32'h393107f7),
	.w5(32'h3ac31af2),
	.w6(32'hb9b5f848),
	.w7(32'h3a8e7414),
	.w8(32'h3a4e4c72),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80cea3),
	.w1(32'hb9b2b39f),
	.w2(32'hba808cb7),
	.w3(32'h3a11dd9a),
	.w4(32'hb897d0f4),
	.w5(32'hba2f7f5d),
	.w6(32'h39ab9191),
	.w7(32'hb9a4ad5d),
	.w8(32'h3b0c5db2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba637e5a),
	.w1(32'hbb4c58ab),
	.w2(32'hbb55eaca),
	.w3(32'hbb282597),
	.w4(32'hbb440885),
	.w5(32'hbb110529),
	.w6(32'hb91d48af),
	.w7(32'hbad10e22),
	.w8(32'hb910788c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39855262),
	.w1(32'hba5362e4),
	.w2(32'hba8483a4),
	.w3(32'h3a0e8081),
	.w4(32'hba725517),
	.w5(32'hba887a72),
	.w6(32'hb9d3bdb5),
	.w7(32'hb9eb5ac9),
	.w8(32'h3ac0a1e4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dc62a),
	.w1(32'h3a4cf422),
	.w2(32'h398675c6),
	.w3(32'h3a95bf0e),
	.w4(32'h39cd47c6),
	.w5(32'h38bf7575),
	.w6(32'h3a97ec1d),
	.w7(32'h3a363494),
	.w8(32'hb725d2b1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ffbe6),
	.w1(32'h38829adb),
	.w2(32'hba96e2e9),
	.w3(32'hba93980f),
	.w4(32'hba08dd95),
	.w5(32'hbb164094),
	.w6(32'h3aae52f7),
	.w7(32'hb9c6d742),
	.w8(32'h3b1899fb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58711e),
	.w1(32'h3b69f55d),
	.w2(32'h3a9a5cc9),
	.w3(32'hbb1eab9c),
	.w4(32'hbbf5113e),
	.w5(32'hba48bde9),
	.w6(32'h3b745ec5),
	.w7(32'h3a8ae712),
	.w8(32'hb8e26cd8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f00cf2),
	.w1(32'hbb1bb1e9),
	.w2(32'hbae865a0),
	.w3(32'hb9aebcb7),
	.w4(32'hbae910ad),
	.w5(32'hbb3a9c55),
	.w6(32'hbafa4320),
	.w7(32'hba85ada2),
	.w8(32'h3a6fdac2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab55335),
	.w1(32'h3a251142),
	.w2(32'h3a5b346e),
	.w3(32'h3b248195),
	.w4(32'h3b2f4361),
	.w5(32'h3b3cee6e),
	.w6(32'hb9949574),
	.w7(32'hb82cfdac),
	.w8(32'h3a84cdfd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87f1a4),
	.w1(32'h380a367b),
	.w2(32'hba318670),
	.w3(32'h3a6eefdd),
	.w4(32'hb818ce7d),
	.w5(32'hba383371),
	.w6(32'h3a81d708),
	.w7(32'h3953316e),
	.w8(32'h39e1932c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12b438),
	.w1(32'hb860bab5),
	.w2(32'hb880d19d),
	.w3(32'h3a5b6b5d),
	.w4(32'h38b5344a),
	.w5(32'hb8b57686),
	.w6(32'h39903907),
	.w7(32'h399a0bcb),
	.w8(32'h3a458991),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed7ed),
	.w1(32'hba3b12d4),
	.w2(32'hba457d90),
	.w3(32'h3ab4eda9),
	.w4(32'hba11d7cd),
	.w5(32'hba29d8ca),
	.w6(32'h37e8af56),
	.w7(32'h3799e8f9),
	.w8(32'h3a85a445),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf40c8),
	.w1(32'h3c1454ed),
	.w2(32'hb9866757),
	.w3(32'hbb951b87),
	.w4(32'h3b856bf3),
	.w5(32'h3a4d650d),
	.w6(32'h3bb41b35),
	.w7(32'hbab303cb),
	.w8(32'hb981ce11),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2489f3),
	.w1(32'h3ad166bd),
	.w2(32'h3adeac3f),
	.w3(32'h3b0782b6),
	.w4(32'h3b63c787),
	.w5(32'h3b769539),
	.w6(32'h3a9ff1ce),
	.w7(32'h3ac85576),
	.w8(32'h3a9152f9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78c4e1),
	.w1(32'h3b049fdf),
	.w2(32'hbb074d4c),
	.w3(32'h39825ef7),
	.w4(32'hba5926c0),
	.w5(32'hbb19b598),
	.w6(32'h3b5de319),
	.w7(32'hbb2665ea),
	.w8(32'hbab55dbe),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab92b1f),
	.w1(32'h3ac64e94),
	.w2(32'hbbdf4893),
	.w3(32'hbb2ef960),
	.w4(32'hbb1ee735),
	.w5(32'hbba6dd3b),
	.w6(32'hbb069980),
	.w7(32'hbbdc4954),
	.w8(32'hbaab222b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1291a),
	.w1(32'h39aa3b8b),
	.w2(32'h3b2870c8),
	.w3(32'h3a6fd670),
	.w4(32'hb9b655b4),
	.w5(32'hba89714b),
	.w6(32'hbad13247),
	.w7(32'h3a50bfb8),
	.w8(32'h3b0337cd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ce1db),
	.w1(32'hb9e73627),
	.w2(32'h3a40f376),
	.w3(32'hbb2e8138),
	.w4(32'h3aea0efa),
	.w5(32'hbb1f5b24),
	.w6(32'hbb3eddc9),
	.w7(32'hbae58ccd),
	.w8(32'h3b3878a3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29ef18),
	.w1(32'hb8d66261),
	.w2(32'h39fe3408),
	.w3(32'h3b770d09),
	.w4(32'h3aad24ff),
	.w5(32'h3ace67a0),
	.w6(32'hb995d62c),
	.w7(32'h397c0700),
	.w8(32'hbbd4cbfe),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc432c),
	.w1(32'hb9b50810),
	.w2(32'hbb8a04d4),
	.w3(32'hbbde5071),
	.w4(32'hbb9621a6),
	.w5(32'hbba60018),
	.w6(32'hbb33e2e3),
	.w7(32'hbb784f8a),
	.w8(32'hba8ac165),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe758d),
	.w1(32'hba29a622),
	.w2(32'hba45ee04),
	.w3(32'hbb84944b),
	.w4(32'hbb999417),
	.w5(32'hbb64a6d7),
	.w6(32'hbaeea769),
	.w7(32'h3a938080),
	.w8(32'hba0deecc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d83e38),
	.w1(32'hbb1835e7),
	.w2(32'hbb09f20c),
	.w3(32'hbaf784db),
	.w4(32'hbaf261fc),
	.w5(32'hbb561198),
	.w6(32'h39e279be),
	.w7(32'hbaa58bc1),
	.w8(32'h3a4cb24d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f9434),
	.w1(32'hba97b9ce),
	.w2(32'hbaa41441),
	.w3(32'h3b154616),
	.w4(32'h398aecc8),
	.w5(32'hba405984),
	.w6(32'hb9418327),
	.w7(32'hb914d2f9),
	.w8(32'hbb01d355),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab00017),
	.w1(32'h39ddebd2),
	.w2(32'h3b12a038),
	.w3(32'hbb6ac301),
	.w4(32'hbb5ee1c5),
	.w5(32'h3a08e5b7),
	.w6(32'hbb5185a4),
	.w7(32'hbb3633a1),
	.w8(32'h3a03abbe),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule