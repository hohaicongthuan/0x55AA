module layer_10_featuremap_470(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dcec3),
	.w1(32'hb9cf34c5),
	.w2(32'hba21b019),
	.w3(32'h38ebcbfb),
	.w4(32'hb98ff559),
	.w5(32'hba60bbba),
	.w6(32'hb9e80720),
	.w7(32'h3a2346c3),
	.w8(32'h398492a3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26faec),
	.w1(32'hba520bd9),
	.w2(32'h39e6bfd9),
	.w3(32'hba769f6b),
	.w4(32'hbae964f3),
	.w5(32'h3a50bf31),
	.w6(32'hba8e2fd0),
	.w7(32'hbb1523cc),
	.w8(32'hb91f23a2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e97daa),
	.w1(32'h3a17551b),
	.w2(32'h39b12628),
	.w3(32'hba1a17fe),
	.w4(32'h3a9ecc6b),
	.w5(32'hb9d87b2d),
	.w6(32'hb9b178c3),
	.w7(32'h39488c28),
	.w8(32'hb97439d7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b195652),
	.w1(32'h3ad6308f),
	.w2(32'h3af5d45d),
	.w3(32'h39bdc822),
	.w4(32'h3a13b7e9),
	.w5(32'h3ac159b1),
	.w6(32'h397b64e7),
	.w7(32'hba8478c6),
	.w8(32'h3a1f4f7b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f1f0b3),
	.w1(32'hb9a2f3ba),
	.w2(32'h38eadd6c),
	.w3(32'h396f5165),
	.w4(32'hba5a9aaa),
	.w5(32'hb94c0257),
	.w6(32'hb8b94376),
	.w7(32'hba13cd33),
	.w8(32'hb7b8e2d4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb468d68e),
	.w1(32'h39796e48),
	.w2(32'h3b099a23),
	.w3(32'hb9ff0c17),
	.w4(32'h3b0ad1f9),
	.w5(32'h3bb7442f),
	.w6(32'hb97f6d77),
	.w7(32'h3ab6a70e),
	.w8(32'h3b5e1881),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae46617),
	.w1(32'hbb0a3805),
	.w2(32'hbb06dbee),
	.w3(32'h3b2b23ac),
	.w4(32'hbb16d9be),
	.w5(32'hbb8ea4c8),
	.w6(32'h3b484caa),
	.w7(32'hba8c04e0),
	.w8(32'hbb0189dc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a3a7b),
	.w1(32'hba93132e),
	.w2(32'hbb9109be),
	.w3(32'h390795a3),
	.w4(32'h3a8fa3fd),
	.w5(32'hbb0f73d8),
	.w6(32'hbb59960a),
	.w7(32'hbaf01e04),
	.w8(32'hbb93cc95),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f1299),
	.w1(32'h3a1fbc69),
	.w2(32'h3a9da5e8),
	.w3(32'hba56fee3),
	.w4(32'h37bfec10),
	.w5(32'h3999aa01),
	.w6(32'hba48395e),
	.w7(32'hb7c9a6c6),
	.w8(32'hba57349f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22b890),
	.w1(32'hbaeb596e),
	.w2(32'hbb60e1b4),
	.w3(32'hbb133bd6),
	.w4(32'hba87ed96),
	.w5(32'hbb70f82e),
	.w6(32'hbb33b716),
	.w7(32'hbb08bd52),
	.w8(32'hbb947051),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4dd665),
	.w1(32'hb9ea36d8),
	.w2(32'hba0622b3),
	.w3(32'hb9840bd4),
	.w4(32'hba0e395d),
	.w5(32'hb98ddaf1),
	.w6(32'hb8ff0ad8),
	.w7(32'hba10e718),
	.w8(32'hb8fd2ada),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f8579),
	.w1(32'hbadf8cdb),
	.w2(32'hbb3ceeaf),
	.w3(32'h3b43efc0),
	.w4(32'hbace899f),
	.w5(32'hbb841bc0),
	.w6(32'h3b2925ac),
	.w7(32'hba4e5042),
	.w8(32'hbb618f66),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b04eb),
	.w1(32'hbb3da639),
	.w2(32'hbb54ae87),
	.w3(32'hbb544f0a),
	.w4(32'hbb074916),
	.w5(32'hbaad25f2),
	.w6(32'hbb77c5f2),
	.w7(32'hbb94fbf8),
	.w8(32'hbba4b19e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3be2a4),
	.w1(32'hba03f1dc),
	.w2(32'hb91407af),
	.w3(32'h3a63effc),
	.w4(32'hba04d493),
	.w5(32'hb8541b73),
	.w6(32'h392a1c9a),
	.w7(32'hba16a3df),
	.w8(32'h3a81411e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4ab9d),
	.w1(32'h38b88e4d),
	.w2(32'h388a6422),
	.w3(32'hb9e51d7b),
	.w4(32'hbab2cf9a),
	.w5(32'h3a75070c),
	.w6(32'h38b6f165),
	.w7(32'hbabe4b01),
	.w8(32'hba078c3a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4de04a),
	.w1(32'hbb118526),
	.w2(32'hbbb9a351),
	.w3(32'hba9b9b21),
	.w4(32'hbabe4b04),
	.w5(32'hbb7d73f7),
	.w6(32'hba89b728),
	.w7(32'hbafd0a6a),
	.w8(32'hbb93490d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f6d68),
	.w1(32'hbad71d26),
	.w2(32'hbaa4e769),
	.w3(32'h39f9f723),
	.w4(32'hbaf7188b),
	.w5(32'hba9e7278),
	.w6(32'hb822564f),
	.w7(32'hbaf1d0c7),
	.w8(32'hbade49f8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3883c4),
	.w1(32'hbb82e727),
	.w2(32'hbbe0957c),
	.w3(32'h3a83b54e),
	.w4(32'hbb1b0a05),
	.w5(32'hbbb79b1a),
	.w6(32'hba414a3e),
	.w7(32'hbb33f242),
	.w8(32'hbbe55877),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab97fb9),
	.w1(32'hbb86471c),
	.w2(32'hbb9988cb),
	.w3(32'hbac65207),
	.w4(32'hbb72e0ea),
	.w5(32'hbb8e353c),
	.w6(32'hbaa4059b),
	.w7(32'hbb89af8e),
	.w8(32'hbbd7c7f8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c35c5),
	.w1(32'hbae609bd),
	.w2(32'hba16b248),
	.w3(32'hbaf41f06),
	.w4(32'hba7a0d27),
	.w5(32'hba99aeaa),
	.w6(32'hbaa6e037),
	.w7(32'h390c30d0),
	.w8(32'hbb1e106b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac05fef),
	.w1(32'h3a9491eb),
	.w2(32'h3b175661),
	.w3(32'hbac32825),
	.w4(32'h3ab40fb9),
	.w5(32'h3b19de82),
	.w6(32'hba809eb4),
	.w7(32'h3a876518),
	.w8(32'h3a896d3d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9499894),
	.w1(32'hbb1ff0f7),
	.w2(32'hba653cf7),
	.w3(32'hba316c0b),
	.w4(32'hbb5fad21),
	.w5(32'hbb157cb7),
	.w6(32'hb9c536f9),
	.w7(32'hbb41458a),
	.w8(32'hbb172aa9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb053e71),
	.w1(32'hbae6396c),
	.w2(32'hbb9c1c07),
	.w3(32'hbb5fa558),
	.w4(32'hb78f78d1),
	.w5(32'hbaa5ba43),
	.w6(32'hba854bec),
	.w7(32'hbb051c67),
	.w8(32'hbb979372),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7de15),
	.w1(32'hba254c99),
	.w2(32'hbb36b743),
	.w3(32'hb9a6de0b),
	.w4(32'hbac57dbb),
	.w5(32'hbb2b6736),
	.w6(32'hbaee5ba7),
	.w7(32'hb95e6e1e),
	.w8(32'hbad533a1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35ae54),
	.w1(32'hba6818cf),
	.w2(32'hbb5dfc38),
	.w3(32'hbb9e76df),
	.w4(32'hbabe4b63),
	.w5(32'hbb6d2f2a),
	.w6(32'hbb6123d6),
	.w7(32'hba5d815c),
	.w8(32'hbaf55f13),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80caa7),
	.w1(32'hba481509),
	.w2(32'hbb5e17c5),
	.w3(32'hbb862913),
	.w4(32'hba5bceee),
	.w5(32'hbb7b3733),
	.w6(32'hbb883915),
	.w7(32'hba8fdb41),
	.w8(32'hbb12cf48),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27deb4),
	.w1(32'h39b14265),
	.w2(32'hb97e1a2f),
	.w3(32'hbb396d4d),
	.w4(32'h35a31bf4),
	.w5(32'hb9e26bae),
	.w6(32'hbaea3172),
	.w7(32'hb910b0c9),
	.w8(32'h3a12d1eb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f9daf),
	.w1(32'h3a1558e5),
	.w2(32'h39472fab),
	.w3(32'h3a9c4786),
	.w4(32'h3a7d7ae7),
	.w5(32'hb8585405),
	.w6(32'h3a05480f),
	.w7(32'h3ac6078e),
	.w8(32'h3a2e026c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86e5e4),
	.w1(32'hba6c0c77),
	.w2(32'hbb057324),
	.w3(32'hb9f1411b),
	.w4(32'hbaf7dbeb),
	.w5(32'hbae49603),
	.w6(32'hb99d4764),
	.w7(32'hb9951c23),
	.w8(32'hb9952151),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94fb7f),
	.w1(32'h3b6ddf90),
	.w2(32'h3b618100),
	.w3(32'hbb1052f9),
	.w4(32'h3ad8ea56),
	.w5(32'h3aaa83c8),
	.w6(32'hbaa12451),
	.w7(32'h39fc1d6d),
	.w8(32'h39e02dd0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8564f1),
	.w1(32'hba55012b),
	.w2(32'h399c2f72),
	.w3(32'hb9927e70),
	.w4(32'hb9a86e45),
	.w5(32'h3918fe75),
	.w6(32'hba33d25a),
	.w7(32'hb8b8377c),
	.w8(32'hba145e25),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79b27b),
	.w1(32'hb6a01b55),
	.w2(32'h3a00faf3),
	.w3(32'h392a1e5e),
	.w4(32'hb97e4665),
	.w5(32'h3962ac22),
	.w6(32'hba1772ea),
	.w7(32'hba87adbe),
	.w8(32'hb82eb75b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a949d46),
	.w1(32'h39d587cc),
	.w2(32'hba8741ce),
	.w3(32'hb869d04d),
	.w4(32'h3a96794e),
	.w5(32'hba2e2573),
	.w6(32'hba098e6f),
	.w7(32'h3a90fd86),
	.w8(32'hb93880f8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27d4cd),
	.w1(32'hba84d4a4),
	.w2(32'hba419c12),
	.w3(32'h390e6787),
	.w4(32'hb744d0f4),
	.w5(32'h3a0520d6),
	.w6(32'hba6ec11a),
	.w7(32'hba1a2ef4),
	.w8(32'h395cd7f2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbf782),
	.w1(32'h3a0de3ca),
	.w2(32'h3a9fbbe3),
	.w3(32'h3a6673ba),
	.w4(32'hb9d2176d),
	.w5(32'h39e861db),
	.w6(32'hb9f6b3a9),
	.w7(32'h3abc74ed),
	.w8(32'h3abe808f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab23b2d),
	.w1(32'h39d03487),
	.w2(32'h3a4199fd),
	.w3(32'h3a941375),
	.w4(32'h3a150a2e),
	.w5(32'h39f954af),
	.w6(32'h3b02a380),
	.w7(32'hb97d024c),
	.w8(32'h38bdd4ff),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82e598),
	.w1(32'hba8bdaae),
	.w2(32'hbbfc0d3c),
	.w3(32'hbaf45b68),
	.w4(32'h3af76ac1),
	.w5(32'hbba59bb8),
	.w6(32'hbbcfe91e),
	.w7(32'h3a913454),
	.w8(32'hbb795d1d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0a4e3),
	.w1(32'h3bd8e872),
	.w2(32'h3bdfe28f),
	.w3(32'h3882ba06),
	.w4(32'h3bb8ddde),
	.w5(32'h3c0b9c0e),
	.w6(32'hbafc28a9),
	.w7(32'h3ba30f00),
	.w8(32'h3c0219b4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49f099),
	.w1(32'h3b5e4aa3),
	.w2(32'h3ba9f45e),
	.w3(32'hbae312e6),
	.w4(32'h3b0a5318),
	.w5(32'h3be38b78),
	.w6(32'hba09d5d4),
	.w7(32'h3b9690e1),
	.w8(32'h3be2731d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa034c),
	.w1(32'h3abd557b),
	.w2(32'h3a50f4f7),
	.w3(32'hb9c40f35),
	.w4(32'h3b3dd7cb),
	.w5(32'h3b21520f),
	.w6(32'h3abf40eb),
	.w7(32'h3b1d7298),
	.w8(32'h3b1117a3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ec315),
	.w1(32'h3a8a7655),
	.w2(32'hba2dcb35),
	.w3(32'hb9c0fe3f),
	.w4(32'hbb081a5c),
	.w5(32'hbaad2624),
	.w6(32'h39191f07),
	.w7(32'hbb037cf2),
	.w8(32'hb9fce85a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d6bce),
	.w1(32'hbac311af),
	.w2(32'h38a31fa0),
	.w3(32'hba9f4ff4),
	.w4(32'hbafd148f),
	.w5(32'h3a5f4619),
	.w6(32'hba203bf1),
	.w7(32'hbb0e0556),
	.w8(32'hbab207e7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a846fbb),
	.w1(32'h3ab20a74),
	.w2(32'h3a35211c),
	.w3(32'h39e729cc),
	.w4(32'h3abd4eb5),
	.w5(32'h3ac866a8),
	.w6(32'h39f46eb4),
	.w7(32'h39f1ef78),
	.w8(32'h3a9c5ffc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e49861),
	.w1(32'hbaa070ed),
	.w2(32'hbbf7c7be),
	.w3(32'hb9ccc252),
	.w4(32'h3aa9c4a7),
	.w5(32'hbb8cbe47),
	.w6(32'h3aa62f9d),
	.w7(32'h389e4b63),
	.w8(32'hbbdd6b5b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a48b1),
	.w1(32'hba76c893),
	.w2(32'hbae904db),
	.w3(32'hba9ca212),
	.w4(32'hba21c79e),
	.w5(32'hba6c19e7),
	.w6(32'hbaa9551d),
	.w7(32'hbac51349),
	.w8(32'hbb1bbe8e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4911d3),
	.w1(32'hba561056),
	.w2(32'hbb3f703a),
	.w3(32'hbb1dbece),
	.w4(32'hbac65c46),
	.w5(32'hbb1a79b2),
	.w6(32'hbb381d45),
	.w7(32'hbb00a489),
	.w8(32'hbb3d0fdd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b3ada),
	.w1(32'hba02c3e2),
	.w2(32'hbac758ac),
	.w3(32'hbae7635d),
	.w4(32'h38c745eb),
	.w5(32'hba37437c),
	.w6(32'hbae99ae0),
	.w7(32'hb896326d),
	.w8(32'hb98d92a1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52405c),
	.w1(32'hbb8d650d),
	.w2(32'hbbee8b12),
	.w3(32'h3adb7b77),
	.w4(32'hbb804764),
	.w5(32'hbbe9e8dd),
	.w6(32'h3969fcf0),
	.w7(32'hbb9fb612),
	.w8(32'hbc1c4af8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35750dce),
	.w1(32'h3a56b87f),
	.w2(32'h3b17b2f8),
	.w3(32'hb99f4911),
	.w4(32'h399dddaf),
	.w5(32'h3accc0a5),
	.w6(32'h3a1419cc),
	.w7(32'h3930f70e),
	.w8(32'h3b0842f6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04fb0c),
	.w1(32'h3a558f11),
	.w2(32'h3a27bd85),
	.w3(32'h39873c87),
	.w4(32'h3a2348d0),
	.w5(32'h389430db),
	.w6(32'h396a8de0),
	.w7(32'h375b202b),
	.w8(32'h3a3eb04f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cc545),
	.w1(32'hba09ecea),
	.w2(32'hba7ddbe4),
	.w3(32'h3a3bfcf2),
	.w4(32'hbb0ee5c7),
	.w5(32'hba79bbd9),
	.w6(32'h3a351c50),
	.w7(32'hbab8e1b0),
	.w8(32'hbafde05b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4052e1),
	.w1(32'hba4a82e8),
	.w2(32'hbac13fe9),
	.w3(32'hbb3d0da8),
	.w4(32'hba296426),
	.w5(32'hbb389e4b),
	.w6(32'hbafab844),
	.w7(32'hba9e0895),
	.w8(32'hbb3cdd13),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c4e18a),
	.w1(32'hb97d27f3),
	.w2(32'hba1225a8),
	.w3(32'h3944651a),
	.w4(32'h3a317678),
	.w5(32'h39707796),
	.w6(32'hb99d2a7f),
	.w7(32'h3a95fdf4),
	.w8(32'h3a4e6023),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa99930),
	.w1(32'hbb35c4d2),
	.w2(32'hbbdf988f),
	.w3(32'h3b1bade0),
	.w4(32'hba387e07),
	.w5(32'hbb9d7a5f),
	.w6(32'h3b4b53e6),
	.w7(32'hba290654),
	.w8(32'hbbafaed4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec8e24),
	.w1(32'hb9049bf5),
	.w2(32'hbab482fd),
	.w3(32'hb9ebeabc),
	.w4(32'h39ae8a0f),
	.w5(32'hba4fb309),
	.w6(32'h38a1eaeb),
	.w7(32'hb9a0ba77),
	.w8(32'hbac95fcb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d339a0),
	.w1(32'h380bef00),
	.w2(32'hb760f9d5),
	.w3(32'hba664f27),
	.w4(32'h39d5dfb6),
	.w5(32'h3ab73590),
	.w6(32'hba927d5a),
	.w7(32'h3a5073c7),
	.w8(32'h3ae27292),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09c087),
	.w1(32'h368cbacf),
	.w2(32'hba4a9c83),
	.w3(32'hba9d3030),
	.w4(32'hb9bef97a),
	.w5(32'hbaf4b430),
	.w6(32'hba4e4fc5),
	.w7(32'hba590b09),
	.w8(32'hbad2b1a9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99731b),
	.w1(32'hb91fa435),
	.w2(32'h3b1d6400),
	.w3(32'hbb071447),
	.w4(32'hba801dab),
	.w5(32'h3b86aa0e),
	.w6(32'hbad22658),
	.w7(32'hbb0f502f),
	.w8(32'h3b223d90),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac53a0c),
	.w1(32'h3b08593f),
	.w2(32'hba642ebe),
	.w3(32'h3b0c5969),
	.w4(32'h3afeb096),
	.w5(32'hba1c8cab),
	.w6(32'h3b2bd236),
	.w7(32'h3adaa310),
	.w8(32'hba51549e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b438b9),
	.w1(32'hbb1ea302),
	.w2(32'hbb09712b),
	.w3(32'h37ca20ca),
	.w4(32'hba22f13d),
	.w5(32'hbb126356),
	.w6(32'h398ad60f),
	.w7(32'hbaa94518),
	.w8(32'hbb2c50c6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1db967),
	.w1(32'hb82b0dc3),
	.w2(32'hbb19fe53),
	.w3(32'hbb843b1e),
	.w4(32'h38c66cd2),
	.w5(32'hbaf80812),
	.w6(32'hbbb03a68),
	.w7(32'hba9a7dcb),
	.w8(32'hbb89fb0a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cebfb),
	.w1(32'hba07a2bc),
	.w2(32'hbb84d18a),
	.w3(32'h3a5d5759),
	.w4(32'h37ee8c52),
	.w5(32'hbb49794f),
	.w6(32'h39deff93),
	.w7(32'hbac7526c),
	.w8(32'hbb8d0f01),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937896c),
	.w1(32'h3a0fb036),
	.w2(32'hba81273f),
	.w3(32'hbae758a0),
	.w4(32'h390359bc),
	.w5(32'hba1c360b),
	.w6(32'hba0578b9),
	.w7(32'h3a4a196f),
	.w8(32'h3916ee35),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9688a30),
	.w1(32'hba2e4294),
	.w2(32'hbabf4494),
	.w3(32'hbac0a196),
	.w4(32'hbac4f9d7),
	.w5(32'hbb47b36d),
	.w6(32'hba5c863b),
	.w7(32'hbadbc79b),
	.w8(32'hbb311a06),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d47fcc),
	.w1(32'h3af309f8),
	.w2(32'h3ac6221c),
	.w3(32'hbad26fe7),
	.w4(32'h3af4f304),
	.w5(32'h3a541ea0),
	.w6(32'hba4c39c9),
	.w7(32'h3b0ade48),
	.w8(32'h3b0c294b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49a1e7),
	.w1(32'h3a7a1827),
	.w2(32'h3a69dc9c),
	.w3(32'h39a72996),
	.w4(32'h3a0dc794),
	.w5(32'h3a65c3da),
	.w6(32'h3a54993a),
	.w7(32'h3ae0f184),
	.w8(32'h3adedcd9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a340b24),
	.w1(32'hbb7801db),
	.w2(32'hbbcfe7ca),
	.w3(32'h3b70f441),
	.w4(32'hbb2c1fc6),
	.w5(32'hbb8dbd24),
	.w6(32'h3b2d532f),
	.w7(32'hbb18941e),
	.w8(32'hbb9dbb8e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc250a),
	.w1(32'h3b10c677),
	.w2(32'hb90799ad),
	.w3(32'hbacda475),
	.w4(32'h3b0638f4),
	.w5(32'hb95bf448),
	.w6(32'hbad176d2),
	.w7(32'h3a38472f),
	.w8(32'hbb99867f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad81ef8),
	.w1(32'hbaa8fa31),
	.w2(32'hbb766f41),
	.w3(32'h39d74cd5),
	.w4(32'hba711519),
	.w5(32'hbafceec6),
	.w6(32'h3a2cc2e6),
	.w7(32'hba8a6409),
	.w8(32'hbb75267d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72a5c6),
	.w1(32'hbaf8ebcb),
	.w2(32'hbc4db70c),
	.w3(32'hbb3b6c0d),
	.w4(32'h3b82d615),
	.w5(32'hbba69eac),
	.w6(32'hbb789a4c),
	.w7(32'hbb88bf6b),
	.w8(32'hbae76d0f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8ad23),
	.w1(32'hbb895fbb),
	.w2(32'hbc157c16),
	.w3(32'h3a4cea49),
	.w4(32'hbc2f6271),
	.w5(32'hbb65fe2f),
	.w6(32'hbb2ba83c),
	.w7(32'hbc4ce5b1),
	.w8(32'hbc50c39e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d2fbc),
	.w1(32'h3b96789c),
	.w2(32'hba859c36),
	.w3(32'hbc030761),
	.w4(32'hbbb1e82b),
	.w5(32'hbafeeeb7),
	.w6(32'hbc34c5e6),
	.w7(32'hbc101fa8),
	.w8(32'hbbfeabcc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdae86f),
	.w1(32'hba40c81a),
	.w2(32'hbc0a15f4),
	.w3(32'hbb370adf),
	.w4(32'h3b090ef2),
	.w5(32'hbbf84483),
	.w6(32'h3a827d68),
	.w7(32'h3b2619cc),
	.w8(32'hbc03f86f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95f158),
	.w1(32'h3b97ba75),
	.w2(32'hba99c20a),
	.w3(32'hba69eacc),
	.w4(32'h3bd05fd4),
	.w5(32'hbb5e7999),
	.w6(32'hbb7f62e8),
	.w7(32'h39ce23cf),
	.w8(32'hbb85782d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1d669),
	.w1(32'h3c8119f2),
	.w2(32'h3a946b64),
	.w3(32'h3b0448f4),
	.w4(32'h3b8a390f),
	.w5(32'hba7a7b1b),
	.w6(32'h3a9713ee),
	.w7(32'hbba0489d),
	.w8(32'h3b0ec1d3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa23820),
	.w1(32'h3965eebb),
	.w2(32'hba039432),
	.w3(32'h3b1d6175),
	.w4(32'hbb90786f),
	.w5(32'hbb209f8d),
	.w6(32'hbb936ed8),
	.w7(32'hbb8656e2),
	.w8(32'hbbe35764),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4c5f4),
	.w1(32'h3c39b25d),
	.w2(32'h3b16320e),
	.w3(32'hbb4b0af6),
	.w4(32'h3c6641bf),
	.w5(32'hbc28f10f),
	.w6(32'hbbaa3fb3),
	.w7(32'h3c2943d1),
	.w8(32'hbb3faef8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd127a),
	.w1(32'hbbaaf9d8),
	.w2(32'h3b1980c1),
	.w3(32'h3c604659),
	.w4(32'hbc977e24),
	.w5(32'h3cb7198e),
	.w6(32'h3ae121ea),
	.w7(32'hbbb83bd5),
	.w8(32'hbc5452d6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb341c49),
	.w1(32'h39f7f7f3),
	.w2(32'h3a45dbef),
	.w3(32'h3bfc807c),
	.w4(32'hbc0a30e8),
	.w5(32'hbc4733c7),
	.w6(32'hbb12010b),
	.w7(32'hbb47412b),
	.w8(32'hbbe5547b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2454a1),
	.w1(32'hbb83cd5f),
	.w2(32'hbbe91c34),
	.w3(32'h3b59f804),
	.w4(32'hbc1ab346),
	.w5(32'hbb58427c),
	.w6(32'hbb0377dd),
	.w7(32'hbc44c4e5),
	.w8(32'hbc60e087),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d04ea),
	.w1(32'h3c7aaeb4),
	.w2(32'h3c4d7cc7),
	.w3(32'hbaa22fb5),
	.w4(32'h3c9b749e),
	.w5(32'hbc14f66e),
	.w6(32'hbbbba1d6),
	.w7(32'h3c52d2fc),
	.w8(32'h3b69504d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b0af9),
	.w1(32'hbc3ed639),
	.w2(32'h3c21ea7d),
	.w3(32'h3b5a1f06),
	.w4(32'hbccfff4c),
	.w5(32'h3c584dd4),
	.w6(32'h3c2f026b),
	.w7(32'hbcac2b6b),
	.w8(32'hbc27ae57),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c050af1),
	.w1(32'hbb17066e),
	.w2(32'h3b88baf6),
	.w3(32'h3cbb27a6),
	.w4(32'h3ad25c90),
	.w5(32'hbaf5ac9e),
	.w6(32'h3be7812a),
	.w7(32'hbb16a24c),
	.w8(32'hbb80d893),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a185231),
	.w1(32'h3945fb00),
	.w2(32'hbb6d401b),
	.w3(32'hba2282a2),
	.w4(32'h3b0ab1e1),
	.w5(32'hbb65fbfa),
	.w6(32'hbb20dc85),
	.w7(32'hbb738ce7),
	.w8(32'hbb850728),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc043f10),
	.w1(32'hbbe3c67f),
	.w2(32'hbbfddf58),
	.w3(32'hbc636431),
	.w4(32'hbc679e40),
	.w5(32'h3ba24b78),
	.w6(32'hb8e5e6e5),
	.w7(32'h3a00654c),
	.w8(32'hbc2ca52d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8c81),
	.w1(32'h3c6681ee),
	.w2(32'h3b9a1cd2),
	.w3(32'hbb0fb33d),
	.w4(32'hbc0a89c8),
	.w5(32'h3bee02ca),
	.w6(32'hbc0a8f3b),
	.w7(32'hbb90ec88),
	.w8(32'h3a8e3bd2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55a8e3),
	.w1(32'hbb8d24bb),
	.w2(32'hbc1dfae1),
	.w3(32'hbc4c342c),
	.w4(32'h3ba9ea96),
	.w5(32'hbbbf5b80),
	.w6(32'hbbd31294),
	.w7(32'h3c42aa73),
	.w8(32'h3ad4ee14),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51d442),
	.w1(32'h3bacaeca),
	.w2(32'h3b9f0e2e),
	.w3(32'hbc4fb8f2),
	.w4(32'h3b5bb8cb),
	.w5(32'hbc8e7346),
	.w6(32'hbc1dce53),
	.w7(32'h3bc7dfa2),
	.w8(32'hbb2166c5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd96a4d),
	.w1(32'h3afc18ab),
	.w2(32'hbb941596),
	.w3(32'hbbded992),
	.w4(32'hbab08649),
	.w5(32'hbc01b102),
	.w6(32'h39d1b405),
	.w7(32'hbaecddcb),
	.w8(32'h3a4001cf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84981e),
	.w1(32'hbbb4b85d),
	.w2(32'hbb19bc5c),
	.w3(32'h3ba44440),
	.w4(32'hb96d48e7),
	.w5(32'h3c91acec),
	.w6(32'h3b9b9f9a),
	.w7(32'hbb9f8cb7),
	.w8(32'h3bc9c75f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d4f57),
	.w1(32'h3b03ef8b),
	.w2(32'h3ba19433),
	.w3(32'h3ab57b02),
	.w4(32'h3a0bbeb1),
	.w5(32'h3beb10dd),
	.w6(32'h3b80d93b),
	.w7(32'h3ae1a3d6),
	.w8(32'h3af47f90),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aacc7),
	.w1(32'hbb490848),
	.w2(32'hbba3d418),
	.w3(32'h3a1be633),
	.w4(32'h3b0be1c1),
	.w5(32'h3bb37345),
	.w6(32'h3bb0864c),
	.w7(32'h3b9acc33),
	.w8(32'h3c99d60c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8ec64),
	.w1(32'h3bff55b9),
	.w2(32'h3c0fa9d5),
	.w3(32'h3ab4a04c),
	.w4(32'h3c0d9302),
	.w5(32'h3b05c228),
	.w6(32'h3c0e8393),
	.w7(32'h3bd721c6),
	.w8(32'h3c14727c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24c019),
	.w1(32'hbbc555bf),
	.w2(32'hbb816b6a),
	.w3(32'hbbb6bc1c),
	.w4(32'h3ad0dea5),
	.w5(32'hbbc08425),
	.w6(32'hbacc8a92),
	.w7(32'hbbcb52e6),
	.w8(32'hbb3874f7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b136f4b),
	.w1(32'hbb041f24),
	.w2(32'hba78eb14),
	.w3(32'hb9be6177),
	.w4(32'h3ba23efc),
	.w5(32'hb9d8b5dd),
	.w6(32'hbaa3ba4e),
	.w7(32'h3a9b0c69),
	.w8(32'h3bed7777),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14b18b),
	.w1(32'h3a2f43d8),
	.w2(32'hbc17f3d3),
	.w3(32'hbb16df2a),
	.w4(32'h3c7a25eb),
	.w5(32'h3ac8d0d8),
	.w6(32'hbb8c4bba),
	.w7(32'h3c00a1c3),
	.w8(32'h3a724cc6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc143467),
	.w1(32'hba57b66c),
	.w2(32'h3a882093),
	.w3(32'hbcad38ec),
	.w4(32'hbc4abe55),
	.w5(32'hbaf793d0),
	.w6(32'hbbea310d),
	.w7(32'hbc2d2c9a),
	.w8(32'hbc15daea),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da998),
	.w1(32'hbbcb721c),
	.w2(32'hbc2d8c7c),
	.w3(32'h3b617427),
	.w4(32'hbace48bf),
	.w5(32'hbbda70a5),
	.w6(32'h3ac08ab0),
	.w7(32'hbb99221b),
	.w8(32'hbbcce2b0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb600688),
	.w1(32'h3b087e90),
	.w2(32'h3bdd9528),
	.w3(32'hbaac03b1),
	.w4(32'h3bb33de6),
	.w5(32'h3c837960),
	.w6(32'hbc2ce483),
	.w7(32'hbb59f70a),
	.w8(32'h3bed01d0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a96b8),
	.w1(32'h3bb40898),
	.w2(32'h3b907bce),
	.w3(32'hbc090d29),
	.w4(32'h3a68f23a),
	.w5(32'h3c1e9cf4),
	.w6(32'hbc00636a),
	.w7(32'h3b62b46a),
	.w8(32'hbbf37473),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a291cdd),
	.w1(32'h3c3ff652),
	.w2(32'h3c19a432),
	.w3(32'hbae022d9),
	.w4(32'h3c58f690),
	.w5(32'hb9c79533),
	.w6(32'h3c206ac4),
	.w7(32'h3c276d52),
	.w8(32'h3ca74e41),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0909b),
	.w1(32'hbb1ce82d),
	.w2(32'hbc21ddc0),
	.w3(32'hbbfee4e7),
	.w4(32'h39d12799),
	.w5(32'h3c9f6470),
	.w6(32'h3974acc7),
	.w7(32'hbbda07fe),
	.w8(32'hbb42c2cb),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb667522),
	.w1(32'h3bb7714c),
	.w2(32'hbba7a7d2),
	.w3(32'h3b78f625),
	.w4(32'h3c06ee34),
	.w5(32'hbc02363c),
	.w6(32'hbb979f08),
	.w7(32'h3c5bf3fd),
	.w8(32'h3a0e278b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4474d),
	.w1(32'hbc54de79),
	.w2(32'hbbb52829),
	.w3(32'hbb8bc350),
	.w4(32'hbc8bee3c),
	.w5(32'h3b5299d7),
	.w6(32'hba865cd2),
	.w7(32'hbc2eb822),
	.w8(32'hbc34d272),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ece1d),
	.w1(32'h3ba5a91e),
	.w2(32'hbb826dbb),
	.w3(32'h3bbf0f80),
	.w4(32'h3beb728f),
	.w5(32'hbbf8c059),
	.w6(32'hb99516df),
	.w7(32'hb979ce2a),
	.w8(32'hbbe3302c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96339c7),
	.w1(32'hbaa5fb27),
	.w2(32'h3b94aa27),
	.w3(32'h3af4a88d),
	.w4(32'hbc0f346d),
	.w5(32'hbc588a68),
	.w6(32'h3aa8e553),
	.w7(32'hbb8822b9),
	.w8(32'hbbee0eb7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7058e5),
	.w1(32'hbb81f4b2),
	.w2(32'h3bd80367),
	.w3(32'h3c13534a),
	.w4(32'hbc5d3be5),
	.w5(32'h3c550ff3),
	.w6(32'h3b7065a3),
	.w7(32'hbc41dd32),
	.w8(32'hbbbb7637),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb763c81),
	.w1(32'h3b13e11a),
	.w2(32'hbc10aadb),
	.w3(32'h3c276e1f),
	.w4(32'h3be02e89),
	.w5(32'h3b76c74e),
	.w6(32'hbb4d518d),
	.w7(32'h3a44e476),
	.w8(32'hbc31f5a3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16bced),
	.w1(32'hb9a43736),
	.w2(32'hbc2e0275),
	.w3(32'hbc67607f),
	.w4(32'h3c1d01df),
	.w5(32'hbb354ee5),
	.w6(32'hbc2d84b9),
	.w7(32'h3a3a4e53),
	.w8(32'hbb9645d0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd49f9),
	.w1(32'h393c8f72),
	.w2(32'hbbc2b4b1),
	.w3(32'hbbd5ef66),
	.w4(32'h3c13e07d),
	.w5(32'h3bfd8cdc),
	.w6(32'hbbbc48c7),
	.w7(32'h3b99ded8),
	.w8(32'h3b7088e7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4c893),
	.w1(32'h363a8993),
	.w2(32'h3aa6bc6f),
	.w3(32'hbc392c67),
	.w4(32'hbb594947),
	.w5(32'h3afdccf9),
	.w6(32'hbb920f23),
	.w7(32'h3bbe53d5),
	.w8(32'h3b56ce73),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810609),
	.w1(32'h3b85e1d2),
	.w2(32'hba3707e8),
	.w3(32'h39b237a6),
	.w4(32'hbb8f0d31),
	.w5(32'h3cf74511),
	.w6(32'hbba35a4b),
	.w7(32'hbc4fe5f5),
	.w8(32'h3b872378),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1372ec),
	.w1(32'h3b18c7fb),
	.w2(32'h3a1ad14a),
	.w3(32'hbbabf776),
	.w4(32'h3be55c73),
	.w5(32'h3a58d776),
	.w6(32'hbb4637c6),
	.w7(32'h3b634438),
	.w8(32'hbb6a6acf),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba607a4),
	.w1(32'hbb499004),
	.w2(32'hbc23f8cb),
	.w3(32'h3a59b0fb),
	.w4(32'hbc3ef46d),
	.w5(32'hbc734523),
	.w6(32'h3b1f83fa),
	.w7(32'hbb843ea4),
	.w8(32'hbb2c352d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0920d),
	.w1(32'h3c10f2fa),
	.w2(32'hbbec3a29),
	.w3(32'h3bc459f5),
	.w4(32'h3d00cfc1),
	.w5(32'hbcc1338c),
	.w6(32'hbab77af3),
	.w7(32'h3cbf9f9f),
	.w8(32'h3a88337b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd62a34),
	.w1(32'h39ee6b99),
	.w2(32'hbbaa2acd),
	.w3(32'hbbb63261),
	.w4(32'hbc1a0b84),
	.w5(32'hbc2c1f67),
	.w6(32'hbc1d46f4),
	.w7(32'hbb382b89),
	.w8(32'hbc36afde),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb25e3a),
	.w1(32'hbb1afb12),
	.w2(32'h3b21474e),
	.w3(32'hbbaca254),
	.w4(32'hba09e343),
	.w5(32'hbc1dfd5b),
	.w6(32'hbc464138),
	.w7(32'h3bb64e7d),
	.w8(32'hbc3e2819),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e9518),
	.w1(32'hbbd56d5a),
	.w2(32'h3baeaee0),
	.w3(32'h3c7b2be2),
	.w4(32'hbc32ef72),
	.w5(32'h3b1f6582),
	.w6(32'h3bdd60bf),
	.w7(32'hbbb73751),
	.w8(32'hbab2bcff),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cf7c5),
	.w1(32'hbad8c0fc),
	.w2(32'hbbed032f),
	.w3(32'h3b6cc358),
	.w4(32'hbb58222a),
	.w5(32'hbb946b0c),
	.w6(32'hbb28d3d0),
	.w7(32'hbb8eada0),
	.w8(32'hbad50cbd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f59e3),
	.w1(32'hbb6e89e6),
	.w2(32'hbc15e8f4),
	.w3(32'hbc093e9d),
	.w4(32'h3c589e7c),
	.w5(32'hbbe6cbf9),
	.w6(32'h3b3f967b),
	.w7(32'h3bb668b5),
	.w8(32'hbc2374b0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54f28c),
	.w1(32'hbb80fece),
	.w2(32'hb99961b4),
	.w3(32'hbc607caa),
	.w4(32'h3c10a4bd),
	.w5(32'hbc91689b),
	.w6(32'hbc021d74),
	.w7(32'hba946da0),
	.w8(32'hbbec6388),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa88d27),
	.w1(32'h3b41698f),
	.w2(32'hba8ba54f),
	.w3(32'h3c84701f),
	.w4(32'h3c328af1),
	.w5(32'hb9b3457a),
	.w6(32'h3b0bfcc6),
	.w7(32'hbb0a4474),
	.w8(32'hbacb8116),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e257b),
	.w1(32'hbb80461d),
	.w2(32'h3b4bbe1a),
	.w3(32'h3913a339),
	.w4(32'hbb9fbd10),
	.w5(32'hbbe06e25),
	.w6(32'hbb68c6b9),
	.w7(32'hbc1d0689),
	.w8(32'hbb65846b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc21827),
	.w1(32'h3bc6421f),
	.w2(32'h3b5d3bdb),
	.w3(32'hbc1f7fa4),
	.w4(32'hbc094d49),
	.w5(32'h3cb94837),
	.w6(32'hbbdfcafb),
	.w7(32'hbc38c42b),
	.w8(32'h3a773881),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cc0c3),
	.w1(32'hbb5c6157),
	.w2(32'hba532dce),
	.w3(32'h3b893dc3),
	.w4(32'hbc2429b0),
	.w5(32'h3c3b7929),
	.w6(32'h3bb2373b),
	.w7(32'hbb04ccee),
	.w8(32'hbbef6984),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f16fe),
	.w1(32'h3c149f09),
	.w2(32'hbb91ee56),
	.w3(32'h3a08fc30),
	.w4(32'h3bdc8293),
	.w5(32'hbbccd259),
	.w6(32'h3aed14ee),
	.w7(32'h3a678066),
	.w8(32'hbaf1853c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38483a66),
	.w1(32'hbc099edf),
	.w2(32'h3ae1547d),
	.w3(32'h3beee224),
	.w4(32'hbc53238b),
	.w5(32'h3bbd1e69),
	.w6(32'h385b30ea),
	.w7(32'hbc69fb2f),
	.w8(32'hbb22b16f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1253f),
	.w1(32'h3bb4df3c),
	.w2(32'hbb01c990),
	.w3(32'hbb6f2c86),
	.w4(32'hbb51467c),
	.w5(32'h38985085),
	.w6(32'h3c0e3bd3),
	.w7(32'hbb9e42e5),
	.w8(32'h3bd930a3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6e730),
	.w1(32'h3c60e45c),
	.w2(32'hbb888023),
	.w3(32'h3b87e148),
	.w4(32'h3d11f181),
	.w5(32'h39f2bebf),
	.w6(32'hb946fcca),
	.w7(32'h3c8f165a),
	.w8(32'h3c868635),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24ab91),
	.w1(32'hbbbabc7e),
	.w2(32'hbc0b08f5),
	.w3(32'hbcf05895),
	.w4(32'hbbd9b511),
	.w5(32'hbbab820e),
	.w6(32'hbbf92c57),
	.w7(32'hbbe6aeb0),
	.w8(32'hbb83da97),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d7e0d),
	.w1(32'h3bc98815),
	.w2(32'hbb99dca9),
	.w3(32'h3aa6c6fb),
	.w4(32'h3ca126d1),
	.w5(32'h39616c57),
	.w6(32'hbac29aa1),
	.w7(32'h3b839b9b),
	.w8(32'h3b6f9132),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fa2bf),
	.w1(32'h3baf4f77),
	.w2(32'hbc293399),
	.w3(32'hbb8a7747),
	.w4(32'h3be6bc93),
	.w5(32'hbc623be6),
	.w6(32'h3a2b3f5c),
	.w7(32'hbb1837ab),
	.w8(32'hbb51a5bb),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe44e36),
	.w1(32'h3b6af4f5),
	.w2(32'h3bec5a54),
	.w3(32'hbc6ff5d1),
	.w4(32'h3c05aa04),
	.w5(32'h3c62be28),
	.w6(32'hbb6cb0a7),
	.w7(32'h3b30b0eb),
	.w8(32'h3be09a86),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d462b),
	.w1(32'hbb74be78),
	.w2(32'hbae45017),
	.w3(32'h3b808e2a),
	.w4(32'hbc02a2ab),
	.w5(32'h3bdec053),
	.w6(32'hb9e979a1),
	.w7(32'hbbe7d305),
	.w8(32'h39083f39),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb998820),
	.w1(32'hbb2d8019),
	.w2(32'h39bb1083),
	.w3(32'h3baf7b8c),
	.w4(32'hbba13091),
	.w5(32'h3ba35393),
	.w6(32'h3b2ac084),
	.w7(32'h39f29a25),
	.w8(32'hbaeac824),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fc855),
	.w1(32'hbbf00649),
	.w2(32'hb88a952e),
	.w3(32'h3b197b5f),
	.w4(32'hba5b91ee),
	.w5(32'h3b4a019c),
	.w6(32'h3b5dc22c),
	.w7(32'hbbe93665),
	.w8(32'h3bd1b534),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e6d4a),
	.w1(32'h3be271b0),
	.w2(32'hbc2a4a96),
	.w3(32'h3a8e7a26),
	.w4(32'h3c0a5b5e),
	.w5(32'hbc07a4c7),
	.w6(32'hb9f6a85e),
	.w7(32'h3b330fcb),
	.w8(32'hbbdceb41),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccae07),
	.w1(32'h3a56cb01),
	.w2(32'hbc2afd31),
	.w3(32'hbbdd71bb),
	.w4(32'h3bb6f067),
	.w5(32'hbbc64c62),
	.w6(32'hbaf04160),
	.w7(32'hbae68598),
	.w8(32'hbb5a3112),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4057d9),
	.w1(32'h3ad11b9a),
	.w2(32'hbb3a8fdd),
	.w3(32'hba5808a7),
	.w4(32'hbbf15e84),
	.w5(32'h3b2244b3),
	.w6(32'hbaf51ef4),
	.w7(32'hbc04cdad),
	.w8(32'hbbd2488f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a812966),
	.w1(32'hbbd07f50),
	.w2(32'h3bef5aa2),
	.w3(32'h39ff7fba),
	.w4(32'hbc710ab3),
	.w5(32'h388f51cd),
	.w6(32'hbb56ca30),
	.w7(32'hbc29121d),
	.w8(32'hbbe73f08),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f06ed),
	.w1(32'hbb88bd7c),
	.w2(32'hbb5b99b4),
	.w3(32'h3cd7af0b),
	.w4(32'hbc79fca2),
	.w5(32'h3c00a023),
	.w6(32'h3c2a4d30),
	.w7(32'hbb99f246),
	.w8(32'hbc67ab0b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2cf93),
	.w1(32'hbacb6daa),
	.w2(32'h3b74bb8e),
	.w3(32'h3c008a9f),
	.w4(32'h3c1fb24a),
	.w5(32'hbb335b47),
	.w6(32'hbaa73c05),
	.w7(32'h3c1b89c4),
	.w8(32'h3c0d3c51),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10bb7a),
	.w1(32'hbc04032a),
	.w2(32'hbbc62880),
	.w3(32'h3b2ac3ac),
	.w4(32'hbc8a6be1),
	.w5(32'h3cad006a),
	.w6(32'hba077321),
	.w7(32'hbc11049a),
	.w8(32'hbc8226cf),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86bfb4),
	.w1(32'hbc29b84d),
	.w2(32'hbbc7c409),
	.w3(32'hbbfe5c80),
	.w4(32'hbcb6e144),
	.w5(32'h3bf6c994),
	.w6(32'hbc871351),
	.w7(32'hbc8fe7bb),
	.w8(32'hbc8e4d31),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8c7e7),
	.w1(32'h3b191bdc),
	.w2(32'hba1d7fde),
	.w3(32'hbb7e8723),
	.w4(32'hbc079d40),
	.w5(32'h3ab607fa),
	.w6(32'hbbc398cd),
	.w7(32'hbb13a0e3),
	.w8(32'hbc038809),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36a854),
	.w1(32'h3c669b69),
	.w2(32'hbaa2a81c),
	.w3(32'h3b1e57d6),
	.w4(32'h3d065e02),
	.w5(32'hbc314b5e),
	.w6(32'h3b6434c2),
	.w7(32'h3cf20040),
	.w8(32'h3c4902c5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e3730),
	.w1(32'hbb026f37),
	.w2(32'h3b2d864a),
	.w3(32'hbc4baca4),
	.w4(32'hbc173806),
	.w5(32'h3c8510a6),
	.w6(32'hbc803923),
	.w7(32'hbbefa615),
	.w8(32'hbb89a169),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dcc81),
	.w1(32'hbc385c21),
	.w2(32'hbbd60433),
	.w3(32'h3c406ed0),
	.w4(32'hbc00b8ca),
	.w5(32'h3c8ae848),
	.w6(32'hb9efae2d),
	.w7(32'hb939ffa6),
	.w8(32'hbc3fc908),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42cae7),
	.w1(32'hba948421),
	.w2(32'h3c36d1a1),
	.w3(32'hbc3d179d),
	.w4(32'hbbcc13e8),
	.w5(32'h3bdb1307),
	.w6(32'hbbcd4d31),
	.w7(32'hbc479ed4),
	.w8(32'hbb9e20b1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6366e),
	.w1(32'hbaca22d1),
	.w2(32'h3b6376dd),
	.w3(32'h3c9f1231),
	.w4(32'hbc09b25e),
	.w5(32'h3c8739e2),
	.w6(32'h3ab1df3b),
	.w7(32'hbb9c9254),
	.w8(32'h3a12b7d1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac16f2),
	.w1(32'h3c1c82ad),
	.w2(32'h3b99e9ee),
	.w3(32'hbcb7bd63),
	.w4(32'h3aae2e37),
	.w5(32'h3b800c4b),
	.w6(32'hbc6ce2d7),
	.w7(32'h3bc13c58),
	.w8(32'hbbb28301),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fa2ab),
	.w1(32'hbbb410ae),
	.w2(32'hbb97e56f),
	.w3(32'h3c718379),
	.w4(32'h3ad871ef),
	.w5(32'h3bd28da5),
	.w6(32'hbb0288f8),
	.w7(32'hbae7984d),
	.w8(32'hbb946fa4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac35a81),
	.w1(32'h397c0ebc),
	.w2(32'hbbca1cb7),
	.w3(32'h3c0bf95d),
	.w4(32'hbc1239ae),
	.w5(32'hbbf6968c),
	.w6(32'h3bdddc46),
	.w7(32'hbc69b737),
	.w8(32'h3ab38d89),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba268bb5),
	.w1(32'h3c57833b),
	.w2(32'h3b98faac),
	.w3(32'hbb4bcc86),
	.w4(32'h3c7dfe8f),
	.w5(32'h3c98fc9f),
	.w6(32'h3b6f2806),
	.w7(32'h3bb71627),
	.w8(32'h3cd77187),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb5e56),
	.w1(32'h3b63cb50),
	.w2(32'h3aea6921),
	.w3(32'hbaf69f8c),
	.w4(32'hbbea3fd3),
	.w5(32'hbb9640aa),
	.w6(32'h3a92ab0e),
	.w7(32'hbbf74aa9),
	.w8(32'hbb045467),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb26889),
	.w1(32'h3be07f43),
	.w2(32'hbbae30de),
	.w3(32'h3b1f4bc4),
	.w4(32'h3bc054f6),
	.w5(32'h3b492cad),
	.w6(32'hbb9b0ca1),
	.w7(32'h3ad70fbe),
	.w8(32'h3b957338),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc8e52),
	.w1(32'h3bd6abe5),
	.w2(32'h3b9cbc1f),
	.w3(32'h3be73c3f),
	.w4(32'h3af11977),
	.w5(32'hbb3baade),
	.w6(32'h3c616237),
	.w7(32'h3bccf8f8),
	.w8(32'hbbacb1e5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca7349),
	.w1(32'hbbdd6a2f),
	.w2(32'h3c9d46ce),
	.w3(32'h3b10618c),
	.w4(32'hbcea6369),
	.w5(32'h3cdc05c4),
	.w6(32'hbc3b419e),
	.w7(32'hbcc16c14),
	.w8(32'hba620990),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ac456),
	.w1(32'hbbb5c6f8),
	.w2(32'h3988478a),
	.w3(32'h3ce49104),
	.w4(32'hb997ab44),
	.w5(32'h3b9bd863),
	.w6(32'h3c4a46f9),
	.w7(32'h3c20db0b),
	.w8(32'hba9d1bcd),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4089c),
	.w1(32'hbc13118a),
	.w2(32'hbbab18ea),
	.w3(32'h3c87698e),
	.w4(32'hbb444d3d),
	.w5(32'hbb09a6aa),
	.w6(32'h3bd45624),
	.w7(32'hbaa93cca),
	.w8(32'hbc03e84b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98acfd0),
	.w1(32'hbb7916e9),
	.w2(32'hbc0802b3),
	.w3(32'hbb107787),
	.w4(32'hbacc8c72),
	.w5(32'hbc418b58),
	.w6(32'hbb7521d4),
	.w7(32'hbaaca078),
	.w8(32'hb9af4f66),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc85adc),
	.w1(32'h3a5027f4),
	.w2(32'hbae5ac87),
	.w3(32'hbba1f6bf),
	.w4(32'h3b1d2038),
	.w5(32'hbabeb995),
	.w6(32'h39cc4b97),
	.w7(32'h3b1b727d),
	.w8(32'hba98e407),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5872a1),
	.w1(32'hbc24b115),
	.w2(32'h3bca81af),
	.w3(32'h3b2c29ce),
	.w4(32'hbc67aa41),
	.w5(32'hbb8114db),
	.w6(32'h3b8cc335),
	.w7(32'hbc0b4eeb),
	.w8(32'hbbb7581b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398027d6),
	.w1(32'h3bda2bb3),
	.w2(32'hbabedc56),
	.w3(32'hbb0d11ba),
	.w4(32'h3c32064e),
	.w5(32'hbc649c74),
	.w6(32'hbb8dc8b3),
	.w7(32'h3bd3ef76),
	.w8(32'hbb96d9b9),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5d124),
	.w1(32'h3b1bb4a0),
	.w2(32'hb8e15942),
	.w3(32'hbba2e3ee),
	.w4(32'hbbb3b914),
	.w5(32'h3b9b9a4b),
	.w6(32'hbbaff928),
	.w7(32'hba79eea9),
	.w8(32'hbafa436c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cca51),
	.w1(32'hbb067345),
	.w2(32'h3b89d243),
	.w3(32'hbc2dd978),
	.w4(32'hbb5d2df7),
	.w5(32'h3b8d2fd3),
	.w6(32'hbc1f760b),
	.w7(32'h3bcd9eae),
	.w8(32'hbc1425ed),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8744b1),
	.w1(32'h38c48e15),
	.w2(32'hbc34059a),
	.w3(32'h3c029e5f),
	.w4(32'h3cca9dff),
	.w5(32'h3beac1ec),
	.w6(32'h3b1a2993),
	.w7(32'h3c4ab64c),
	.w8(32'h3bda7742),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc24dc2),
	.w1(32'h3b28857e),
	.w2(32'hbbfe02b4),
	.w3(32'hbc9eed92),
	.w4(32'h3c91a935),
	.w5(32'h3b28db7b),
	.w6(32'hbbf813ed),
	.w7(32'h3c1b26fa),
	.w8(32'hb90ab376),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07cb62),
	.w1(32'hbb0942d4),
	.w2(32'hbc370f67),
	.w3(32'hbbf3e0f0),
	.w4(32'h3b189375),
	.w5(32'hbc564a45),
	.w6(32'hbbe24bcc),
	.w7(32'h3b8bbb60),
	.w8(32'hbb61cc5b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28aec4),
	.w1(32'hbaa3a8c6),
	.w2(32'h3b5eafb5),
	.w3(32'h3be67a0a),
	.w4(32'hbc42f6da),
	.w5(32'h3c4d5374),
	.w6(32'h3aa0a834),
	.w7(32'hbc227868),
	.w8(32'hbbf0d747),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cc6d1),
	.w1(32'h3ab764c7),
	.w2(32'hbb8745e6),
	.w3(32'h3bcf8f2a),
	.w4(32'h39df9a8a),
	.w5(32'h3c17cae8),
	.w6(32'hbb199a62),
	.w7(32'h3bc61f49),
	.w8(32'hbb9afda1),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2f0bb),
	.w1(32'hba0b9d26),
	.w2(32'hbc3d8325),
	.w3(32'hbb20b2ce),
	.w4(32'h3c9dde96),
	.w5(32'hbc17a433),
	.w6(32'hbb94e74c),
	.w7(32'h3bd5155b),
	.w8(32'h3c300480),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f2225),
	.w1(32'h3a69d4a3),
	.w2(32'hbc464eb9),
	.w3(32'hbca9fc24),
	.w4(32'hbb64ae34),
	.w5(32'hbc37fcf1),
	.w6(32'hbc06d482),
	.w7(32'hbb3ab279),
	.w8(32'hbc58b32d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6e1db),
	.w1(32'hbc68d7c9),
	.w2(32'hbc3eebad),
	.w3(32'hbbcab929),
	.w4(32'hbc8ebcfc),
	.w5(32'hbbc0b134),
	.w6(32'hbad996fb),
	.w7(32'hbc7338c1),
	.w8(32'hbc880e42),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0d875),
	.w1(32'h3b6bdaa9),
	.w2(32'hba2dc552),
	.w3(32'hbba56c9b),
	.w4(32'h3885bbcd),
	.w5(32'hbc576701),
	.w6(32'hbb656192),
	.w7(32'h3b8a23e6),
	.w8(32'hbb9ac490),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e9fbfe),
	.w1(32'hbc1cf695),
	.w2(32'hbb82bacf),
	.w3(32'hbb7e2adb),
	.w4(32'h3aaa43d6),
	.w5(32'h3be96992),
	.w6(32'hbbf62737),
	.w7(32'hbb92ce35),
	.w8(32'h3ba9eafa),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc212004),
	.w1(32'h3b4b986b),
	.w2(32'h3bc41c1a),
	.w3(32'hbc769f3e),
	.w4(32'h3b78bd1f),
	.w5(32'hbbc18daa),
	.w6(32'hbc2a760b),
	.w7(32'hb906035c),
	.w8(32'hbaed6d0f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1dbb4),
	.w1(32'h3b63a1ff),
	.w2(32'h3a5b005a),
	.w3(32'h3b516da0),
	.w4(32'h3c47e9a5),
	.w5(32'hbbefea99),
	.w6(32'h3bacabc0),
	.w7(32'hb8ad03a8),
	.w8(32'hbb477611),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98bf47),
	.w1(32'h3a91c150),
	.w2(32'h3aeb1514),
	.w3(32'h3b60f543),
	.w4(32'h3c605d84),
	.w5(32'hbc9e3235),
	.w6(32'hbb4bdd50),
	.w7(32'h3bdee62f),
	.w8(32'hbbd63a55),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39493b68),
	.w1(32'hbc8c2432),
	.w2(32'hbc4d7359),
	.w3(32'h3cde4446),
	.w4(32'hbca30170),
	.w5(32'hbb918252),
	.w6(32'h3bccd0a5),
	.w7(32'hbc88138b),
	.w8(32'hbc5361fa),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2554dd),
	.w1(32'h3ba8ad08),
	.w2(32'h3b98e066),
	.w3(32'hbc05acf4),
	.w4(32'h3b376b89),
	.w5(32'h3b5e4eb2),
	.w6(32'hbc27aa73),
	.w7(32'hbb91da93),
	.w8(32'h3a2af600),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ac669),
	.w1(32'h3b5fa21f),
	.w2(32'h3c24229c),
	.w3(32'hbb9fe829),
	.w4(32'h3ad1fcc5),
	.w5(32'hbc3b52f1),
	.w6(32'h381270cc),
	.w7(32'h3baea7c2),
	.w8(32'h3b296db2),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c661ed),
	.w1(32'hbbc4cd23),
	.w2(32'hbc6a7947),
	.w3(32'hbbbedf5d),
	.w4(32'hbb86daf6),
	.w5(32'hbab2ce41),
	.w6(32'hbc216e6a),
	.w7(32'h38e0d4f8),
	.w8(32'hbc3a7d3d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb092f56),
	.w1(32'hbb3d9ffa),
	.w2(32'hbc1bc31f),
	.w3(32'hbbd6897f),
	.w4(32'h3b53507b),
	.w5(32'hbb4b010d),
	.w6(32'hbc311c27),
	.w7(32'h3bc57ef0),
	.w8(32'hbb5bbb7d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb257c9d),
	.w1(32'hbb9f53d8),
	.w2(32'h3c662cd2),
	.w3(32'hbbc8f912),
	.w4(32'hbcaf4f16),
	.w5(32'h3c9c8978),
	.w6(32'hbbe2eea2),
	.w7(32'hbc20a532),
	.w8(32'h3b1267e0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c723424),
	.w1(32'h3b4237ff),
	.w2(32'hbc9e0929),
	.w3(32'h3d0f278b),
	.w4(32'h3bbf980f),
	.w5(32'hbc310351),
	.w6(32'h3cc1b906),
	.w7(32'hbb0a3740),
	.w8(32'hbbfbd3de),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b53f7),
	.w1(32'hbb60b91f),
	.w2(32'hbc55a60b),
	.w3(32'hbc35b183),
	.w4(32'hbaceced5),
	.w5(32'hbc0a37cb),
	.w6(32'hbc263abc),
	.w7(32'hbbbdb33d),
	.w8(32'hbb1b66a6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac48dd2),
	.w1(32'hbc2837cc),
	.w2(32'hbc0ea4c6),
	.w3(32'hbb16ee91),
	.w4(32'hbba63fcf),
	.w5(32'hbc48a195),
	.w6(32'hbbf51bbe),
	.w7(32'hbc0323b6),
	.w8(32'hbc3062c4),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5657df),
	.w1(32'h3c329dd9),
	.w2(32'h3b9a95bb),
	.w3(32'hba47c353),
	.w4(32'h3c2b6747),
	.w5(32'h3c3e0b4d),
	.w6(32'hbc8582e2),
	.w7(32'h3b4f599c),
	.w8(32'h3cc331e1),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfda34),
	.w1(32'hb9ba7eca),
	.w2(32'h3b8a915d),
	.w3(32'hbb5a2f3d),
	.w4(32'hbb67e887),
	.w5(32'h3be157ac),
	.w6(32'h3b4f2d04),
	.w7(32'h3b6e5e00),
	.w8(32'hbb192b14),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e576c),
	.w1(32'hbba89a38),
	.w2(32'hbc54ceb1),
	.w3(32'h3bb51f04),
	.w4(32'h3c415068),
	.w5(32'hbb1f887e),
	.w6(32'h3b51e212),
	.w7(32'h3a122e84),
	.w8(32'h37b9dc27),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7957ef),
	.w1(32'hbbcfc40c),
	.w2(32'h3c2b89c8),
	.w3(32'hbc5c73aa),
	.w4(32'hbc24bcc0),
	.w5(32'hbad99a67),
	.w6(32'hbc2dc5ae),
	.w7(32'hbb312334),
	.w8(32'h3b5a1122),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c276db1),
	.w1(32'h3bfaf800),
	.w2(32'h3c291389),
	.w3(32'h3c95a2b5),
	.w4(32'h3c042894),
	.w5(32'h3aaaea0b),
	.w6(32'h3c2549ce),
	.w7(32'h3bbed599),
	.w8(32'h3b17db39),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde8ed6),
	.w1(32'h3b85ac46),
	.w2(32'hbc01cabd),
	.w3(32'h3beb1dd5),
	.w4(32'h3c4e87e8),
	.w5(32'hbb2057b9),
	.w6(32'h3b449fc1),
	.w7(32'h3c845c67),
	.w8(32'hba28350c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00cc43),
	.w1(32'hb964be31),
	.w2(32'hbae48239),
	.w3(32'hbc87cb74),
	.w4(32'h3ac40b40),
	.w5(32'hbc806bfd),
	.w6(32'hbba5f5bc),
	.w7(32'h3b31a99d),
	.w8(32'hbab21ec6),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b8cd3),
	.w1(32'h3a486d0a),
	.w2(32'hbb4d02bb),
	.w3(32'h3a4a99b9),
	.w4(32'h3b8234d9),
	.w5(32'h3b63e8da),
	.w6(32'hbb2b9002),
	.w7(32'hbb614059),
	.w8(32'hbb09d016),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfd473),
	.w1(32'hbca47150),
	.w2(32'hbb943226),
	.w3(32'hbb909f6e),
	.w4(32'hbc04068e),
	.w5(32'h3b263947),
	.w6(32'h39c5f0a9),
	.w7(32'hbc85cc11),
	.w8(32'h3b598592),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba914e1),
	.w1(32'hbc1d206b),
	.w2(32'h3b985e9d),
	.w3(32'hbc0a3621),
	.w4(32'hbc2fea9d),
	.w5(32'h3b999161),
	.w6(32'hbbbd76fa),
	.w7(32'hbc28f201),
	.w8(32'hbaa2c51c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c026a12),
	.w1(32'h3abf4946),
	.w2(32'hbb8f553a),
	.w3(32'h3c0dac49),
	.w4(32'hba6cc2d2),
	.w5(32'hbb9d4fac),
	.w6(32'h3b97f6f1),
	.w7(32'hbb8cb16e),
	.w8(32'hbbec0762),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd46ec),
	.w1(32'hbb8fcc2b),
	.w2(32'hbb3051f0),
	.w3(32'hbbe53bc1),
	.w4(32'hbb0fd31c),
	.w5(32'hbaf883d4),
	.w6(32'hbb3b06ef),
	.w7(32'hb962e9f9),
	.w8(32'hbb8f4aa3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2621b9),
	.w1(32'hbc1094d7),
	.w2(32'hbaa830bc),
	.w3(32'hbb8553e4),
	.w4(32'hbb379a38),
	.w5(32'h3afe232c),
	.w6(32'hbb458aaa),
	.w7(32'hbbf886dc),
	.w8(32'hbabe3ddf),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf4efd),
	.w1(32'hbb99dbc4),
	.w2(32'h3965a624),
	.w3(32'h3c94b38e),
	.w4(32'hba37c007),
	.w5(32'h3ab9f7a1),
	.w6(32'h3c5bdc6d),
	.w7(32'hb9dfe3ac),
	.w8(32'h3a17e7b7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b177200),
	.w1(32'hbaacaa56),
	.w2(32'hbb21be1b),
	.w3(32'h3b0b36d2),
	.w4(32'hbbb907e2),
	.w5(32'hbb8fc2d1),
	.w6(32'hbb9f80ae),
	.w7(32'hbc2f25a5),
	.w8(32'hbc0e4919),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2135ab),
	.w1(32'hbb6bb775),
	.w2(32'h394cc35c),
	.w3(32'hbaa9eff2),
	.w4(32'hba64bd4a),
	.w5(32'h3af85264),
	.w6(32'hbb5330cd),
	.w7(32'hbb3b5043),
	.w8(32'hbb2a3b29),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cf703),
	.w1(32'h3ba7aa8f),
	.w2(32'h3a1372f1),
	.w3(32'hbb10c620),
	.w4(32'h3ba6f9e6),
	.w5(32'hbc164b25),
	.w6(32'hbb879130),
	.w7(32'h3bb72c05),
	.w8(32'hbb822f5a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3487b5),
	.w1(32'hba7d96a4),
	.w2(32'h3abc1ccc),
	.w3(32'h3b0140eb),
	.w4(32'hbbed7d9a),
	.w5(32'h3af4e498),
	.w6(32'h39aaa195),
	.w7(32'hb97c8e23),
	.w8(32'h3b93bcb6),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd8c43),
	.w1(32'h3bb22a10),
	.w2(32'h378af072),
	.w3(32'h3ad124ce),
	.w4(32'h3786d355),
	.w5(32'h39c48756),
	.w6(32'hbb8a32f3),
	.w7(32'h3a980f17),
	.w8(32'hba921a74),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb670a60),
	.w1(32'hbb761e04),
	.w2(32'hbbe674ae),
	.w3(32'h3ab60744),
	.w4(32'h3b0d1d2b),
	.w5(32'hbb29bd1d),
	.w6(32'h3b97189f),
	.w7(32'hbb07ecf5),
	.w8(32'hba8df184),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03b370),
	.w1(32'h3c044a36),
	.w2(32'h3b753d7c),
	.w3(32'h3b83a2f0),
	.w4(32'h3c36e8ef),
	.w5(32'h3a2ea4ad),
	.w6(32'hbbd9dca5),
	.w7(32'h3c4fe494),
	.w8(32'h3c081ce6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad729f7),
	.w1(32'hbb66caae),
	.w2(32'hba697348),
	.w3(32'h3b1e5752),
	.w4(32'hba95987c),
	.w5(32'h3ba9c3bf),
	.w6(32'h3be74523),
	.w7(32'hba04ecc2),
	.w8(32'h3afeec2d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985cfa4),
	.w1(32'h3b6ef0d5),
	.w2(32'h3b246cd6),
	.w3(32'hb8b36099),
	.w4(32'hbaa5d4c9),
	.w5(32'h3b516b3c),
	.w6(32'hbb0f144d),
	.w7(32'hbb27072a),
	.w8(32'hba7a5585),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b359b58),
	.w1(32'h3b5343b2),
	.w2(32'h3a8aba5a),
	.w3(32'h3b1d12bb),
	.w4(32'h3b99542a),
	.w5(32'h3b756edd),
	.w6(32'hbaf7e511),
	.w7(32'h3b32435b),
	.w8(32'hbc1c2a74),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe4f07),
	.w1(32'hbbdc273d),
	.w2(32'hbbb63f59),
	.w3(32'hbbac46e2),
	.w4(32'hbb4afdd7),
	.w5(32'hbad22cca),
	.w6(32'hbb86e34c),
	.w7(32'hbb133629),
	.w8(32'hbb6040f7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3a67c),
	.w1(32'hbb19512a),
	.w2(32'h3c1b6605),
	.w3(32'hbba66091),
	.w4(32'h3a976f9b),
	.w5(32'h3c9c80f0),
	.w6(32'hbbc2ce73),
	.w7(32'h3bccc1a0),
	.w8(32'hbb007058),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5b765),
	.w1(32'hbbcba997),
	.w2(32'hbc18447f),
	.w3(32'h3aeab1a6),
	.w4(32'hbbe3d6ee),
	.w5(32'hbc25a06e),
	.w6(32'hbb1cf2f0),
	.w7(32'hbb9b6cb4),
	.w8(32'hbbbebd7e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba57f37),
	.w1(32'hbc015b13),
	.w2(32'hbc0617f5),
	.w3(32'hbbb89bac),
	.w4(32'hbc1ea5c7),
	.w5(32'hbc18d0b3),
	.w6(32'hbb37b876),
	.w7(32'hbba6e028),
	.w8(32'hbb1c12f3),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a29b),
	.w1(32'h3abe3dd3),
	.w2(32'h3a4b2ebb),
	.w3(32'h3b47b98b),
	.w4(32'h3b848a35),
	.w5(32'hbc068e79),
	.w6(32'hbb9c1332),
	.w7(32'h3a6d8002),
	.w8(32'hb9f413cc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081b13),
	.w1(32'h3bc8dad1),
	.w2(32'h3b3b345c),
	.w3(32'hbaaec1ea),
	.w4(32'h3c931d76),
	.w5(32'h3c39e940),
	.w6(32'hba98a102),
	.w7(32'h3bdaa98c),
	.w8(32'h3c1b3121),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9666c),
	.w1(32'hbabb4b82),
	.w2(32'hbb8a0519),
	.w3(32'hb9f64ccf),
	.w4(32'h3b103a20),
	.w5(32'hbbd4681f),
	.w6(32'hbb888923),
	.w7(32'hbb2fadd7),
	.w8(32'hbba3d745),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbefd4),
	.w1(32'hba01a8b7),
	.w2(32'hba6b1dbb),
	.w3(32'hba7d6192),
	.w4(32'hbad51bb7),
	.w5(32'h386e9216),
	.w6(32'h3b881d71),
	.w7(32'h3b04c895),
	.w8(32'hbae26401),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb212c36),
	.w1(32'h3a8a3e7d),
	.w2(32'h3b8ce73a),
	.w3(32'h3a95eed1),
	.w4(32'hbba2ea63),
	.w5(32'h3b91cb3c),
	.w6(32'hbb9f1b49),
	.w7(32'h3b2f9057),
	.w8(32'h3b808d1c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93269d),
	.w1(32'hbbb6d785),
	.w2(32'hba812ae5),
	.w3(32'hbb94add0),
	.w4(32'hbb41e8ef),
	.w5(32'h3bbb9af4),
	.w6(32'hbbb06b82),
	.w7(32'hbb33ba53),
	.w8(32'h3aa57661),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aa8fd),
	.w1(32'hbba2e52d),
	.w2(32'h3ae82b9c),
	.w3(32'hb9c6d7ad),
	.w4(32'hbb088e3f),
	.w5(32'h3980c274),
	.w6(32'hbb58be98),
	.w7(32'hbbfd62fe),
	.w8(32'hbbab2d18),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a057c59),
	.w1(32'hbb4b28a7),
	.w2(32'h3bc3b0f3),
	.w3(32'h3a712196),
	.w4(32'hbb94b010),
	.w5(32'h379591c0),
	.w6(32'hbc315613),
	.w7(32'hbb9a90f8),
	.w8(32'hbbdf8dab),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89b898),
	.w1(32'hbaf43ca3),
	.w2(32'hba364118),
	.w3(32'h3b07fcd6),
	.w4(32'hbbe3514e),
	.w5(32'h3c06523c),
	.w6(32'hbafd9f69),
	.w7(32'hbb924dce),
	.w8(32'h3b2e2ac6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb988532),
	.w1(32'h3c23ba4d),
	.w2(32'h3c46b3c0),
	.w3(32'h37c65a6d),
	.w4(32'h3ca60790),
	.w5(32'h3cb0208d),
	.w6(32'hba4b758b),
	.w7(32'h3c8e1dfe),
	.w8(32'h3c903929),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cc7e7),
	.w1(32'hbb528c6c),
	.w2(32'h3bb86986),
	.w3(32'h3b8eff61),
	.w4(32'h3ba93078),
	.w5(32'hb91fd39c),
	.w6(32'h3b3dc80b),
	.w7(32'hbb6f368c),
	.w8(32'h3abf5a7b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb14af4),
	.w1(32'h3c35edff),
	.w2(32'h3bce8529),
	.w3(32'h3c3210fc),
	.w4(32'h3bcb3fc5),
	.w5(32'h3c857c3b),
	.w6(32'h3c57db70),
	.w7(32'hbb274212),
	.w8(32'h3bd344ca),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57968c),
	.w1(32'hbb587f13),
	.w2(32'hbb1b5c17),
	.w3(32'hbb113332),
	.w4(32'h39c90d37),
	.w5(32'hbbc7e4d8),
	.w6(32'h3bd4b07c),
	.w7(32'hbb8efa7f),
	.w8(32'hbb810c3e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f77b4),
	.w1(32'hbaf67fc7),
	.w2(32'h3b01cdc6),
	.w3(32'hbb3afaed),
	.w4(32'hbba142f9),
	.w5(32'h3c2c3734),
	.w6(32'hbb059a7d),
	.w7(32'hbb6f24bf),
	.w8(32'h3b97fe54),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e7179),
	.w1(32'h39979c27),
	.w2(32'hbb970fd6),
	.w3(32'hbb6280c6),
	.w4(32'hba4b3193),
	.w5(32'hbb15a6f0),
	.w6(32'hba81bb84),
	.w7(32'hba3cd7ac),
	.w8(32'hbc1bce8b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaad9bc),
	.w1(32'hbb35984d),
	.w2(32'h3b3fbda0),
	.w3(32'h3badc19a),
	.w4(32'hb9f0631f),
	.w5(32'h3c2129d3),
	.w6(32'hb98ef673),
	.w7(32'h38b69aa1),
	.w8(32'h3b3867a5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea7a1b),
	.w1(32'hb8a7c2b4),
	.w2(32'hba8f398e),
	.w3(32'h3b1db2ee),
	.w4(32'hba90cfc2),
	.w5(32'hba115370),
	.w6(32'h3b5a09a4),
	.w7(32'hbc426781),
	.w8(32'hbbc10f7e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b064f92),
	.w1(32'hbbaa2888),
	.w2(32'hba9102c3),
	.w3(32'hba62a07d),
	.w4(32'hbae05370),
	.w5(32'h3b55e3d4),
	.w6(32'h3a567210),
	.w7(32'hbb1e3a95),
	.w8(32'h3b56ae83),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47159a),
	.w1(32'h3b38c3d9),
	.w2(32'hbb0542ad),
	.w3(32'h3b5c2536),
	.w4(32'h3ac0da4f),
	.w5(32'h3b5276df),
	.w6(32'h3bb1c3eb),
	.w7(32'hb97175d4),
	.w8(32'h36fa6eae),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb211170),
	.w1(32'hbb8676eb),
	.w2(32'hbbf07f96),
	.w3(32'hbb98e87d),
	.w4(32'hbba5f6a6),
	.w5(32'hbb591cab),
	.w6(32'hbc117225),
	.w7(32'hbbd5f099),
	.w8(32'hbb034a80),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b05698),
	.w1(32'hba86d097),
	.w2(32'h3afcaf99),
	.w3(32'hbb3a0aab),
	.w4(32'h3bb7fede),
	.w5(32'h3c41abff),
	.w6(32'hbb0d3850),
	.w7(32'hbb35a2b9),
	.w8(32'h3c17aecb),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab18da1),
	.w1(32'h3af66430),
	.w2(32'h3a6f46cf),
	.w3(32'h3b87c17d),
	.w4(32'h3993233f),
	.w5(32'hbbcb6955),
	.w6(32'h3c0c111a),
	.w7(32'hbab03adb),
	.w8(32'h3a0ca72b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bbb97),
	.w1(32'hb8c60693),
	.w2(32'h3bcefc21),
	.w3(32'hbabba44a),
	.w4(32'h3b9fe8da),
	.w5(32'h3bb6be6c),
	.w6(32'hbb8a83c0),
	.w7(32'h3ba5b149),
	.w8(32'hba24d7ba),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4edbda),
	.w1(32'h3a5369aa),
	.w2(32'h3a386d27),
	.w3(32'h3b8d5602),
	.w4(32'h3a804d5d),
	.w5(32'h3c5c81b9),
	.w6(32'h3ba305a8),
	.w7(32'hb8c59a78),
	.w8(32'h3c579359),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7546e6),
	.w1(32'hbc098dd4),
	.w2(32'hbb7f0ac5),
	.w3(32'hba045808),
	.w4(32'hbbe0da5e),
	.w5(32'h3b4277fc),
	.w6(32'h3b08d960),
	.w7(32'hbb224d71),
	.w8(32'hba87b45e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6260a),
	.w1(32'hbc16e6f7),
	.w2(32'hbba219b6),
	.w3(32'h3bb85326),
	.w4(32'hbbb47ee5),
	.w5(32'h3ac00c40),
	.w6(32'hbb5906e6),
	.w7(32'hbb76ea2e),
	.w8(32'hbc094afc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e704),
	.w1(32'hbc293641),
	.w2(32'hb72b5f51),
	.w3(32'h3a66d9ab),
	.w4(32'hbc61313e),
	.w5(32'h3b127a30),
	.w6(32'hbb823ea9),
	.w7(32'hbc1b6372),
	.w8(32'hbba3bbf1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96958d),
	.w1(32'hbaecae7b),
	.w2(32'hbaa47922),
	.w3(32'h3c37576f),
	.w4(32'hbb7c4fd4),
	.w5(32'h3b38a9c6),
	.w6(32'h3ba6c7e8),
	.w7(32'hbb4cee98),
	.w8(32'hbae1b3f1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b8d26),
	.w1(32'hbb8da6c2),
	.w2(32'h3b902e2e),
	.w3(32'h3a40f08c),
	.w4(32'hbbfa533d),
	.w5(32'h3aae41d1),
	.w6(32'h3aebda56),
	.w7(32'hbbf641a0),
	.w8(32'hba7f9fd3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7733f9),
	.w1(32'hbbd14faa),
	.w2(32'hbb8b6b01),
	.w3(32'h3b1021cc),
	.w4(32'hbae460b0),
	.w5(32'h38ec8336),
	.w6(32'hb99caf36),
	.w7(32'h3a2bd862),
	.w8(32'h3a9d7cf6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d43ef8),
	.w1(32'h3b05343b),
	.w2(32'h3b6176d1),
	.w3(32'hbb168f66),
	.w4(32'hbbd5a258),
	.w5(32'hbb0868d1),
	.w6(32'hbb849f84),
	.w7(32'hbb40a47b),
	.w8(32'hbb17d707),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9a287),
	.w1(32'hbb80630b),
	.w2(32'hbb199917),
	.w3(32'h3bfbb454),
	.w4(32'hbb70b036),
	.w5(32'h3a29331f),
	.w6(32'h3b07d338),
	.w7(32'hbbf03b7c),
	.w8(32'hbb53c8d3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ceb5c),
	.w1(32'h3ba69fad),
	.w2(32'hba692487),
	.w3(32'hbbabfc31),
	.w4(32'h3b55caa5),
	.w5(32'hbc247f52),
	.w6(32'hbb822abd),
	.w7(32'h3b7341b3),
	.w8(32'hbaa6fefd),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8a40b),
	.w1(32'hbb2aed89),
	.w2(32'hba6f1a38),
	.w3(32'hbb85c1ed),
	.w4(32'h3c1f145e),
	.w5(32'h3c2198a1),
	.w6(32'h3a19284e),
	.w7(32'hbbf2d9d1),
	.w8(32'hbaee360d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba293d8),
	.w1(32'h3a9921e3),
	.w2(32'hbbc7bb21),
	.w3(32'h3c0a964a),
	.w4(32'hbaeedb55),
	.w5(32'hbb9a17da),
	.w6(32'h3b9f8873),
	.w7(32'hbb8dccd5),
	.w8(32'hbbaf2630),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2e4a1),
	.w1(32'hbb92700f),
	.w2(32'h3ba41a3d),
	.w3(32'hbb1579a8),
	.w4(32'hbb9ba2a8),
	.w5(32'h3c179e37),
	.w6(32'hbb105ab3),
	.w7(32'hbb46dbc0),
	.w8(32'h3ba15166),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b732f67),
	.w1(32'hbb4d013f),
	.w2(32'hbacafa76),
	.w3(32'h3a9a5f0e),
	.w4(32'hbac6c0bf),
	.w5(32'hbb5817b9),
	.w6(32'h3aff2981),
	.w7(32'h371798e1),
	.w8(32'hbb414f12),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372ffc23),
	.w1(32'hbb12dacd),
	.w2(32'hbc06d25a),
	.w3(32'hbb5fac69),
	.w4(32'hbb140ac2),
	.w5(32'hbac01f6b),
	.w6(32'hbb51e4fa),
	.w7(32'hbb473a5c),
	.w8(32'hbbc892d6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6c48a),
	.w1(32'h3bdf64d4),
	.w2(32'h3ba87b01),
	.w3(32'h3b8303e5),
	.w4(32'hbb9b6c36),
	.w5(32'hbbf1ca16),
	.w6(32'h3b69d4b2),
	.w7(32'hbad48b09),
	.w8(32'hbbd12d9a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab22c39),
	.w1(32'h3a213d8d),
	.w2(32'hb8afcd76),
	.w3(32'hbbeecd93),
	.w4(32'h3b228652),
	.w5(32'h3b146bad),
	.w6(32'hbbeb7c64),
	.w7(32'hba9f6915),
	.w8(32'hbbb59bd6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule