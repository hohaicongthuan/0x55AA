module layer_10_featuremap_126(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376a4fe3),
	.w1(32'h36c53f67),
	.w2(32'h36d0b16b),
	.w3(32'h369ed8ad),
	.w4(32'hb590ea06),
	.w5(32'h360cb941),
	.w6(32'hb695cf3a),
	.w7(32'hb76991e8),
	.w8(32'hb696c7e0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff81ab),
	.w1(32'hb937dbac),
	.w2(32'hbaa70d7a),
	.w3(32'hbb386e42),
	.w4(32'hb939d035),
	.w5(32'hba65d476),
	.w6(32'hbb253eac),
	.w7(32'hba6761ab),
	.w8(32'hbae8c713),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362bd60f),
	.w1(32'h36209658),
	.w2(32'h364caa73),
	.w3(32'h36cabab7),
	.w4(32'h36ba54a8),
	.w5(32'h36590858),
	.w6(32'h368a91d4),
	.w7(32'h367b2efd),
	.w8(32'h368cbb4e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c5cfd),
	.w1(32'h3a75eac9),
	.w2(32'h3a1098c3),
	.w3(32'hb8e05ecf),
	.w4(32'h3a7edd37),
	.w5(32'h3898284f),
	.w6(32'h393b0ab6),
	.w7(32'h3a22d567),
	.w8(32'h39f94482),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3770eec9),
	.w1(32'hb887a199),
	.w2(32'hb9902ded),
	.w3(32'h388139b4),
	.w4(32'hb824d0c2),
	.w5(32'hb963b99b),
	.w6(32'h38c423e0),
	.w7(32'h37c705b5),
	.w8(32'hb8e76528),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368cb905),
	.w1(32'h368bc7e6),
	.w2(32'h379cae05),
	.w3(32'h3664f3de),
	.w4(32'h3750971e),
	.w5(32'h3791f4ce),
	.w6(32'hb62a39c3),
	.w7(32'hb68640b0),
	.w8(32'h352cc222),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b727dbe),
	.w1(32'hbad978ee),
	.w2(32'hbb4768d3),
	.w3(32'h3b7b5da8),
	.w4(32'hbacf81d9),
	.w5(32'hbb496bbb),
	.w6(32'h3bb46b2d),
	.w7(32'h3aa6ecc4),
	.w8(32'hbb16dd7f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb617484),
	.w1(32'hbb0a35a5),
	.w2(32'hbb8d72fe),
	.w3(32'h3b707d1e),
	.w4(32'hba8ad3af),
	.w5(32'hbb5b0a76),
	.w6(32'h3b9eb0ac),
	.w7(32'hbaa8a967),
	.w8(32'hbbbcd015),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38578d25),
	.w1(32'hb8679edf),
	.w2(32'hb974dd9f),
	.w3(32'h39e026ba),
	.w4(32'h393c72a2),
	.w5(32'h3906d314),
	.w6(32'h39e92ef0),
	.w7(32'h39bc6cbf),
	.w8(32'hb8cfc4c0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4175af),
	.w1(32'hbae11036),
	.w2(32'hbb8c0f61),
	.w3(32'h39113e7f),
	.w4(32'hba01441c),
	.w5(32'hbb098346),
	.w6(32'h3b57d028),
	.w7(32'h39aa367e),
	.w8(32'hbb3ef5db),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df543d),
	.w1(32'hb9dd1962),
	.w2(32'hba60c6ae),
	.w3(32'hb8179083),
	.w4(32'hb98d4a36),
	.w5(32'hba293c8f),
	.w6(32'hb8cd45a7),
	.w7(32'hb978f42f),
	.w8(32'hba257398),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad74a6),
	.w1(32'h3b1c794a),
	.w2(32'hbb98496c),
	.w3(32'h3bb0a332),
	.w4(32'h3aecede1),
	.w5(32'hbbb886f5),
	.w6(32'h3c162d5f),
	.w7(32'h3b60d297),
	.w8(32'hbb6dbd86),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b301c9c),
	.w1(32'hbaf9da51),
	.w2(32'hbbde276e),
	.w3(32'h3b96793e),
	.w4(32'hba2d43fa),
	.w5(32'hbb8c0fc4),
	.w6(32'h3b7a0371),
	.w7(32'hbb1554f1),
	.w8(32'hbbb64e82),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8797d36),
	.w1(32'hbb35d6b6),
	.w2(32'hbad794f0),
	.w3(32'hba2d974c),
	.w4(32'hbb427d21),
	.w5(32'hbab0b486),
	.w6(32'hb948d218),
	.w7(32'hbb2b95f9),
	.w8(32'hbabb8927),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7583f2),
	.w1(32'h3aa8b3b9),
	.w2(32'h3a8774e3),
	.w3(32'hbafd46c8),
	.w4(32'h3a82bddf),
	.w5(32'h39a44fdc),
	.w6(32'hba57840e),
	.w7(32'h3a827f50),
	.w8(32'hb9995933),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ded6e),
	.w1(32'hbb9fb0a5),
	.w2(32'hbc17b813),
	.w3(32'hbb545679),
	.w4(32'hbb29c5e4),
	.w5(32'hbba91fd2),
	.w6(32'hba7adac1),
	.w7(32'hbb6ef9ca),
	.w8(32'hbbcb05e9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3802a5bb),
	.w1(32'hb9098e7e),
	.w2(32'hb9307c00),
	.w3(32'h3917397e),
	.w4(32'h3833b8d2),
	.w5(32'hb88752de),
	.w6(32'h391dea21),
	.w7(32'hb8196ade),
	.w8(32'hb8b4cab0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24002e),
	.w1(32'hbbb8e149),
	.w2(32'hbc0c3fc0),
	.w3(32'h3b9c4ed7),
	.w4(32'hbba4b3f7),
	.w5(32'hbba7f74f),
	.w6(32'h3bc6719a),
	.w7(32'hbb2cb828),
	.w8(32'hbbccab04),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07dfa9),
	.w1(32'hbb17c00b),
	.w2(32'hbb890cc5),
	.w3(32'h3b1c348d),
	.w4(32'hbaca5740),
	.w5(32'hbb306267),
	.w6(32'h3b2adb64),
	.w7(32'hbb06f5b5),
	.w8(32'hbb854bbb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e3134e),
	.w1(32'h391280ab),
	.w2(32'hb7971e11),
	.w3(32'hb82405a0),
	.w4(32'h39647c5a),
	.w5(32'h38710717),
	.w6(32'hb898fe82),
	.w7(32'h392ef0a3),
	.w8(32'hb5e61edc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970ff31),
	.w1(32'hb741254a),
	.w2(32'hb8170ac3),
	.w3(32'h399259b2),
	.w4(32'h38e80988),
	.w5(32'h38840078),
	.w6(32'h393024ca),
	.w7(32'h393b0bb8),
	.w8(32'h391d256b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9080ae9),
	.w1(32'h3ab36873),
	.w2(32'h3a120124),
	.w3(32'hba004498),
	.w4(32'h3aa31b45),
	.w5(32'hb88c284e),
	.w6(32'hba2933d7),
	.w7(32'h3a02ee2b),
	.w8(32'hb9fd3623),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9233a0),
	.w1(32'hbc11cd08),
	.w2(32'hbc574475),
	.w3(32'hbb0d2e11),
	.w4(32'hba2823e9),
	.w5(32'hbc16570e),
	.w6(32'h3b808505),
	.w7(32'hbaa5f56a),
	.w8(32'hbbcfd7da),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60c2aa),
	.w1(32'h3a81a32d),
	.w2(32'h37308132),
	.w3(32'hbad77349),
	.w4(32'h3a604ea4),
	.w5(32'h39262a49),
	.w6(32'hb5e38332),
	.w7(32'h3a880ba9),
	.w8(32'hb9e7dc38),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22db8e),
	.w1(32'h3b6a7f36),
	.w2(32'h3b3389d1),
	.w3(32'hbb6540b9),
	.w4(32'h3b627b4b),
	.w5(32'h3a161bda),
	.w6(32'hbb9c1fcc),
	.w7(32'h3afabe76),
	.w8(32'hb64b5364),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c31458),
	.w1(32'h38f94840),
	.w2(32'h3906d93c),
	.w3(32'h394a1e3b),
	.w4(32'h39e014ce),
	.w5(32'h3a07b614),
	.w6(32'h38200b61),
	.w7(32'h39bf089c),
	.w8(32'h39cab803),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dd5bb3),
	.w1(32'h38487e1f),
	.w2(32'h384ba1a1),
	.w3(32'h368756b5),
	.w4(32'h37fe4a5a),
	.w5(32'h38001c92),
	.w6(32'hb83f4dde),
	.w7(32'hb7720f59),
	.w8(32'h378eab01),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a120191),
	.w1(32'h3ba20ac8),
	.w2(32'h3a899074),
	.w3(32'h3a6bdec4),
	.w4(32'h3ba8140f),
	.w5(32'h3b098a38),
	.w6(32'h3970e236),
	.w7(32'h3b76e8b9),
	.w8(32'hb9e44768),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28094e),
	.w1(32'h3a3b95a1),
	.w2(32'hb8e2ad0e),
	.w3(32'h392e4df8),
	.w4(32'h39d14836),
	.w5(32'h382c80e9),
	.w6(32'h35b38c62),
	.w7(32'h38009673),
	.w8(32'hb8c49fcb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ab2d4),
	.w1(32'h3bb26394),
	.w2(32'h3bcce481),
	.w3(32'hbb5df7ea),
	.w4(32'h3b8ee87a),
	.w5(32'h3bb384c8),
	.w6(32'hbb825af1),
	.w7(32'h3b0e94a2),
	.w8(32'h3b3a882a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371006be),
	.w1(32'h36ee36b7),
	.w2(32'h35cc8ef4),
	.w3(32'h3594b1ad),
	.w4(32'h363131a9),
	.w5(32'hb6a5c4e8),
	.w6(32'hb712b21e),
	.w7(32'hb653d279),
	.w8(32'hb6e17479),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3810285f),
	.w1(32'hb776a31c),
	.w2(32'hb4a6ade2),
	.w3(32'h36a2d200),
	.w4(32'hb81e3b75),
	.w5(32'hb820946d),
	.w6(32'h3780cefa),
	.w7(32'hb72b50a4),
	.w8(32'h3607fea4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38410e94),
	.w1(32'hba730158),
	.w2(32'hbae3a43c),
	.w3(32'h382d10b4),
	.w4(32'hba3f8a37),
	.w5(32'hbab499ac),
	.w6(32'h3a66d303),
	.w7(32'hb9cccccb),
	.w8(32'hbad2d779),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa69b4),
	.w1(32'h3a0a31f3),
	.w2(32'hba02ef73),
	.w3(32'hbace3111),
	.w4(32'h3a33fe60),
	.w5(32'hba62eada),
	.w6(32'hbac02c75),
	.w7(32'hb9b6e2aa),
	.w8(32'hbaa303af),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18904f),
	.w1(32'hb710ab0a),
	.w2(32'hba3ba0a9),
	.w3(32'h37ee08b6),
	.w4(32'h39463f3b),
	.w5(32'hb9a45df4),
	.w6(32'h39f0ec79),
	.w7(32'h37f77c39),
	.w8(32'hba28438e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8df1ac),
	.w1(32'h39ebc2f2),
	.w2(32'hbb19d151),
	.w3(32'h3b3b624a),
	.w4(32'h39c5088b),
	.w5(32'hbaee2708),
	.w6(32'h3b7611f8),
	.w7(32'h3ad8a908),
	.w8(32'hba8fc4f6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42358a),
	.w1(32'h3bceba9a),
	.w2(32'hbc4520bf),
	.w3(32'hbb845760),
	.w4(32'h3bc2d57f),
	.w5(32'hbc55a889),
	.w6(32'h3b0519cb),
	.w7(32'h3c20bd5d),
	.w8(32'hbbee82c6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bcea5),
	.w1(32'h3c4a63d5),
	.w2(32'h3c04d9dc),
	.w3(32'hbbd6e8a7),
	.w4(32'h3c41a7b3),
	.w5(32'h3bb9c1e6),
	.w6(32'hbba625be),
	.w7(32'h3c0e2065),
	.w8(32'h3b9298fa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1cf34),
	.w1(32'h3b9ba35a),
	.w2(32'h3b838c6f),
	.w3(32'hbbcd1cec),
	.w4(32'h3bad9543),
	.w5(32'h3bb15d02),
	.w6(32'hbb226c5c),
	.w7(32'h3bec8f19),
	.w8(32'h3bf5b52f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abfeee),
	.w1(32'h3b1f7b2c),
	.w2(32'h3ac1bad5),
	.w3(32'hba1d602c),
	.w4(32'h3b333d77),
	.w5(32'h3a8153cf),
	.w6(32'hb950392e),
	.w7(32'h3b341199),
	.w8(32'h3a5a0a47),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906fd41),
	.w1(32'h38bcd934),
	.w2(32'h38e9c017),
	.w3(32'h38995bbb),
	.w4(32'h3896b1ef),
	.w5(32'h38b79d15),
	.w6(32'h3815c292),
	.w7(32'h36b996d9),
	.w8(32'h3816369b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e504d2),
	.w1(32'h390edfe6),
	.w2(32'h388bba16),
	.w3(32'hb817ad63),
	.w4(32'h38b65864),
	.w5(32'h3854d10a),
	.w6(32'hb8644b8d),
	.w7(32'h37c97893),
	.w8(32'h365001a1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d2dad),
	.w1(32'hba1e8687),
	.w2(32'h3837866f),
	.w3(32'hb8d838f7),
	.w4(32'hb95987d4),
	.w5(32'h3a8a2ff1),
	.w6(32'h39512478),
	.w7(32'h3a0c71cd),
	.w8(32'h39ccc011),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65c356),
	.w1(32'hbb0df17c),
	.w2(32'hbb9e6759),
	.w3(32'h3b5bd1c5),
	.w4(32'h3aa89a65),
	.w5(32'hba227d72),
	.w6(32'h3b9a4325),
	.w7(32'h3add8a1f),
	.w8(32'hbb32933b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d86c5),
	.w1(32'h3b03a440),
	.w2(32'h3ac24ee9),
	.w3(32'hbb4d8e2c),
	.w4(32'h3b162ba4),
	.w5(32'h3a662290),
	.w6(32'hbb62f21f),
	.w7(32'h39fb6b25),
	.w8(32'hba1106cd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11d792),
	.w1(32'h3a2a06e8),
	.w2(32'hba036da0),
	.w3(32'hba85ccfd),
	.w4(32'h3b00ae92),
	.w5(32'hb9cadc96),
	.w6(32'hbad687e5),
	.w7(32'h3981033e),
	.w8(32'hbb3fb7e1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d50f7),
	.w1(32'hb99620e6),
	.w2(32'hbb2f5e5e),
	.w3(32'hbb659deb),
	.w4(32'h3933dbcb),
	.w5(32'hbac05a8b),
	.w6(32'hba8e4fc6),
	.w7(32'h3a705906),
	.w8(32'hba519ffa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeec984),
	.w1(32'hbb924435),
	.w2(32'hbc303ef4),
	.w3(32'h3be6421f),
	.w4(32'hbb0ca44e),
	.w5(32'hbbdf460f),
	.w6(32'h3c2ee794),
	.w7(32'h3a4ff477),
	.w8(32'hbb93b5f9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3855ddce),
	.w1(32'hb699864d),
	.w2(32'h387cb340),
	.w3(32'hb7851bd8),
	.w4(32'hb78db00d),
	.w5(32'h388a63b2),
	.w6(32'hb8702025),
	.w7(32'hb79ad177),
	.w8(32'h38174388),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39339af3),
	.w1(32'h3983a31a),
	.w2(32'h39327071),
	.w3(32'h391ee72c),
	.w4(32'h39cb25d3),
	.w5(32'h39fa3097),
	.w6(32'h3985cdeb),
	.w7(32'h39832c60),
	.w8(32'h394aeb59),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987fde0),
	.w1(32'hb9839111),
	.w2(32'hb8805aa4),
	.w3(32'hb98891e4),
	.w4(32'hb932b475),
	.w5(32'h37fde1de),
	.w6(32'hb95901e0),
	.w7(32'hb8cbd142),
	.w8(32'h38809fe3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa95754),
	.w1(32'hba8d2a55),
	.w2(32'hbb2b4bd4),
	.w3(32'h3a5ae0b7),
	.w4(32'hb81614ac),
	.w5(32'hbac0deb1),
	.w6(32'h3a017f9f),
	.w7(32'hb9649456),
	.w8(32'hbab10b35),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba934de8),
	.w1(32'hba9096e6),
	.w2(32'hbae32d7f),
	.w3(32'hba5f610a),
	.w4(32'hba6eb82d),
	.w5(32'hbaa571d8),
	.w6(32'hb9d53e14),
	.w7(32'hb9c0c4f8),
	.w8(32'hba841328),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a193cb7),
	.w1(32'hbb9b21e5),
	.w2(32'hbc04638a),
	.w3(32'h3b2ed104),
	.w4(32'hbb6c1e2c),
	.w5(32'hbbb0e8ba),
	.w6(32'h3be5dff9),
	.w7(32'hba87e405),
	.w8(32'hbbacc135),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e50a19),
	.w1(32'hb9ff8708),
	.w2(32'hba254b49),
	.w3(32'hb9067f1f),
	.w4(32'hba19629a),
	.w5(32'hba055ef7),
	.w6(32'hb8d28905),
	.w7(32'hb9e537c0),
	.w8(32'hbab66993),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c9d9d2),
	.w1(32'h39213054),
	.w2(32'hb755e64a),
	.w3(32'hb81d9cd7),
	.w4(32'h395c08cf),
	.w5(32'h38647da6),
	.w6(32'hb8b348f1),
	.w7(32'h387f9e40),
	.w8(32'h3714b56f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4ad66a8),
	.w1(32'h378791fb),
	.w2(32'hb6ba58cf),
	.w3(32'h35949825),
	.w4(32'h379ea11e),
	.w5(32'hb7d2a0ef),
	.w6(32'hb784922a),
	.w7(32'h347382a4),
	.w8(32'hb8080174),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94884b1),
	.w1(32'h38f8ad3b),
	.w2(32'h39f6d9aa),
	.w3(32'hb8bdb33b),
	.w4(32'h3880f5bc),
	.w5(32'h39d76336),
	.w6(32'hb96912e5),
	.w7(32'h38b320c2),
	.w8(32'h3a191dc7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d55928),
	.w1(32'h39eea3be),
	.w2(32'hb914197e),
	.w3(32'h38c15ea4),
	.w4(32'h39c9e42a),
	.w5(32'hb8c3e60c),
	.w6(32'hb8be307e),
	.w7(32'h39a602e6),
	.w8(32'hb71babf8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b66d3d),
	.w1(32'hb9e09397),
	.w2(32'hb90a4cb1),
	.w3(32'hb81788a3),
	.w4(32'hb992e784),
	.w5(32'h387c38fa),
	.w6(32'h38514576),
	.w7(32'hba1774a1),
	.w8(32'hb92de32c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d2320),
	.w1(32'hbb510a3a),
	.w2(32'hbb8a963a),
	.w3(32'h3b16c8d2),
	.w4(32'hbb194bd4),
	.w5(32'hbb602d0f),
	.w6(32'h3afecc5e),
	.w7(32'hbb0ff624),
	.w8(32'hbb769ae5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c7e2f),
	.w1(32'hbb459477),
	.w2(32'hbb811cba),
	.w3(32'hb9b47723),
	.w4(32'h3a717b29),
	.w5(32'hbaac9ace),
	.w6(32'h3a8d0a23),
	.w7(32'hb9114d9b),
	.w8(32'hbb1cbeb0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb780d60e),
	.w1(32'hb6b640ce),
	.w2(32'h36a19168),
	.w3(32'hb8632d1a),
	.w4(32'hb82a920f),
	.w5(32'h36f9df58),
	.w6(32'hb89a011c),
	.w7(32'hb8811af9),
	.w8(32'hb7ab06b0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3704d4f3),
	.w1(32'h37ccd679),
	.w2(32'h38361a36),
	.w3(32'h369a11bc),
	.w4(32'h37e06535),
	.w5(32'h3849f348),
	.w6(32'hb6751808),
	.w7(32'h37960e13),
	.w8(32'h3833ecba),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84aa484),
	.w1(32'hb8202fd7),
	.w2(32'hb7df7e12),
	.w3(32'hb8986fa3),
	.w4(32'hb83bd485),
	.w5(32'hb835bc24),
	.w6(32'hb8735563),
	.w7(32'hb827cfa4),
	.w8(32'hb7a5a178),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5d394fc),
	.w1(32'h3707f131),
	.w2(32'h37cf9bac),
	.w3(32'h3799a475),
	.w4(32'h36839aba),
	.w5(32'h37290e7f),
	.w6(32'hb6e72d21),
	.w7(32'hb71e95a6),
	.w8(32'h376271af),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b385f2b),
	.w1(32'hbc027a56),
	.w2(32'hbc5fbf0e),
	.w3(32'hbb64a9d0),
	.w4(32'hbc014b35),
	.w5(32'hbc0cb02b),
	.w6(32'h3bab2a56),
	.w7(32'hbb2a316d),
	.w8(32'hbc137bda),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f0fc46),
	.w1(32'hbb008943),
	.w2(32'hbbb05394),
	.w3(32'h3b7374e7),
	.w4(32'h37bc3ddd),
	.w5(32'hbba8815c),
	.w6(32'hbae656e9),
	.w7(32'hbb3d6912),
	.w8(32'hbc2a0593),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad60623),
	.w1(32'hbbc6f211),
	.w2(32'hbbf29425),
	.w3(32'hba0d45ad),
	.w4(32'hbb88b480),
	.w5(32'hbbd8b3ba),
	.w6(32'h3990f673),
	.w7(32'hbb2ade1b),
	.w8(32'hbbdbb99b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8cb97),
	.w1(32'h3bbe310b),
	.w2(32'h3bc79e46),
	.w3(32'hbb894e20),
	.w4(32'h3be04ca1),
	.w5(32'h3a00fe47),
	.w6(32'hbbad1c58),
	.w7(32'h3b253e48),
	.w8(32'h3ab84d8f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385fe908),
	.w1(32'h380d570e),
	.w2(32'h37e93394),
	.w3(32'h38bcdfd3),
	.w4(32'h380d0160),
	.w5(32'h37f603a7),
	.w6(32'h3839aef2),
	.w7(32'h37c38e75),
	.w8(32'h37edd4a0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb611b2a6),
	.w1(32'hb7379d77),
	.w2(32'h38311508),
	.w3(32'hb7a6f8d5),
	.w4(32'hb4f55356),
	.w5(32'h38636f3d),
	.w6(32'hb7ec8832),
	.w7(32'hb6bc430d),
	.w8(32'h3830817c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f14db),
	.w1(32'h3781bd47),
	.w2(32'h382dc69d),
	.w3(32'h3801d5b6),
	.w4(32'h384dcd85),
	.w5(32'h3892eb8f),
	.w6(32'hb717bc91),
	.w7(32'h366c7a71),
	.w8(32'h37f25a34),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65ebc8),
	.w1(32'hbac0c458),
	.w2(32'hbb3018ce),
	.w3(32'h3aec7d6c),
	.w4(32'hba85f445),
	.w5(32'hbadf9e99),
	.w6(32'h3aa52811),
	.w7(32'hbaaa0ef6),
	.w8(32'hbb2721b5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ca73e1),
	.w1(32'h355a2046),
	.w2(32'h3722c290),
	.w3(32'h382a088c),
	.w4(32'h36cca0c6),
	.w5(32'h37b2e385),
	.w6(32'h381d96a2),
	.w7(32'h36d69b42),
	.w8(32'h372c84e7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c57a6c),
	.w1(32'hbb52e72d),
	.w2(32'hbbb1666c),
	.w3(32'hba966284),
	.w4(32'hbb6bdfd0),
	.w5(32'hbb984d41),
	.w6(32'h3b477d3a),
	.w7(32'hb930bd1d),
	.w8(32'hbb3695bd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b898b1d),
	.w1(32'h3984dc46),
	.w2(32'hbbe2d8ac),
	.w3(32'h3bd07715),
	.w4(32'h3980636f),
	.w5(32'hbbf12e81),
	.w6(32'h3ba59c19),
	.w7(32'h3abb7d22),
	.w8(32'hbbbb0a77),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b8d46),
	.w1(32'h3b637cb8),
	.w2(32'hb9ac5b97),
	.w3(32'h3a69d381),
	.w4(32'h3b85765c),
	.w5(32'hb99ad233),
	.w6(32'hb8c1967f),
	.w7(32'h3b2661f4),
	.w8(32'hba63e39b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c71faa),
	.w1(32'hbac3d044),
	.w2(32'hbb5e5f9f),
	.w3(32'h390c832a),
	.w4(32'hbabcd8f4),
	.w5(32'hbb28505c),
	.w6(32'h3a705126),
	.w7(32'hba962f4a),
	.w8(32'hbb3850da),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f9ba9),
	.w1(32'h396dbc00),
	.w2(32'hbb69751f),
	.w3(32'hb9d3c63f),
	.w4(32'hb9b2e1ee),
	.w5(32'hbae219b9),
	.w6(32'h3ad32481),
	.w7(32'h3a88460a),
	.w8(32'hbb687e7b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61674b),
	.w1(32'hb9062d7d),
	.w2(32'hba1a4b82),
	.w3(32'hbaa4d0da),
	.w4(32'h3a0df61b),
	.w5(32'hb984d0ab),
	.w6(32'hba3bd24c),
	.w7(32'hb906e00d),
	.w8(32'hba5f93a1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fa88b),
	.w1(32'hbaf5c62e),
	.w2(32'hbb802bbf),
	.w3(32'h3adc8908),
	.w4(32'hbacf0219),
	.w5(32'hbb2b7856),
	.w6(32'h3b13a2e6),
	.w7(32'hbab60477),
	.w8(32'hbb4c24a3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ed2e71),
	.w1(32'h36f0ab92),
	.w2(32'h36158a08),
	.w3(32'h36e07cc0),
	.w4(32'h369930c7),
	.w5(32'h3412d221),
	.w6(32'h374e913c),
	.w7(32'h364b0a97),
	.w8(32'hb68487e4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38274dad),
	.w1(32'hb7d9b966),
	.w2(32'hb821d66b),
	.w3(32'h362e0fa7),
	.w4(32'hb776355d),
	.w5(32'hb82999d3),
	.w6(32'h33f966c8),
	.w7(32'hb81028e6),
	.w8(32'hb7cbb165),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f60bfb),
	.w1(32'hb525362e),
	.w2(32'hb5cbd786),
	.w3(32'hb8e41dc9),
	.w4(32'h3860374b),
	.w5(32'h375ccfd8),
	.w6(32'h37c7c0e9),
	.w7(32'h38e0b568),
	.w8(32'h3732c017),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98da828),
	.w1(32'h3a086db8),
	.w2(32'h3aadc8c3),
	.w3(32'hb975a155),
	.w4(32'h3a212aee),
	.w5(32'h3a9ae257),
	.w6(32'hb92eb751),
	.w7(32'h3a1b6a0b),
	.w8(32'h3aa296d6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02db51),
	.w1(32'h3b815cd8),
	.w2(32'h3ab36f94),
	.w3(32'hbb841ade),
	.w4(32'h3b032082),
	.w5(32'hba791b51),
	.w6(32'hbb527da1),
	.w7(32'h3a508da7),
	.w8(32'hba5813dd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a007090),
	.w1(32'h3a5b51bb),
	.w2(32'h38fc7ad1),
	.w3(32'h3a123e3e),
	.w4(32'h3a6a5998),
	.w5(32'hb948f658),
	.w6(32'h39b3fab3),
	.w7(32'h3a39104f),
	.w8(32'hb94e8776),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8330a4),
	.w1(32'h38877a83),
	.w2(32'hb91d9024),
	.w3(32'hbb2376ad),
	.w4(32'h3a5d0a45),
	.w5(32'hba04f3b1),
	.w6(32'hbb7372ac),
	.w7(32'hb93ebf76),
	.w8(32'hbb470173),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca2e33),
	.w1(32'hbbe8394c),
	.w2(32'hbc019ecc),
	.w3(32'hb8dea78f),
	.w4(32'hbbe87661),
	.w5(32'hbbcc83ef),
	.w6(32'h3b049b9f),
	.w7(32'hbb0dbf9e),
	.w8(32'hbb846d63),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f2b19),
	.w1(32'h3b51c9b9),
	.w2(32'h3b18576a),
	.w3(32'hbb53d2e0),
	.w4(32'h3b2215be),
	.w5(32'h3b1611b6),
	.w6(32'hba77152a),
	.w7(32'h3b8caca7),
	.w8(32'h3b63ce08),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83b03d),
	.w1(32'hbb33033b),
	.w2(32'hbc78808c),
	.w3(32'h3b20f95a),
	.w4(32'h38ad5f85),
	.w5(32'hbc2300c8),
	.w6(32'h3c0ddc51),
	.w7(32'h3b0806b7),
	.w8(32'hbc158078),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa137cc),
	.w1(32'h3ba87448),
	.w2(32'h3bc958ed),
	.w3(32'h3a254256),
	.w4(32'h3b98b22b),
	.w5(32'h3bb4b78f),
	.w6(32'h3975ae64),
	.w7(32'h3b8c47e6),
	.w8(32'h3ba11087),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26301a),
	.w1(32'hbb2de650),
	.w2(32'hbbd4e747),
	.w3(32'hb9b08f81),
	.w4(32'hbaf1cf56),
	.w5(32'hbb75c5ee),
	.w6(32'h3a43b87a),
	.w7(32'hbb27b3e4),
	.w8(32'hbbe18705),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e809c),
	.w1(32'hbae24555),
	.w2(32'hbb0a6cdf),
	.w3(32'hbb332f42),
	.w4(32'hbae0cd13),
	.w5(32'hbb0c7852),
	.w6(32'hbb13627f),
	.w7(32'hb979becf),
	.w8(32'hbb3f9eea),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebdd6a),
	.w1(32'h3bb184a8),
	.w2(32'h3b8ecc7a),
	.w3(32'hbaf63288),
	.w4(32'h3b9495dc),
	.w5(32'h3b768b10),
	.w6(32'hba97dc7c),
	.w7(32'h3b831903),
	.w8(32'h3ac838bc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e2a0c),
	.w1(32'h355cb5a3),
	.w2(32'h3935e839),
	.w3(32'hb82fcef1),
	.w4(32'h38ca865e),
	.w5(32'h39384e1a),
	.w6(32'hb98464ca),
	.w7(32'hb92cfd88),
	.w8(32'hb867d7b5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b6c29),
	.w1(32'hbb33bbfb),
	.w2(32'hbb93e836),
	.w3(32'h39e9344b),
	.w4(32'hbacecb2b),
	.w5(32'hbb281a79),
	.w6(32'h3b1513cc),
	.w7(32'hba843ad7),
	.w8(32'hbb6925e7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58700a),
	.w1(32'hbb849b2b),
	.w2(32'hbc085b0c),
	.w3(32'hbb432af6),
	.w4(32'hbb833408),
	.w5(32'hbbf621b3),
	.w6(32'h3bb464eb),
	.w7(32'h3a13b461),
	.w8(32'hbb702948),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb729b6a),
	.w1(32'hbb296642),
	.w2(32'hbc3d00d3),
	.w3(32'h3b66e030),
	.w4(32'h3bce0a4c),
	.w5(32'hbc63223a),
	.w6(32'h3acb272e),
	.w7(32'h3b3bbefe),
	.w8(32'hbbf6b590),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dc2af),
	.w1(32'h3c19aa2c),
	.w2(32'h3b9e4fa0),
	.w3(32'hbbcebada),
	.w4(32'h3c25bd3b),
	.w5(32'h3bf4a6e9),
	.w6(32'hbb4f7275),
	.w7(32'h3c2f4895),
	.w8(32'h3bf6dca0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfb832),
	.w1(32'h3b631099),
	.w2(32'h3b55743f),
	.w3(32'hbb1d1a04),
	.w4(32'h3b71d2eb),
	.w5(32'h3b30a96a),
	.w6(32'hbb5cf8b6),
	.w7(32'h3b202273),
	.w8(32'h3a60c1ee),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2da6dd),
	.w1(32'hbb509291),
	.w2(32'hbc3b0f1f),
	.w3(32'hbb556a6e),
	.w4(32'hba9a5151),
	.w5(32'hbc0e47b6),
	.w6(32'h3b86a31a),
	.w7(32'h3b0676fa),
	.w8(32'hbbb9d115),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98723e1),
	.w1(32'hb9185cdc),
	.w2(32'h37f24cd1),
	.w3(32'h378a1ac8),
	.w4(32'h3984a353),
	.w5(32'h3a0287ef),
	.w6(32'h38cc5427),
	.w7(32'h3901ac3b),
	.w8(32'h38fa5372),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95741a8),
	.w1(32'h38b0baf2),
	.w2(32'hbc1758d3),
	.w3(32'hb9bf55da),
	.w4(32'h3a8db755),
	.w5(32'hbbffae98),
	.w6(32'h3a702050),
	.w7(32'h3bb2367f),
	.w8(32'hbba256d9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ca518),
	.w1(32'h3bdabd8d),
	.w2(32'hbaf0267a),
	.w3(32'h3bfaebc4),
	.w4(32'h3bba974f),
	.w5(32'hbaa52ac0),
	.w6(32'h3c35ef8e),
	.w7(32'h3baa1336),
	.w8(32'hb9a3e7a9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68806af),
	.w1(32'h38c12661),
	.w2(32'hb80a7168),
	.w3(32'hb85d51e0),
	.w4(32'h3901fa31),
	.w5(32'h36c2789c),
	.w6(32'hb866a621),
	.w7(32'h38cc41d6),
	.w8(32'h3796abce),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ab60f),
	.w1(32'hba4488a1),
	.w2(32'hbb0cffa8),
	.w3(32'hb8eb49a2),
	.w4(32'hb918c7cd),
	.w5(32'hbb1c4f38),
	.w6(32'hba9a59dd),
	.w7(32'hba5af168),
	.w8(32'hbac92ca3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a820956),
	.w1(32'h3a0cc7cc),
	.w2(32'hbb2b898a),
	.w3(32'h3b57e865),
	.w4(32'h3b4c5c2d),
	.w5(32'h3971bf88),
	.w6(32'h3b8cb965),
	.w7(32'h3b2427fc),
	.w8(32'hba5162b1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92f917),
	.w1(32'h3b8281a0),
	.w2(32'h3b6e49d5),
	.w3(32'hba7abaaa),
	.w4(32'h3b8089a8),
	.w5(32'h3b490798),
	.w6(32'hbab543e5),
	.w7(32'h3b2945a1),
	.w8(32'h3afd5d79),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb763864),
	.w1(32'h3a5d938e),
	.w2(32'h3b43d6db),
	.w3(32'hbb1c6bee),
	.w4(32'h3ab1a3a4),
	.w5(32'h3b928f1f),
	.w6(32'hb90ab2bf),
	.w7(32'h3b72f232),
	.w8(32'h3bb38eab),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabff3bd),
	.w1(32'h3a5de778),
	.w2(32'h3990802d),
	.w3(32'hba23f822),
	.w4(32'h3aa6cde5),
	.w5(32'h3a1c84a7),
	.w6(32'hba3f606a),
	.w7(32'h3a4fddc3),
	.w8(32'hba98c3bf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987b05b),
	.w1(32'h3aa8f1c2),
	.w2(32'hbab7db82),
	.w3(32'h3b172962),
	.w4(32'h3b57bc7a),
	.w5(32'hbb39baf5),
	.w6(32'hb8e6e580),
	.w7(32'h3b289f16),
	.w8(32'hbb4ad5f6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec9930),
	.w1(32'hbbc32002),
	.w2(32'hbc0457ca),
	.w3(32'hbb413c3e),
	.w4(32'hbb625876),
	.w5(32'hbba63f23),
	.w6(32'hbab0edbc),
	.w7(32'hbb8e3c89),
	.w8(32'hbbd08e36),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988b411),
	.w1(32'h3a839650),
	.w2(32'h3a2790d5),
	.w3(32'hb9f28521),
	.w4(32'h3a96ee0d),
	.w5(32'h3a281d5c),
	.w6(32'hb98b89e9),
	.w7(32'h3a88106c),
	.w8(32'h391294e7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3841ac2e),
	.w1(32'h378bda98),
	.w2(32'h37611c52),
	.w3(32'h383ed598),
	.w4(32'h38425cdb),
	.w5(32'h37e314c6),
	.w6(32'h36a9cc72),
	.w7(32'hb78e548d),
	.w8(32'h37a9949a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fbad8b),
	.w1(32'hb9dec9ab),
	.w2(32'hbab1d929),
	.w3(32'hb95b8492),
	.w4(32'hb9ae269b),
	.w5(32'hba94c5c1),
	.w6(32'hb951b04c),
	.w7(32'hba4a21ac),
	.w8(32'hba8f6174),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f68f62),
	.w1(32'h364db880),
	.w2(32'h37b2d198),
	.w3(32'hb7a68494),
	.w4(32'hb80793e0),
	.w5(32'h37bf1946),
	.w6(32'hb66b4150),
	.w7(32'hb7382d82),
	.w8(32'h3792f75f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf0d88),
	.w1(32'hb7ee127a),
	.w2(32'hb94cae0b),
	.w3(32'hb82d0e9f),
	.w4(32'hb8a9c0eb),
	.w5(32'hb8fcffa0),
	.w6(32'hb8d93385),
	.w7(32'hb814218c),
	.w8(32'h390f37ff),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a502f),
	.w1(32'h3a93760a),
	.w2(32'h3a53ea11),
	.w3(32'hba9137be),
	.w4(32'h3abc05ab),
	.w5(32'h3a0eca6c),
	.w6(32'hba959996),
	.w7(32'h399be4b0),
	.w8(32'hba4ca149),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98122af),
	.w1(32'hb99a17aa),
	.w2(32'hba4b923d),
	.w3(32'hb6b2ad94),
	.w4(32'hb949388d),
	.w5(32'hba2f101a),
	.w6(32'hb8f8b941),
	.w7(32'hb9b62c09),
	.w8(32'hba07218c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f9378),
	.w1(32'hb8eb4944),
	.w2(32'hbb499d78),
	.w3(32'h3a88c821),
	.w4(32'hba7a7866),
	.w5(32'hbaf81ce0),
	.w6(32'h3b34fb26),
	.w7(32'h3906621f),
	.w8(32'hba8eae0f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e3cb7),
	.w1(32'h3b2f6689),
	.w2(32'hb99b5030),
	.w3(32'hb8f84bf7),
	.w4(32'h3b39d737),
	.w5(32'h3a0fc599),
	.w6(32'hba4cbdce),
	.w7(32'h3b11c35d),
	.w8(32'hbad1b45b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a8fe4e),
	.w1(32'h34b7d558),
	.w2(32'hb890ed76),
	.w3(32'h38dfbcfb),
	.w4(32'hb9322416),
	.w5(32'hb8682285),
	.w6(32'h39166843),
	.w7(32'hb917a70f),
	.w8(32'h37ce38bd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7826e98),
	.w1(32'hb916ecf1),
	.w2(32'hb9398df6),
	.w3(32'h39288567),
	.w4(32'h388ce070),
	.w5(32'hb896ca46),
	.w6(32'h38e48f0b),
	.w7(32'hb7100022),
	.w8(32'hb8ed9a31),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ea9059),
	.w1(32'h3742744c),
	.w2(32'h362bf547),
	.w3(32'h3791d500),
	.w4(32'hb50837ee),
	.w5(32'h358281c6),
	.w6(32'h374836f3),
	.w7(32'hb7022d17),
	.w8(32'hb6d6b5b4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecd203),
	.w1(32'h3957a4d5),
	.w2(32'hb99dc46a),
	.w3(32'hb853ded4),
	.w4(32'h39ceb38a),
	.w5(32'hb9794fed),
	.w6(32'h398bce6d),
	.w7(32'h3a2a364d),
	.w8(32'h37b3da00),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e01f7),
	.w1(32'hbafadc4b),
	.w2(32'hbb9fb24c),
	.w3(32'h3c08311d),
	.w4(32'hbaea6a66),
	.w5(32'hbb84b522),
	.w6(32'h3b227dfd),
	.w7(32'h3a913077),
	.w8(32'hbb9fd730),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962c398),
	.w1(32'hbb2a8bad),
	.w2(32'hbb91af68),
	.w3(32'h3ab96964),
	.w4(32'hbaf52e4c),
	.w5(32'hbb1423ce),
	.w6(32'h3b6a798a),
	.w7(32'hba28693c),
	.w8(32'hbb57e305),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55ff28),
	.w1(32'hb94960e2),
	.w2(32'hba90b62d),
	.w3(32'h39968374),
	.w4(32'hb979a439),
	.w5(32'hba46f65b),
	.w6(32'h3a859ba6),
	.w7(32'h39481a3f),
	.w8(32'hb9a2f2f2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d03b3e),
	.w1(32'hbab8616f),
	.w2(32'hbb151765),
	.w3(32'h3a57272b),
	.w4(32'hba2db9c3),
	.w5(32'hbaf8525e),
	.w6(32'h3a80cdb6),
	.w7(32'hba0a6b2d),
	.w8(32'hbb1b46ac),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc4e3b),
	.w1(32'h3a513a3b),
	.w2(32'hb96ae368),
	.w3(32'hba0bca45),
	.w4(32'h39983cc0),
	.w5(32'h39e348c4),
	.w6(32'hb921f7be),
	.w7(32'h3a40c43a),
	.w8(32'hb97d5b12),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb869e25f),
	.w1(32'hbaa0077e),
	.w2(32'hbaf862ce),
	.w3(32'h38b04c3e),
	.w4(32'hba04cbe8),
	.w5(32'hba71310d),
	.w6(32'h39cdbbf3),
	.w7(32'hba07d564),
	.w8(32'hbacd6f48),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d321f),
	.w1(32'hbb43de6b),
	.w2(32'hbb618416),
	.w3(32'hbba0bd6d),
	.w4(32'hbb00758b),
	.w5(32'hbb56eafc),
	.w6(32'hbb7a6194),
	.w7(32'hbad6e5bc),
	.w8(32'hbb6c12bd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada5db2),
	.w1(32'hbb85c8eb),
	.w2(32'hbc0c93ee),
	.w3(32'h3b02364c),
	.w4(32'hbb967d4b),
	.w5(32'hbbb908fb),
	.w6(32'h3bdb6a71),
	.w7(32'hbaa4fe0c),
	.w8(32'hbba26fc3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab176ce),
	.w1(32'h3b5ba4c5),
	.w2(32'h3b0e2f58),
	.w3(32'hbafdfb83),
	.w4(32'h3b4a1db0),
	.w5(32'h3ad54a8a),
	.w6(32'hbace71ce),
	.w7(32'h3b1b5a4e),
	.w8(32'h39d8cf25),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c166fd),
	.w1(32'hba71d364),
	.w2(32'hbb8fc9f0),
	.w3(32'h3a839ae7),
	.w4(32'hbb1a3db8),
	.w5(32'hbba94d5e),
	.w6(32'h3ad4deb1),
	.w7(32'hb951c978),
	.w8(32'hbb530618),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7aa0a2),
	.w1(32'hbb849f2b),
	.w2(32'hbb999641),
	.w3(32'h3adcc4e6),
	.w4(32'hbaf0165e),
	.w5(32'hbb7616e9),
	.w6(32'h3b9c7d17),
	.w7(32'h37b2b950),
	.w8(32'hbac50931),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85d9dd),
	.w1(32'h3b09c26c),
	.w2(32'hba431d36),
	.w3(32'h3a2cba1f),
	.w4(32'h3b4a274f),
	.w5(32'hba9661f1),
	.w6(32'hba2fb511),
	.w7(32'h3afe72aa),
	.w8(32'hbafb3dca),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0a812),
	.w1(32'hba23ac16),
	.w2(32'hbb61c3d9),
	.w3(32'h393370c7),
	.w4(32'h39f5a87a),
	.w5(32'hba93c535),
	.w6(32'h3b27d1be),
	.w7(32'h3a68453d),
	.w8(32'hbafee5b6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e842e),
	.w1(32'h39238e3f),
	.w2(32'hb9495e38),
	.w3(32'hb92ee66c),
	.w4(32'h394095ee),
	.w5(32'hb997cada),
	.w6(32'hb8f16e1f),
	.w7(32'h38a07442),
	.w8(32'hb9f61fc0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7dd7f),
	.w1(32'h3c092227),
	.w2(32'h3be6684f),
	.w3(32'hbb040428),
	.w4(32'h3bfc3909),
	.w5(32'h3bd59e37),
	.w6(32'hb831bbda),
	.w7(32'h3bf25844),
	.w8(32'h3ba6d314),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7598f),
	.w1(32'h39d480a5),
	.w2(32'hba09925f),
	.w3(32'h3880eb11),
	.w4(32'h39bd9420),
	.w5(32'hb9f9fb4b),
	.w6(32'h394d14ff),
	.w7(32'h39da82f8),
	.w8(32'hb9e99167),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3816849b),
	.w1(32'hb7a9d5cc),
	.w2(32'hb8b2c8a6),
	.w3(32'h3930bfd7),
	.w4(32'h38699009),
	.w5(32'hb82775d4),
	.w6(32'h383779f1),
	.w7(32'hb7dc17c8),
	.w8(32'hb90b4031),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848d0dc),
	.w1(32'h37adc30f),
	.w2(32'h38929027),
	.w3(32'hb853ba05),
	.w4(32'hb683c928),
	.w5(32'h3889a395),
	.w6(32'hb7b240cc),
	.w7(32'h389fe908),
	.w8(32'h38cd1aca),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b038c8c),
	.w1(32'h3b2f7967),
	.w2(32'hbaa2792e),
	.w3(32'h3b0df70d),
	.w4(32'h3b2b1356),
	.w5(32'hbaa38c44),
	.w6(32'h3b25f0e8),
	.w7(32'h3acc91b2),
	.w8(32'h3944e612),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb2678),
	.w1(32'h3b8cc094),
	.w2(32'h3a740f5a),
	.w3(32'hbae8ab2a),
	.w4(32'h3b53215a),
	.w5(32'h39d3afe8),
	.w6(32'hba49904a),
	.w7(32'h3b54439f),
	.w8(32'hba0559f3),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28c531),
	.w1(32'hb984d559),
	.w2(32'hbb95e237),
	.w3(32'h3b83a6c0),
	.w4(32'h3a6651e5),
	.w5(32'hbb576570),
	.w6(32'h3b777623),
	.w7(32'hb914a40a),
	.w8(32'hbb6d0a36),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3711ab65),
	.w1(32'h363f138c),
	.w2(32'h37aff0fd),
	.w3(32'h3647faf9),
	.w4(32'h35f8ba79),
	.w5(32'h37d3b7c0),
	.w6(32'hb777a59e),
	.w7(32'hb7d04e0d),
	.w8(32'h37156cf9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392cb58e),
	.w1(32'hbb107bba),
	.w2(32'hbb85611b),
	.w3(32'hbaee938a),
	.w4(32'hbab0064b),
	.w5(32'hbaffdea5),
	.w6(32'h3aed4b55),
	.w7(32'hb8ef0932),
	.w8(32'hbb1774ce),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f87f1),
	.w1(32'h3a6f48ed),
	.w2(32'h39dbef3d),
	.w3(32'hba3e800d),
	.w4(32'h3ab065b1),
	.w5(32'h3a938de3),
	.w6(32'h396f0c94),
	.w7(32'h3ad020f5),
	.w8(32'h3a4bb390),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b409527),
	.w1(32'hbb0c299a),
	.w2(32'hbc128637),
	.w3(32'h3afdffee),
	.w4(32'hbac350d9),
	.w5(32'hbbb01807),
	.w6(32'h3b8bce4d),
	.w7(32'hb9a1e584),
	.w8(32'hbb65f79a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacf230),
	.w1(32'h3a87278e),
	.w2(32'h3abc87f9),
	.w3(32'hbae18d04),
	.w4(32'h3b50cc9b),
	.w5(32'h3b57537c),
	.w6(32'hbad227cb),
	.w7(32'h3b2be243),
	.w8(32'h38fc6959),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3117a),
	.w1(32'hba7c7be0),
	.w2(32'hbae71b80),
	.w3(32'hbad66fa5),
	.w4(32'hb996b353),
	.w5(32'hbaa472d1),
	.w6(32'hba9f1e7c),
	.w7(32'hba1f70f8),
	.w8(32'hbab0cad4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad64ca),
	.w1(32'h39831cab),
	.w2(32'h377a1185),
	.w3(32'hb94b4706),
	.w4(32'h3926e7c4),
	.w5(32'h38e150a0),
	.w6(32'hb9629c60),
	.w7(32'h39036fb2),
	.w8(32'h3812e131),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dc2ce),
	.w1(32'h3b3ea88a),
	.w2(32'h3b33b419),
	.w3(32'hbafd4453),
	.w4(32'h3b395e59),
	.w5(32'h3b118431),
	.w6(32'hbb146c60),
	.w7(32'h3ac9dfb6),
	.w8(32'h3aa20b82),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40946d),
	.w1(32'h39ff2dcc),
	.w2(32'hba517c67),
	.w3(32'hbb94d655),
	.w4(32'hb9523b5d),
	.w5(32'hba5559d4),
	.w6(32'hbb6731f7),
	.w7(32'hb994cb91),
	.w8(32'hba8f7c7b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf5153),
	.w1(32'h3b29eefc),
	.w2(32'h3ac93abe),
	.w3(32'hba906671),
	.w4(32'h3b12595f),
	.w5(32'h3ad1a193),
	.w6(32'hba58652e),
	.w7(32'h3b0c63a8),
	.w8(32'h3a9fca8c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1aec9a),
	.w1(32'hba4f1e07),
	.w2(32'hbb1754db),
	.w3(32'h38eaed22),
	.w4(32'hba9fbbe1),
	.w5(32'hbaf3b7fb),
	.w6(32'h3a3d4ec0),
	.w7(32'hba146c0a),
	.w8(32'hba9d73ff),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8a4e9),
	.w1(32'hb969c06a),
	.w2(32'hb9a6584b),
	.w3(32'hb9b85c7f),
	.w4(32'hb96682ce),
	.w5(32'hb9c6b666),
	.w6(32'hb9877ce4),
	.w7(32'hb9ab6910),
	.w8(32'hb9ae63e5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aced30d),
	.w1(32'hbaaeb34c),
	.w2(32'hbb4a9541),
	.w3(32'h3af6d00d),
	.w4(32'h3a2eb9b3),
	.w5(32'hbaaf6b1d),
	.w6(32'h3b4ce35f),
	.w7(32'h3a57f8fc),
	.w8(32'hbb0c56df),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f4a87),
	.w1(32'h3a622b28),
	.w2(32'hb9771851),
	.w3(32'h3a2f2e6c),
	.w4(32'h39dad25c),
	.w5(32'hb80449f8),
	.w6(32'h3aacd4b8),
	.w7(32'h3a5e6c12),
	.w8(32'h39fe950b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1de827),
	.w1(32'h3a787149),
	.w2(32'h3aebcf8b),
	.w3(32'hba5c5076),
	.w4(32'h3a833ab8),
	.w5(32'h3ae10805),
	.w6(32'hbaf4cb90),
	.w7(32'hb9aa72aa),
	.w8(32'hba197f32),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8693c),
	.w1(32'hb882a959),
	.w2(32'hb95b45b7),
	.w3(32'h394db4da),
	.w4(32'hb87430b2),
	.w5(32'hb9746411),
	.w6(32'h396332fe),
	.w7(32'h3825bcd5),
	.w8(32'hb92130e6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56108f),
	.w1(32'h3ad8411f),
	.w2(32'h396fb622),
	.w3(32'h3b9a3329),
	.w4(32'hb995c0d0),
	.w5(32'hbab85abb),
	.w6(32'h3b86514d),
	.w7(32'h393f4716),
	.w8(32'hba8d17d1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37077f47),
	.w1(32'h37ada7b4),
	.w2(32'h372c346e),
	.w3(32'h36d7b30c),
	.w4(32'h375e8924),
	.w5(32'hb6d793a8),
	.w6(32'hb73f98cb),
	.w7(32'hb7c6609c),
	.w8(32'hb821ab32),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9377461),
	.w1(32'hb9a7fc95),
	.w2(32'hb9c031d7),
	.w3(32'hb8b43337),
	.w4(32'hb97e8564),
	.w5(32'hb9c299c7),
	.w6(32'hb8473308),
	.w7(32'hb9576a6a),
	.w8(32'hb96cc398),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f9c84),
	.w1(32'h3adace52),
	.w2(32'h3acc44e1),
	.w3(32'hbb6f33c7),
	.w4(32'h3afb6706),
	.w5(32'h3b0ba0e6),
	.w6(32'hbb5d789f),
	.w7(32'h3a93d480),
	.w8(32'h39b09161),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a085ed1),
	.w1(32'h3b28e588),
	.w2(32'hbb33a2de),
	.w3(32'h3b5b23eb),
	.w4(32'h3b90fb9c),
	.w5(32'h371d10cd),
	.w6(32'h3b8957c9),
	.w7(32'h3b82b132),
	.w8(32'hbad1c8ea),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5779e4),
	.w1(32'h3a2ac8d3),
	.w2(32'hba355a85),
	.w3(32'h3a5ed1a2),
	.w4(32'h3a41cbca),
	.w5(32'hba1005b3),
	.w6(32'h3a0e6d5d),
	.w7(32'h3a528aa7),
	.w8(32'hba08928e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fe94f),
	.w1(32'h3aca1356),
	.w2(32'h3aca16f9),
	.w3(32'hbaf3aabd),
	.w4(32'h3ae2ae81),
	.w5(32'h3ab53251),
	.w6(32'hbb1d9aa5),
	.w7(32'h3a4f8771),
	.w8(32'hb89b6ff0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a830a0f),
	.w1(32'h3a858302),
	.w2(32'hb9e3c89d),
	.w3(32'h39718dca),
	.w4(32'h3a7b1174),
	.w5(32'h3a6332ce),
	.w6(32'h3a02c17c),
	.w7(32'h3a7b264e),
	.w8(32'h3a1fcb82),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac465e),
	.w1(32'hbb1254a3),
	.w2(32'hbbeaa326),
	.w3(32'h3ac9d84e),
	.w4(32'hba8d9fa4),
	.w5(32'hbb9d47cc),
	.w6(32'h3b0e4767),
	.w7(32'hba3fbf37),
	.w8(32'hbb9b861d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a710f93),
	.w1(32'hba8f6079),
	.w2(32'hbb88c221),
	.w3(32'h39bb9e8c),
	.w4(32'hbacb0053),
	.w5(32'hbb588916),
	.w6(32'h3ab0b524),
	.w7(32'hb98993fe),
	.w8(32'hbb1a0679),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba483e06),
	.w1(32'hbb7d5e59),
	.w2(32'hbb81ce5a),
	.w3(32'hba320ad1),
	.w4(32'hbb551a3a),
	.w5(32'hbb196be2),
	.w6(32'h39e3d3b4),
	.w7(32'hbb347106),
	.w8(32'hbb82d05f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a27c0),
	.w1(32'hb8a93422),
	.w2(32'h387ceb3d),
	.w3(32'h383b702d),
	.w4(32'hb904a56b),
	.w5(32'h388b9b3c),
	.w6(32'h3864f952),
	.w7(32'hb819d774),
	.w8(32'h37ce1f9b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90b719),
	.w1(32'hbad01462),
	.w2(32'hbb41ba07),
	.w3(32'hbb37fb42),
	.w4(32'hbadc352a),
	.w5(32'hbb09343f),
	.w6(32'hba94d5ff),
	.w7(32'hbafb7ba5),
	.w8(32'hbb6544b6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3829944c),
	.w1(32'h37520bea),
	.w2(32'h37d79eb3),
	.w3(32'h3824b5a0),
	.w4(32'h36e117db),
	.w5(32'h377ea131),
	.w6(32'h37b02332),
	.w7(32'h36012599),
	.w8(32'h37992158),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d96bf),
	.w1(32'hba2810c1),
	.w2(32'hba4164e6),
	.w3(32'hb9484597),
	.w4(32'hb9038437),
	.w5(32'hba876aa0),
	.w6(32'h3924c2a3),
	.w7(32'hb9c40b5d),
	.w8(32'hb9e78dff),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b6a95),
	.w1(32'h37d958c3),
	.w2(32'h3887c269),
	.w3(32'hb9b736a9),
	.w4(32'hb91a3b37),
	.w5(32'hb96e9cfb),
	.w6(32'hb9e28e52),
	.w7(32'hb88fad75),
	.w8(32'hba03f2db),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f7ff9),
	.w1(32'hbb164024),
	.w2(32'hbbb136ca),
	.w3(32'hba91dff7),
	.w4(32'hbad70f1d),
	.w5(32'hbb5860f8),
	.w6(32'h39e7dbdc),
	.w7(32'hba72fe31),
	.w8(32'hbb70aad8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71df7e2),
	.w1(32'hb61715fa),
	.w2(32'hb5475205),
	.w3(32'hb7709460),
	.w4(32'h34f31c48),
	.w5(32'hb638ffaa),
	.w6(32'hb7aa99e1),
	.w7(32'hb795ea2a),
	.w8(32'hb70f790c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b9713e),
	.w1(32'h37fc685d),
	.w2(32'h383b52a6),
	.w3(32'hb5e9e9f3),
	.w4(32'h358003d1),
	.w5(32'h354825ce),
	.w6(32'hb6e9f2a6),
	.w7(32'hb817921b),
	.w8(32'hb8b20d5b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c70b52),
	.w1(32'h3916a1bc),
	.w2(32'h39c2568e),
	.w3(32'hba22dc62),
	.w4(32'h39b69e2f),
	.w5(32'h3815818e),
	.w6(32'hbaa6b5eb),
	.w7(32'h39328fdb),
	.w8(32'h390d36ea),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab87032),
	.w1(32'hbb94a74a),
	.w2(32'hbc113c2b),
	.w3(32'hba9494f8),
	.w4(32'hbb8722fe),
	.w5(32'hbbea5e01),
	.w6(32'h3a806032),
	.w7(32'hbb76558a),
	.w8(32'hbbbe63ce),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaf141),
	.w1(32'h3b432b4f),
	.w2(32'hbb8b1087),
	.w3(32'hbb1c6eec),
	.w4(32'h3b40f98c),
	.w5(32'hbb6b0964),
	.w6(32'h3a38f427),
	.w7(32'h3b887c47),
	.w8(32'hbaa64ae4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be5da6),
	.w1(32'hba53c5b1),
	.w2(32'hb9ee4405),
	.w3(32'hb99c1f6b),
	.w4(32'hb953f262),
	.w5(32'hba275809),
	.w6(32'hb9538a89),
	.w7(32'hb900836d),
	.w8(32'hb9c0b56a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b59ab),
	.w1(32'hbc037916),
	.w2(32'hbc2b88e7),
	.w3(32'h3bf07ec2),
	.w4(32'hbbbdb97c),
	.w5(32'hbc19749b),
	.w6(32'h3b31700a),
	.w7(32'hbc368d45),
	.w8(32'hbc676587),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa64e),
	.w1(32'h3b51d48a),
	.w2(32'hbaedd676),
	.w3(32'hbbfc07b3),
	.w4(32'h3b4290b5),
	.w5(32'h3aaa4da6),
	.w6(32'hbb909454),
	.w7(32'h3b1ff0b5),
	.w8(32'hba87aaff),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac844f5),
	.w1(32'h3a364aff),
	.w2(32'hbb0a308c),
	.w3(32'h398308bc),
	.w4(32'h38b78759),
	.w5(32'hbad862b5),
	.w6(32'h3a8918cc),
	.w7(32'h3aa83afc),
	.w8(32'hba8c2495),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3714faf7),
	.w1(32'hb872487b),
	.w2(32'hb7fd6e9f),
	.w3(32'hb76ddf43),
	.w4(32'hb75db526),
	.w5(32'hb78792f6),
	.w6(32'hb7a8fbdb),
	.w7(32'hb8416698),
	.w8(32'hb7f07825),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77531a8),
	.w1(32'hb800a236),
	.w2(32'hb82ea8c7),
	.w3(32'hb88ca69a),
	.w4(32'hb842d843),
	.w5(32'h3805094c),
	.w6(32'hb83d397a),
	.w7(32'hb7f4885e),
	.w8(32'h37cf5dd0),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cc0b69),
	.w1(32'hb6c33453),
	.w2(32'h36d989ea),
	.w3(32'h36c4eb20),
	.w4(32'hb67d948e),
	.w5(32'h36fa8820),
	.w6(32'h37500ddd),
	.w7(32'hb4f3da9e),
	.w8(32'h3734b9f0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ed19f),
	.w1(32'h3a947485),
	.w2(32'hbaf91c31),
	.w3(32'h3ab14be0),
	.w4(32'h3aba421c),
	.w5(32'hba924d2d),
	.w6(32'h3b63a7f7),
	.w7(32'h3b33168f),
	.w8(32'h391f471c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3973e0),
	.w1(32'hb9d4c65d),
	.w2(32'hbb11f9b9),
	.w3(32'hb99361b4),
	.w4(32'h3980bc1e),
	.w5(32'hba83bfc1),
	.w6(32'h3a755796),
	.w7(32'h3b033674),
	.w8(32'hba776c69),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39987813),
	.w1(32'h3b3c13f1),
	.w2(32'hb9877e2d),
	.w3(32'hb92f7780),
	.w4(32'h3b6783bd),
	.w5(32'hba04ee0d),
	.w6(32'hbae60512),
	.w7(32'h3ae45c53),
	.w8(32'hbad52bda),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e4b97),
	.w1(32'h3a12fefa),
	.w2(32'h39d317e6),
	.w3(32'h38345ff5),
	.w4(32'h3a55ed39),
	.w5(32'h3a1f67c2),
	.w6(32'hb99c906f),
	.w7(32'h3a014d41),
	.w8(32'h395a60f0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35b29c),
	.w1(32'hbb104c04),
	.w2(32'hbba16808),
	.w3(32'h3b3ea913),
	.w4(32'hb83ad88c),
	.w5(32'hbb3e152e),
	.w6(32'h3b714960),
	.w7(32'hb9a67a42),
	.w8(32'hbb63e2da),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e04c4d),
	.w1(32'h3b08d73f),
	.w2(32'hbb1b53b1),
	.w3(32'h3b1b5293),
	.w4(32'h3afe4dbd),
	.w5(32'hbb2587a7),
	.w6(32'h3af73615),
	.w7(32'h3a80a5a1),
	.w8(32'hbacba379),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b16d45),
	.w1(32'h37491a5e),
	.w2(32'h380696f1),
	.w3(32'h3751a149),
	.w4(32'h37089fa0),
	.w5(32'h37c2ee12),
	.w6(32'h35dbaf93),
	.w7(32'hb622117d),
	.w8(32'h378d5f80),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cf3eb),
	.w1(32'hbb2976ed),
	.w2(32'hbb82510f),
	.w3(32'hbaff33af),
	.w4(32'hba867023),
	.w5(32'hbb07ee4a),
	.w6(32'hb9845060),
	.w7(32'hb9e8d74a),
	.w8(32'hbafe3259),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f9d02d),
	.w1(32'h3804954b),
	.w2(32'h389c7060),
	.w3(32'h36aaaf5a),
	.w4(32'h37af5a60),
	.w5(32'h38887a7b),
	.w6(32'hb78909b7),
	.w7(32'hb6b3ce15),
	.w8(32'h3832b3b5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b96b4),
	.w1(32'h3b33338b),
	.w2(32'hbb3d2df6),
	.w3(32'h3bae213c),
	.w4(32'h3a4acb17),
	.w5(32'hbab134e3),
	.w6(32'h3ba49659),
	.w7(32'h39ed466b),
	.w8(32'hbac63eb1),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa27dff),
	.w1(32'h3b7052de),
	.w2(32'h3a3d9bda),
	.w3(32'hbb379ece),
	.w4(32'h3b2c2adc),
	.w5(32'hba82bb60),
	.w6(32'hbb59269b),
	.w7(32'h3a186a06),
	.w8(32'hbb16569a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafba1bc),
	.w1(32'h3a89c412),
	.w2(32'hb8ea40b8),
	.w3(32'hbb149e9e),
	.w4(32'h3abc17a6),
	.w5(32'hb822c302),
	.w6(32'hbaddd8eb),
	.w7(32'h3a88fdd0),
	.w8(32'hb9b04239),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390712f0),
	.w1(32'h39a045f4),
	.w2(32'hba5e01d2),
	.w3(32'h39b7ba8f),
	.w4(32'h38773257),
	.w5(32'hba3109f7),
	.w6(32'h39a8e3b4),
	.w7(32'h3943d2a2),
	.w8(32'hba19880f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb234cd1),
	.w1(32'h3b1b8ba0),
	.w2(32'h3a61f618),
	.w3(32'hbb7f468b),
	.w4(32'h3b259998),
	.w5(32'h3a6befa4),
	.w6(32'hbb5caa3d),
	.w7(32'h3b0dc624),
	.w8(32'hb8120f82),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152971),
	.w1(32'hba5e8019),
	.w2(32'hbb29f169),
	.w3(32'h3ab15b3c),
	.w4(32'hba2fa846),
	.w5(32'hba885577),
	.w6(32'h3b102b35),
	.w7(32'hb9b749d5),
	.w8(32'hbb146957),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95fe29),
	.w1(32'h3a87ba53),
	.w2(32'hbb40d8f8),
	.w3(32'h3bd63adb),
	.w4(32'h3acb90c3),
	.w5(32'hbb398841),
	.w6(32'h3b97403a),
	.w7(32'h3aa61903),
	.w8(32'hbb2d31d9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380c6bc1),
	.w1(32'h3758bb1c),
	.w2(32'h37b166a4),
	.w3(32'h377e20f5),
	.w4(32'hb63b7c7a),
	.w5(32'h377d307c),
	.w6(32'h3777734e),
	.w7(32'hb70ec51d),
	.w8(32'h3741b828),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3700f6db),
	.w1(32'hb8881b50),
	.w2(32'hb8e5211f),
	.w3(32'hb84efb2c),
	.w4(32'hb8a98550),
	.w5(32'hb8ee1109),
	.w6(32'hb8427104),
	.w7(32'hb91dd7f1),
	.w8(32'hb91a858f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1651b7),
	.w1(32'h3a344026),
	.w2(32'hbb891aee),
	.w3(32'h3b4d650b),
	.w4(32'h3b27a16b),
	.w5(32'hbb873188),
	.w6(32'h3b02b375),
	.w7(32'h3a6d8823),
	.w8(32'hbbbdb059),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab765ee),
	.w1(32'hbaab68ea),
	.w2(32'hbb4d5a3a),
	.w3(32'h3a7fd8aa),
	.w4(32'h3a2283b8),
	.w5(32'hbb0645b2),
	.w6(32'h3aa74c31),
	.w7(32'h39b7ccba),
	.w8(32'hbb92bbf6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ad793),
	.w1(32'h3a6cbb06),
	.w2(32'hb8f1ae54),
	.w3(32'hbb0abb69),
	.w4(32'h3a929382),
	.w5(32'hba195000),
	.w6(32'hba69a809),
	.w7(32'h39fd24ce),
	.w8(32'hbaa92592),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b384d28),
	.w1(32'hbb23783d),
	.w2(32'hbbfa53c6),
	.w3(32'hbb1c0dbd),
	.w4(32'hbb7c6305),
	.w5(32'hbbb991a5),
	.w6(32'h3b43bf5b),
	.w7(32'hb945c0ba),
	.w8(32'hbbbb7ab3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e03baf),
	.w1(32'hb953797a),
	.w2(32'h37f90da5),
	.w3(32'h3a1bcf30),
	.w4(32'h3918e54b),
	.w5(32'h399b9a15),
	.w6(32'hb8bb9d21),
	.w7(32'h3902fefe),
	.w8(32'h3684cf46),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3970e602),
	.w1(32'hba3b0ed8),
	.w2(32'hba6e22b4),
	.w3(32'h3a81a992),
	.w4(32'hb9d4b69a),
	.w5(32'hba1391dc),
	.w6(32'h38c89207),
	.w7(32'hba4a9ce8),
	.w8(32'hba831950),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bc6f6),
	.w1(32'h3be337fe),
	.w2(32'hbbb6172d),
	.w3(32'h3bf607e6),
	.w4(32'h3c247c0e),
	.w5(32'hbb8411e7),
	.w6(32'h3bf65bbd),
	.w7(32'h3c301e6c),
	.w8(32'hbaf87488),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f64d1),
	.w1(32'hbb92732f),
	.w2(32'hbbdc8378),
	.w3(32'h3bd69326),
	.w4(32'hbb4d8c6d),
	.w5(32'hbbe878a2),
	.w6(32'h3bb96993),
	.w7(32'hbb5926b3),
	.w8(32'hbbdfe05a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05699d),
	.w1(32'hba4db5ef),
	.w2(32'hbbd391c1),
	.w3(32'h3afd12e4),
	.w4(32'h3a65cdac),
	.w5(32'hbb98e3a4),
	.w6(32'h3b908c10),
	.w7(32'h3b52409a),
	.w8(32'hbaa5b493),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d60d9),
	.w1(32'h3b573bd9),
	.w2(32'h3b5c689b),
	.w3(32'hbaaa5377),
	.w4(32'h3b352a03),
	.w5(32'h3b1edb06),
	.w6(32'hbaca1ba7),
	.w7(32'h3b1322fb),
	.w8(32'h3af2f5d7),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b6db9),
	.w1(32'h3aabcdba),
	.w2(32'h39c1f2e5),
	.w3(32'hbb7b77e4),
	.w4(32'h3abd146b),
	.w5(32'h3a51895c),
	.w6(32'hbb650ab1),
	.w7(32'hba173e24),
	.w8(32'hba27cecd),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3706eb77),
	.w1(32'h375223b0),
	.w2(32'h37779947),
	.w3(32'h37131f37),
	.w4(32'h37128c53),
	.w5(32'h36d9c383),
	.w6(32'hb65a565b),
	.w7(32'h35cc01d6),
	.w8(32'h36c11304),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d97f38),
	.w1(32'h377f3d2e),
	.w2(32'h37bb1c53),
	.w3(32'h37a86eff),
	.w4(32'h374eae27),
	.w5(32'h37c8b583),
	.w6(32'h371e08de),
	.w7(32'h344f9fa4),
	.w8(32'h37612fa6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc01eb),
	.w1(32'hb9c73ea2),
	.w2(32'hba44f22f),
	.w3(32'hb82f89e7),
	.w4(32'hba0d11d0),
	.w5(32'hba20f567),
	.w6(32'h36779358),
	.w7(32'hba2f32ec),
	.w8(32'hba7a5f20),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371ff74b),
	.w1(32'hb650185c),
	.w2(32'h37d4b6f4),
	.w3(32'h36bb4578),
	.w4(32'hb682cb57),
	.w5(32'h37987d6a),
	.w6(32'h3698dd38),
	.w7(32'hb70ab857),
	.w8(32'h37876a72),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af16895),
	.w1(32'h39863bdf),
	.w2(32'hba7a1b57),
	.w3(32'h3ab952ea),
	.w4(32'hba3bf35d),
	.w5(32'hbaa57bde),
	.w6(32'h3b132bb6),
	.w7(32'hb9d088e6),
	.w8(32'hba90130c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b66c7),
	.w1(32'hbb20b969),
	.w2(32'hbb9cde4c),
	.w3(32'h3af6b740),
	.w4(32'hbaa012d2),
	.w5(32'hbb341aa0),
	.w6(32'h3a29e121),
	.w7(32'hbb18db52),
	.w8(32'hbb9cecb6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabed6f),
	.w1(32'h3a4da4ba),
	.w2(32'hb9195c13),
	.w3(32'hba038b9d),
	.w4(32'h3a9343fc),
	.w5(32'h38a652cb),
	.w6(32'hb930fd3b),
	.w7(32'h3ae32139),
	.w8(32'h38d11575),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3835cf52),
	.w1(32'h37cde683),
	.w2(32'h3759debc),
	.w3(32'h379fe3d9),
	.w4(32'hb4c82bfc),
	.w5(32'hb689737c),
	.w6(32'h3726d8bb),
	.w7(32'h374e83e4),
	.w8(32'hb5a65866),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2bfae),
	.w1(32'hb9122486),
	.w2(32'hbc3d8e4b),
	.w3(32'h3b742487),
	.w4(32'hb710d15d),
	.w5(32'hbc028449),
	.w6(32'h3c07e4c2),
	.w7(32'h3b8be3e8),
	.w8(32'hbb8934a8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb9534),
	.w1(32'hbac8c996),
	.w2(32'hbb1d3e69),
	.w3(32'h3aef1e3b),
	.w4(32'hba1ab25f),
	.w5(32'hbaf2ad82),
	.w6(32'h3ae8313e),
	.w7(32'hba1856e0),
	.w8(32'hbb1baf74),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380bbd87),
	.w1(32'hb789985b),
	.w2(32'h37f5929c),
	.w3(32'h38235b79),
	.w4(32'h367911fb),
	.w5(32'h38d5b667),
	.w6(32'h3861b8a1),
	.w7(32'h38baae90),
	.w8(32'h38e8ea96),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b103246),
	.w1(32'hbae57e0a),
	.w2(32'hbb7cc93a),
	.w3(32'h3b5012af),
	.w4(32'hba02ce18),
	.w5(32'hbb214534),
	.w6(32'h3b81b980),
	.w7(32'h3896ca10),
	.w8(32'hbb05a35a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8125c85),
	.w1(32'hb79d3a9c),
	.w2(32'h37b96ca6),
	.w3(32'hb743df11),
	.w4(32'h38036411),
	.w5(32'h38a1a655),
	.w6(32'h381d1172),
	.w7(32'h386a66af),
	.w8(32'h389b1b9f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f1532),
	.w1(32'hb8943077),
	.w2(32'hb904f349),
	.w3(32'h39951b34),
	.w4(32'h392ef5f3),
	.w5(32'h3895d3e3),
	.w6(32'h3932c307),
	.w7(32'h38719f5f),
	.w8(32'h380ca515),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79b9f8b),
	.w1(32'hb75d9f08),
	.w2(32'h3701c72b),
	.w3(32'hb7a0a7be),
	.w4(32'h3735ba33),
	.w5(32'h3778de4f),
	.w6(32'hb70a1432),
	.w7(32'h36fc257d),
	.w8(32'h370fdded),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387737be),
	.w1(32'hb873033e),
	.w2(32'hb7916940),
	.w3(32'h37da4b59),
	.w4(32'hb8059555),
	.w5(32'h37326ff7),
	.w6(32'h37998acb),
	.w7(32'h37482788),
	.w8(32'h380562ca),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2a42a),
	.w1(32'h3aba55a5),
	.w2(32'h3a82db43),
	.w3(32'hba3a7774),
	.w4(32'h3aa7e48b),
	.w5(32'h39b9729a),
	.w6(32'hba270bd8),
	.w7(32'h3a93e612),
	.w8(32'h3a2792be),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39230ff1),
	.w1(32'hbbd1e4bf),
	.w2(32'hbbfeafd7),
	.w3(32'hbb63f8d0),
	.w4(32'hbb82ee5e),
	.w5(32'hbb7c93ff),
	.w6(32'h3b026f84),
	.w7(32'hbb14d8f7),
	.w8(32'hbb908dbe),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b029a1e),
	.w1(32'hbac37092),
	.w2(32'hbb1f285b),
	.w3(32'h3b027e2d),
	.w4(32'hb9f7dd8f),
	.w5(32'hbaa1e32a),
	.w6(32'h3b264a1d),
	.w7(32'hba52bc1b),
	.w8(32'hbb286abc),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2e004),
	.w1(32'hbb210a77),
	.w2(32'hbb8d03bd),
	.w3(32'h3a8e4f19),
	.w4(32'hbaa5ac54),
	.w5(32'hbaf6caf6),
	.w6(32'h3b7a1384),
	.w7(32'hba5c50fb),
	.w8(32'hbb5a6fb2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384770f7),
	.w1(32'h38948c32),
	.w2(32'hb8b9624d),
	.w3(32'h3802a585),
	.w4(32'h385b3595),
	.w5(32'hb899b2fb),
	.w6(32'hb777dd77),
	.w7(32'h37fc7f2a),
	.w8(32'hb8c66b2f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91df2b3),
	.w1(32'hb96c2927),
	.w2(32'hb9f1b060),
	.w3(32'hb80899ae),
	.w4(32'hb9764b5a),
	.w5(32'hb9ce7f75),
	.w6(32'h3969d757),
	.w7(32'hb91da2a2),
	.w8(32'hb9fef3d3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3727cb3b),
	.w1(32'h36e184db),
	.w2(32'h378017ef),
	.w3(32'h36ea0d55),
	.w4(32'h36e99fb5),
	.w5(32'h374c928a),
	.w6(32'h36d7b5fe),
	.w7(32'hb62a3ccd),
	.w8(32'h3723605a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378cdd00),
	.w1(32'hb78458b8),
	.w2(32'hb78d3892),
	.w3(32'h380ba72f),
	.w4(32'hb65339a7),
	.w5(32'hb74850cc),
	.w6(32'h3781ad51),
	.w7(32'hb7ee08c1),
	.w8(32'hb7d2b817),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbb7c7),
	.w1(32'hbb7805fe),
	.w2(32'hbbb3a2a7),
	.w3(32'hbaea7213),
	.w4(32'hbb252501),
	.w5(32'hbb48c0ff),
	.w6(32'hb9b9689d),
	.w7(32'hbb3c495b),
	.w8(32'hbb9a1f3a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d3d10b),
	.w1(32'h37a297be),
	.w2(32'h3853b2b4),
	.w3(32'h38916341),
	.w4(32'h3899c7d4),
	.w5(32'h38ef7af1),
	.w6(32'h3800c0fa),
	.w7(32'h381834f3),
	.w8(32'h38b8bcc1),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2f96e),
	.w1(32'h399dd777),
	.w2(32'hba82547b),
	.w3(32'h39fd894b),
	.w4(32'hb87c6481),
	.w5(32'hba6fd4a5),
	.w6(32'h3996cbe5),
	.w7(32'hb89e0c5b),
	.w8(32'hba5914db),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939d014),
	.w1(32'h39d1e7bb),
	.w2(32'hbac0a623),
	.w3(32'h397faee3),
	.w4(32'h39bb7952),
	.w5(32'hba8a1a5e),
	.w6(32'h392d2750),
	.w7(32'h39948937),
	.w8(32'hb9e9ecb9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3786f4b8),
	.w1(32'h3757698a),
	.w2(32'h3692d108),
	.w3(32'h341647f7),
	.w4(32'h379c02ee),
	.w5(32'h373fd477),
	.w6(32'hb69d6994),
	.w7(32'h37e71e26),
	.w8(32'h379e7aa4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a404668),
	.w1(32'hba349298),
	.w2(32'hbad9bc18),
	.w3(32'h3ac48165),
	.w4(32'hb90f8751),
	.w5(32'hbacf0703),
	.w6(32'h3af161fb),
	.w7(32'hb9214860),
	.w8(32'hbad56dbc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370b0263),
	.w1(32'hb97af8eb),
	.w2(32'hb9b8b78a),
	.w3(32'hb942ae44),
	.w4(32'hb9aad702),
	.w5(32'hb9711fcb),
	.w6(32'hb774a7a2),
	.w7(32'hb9c39b82),
	.w8(32'hb9d70dc0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04d0d2),
	.w1(32'hbbe5c257),
	.w2(32'hbc3e7177),
	.w3(32'hbb4c0158),
	.w4(32'hbb553c57),
	.w5(32'hbbd479d1),
	.w6(32'hb99cdea6),
	.w7(32'hbb0551f2),
	.w8(32'hbbce31ab),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912d96d),
	.w1(32'h3b16644e),
	.w2(32'h3b00914b),
	.w3(32'h388d2b92),
	.w4(32'hba442794),
	.w5(32'h3a314abb),
	.w6(32'h3abf2b08),
	.w7(32'h3af5ec48),
	.w8(32'h3a838c2e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62af7a),
	.w1(32'h3b83f8a6),
	.w2(32'h3af82172),
	.w3(32'hbadbc6b5),
	.w4(32'hbb011865),
	.w5(32'hbb24ab7f),
	.w6(32'hba5b061d),
	.w7(32'h3a5f1040),
	.w8(32'hbb108cb0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule