module layer_8_featuremap_150(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa469bc),
	.w1(32'h3b194d28),
	.w2(32'h3a6cf73c),
	.w3(32'h3ab92fc4),
	.w4(32'h3b4f9bcc),
	.w5(32'h3b023c51),
	.w6(32'h3a24ea24),
	.w7(32'h3b1b57bc),
	.w8(32'h3addde54),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79e24ac),
	.w1(32'hb8e49e0f),
	.w2(32'h3a9cda95),
	.w3(32'hbab45ccb),
	.w4(32'h3add19ad),
	.w5(32'h3ab06cfe),
	.w6(32'hba7717b0),
	.w7(32'h3a95cc18),
	.w8(32'h3aa191d1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e100d3),
	.w1(32'hba8ff30a),
	.w2(32'hbb16b25d),
	.w3(32'hb9a4f916),
	.w4(32'h3b17cad0),
	.w5(32'h3ac2b6e9),
	.w6(32'h3b16f03a),
	.w7(32'h3b05759f),
	.w8(32'h3a936f47),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4075f),
	.w1(32'hba26ae0a),
	.w2(32'hb988d3c6),
	.w3(32'hb8185a8f),
	.w4(32'hba272a02),
	.w5(32'h38c6c77e),
	.w6(32'hb9b6c5e9),
	.w7(32'h396c2182),
	.w8(32'h39a7b3e5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b824856),
	.w1(32'h3bfeb692),
	.w2(32'h3b440664),
	.w3(32'h3b6090ce),
	.w4(32'h3bc4aa50),
	.w5(32'h3b6100e9),
	.w6(32'hb85d33ef),
	.w7(32'h3b739daa),
	.w8(32'h3b2083b8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0af2b8),
	.w1(32'hbb1391aa),
	.w2(32'hba8ae8d0),
	.w3(32'h3af8c5ae),
	.w4(32'hb96856bb),
	.w5(32'h39e8acf1),
	.w6(32'h3af63f49),
	.w7(32'h3a81b367),
	.w8(32'h3b0b0cd7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920424e),
	.w1(32'hb919a0a1),
	.w2(32'hb9a682e0),
	.w3(32'h3989b9f0),
	.w4(32'hb93fffc5),
	.w5(32'hb8286a91),
	.w6(32'hb937e68c),
	.w7(32'hb9a55202),
	.w8(32'h36d67b1a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2973c1),
	.w1(32'h3a26f06b),
	.w2(32'h38997b60),
	.w3(32'h3c09f9b3),
	.w4(32'h3bf616e9),
	.w5(32'h3b3ef279),
	.w6(32'h3bc77669),
	.w7(32'h3bb5b978),
	.w8(32'h3b261903),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc02025),
	.w1(32'h3c239857),
	.w2(32'h3bbdaa38),
	.w3(32'h3b6ffe8b),
	.w4(32'h3bf6e033),
	.w5(32'h3b9d8d6c),
	.w6(32'h3bb43c14),
	.w7(32'h3c06b2c2),
	.w8(32'h3b2a5b86),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab05b30),
	.w1(32'h3a2e0271),
	.w2(32'hb8dca35a),
	.w3(32'hbac4ac31),
	.w4(32'h3a29a5ad),
	.w5(32'h3a8bdb75),
	.w6(32'h39ea5910),
	.w7(32'h3b684d7f),
	.w8(32'h3992f227),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d56a9),
	.w1(32'h3b9c921b),
	.w2(32'h3b2b4b3e),
	.w3(32'h3a5b6e8c),
	.w4(32'h3b8d08af),
	.w5(32'h3b1eb332),
	.w6(32'h38ce4362),
	.w7(32'h3abfb9b7),
	.w8(32'h3b842a24),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7306e08),
	.w1(32'h3a772c6a),
	.w2(32'h3a776db1),
	.w3(32'h3a166170),
	.w4(32'h3afdee61),
	.w5(32'h3ab6e6ff),
	.w6(32'h3b4e1b08),
	.w7(32'h3b5efe1a),
	.w8(32'h3b384409),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82823fa),
	.w1(32'hb9a3064c),
	.w2(32'hbb39ac1a),
	.w3(32'h3b0962aa),
	.w4(32'hba265117),
	.w5(32'hbaf91f0c),
	.w6(32'h3b4b3877),
	.w7(32'h3b2c23fc),
	.w8(32'h3b0adc83),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2669e6),
	.w1(32'h3a600391),
	.w2(32'hbb1312fc),
	.w3(32'hba7475f1),
	.w4(32'hbb1337df),
	.w5(32'hbbc02af3),
	.w6(32'h39ada317),
	.w7(32'hbb1e35ae),
	.w8(32'hbbcec003),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb652b6),
	.w1(32'hbaecf19c),
	.w2(32'hbbdd0364),
	.w3(32'hb97bb876),
	.w4(32'hbbd35769),
	.w5(32'hbc0d9550),
	.w6(32'hba981122),
	.w7(32'hbbe88760),
	.w8(32'hbc0d81d8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012262),
	.w1(32'hbbd34313),
	.w2(32'h3a8c71bd),
	.w3(32'hbb9dc590),
	.w4(32'h39f9210c),
	.w5(32'h3aab737e),
	.w6(32'hbbebf88f),
	.w7(32'h3a27d3da),
	.w8(32'hb9443182),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e7410),
	.w1(32'hb9d7e418),
	.w2(32'h3bc99f42),
	.w3(32'h39b54402),
	.w4(32'h3b15aa30),
	.w5(32'hbb03e675),
	.w6(32'hb963067e),
	.w7(32'h3be5368b),
	.w8(32'h37d6cf77),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91a438),
	.w1(32'h38ece2cb),
	.w2(32'hbbb6b760),
	.w3(32'hbad3285d),
	.w4(32'h3b0bbd01),
	.w5(32'hbbdb3a46),
	.w6(32'h3a058303),
	.w7(32'h3b1750a2),
	.w8(32'hbb53978f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c163a2f),
	.w1(32'h3bcfbb02),
	.w2(32'hbb1cf3b5),
	.w3(32'h3ab4bb9b),
	.w4(32'h3b8aca0f),
	.w5(32'h3a6962dc),
	.w6(32'hbb748020),
	.w7(32'h3b4e63c6),
	.w8(32'hb9a77b5a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00859a),
	.w1(32'h3be3012a),
	.w2(32'h3c3fd080),
	.w3(32'h3b25e41d),
	.w4(32'h3c611f6b),
	.w5(32'h3beaf53c),
	.w6(32'hbc0da56b),
	.w7(32'hbbb02096),
	.w8(32'hbc1c0145),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f7b5a),
	.w1(32'h3b3d7db9),
	.w2(32'h398b9e8c),
	.w3(32'hb9009fb7),
	.w4(32'h3a23293d),
	.w5(32'h3b607e99),
	.w6(32'hbb645b06),
	.w7(32'hbb016964),
	.w8(32'h3b882266),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beac983),
	.w1(32'hbc655fb5),
	.w2(32'h3c1cba8c),
	.w3(32'hbc2bff9a),
	.w4(32'h3c314d61),
	.w5(32'h3c419954),
	.w6(32'hbc77c325),
	.w7(32'h3c35af0d),
	.w8(32'h3c7aec02),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c677edd),
	.w1(32'h3cacfd79),
	.w2(32'hbb000ba9),
	.w3(32'h3bb9f315),
	.w4(32'h3bed813f),
	.w5(32'hbaa0fb5f),
	.w6(32'h3abdef7a),
	.w7(32'hbbc37499),
	.w8(32'hbc02014f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf68147),
	.w1(32'hbbb9241d),
	.w2(32'hbb97d9b2),
	.w3(32'hbc3e17dd),
	.w4(32'hba964a79),
	.w5(32'hbb03195f),
	.w6(32'hbc77f792),
	.w7(32'hbba19821),
	.w8(32'hbba2c856),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d494d),
	.w1(32'h3aa18d9c),
	.w2(32'hb9c567e8),
	.w3(32'h3ada1167),
	.w4(32'hba0565b7),
	.w5(32'hbb205dc5),
	.w6(32'h3b324408),
	.w7(32'h3b0797be),
	.w8(32'hbb5561c9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf302f3),
	.w1(32'h3c494cf6),
	.w2(32'h3c0a6696),
	.w3(32'h3be2c26f),
	.w4(32'h3c2c5259),
	.w5(32'hbb1d0054),
	.w6(32'hba0548fc),
	.w7(32'h3b3f49cc),
	.w8(32'hbc5985fc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc808d3c),
	.w1(32'hbc0b705c),
	.w2(32'h3b70615a),
	.w3(32'hba0a1a2d),
	.w4(32'hba1a97f1),
	.w5(32'hbb1b9215),
	.w6(32'hbc0de61f),
	.w7(32'hbacaa342),
	.w8(32'hbba911fc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce26678),
	.w1(32'h3cf730b1),
	.w2(32'h3cda03d5),
	.w3(32'h3c56ff7e),
	.w4(32'h3c8635b9),
	.w5(32'h3c75bdb5),
	.w6(32'hbb857a51),
	.w7(32'h3ac1cefe),
	.w8(32'hbb001c59),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c003763),
	.w1(32'h3b5240ea),
	.w2(32'h3c0a66fc),
	.w3(32'h3b8c46d0),
	.w4(32'h3baf741a),
	.w5(32'h3b76eada),
	.w6(32'h3a015c21),
	.w7(32'h3bde87ae),
	.w8(32'h3c13610a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b727487),
	.w1(32'hb991a646),
	.w2(32'h3bf0f044),
	.w3(32'hbb57ec06),
	.w4(32'h3ab0b835),
	.w5(32'h3ba2f133),
	.w6(32'h3b104e6f),
	.w7(32'h3c8ef8f4),
	.w8(32'h3d1b621d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71c9a6),
	.w1(32'h3b776601),
	.w2(32'hbbecd0d5),
	.w3(32'h366c3a91),
	.w4(32'hbc128a2d),
	.w5(32'hbc090eee),
	.w6(32'h3c1cb2a3),
	.w7(32'hbbfa1a0d),
	.w8(32'hbc006039),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f91d1),
	.w1(32'hbb1a8d86),
	.w2(32'h3b9b95c2),
	.w3(32'hbbb0eecf),
	.w4(32'h3b683507),
	.w5(32'hba9fd8fc),
	.w6(32'hbbd49b57),
	.w7(32'hbbcb33a1),
	.w8(32'hbc61620b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2300e8),
	.w1(32'hb804a52a),
	.w2(32'hba2958ef),
	.w3(32'hbbb405a0),
	.w4(32'h3bb51bd8),
	.w5(32'h3aeadb6d),
	.w6(32'hbc6bceb7),
	.w7(32'h3c08078c),
	.w8(32'h3c0fe1f9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd51172),
	.w1(32'hbc181198),
	.w2(32'h3b3dfdf2),
	.w3(32'hbb004eb7),
	.w4(32'h3bf2999b),
	.w5(32'h3a2534bb),
	.w6(32'h3b47ef73),
	.w7(32'h3be1f4ca),
	.w8(32'hbbab34f9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd9a35),
	.w1(32'hbbb8192c),
	.w2(32'h3c49010f),
	.w3(32'hbbde9b8b),
	.w4(32'h3c0d1fb7),
	.w5(32'h3c427127),
	.w6(32'hbbcb994f),
	.w7(32'h3bfefe63),
	.w8(32'h3c1bc32c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b9b09),
	.w1(32'hba30e278),
	.w2(32'h3b1cc7c2),
	.w3(32'hbb4cfdf4),
	.w4(32'hba21c850),
	.w5(32'h3cc4d1f2),
	.w6(32'hbb99d931),
	.w7(32'h3b8b25b5),
	.w8(32'h3ce9d04e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2dbd2),
	.w1(32'hbb5be0a4),
	.w2(32'hbb01f44d),
	.w3(32'h3bcf6b3c),
	.w4(32'h3b419a56),
	.w5(32'h3b9b916e),
	.w6(32'hbb7417c8),
	.w7(32'hbb27a53d),
	.w8(32'h3a9114fe),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babb92c),
	.w1(32'h3bbbf2f4),
	.w2(32'hb7f42bc2),
	.w3(32'h392aaed3),
	.w4(32'h3a849a5b),
	.w5(32'hbbc90d2b),
	.w6(32'h392bb359),
	.w7(32'h3b030885),
	.w8(32'hbbef0b1a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c334d),
	.w1(32'hbc11d53d),
	.w2(32'h3bd0638a),
	.w3(32'hbbcd4c9d),
	.w4(32'h3b779c0b),
	.w5(32'h38c90b22),
	.w6(32'hbc0a69b8),
	.w7(32'h3b8405a1),
	.w8(32'hbaa4998b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93208e),
	.w1(32'h3aaf27e9),
	.w2(32'hba96d9f6),
	.w3(32'hbbc61d0e),
	.w4(32'hbb9a32cd),
	.w5(32'hbc05cc55),
	.w6(32'hbb035277),
	.w7(32'hbb5c19d2),
	.w8(32'hbb9689dc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47c915),
	.w1(32'h3b94f10f),
	.w2(32'h3a6f9005),
	.w3(32'hbc0358a1),
	.w4(32'hbb9d689d),
	.w5(32'h3a1cce07),
	.w6(32'hbbf64732),
	.w7(32'hbb7d3c87),
	.w8(32'hba5dbf32),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30b5f1),
	.w1(32'hbbb02da8),
	.w2(32'h3ba87f58),
	.w3(32'hbbe1cf16),
	.w4(32'h3c2e484e),
	.w5(32'h3cc7421d),
	.w6(32'hbc00f3a2),
	.w7(32'h3bcfaec3),
	.w8(32'h3c9f8523),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74057d),
	.w1(32'hbb3a7a24),
	.w2(32'h3c04226b),
	.w3(32'hbb071801),
	.w4(32'h3b29abfd),
	.w5(32'h3ad6f11e),
	.w6(32'hbb73580b),
	.w7(32'h3be63f46),
	.w8(32'h3c598965),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c114691),
	.w1(32'h3c154b06),
	.w2(32'hb9862cee),
	.w3(32'h3c0539ff),
	.w4(32'h3a3d2d58),
	.w5(32'h3b0a9bfc),
	.w6(32'h3c5f6c95),
	.w7(32'hba70c83e),
	.w8(32'h3ad31f16),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91947c),
	.w1(32'h3b565cda),
	.w2(32'h3bb4db68),
	.w3(32'h3abf9c8a),
	.w4(32'h3bc8250d),
	.w5(32'h39e2e5ec),
	.w6(32'h3a6bf7cf),
	.w7(32'h3c25e656),
	.w8(32'h3bb9dbff),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c7b5a),
	.w1(32'hba10f10d),
	.w2(32'hbbcc0236),
	.w3(32'hbbd1aa91),
	.w4(32'hbb981ca8),
	.w5(32'h3bb9bc44),
	.w6(32'hbaf8c5aa),
	.w7(32'hbc0ca940),
	.w8(32'h3c1e4e31),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd339ec),
	.w1(32'h3bbc4a04),
	.w2(32'hbab987d1),
	.w3(32'h3b96f799),
	.w4(32'hba5a8cb8),
	.w5(32'h3b0078db),
	.w6(32'h3b91bb7f),
	.w7(32'h3b3e6c59),
	.w8(32'h3c3f777b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37d72f),
	.w1(32'h3af44ac3),
	.w2(32'hbaf1f1c3),
	.w3(32'hbab3ff7a),
	.w4(32'h3bc53776),
	.w5(32'hbb3278ba),
	.w6(32'h3960e20f),
	.w7(32'h3a9f2ee2),
	.w8(32'h3aa0a39e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e55c8a),
	.w1(32'h3c2509f6),
	.w2(32'hba215b45),
	.w3(32'h3b9120e5),
	.w4(32'h39d2d4cd),
	.w5(32'hbbd9c53b),
	.w6(32'h3c3ad823),
	.w7(32'hba8847a8),
	.w8(32'hbc362a5d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb983dc1),
	.w1(32'hbc01c305),
	.w2(32'hba8ebebc),
	.w3(32'hbbe5ea1a),
	.w4(32'h3b6907af),
	.w5(32'hbc71c18f),
	.w6(32'hbc2a473c),
	.w7(32'hbaf5dd33),
	.w8(32'hbcb6f1d1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81e3d2),
	.w1(32'h39f1cd6b),
	.w2(32'hb77f41d7),
	.w3(32'h3aca4620),
	.w4(32'hbb1a1f48),
	.w5(32'hbc007277),
	.w6(32'hb9edfe63),
	.w7(32'h3a51432a),
	.w8(32'hbb9298fe),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f6ce2),
	.w1(32'h3b415948),
	.w2(32'h3c02812e),
	.w3(32'h3c2d566a),
	.w4(32'h3cd46841),
	.w5(32'h3ca9779f),
	.w6(32'h3bbef420),
	.w7(32'h3c653b3d),
	.w8(32'h3ca61465),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90d6c1),
	.w1(32'h3af4d761),
	.w2(32'h3b4c717e),
	.w3(32'h3a8b0e3b),
	.w4(32'h3c5c0d1a),
	.w5(32'h3b47c717),
	.w6(32'hbbd295b9),
	.w7(32'h3c1b21a3),
	.w8(32'hbb148682),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fa0f5),
	.w1(32'h3bee0d95),
	.w2(32'h3b072980),
	.w3(32'h3b57e0b9),
	.w4(32'h3af4534b),
	.w5(32'h3b45bfa0),
	.w6(32'h3a990e7d),
	.w7(32'h3aaac813),
	.w8(32'h3ae1e0e1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c6574),
	.w1(32'hb8b7a1a5),
	.w2(32'hbb569e0a),
	.w3(32'hba3858e2),
	.w4(32'hbbfc8495),
	.w5(32'hbb16e2ba),
	.w6(32'hb9c1d191),
	.w7(32'hbc333edb),
	.w8(32'hbbd4b332),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03a226),
	.w1(32'h3b8fbb6c),
	.w2(32'h3b72abf3),
	.w3(32'hbbacfc38),
	.w4(32'h3bc4f888),
	.w5(32'hbab644e7),
	.w6(32'hbc12d9a2),
	.w7(32'h3be22ef6),
	.w8(32'hba6026ff),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93c15a),
	.w1(32'hbb9e731b),
	.w2(32'hbbdd3710),
	.w3(32'hbaa97356),
	.w4(32'hbc33d68c),
	.w5(32'hbc014324),
	.w6(32'hbb2ea16f),
	.w7(32'hbc06e1c5),
	.w8(32'hbb8ff761),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0c327),
	.w1(32'hbc028f9c),
	.w2(32'h3b8b2446),
	.w3(32'hbaaccda9),
	.w4(32'h3b966021),
	.w5(32'hba06b695),
	.w6(32'hbb570264),
	.w7(32'h3c684d98),
	.w8(32'h3c85585b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf4825),
	.w1(32'h3ae94082),
	.w2(32'hb9d80e13),
	.w3(32'h3803831c),
	.w4(32'h3b04bb93),
	.w5(32'h3af5d3c9),
	.w6(32'h3bebdfd1),
	.w7(32'h3a740fbc),
	.w8(32'h3ac9baf1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a69cf),
	.w1(32'h3a23f565),
	.w2(32'h3ab9d7bb),
	.w3(32'hb95e0a21),
	.w4(32'h3b6e8671),
	.w5(32'hbc7bf18c),
	.w6(32'h39a7986c),
	.w7(32'hbc50f87e),
	.w8(32'hbca9f019),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74433d),
	.w1(32'hbc03e4df),
	.w2(32'h3bfb8588),
	.w3(32'hbb0eb0ef),
	.w4(32'h3b64561c),
	.w5(32'h3c8db3ce),
	.w6(32'hbc91b559),
	.w7(32'h3c00e29e),
	.w8(32'h3c96e511),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c879dd7),
	.w1(32'h3b024fbb),
	.w2(32'hbbf9be95),
	.w3(32'h3bd24664),
	.w4(32'hbafd320a),
	.w5(32'hba6597fc),
	.w6(32'h3b87f697),
	.w7(32'hbbcb49b2),
	.w8(32'hbac15526),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac90122),
	.w1(32'h3b8fa404),
	.w2(32'hba0c416c),
	.w3(32'hba911959),
	.w4(32'h3aa39947),
	.w5(32'hbbbce375),
	.w6(32'hba61f814),
	.w7(32'h3a45447c),
	.w8(32'hbbffa457),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0baf5b),
	.w1(32'hbb868d14),
	.w2(32'hbb4f6f50),
	.w3(32'h3af3de95),
	.w4(32'h392d70cc),
	.w5(32'hbb0fb16a),
	.w6(32'hbb9c4200),
	.w7(32'hbaf9c219),
	.w8(32'hbb930398),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95779),
	.w1(32'h390f9051),
	.w2(32'h3c05b875),
	.w3(32'hbb3bb68a),
	.w4(32'h3ba390e3),
	.w5(32'h3c0478e3),
	.w6(32'hbb2b588b),
	.w7(32'h3b4df49a),
	.w8(32'h3bbc42c8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a2ba5),
	.w1(32'h3be599ee),
	.w2(32'h3bc2f5e3),
	.w3(32'h3b538d0b),
	.w4(32'h3beca3a5),
	.w5(32'h3c43c37d),
	.w6(32'hb922459f),
	.w7(32'h3bc17301),
	.w8(32'h3c21d3b5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d1ffa),
	.w1(32'h3b4083f2),
	.w2(32'hbba0b0a3),
	.w3(32'h3b04226f),
	.w4(32'hbb2e9da0),
	.w5(32'hbb93d525),
	.w6(32'h3b678a61),
	.w7(32'hbb9d8508),
	.w8(32'hbc045752),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ba5a9),
	.w1(32'hbc109311),
	.w2(32'hbacec5c8),
	.w3(32'hbba4d799),
	.w4(32'h3ba0d295),
	.w5(32'h3c6b936a),
	.w6(32'hbbb04295),
	.w7(32'h3b2a3c41),
	.w8(32'h3c9e5919),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c914131),
	.w1(32'hbb8a6a87),
	.w2(32'h3b1990bf),
	.w3(32'hbb3c71bf),
	.w4(32'h39955c48),
	.w5(32'hbaa1ae79),
	.w6(32'hbb771655),
	.w7(32'h3af50453),
	.w8(32'hba70a6c6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a581b63),
	.w1(32'h3c33bb1f),
	.w2(32'h3bfeccc9),
	.w3(32'hbb0edc31),
	.w4(32'h3c543a17),
	.w5(32'h3c185256),
	.w6(32'hbb53c061),
	.w7(32'h3c783c76),
	.w8(32'h3c2e3fa6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1556db),
	.w1(32'hbc016589),
	.w2(32'hbb967f12),
	.w3(32'hbbbbfe6a),
	.w4(32'h394ae83b),
	.w5(32'h3983c5d4),
	.w6(32'hbaad9a01),
	.w7(32'hbaaa5e8e),
	.w8(32'h3b708764),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb84f18),
	.w1(32'h3bb3ebfa),
	.w2(32'h3c1d0a3b),
	.w3(32'hbb13cb8c),
	.w4(32'h3c49bf1b),
	.w5(32'h3bb8ca09),
	.w6(32'hbba91922),
	.w7(32'h3bf5f387),
	.w8(32'hbaadb465),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1081fa),
	.w1(32'hbb3ea1ab),
	.w2(32'hbb899c27),
	.w3(32'h39903cd4),
	.w4(32'h3ab222b0),
	.w5(32'h3b195a79),
	.w6(32'hbaead331),
	.w7(32'hbb755426),
	.w8(32'hbb943d2b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba159bfc),
	.w1(32'hba46d806),
	.w2(32'h3bd2b327),
	.w3(32'h3b63a10b),
	.w4(32'h3ba8c78f),
	.w5(32'hbbb95d1a),
	.w6(32'hbb6f7db8),
	.w7(32'h3c278a2e),
	.w8(32'hbb558664),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90a763),
	.w1(32'hba2f7b57),
	.w2(32'hba367865),
	.w3(32'h3adb19de),
	.w4(32'h3b59f32b),
	.w5(32'hbc3273a1),
	.w6(32'hbb9f56f0),
	.w7(32'hba80817d),
	.w8(32'hbc825738),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1a16f),
	.w1(32'h39bcc873),
	.w2(32'h3b64c269),
	.w3(32'hbb063fb8),
	.w4(32'h3b950382),
	.w5(32'hba692705),
	.w6(32'hbbe181d1),
	.w7(32'h3a9e9874),
	.w8(32'h399f96cb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab97da5),
	.w1(32'hbbfb8cb8),
	.w2(32'hbb7ca8ed),
	.w3(32'hbbd5ecc8),
	.w4(32'h398541e7),
	.w5(32'h3c1e7705),
	.w6(32'hbbf3563c),
	.w7(32'hbc04deb2),
	.w8(32'h3b2973e6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf38617),
	.w1(32'h3b128a3e),
	.w2(32'hb9aef0dc),
	.w3(32'h3c0caad5),
	.w4(32'h3b5feecf),
	.w5(32'h3b8c4e2e),
	.w6(32'hba460dad),
	.w7(32'h3b94fb30),
	.w8(32'h3c2bbba5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddbb5c),
	.w1(32'h3ba1a381),
	.w2(32'h3ab56e86),
	.w3(32'hbb462f84),
	.w4(32'h386a0e85),
	.w5(32'h3af94b86),
	.w6(32'h3b992842),
	.w7(32'h3a7c36bd),
	.w8(32'h3b859240),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15574b),
	.w1(32'h3b726e68),
	.w2(32'hb9ae7393),
	.w3(32'hbb7c6264),
	.w4(32'hbc5b35d3),
	.w5(32'hbbba503c),
	.w6(32'h3b49a6bb),
	.w7(32'h3c72253d),
	.w8(32'h39cde84f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d120e7d),
	.w1(32'h3ce1ce48),
	.w2(32'hbc332008),
	.w3(32'h3ab6d342),
	.w4(32'hba8c7d3f),
	.w5(32'h3bd1cd65),
	.w6(32'hbb980c10),
	.w7(32'h3c4e1f94),
	.w8(32'h3c81ba55),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3018d),
	.w1(32'hbb3e1c6d),
	.w2(32'hbb68523c),
	.w3(32'h3b025f9c),
	.w4(32'h3b7af7b8),
	.w5(32'h3c8773df),
	.w6(32'h3a8ea289),
	.w7(32'hbc80ea33),
	.w8(32'hbc8a73c5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1a1cb),
	.w1(32'h3ce496f7),
	.w2(32'hbbc74363),
	.w3(32'hbbcaf9b0),
	.w4(32'h3c1397ac),
	.w5(32'h3b50ac66),
	.w6(32'hbb93e386),
	.w7(32'h3c9b0d89),
	.w8(32'h3bb2529a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ea8ae),
	.w1(32'h3b2fc674),
	.w2(32'h3c67e93c),
	.w3(32'hbbec0f5b),
	.w4(32'h3b849783),
	.w5(32'hbc34c817),
	.w6(32'hbc3fc8ee),
	.w7(32'hbb84c220),
	.w8(32'hbab34c8b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a892969),
	.w1(32'hbb7c3b7c),
	.w2(32'h3b20645a),
	.w3(32'h3b80dbb1),
	.w4(32'h3c9c2363),
	.w5(32'h3b5bc595),
	.w6(32'h3cbd8b5b),
	.w7(32'h3c361adc),
	.w8(32'h3ba5ae8d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b60b8),
	.w1(32'h3c5d39f6),
	.w2(32'hbb86041f),
	.w3(32'hbbc58b9e),
	.w4(32'h3b277b5f),
	.w5(32'hbb91c2ad),
	.w6(32'hbca99c88),
	.w7(32'hba96c511),
	.w8(32'hbb41d649),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cef6001),
	.w1(32'h3c0dabd6),
	.w2(32'hbc762fce),
	.w3(32'hb8d711fc),
	.w4(32'hbc1faa22),
	.w5(32'hbb8b5e95),
	.w6(32'hba67cd3e),
	.w7(32'hbbffdfa4),
	.w8(32'h3c55ab7a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c376a26),
	.w1(32'h3b734269),
	.w2(32'h3b1a80f5),
	.w3(32'h3912929c),
	.w4(32'hbbd9335f),
	.w5(32'hbc217822),
	.w6(32'h3c2d448d),
	.w7(32'hbb5078d1),
	.w8(32'h38f72bb8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb858ea2),
	.w1(32'hbbd66b06),
	.w2(32'hbb712686),
	.w3(32'hbb6cc2b3),
	.w4(32'hbc86bda9),
	.w5(32'hbc1247a2),
	.w6(32'h3b99d09d),
	.w7(32'h3ab963d5),
	.w8(32'h3bbfbfa1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa032e1),
	.w1(32'h3abbb8ae),
	.w2(32'hbbadf4d8),
	.w3(32'hbc241301),
	.w4(32'h3a73729a),
	.w5(32'hbb4d49e5),
	.w6(32'h389cc79d),
	.w7(32'h3cd932c6),
	.w8(32'h3d21d04a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9d661),
	.w1(32'hbc2af3e9),
	.w2(32'h3cd0cc90),
	.w3(32'hbaa6f580),
	.w4(32'h3c501c3f),
	.w5(32'h3bf8280e),
	.w6(32'h3bebe6db),
	.w7(32'hbb80d908),
	.w8(32'hbcf652de),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e3b31),
	.w1(32'hbb5e5088),
	.w2(32'hbb89b063),
	.w3(32'h394789cf),
	.w4(32'hbbc050c0),
	.w5(32'hbcb2ec89),
	.w6(32'h3a857093),
	.w7(32'hbd5941bd),
	.w8(32'hbd207f3a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db6a275),
	.w1(32'h3d0525de),
	.w2(32'h3b4234b9),
	.w3(32'hbcd70095),
	.w4(32'h3b7fb961),
	.w5(32'h3b599f71),
	.w6(32'hbd0327bd),
	.w7(32'h3c02edde),
	.w8(32'hbc397804),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b042054),
	.w1(32'h3c8224f7),
	.w2(32'hbc551d9f),
	.w3(32'h3c03bcc3),
	.w4(32'h3b63bf1f),
	.w5(32'h3aaa692d),
	.w6(32'hbb48fc79),
	.w7(32'h3b52526b),
	.w8(32'h3d07fd1c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e80ae),
	.w1(32'h3c226dcc),
	.w2(32'hbad70a08),
	.w3(32'h3b9d7a72),
	.w4(32'h3ac04c78),
	.w5(32'h3b50fc31),
	.w6(32'h3c55f92c),
	.w7(32'h392de01f),
	.w8(32'h3b9b40a6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26de26),
	.w1(32'h3b0045c5),
	.w2(32'hbbc5aeca),
	.w3(32'h3a4a73b7),
	.w4(32'hbc3474a2),
	.w5(32'h3a9e3156),
	.w6(32'hba127820),
	.w7(32'hbcd91284),
	.w8(32'hbd3ab4e7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d485dbf),
	.w1(32'h3d35dcc3),
	.w2(32'hbc4e5cf7),
	.w3(32'hbbc8e842),
	.w4(32'h3cec25e7),
	.w5(32'h3c6d65f0),
	.w6(32'hbcb85e3f),
	.w7(32'h3c4da58f),
	.w8(32'h3d105b7f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdb6ccc1),
	.w1(32'hbd0cf6ee),
	.w2(32'h3c24c167),
	.w3(32'h3b831c3a),
	.w4(32'hbc6ec283),
	.w5(32'hba05c7a2),
	.w6(32'h3ccc57cc),
	.w7(32'hb91dd588),
	.w8(32'h3c3a5838),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba63539),
	.w1(32'hbc5a4019),
	.w2(32'hbb2ac14e),
	.w3(32'h3c12272c),
	.w4(32'hbb407a8e),
	.w5(32'hbb306938),
	.w6(32'h3c55f897),
	.w7(32'hbaf37798),
	.w8(32'h3bc17c75),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb209b2a),
	.w1(32'hb9eecb37),
	.w2(32'hbc628940),
	.w3(32'hbb93806d),
	.w4(32'hb93d3b76),
	.w5(32'hb9a22e82),
	.w6(32'h3aa2a682),
	.w7(32'h3b7017d3),
	.w8(32'h3bfd2d6d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1388bc),
	.w1(32'h3c5680f7),
	.w2(32'h3b9a8cf1),
	.w3(32'h3aabe7a8),
	.w4(32'hbc03b034),
	.w5(32'hbbe1be57),
	.w6(32'h3c26718b),
	.w7(32'hbc921e9f),
	.w8(32'hbc910ac3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc13c7c),
	.w1(32'h3ca173de),
	.w2(32'hbace82c5),
	.w3(32'hbc827ea7),
	.w4(32'hbac1754f),
	.w5(32'h3c088213),
	.w6(32'hbca5387a),
	.w7(32'h3c6e8637),
	.w8(32'h3ca03880),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc867a21),
	.w1(32'hbc673c10),
	.w2(32'h3c41847a),
	.w3(32'hbb46945f),
	.w4(32'hbc0beb69),
	.w5(32'hbbf0fbd6),
	.w6(32'hbbae529d),
	.w7(32'hbc45b2f6),
	.w8(32'hbcb752e9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c473ef6),
	.w1(32'h3c0db3c5),
	.w2(32'hbc590887),
	.w3(32'hb9ea2216),
	.w4(32'h3c41d60f),
	.w5(32'h3b100d6b),
	.w6(32'hbb97dab0),
	.w7(32'hbbfdf04d),
	.w8(32'hbc108dd6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf98dc4),
	.w1(32'hbc7167ed),
	.w2(32'h3b3b56ec),
	.w3(32'hba846b82),
	.w4(32'h3b4135de),
	.w5(32'h3ad010dd),
	.w6(32'hbbdf487e),
	.w7(32'h3b5af5ee),
	.w8(32'hbc9993ca),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ac635),
	.w1(32'h3c4e30e7),
	.w2(32'h3aaf8ab2),
	.w3(32'h3bf9b1cf),
	.w4(32'h3c26963a),
	.w5(32'h3c09f6bb),
	.w6(32'hbbfe15c2),
	.w7(32'hbc7c850f),
	.w8(32'hbc5f0640),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2d5187),
	.w1(32'hbbc0956d),
	.w2(32'h3c046fbe),
	.w3(32'hbbdb8763),
	.w4(32'hb9ea32b8),
	.w5(32'h3907c515),
	.w6(32'hbcbee114),
	.w7(32'h3c8a531c),
	.w8(32'h3d32f62b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd20ed56),
	.w1(32'hbb251393),
	.w2(32'hbb886000),
	.w3(32'h3b4707a7),
	.w4(32'h3aad4088),
	.w5(32'h3c544541),
	.w6(32'h3c8c902e),
	.w7(32'hbc13085a),
	.w8(32'h3bfd747c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24ad39),
	.w1(32'hbc0ed77f),
	.w2(32'hba812afe),
	.w3(32'h3bdbc813),
	.w4(32'hbb8c2df9),
	.w5(32'hbbd3bd0b),
	.w6(32'h3b2023ee),
	.w7(32'h3b2cb8be),
	.w8(32'hba459a94),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ed4d1),
	.w1(32'h3bafd889),
	.w2(32'hbc254512),
	.w3(32'hb9b68f83),
	.w4(32'h3c3336fd),
	.w5(32'hbbd554ae),
	.w6(32'h3c0ac9d3),
	.w7(32'hbc0cdae8),
	.w8(32'h3b742b05),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c946923),
	.w1(32'h3bdd1bdf),
	.w2(32'h3b8d2404),
	.w3(32'h3a8720a5),
	.w4(32'h3b7f89bb),
	.w5(32'hbb267338),
	.w6(32'h3c2fb082),
	.w7(32'hbc02cff6),
	.w8(32'hbc7f4742),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c499f66),
	.w1(32'h3c9857ea),
	.w2(32'h3a3b2a56),
	.w3(32'h3b966242),
	.w4(32'h3c09a7a4),
	.w5(32'h3c21375d),
	.w6(32'hbc16aa60),
	.w7(32'h3cc24b24),
	.w8(32'h3cd7907f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd5696),
	.w1(32'hbc858a91),
	.w2(32'h3cd6f022),
	.w3(32'hbaaca16a),
	.w4(32'hbbde9004),
	.w5(32'hbb9e1153),
	.w6(32'h3b199e70),
	.w7(32'hbcd4c0ab),
	.w8(32'hbd46636d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8bca12),
	.w1(32'h3c88df79),
	.w2(32'h3c3d87a3),
	.w3(32'hbc159e0f),
	.w4(32'hbcfb3f86),
	.w5(32'hbc9bd2e1),
	.w6(32'hbd0fd2ed),
	.w7(32'hbcd43870),
	.w8(32'hbcd9ec0b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09f4b3),
	.w1(32'h3cbdf0f1),
	.w2(32'hbc4c3db2),
	.w3(32'hbcb9bc23),
	.w4(32'hbc586575),
	.w5(32'h3bd499b8),
	.w6(32'hbc1dc8c5),
	.w7(32'h3c72eb6c),
	.w8(32'h3d04fd56),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0001c5),
	.w1(32'hbc9e7326),
	.w2(32'h3c7c2bbb),
	.w3(32'h3c07d0c8),
	.w4(32'hbc0c1372),
	.w5(32'h3a5a9afc),
	.w6(32'h3c9e04dd),
	.w7(32'h3c1da7a6),
	.w8(32'h3c67b4d1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5b5d2),
	.w1(32'h37a15952),
	.w2(32'hbb99a8e1),
	.w3(32'h37b8e236),
	.w4(32'hbb27574c),
	.w5(32'h3c3e9dbe),
	.w6(32'hbc82da90),
	.w7(32'hbbf49ba9),
	.w8(32'hbba5de0b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe3599),
	.w1(32'hbbd5f12f),
	.w2(32'hbb866c98),
	.w3(32'hbb9ec61d),
	.w4(32'hb9cc7bd2),
	.w5(32'h3ba8771f),
	.w6(32'h3a2f27be),
	.w7(32'hbb53b96d),
	.w8(32'h3bf29730),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba524cf),
	.w1(32'hbb98debe),
	.w2(32'hba73bb48),
	.w3(32'h3a509606),
	.w4(32'hbbd4e689),
	.w5(32'hbc385c2d),
	.w6(32'h3acfcb7c),
	.w7(32'h3b955820),
	.w8(32'hbc0d7f96),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf70b12),
	.w1(32'hbb61b4ec),
	.w2(32'h3c061d72),
	.w3(32'h3ae1d64c),
	.w4(32'hbc08e5fb),
	.w5(32'hbc3dbefe),
	.w6(32'hbc9209c8),
	.w7(32'hbc5e6f45),
	.w8(32'hbc4cffe8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0644ee),
	.w1(32'h3b8b045d),
	.w2(32'hbc5593c5),
	.w3(32'hbc1f45e3),
	.w4(32'h3c080b7d),
	.w5(32'h3bc3586c),
	.w6(32'hbba5980f),
	.w7(32'hbc056e31),
	.w8(32'hbc505c65),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3013a6),
	.w1(32'hbacc2654),
	.w2(32'h3c3d7d92),
	.w3(32'hbbe95d21),
	.w4(32'hbb1c9b83),
	.w5(32'h3af9e16c),
	.w6(32'hbc17c1ba),
	.w7(32'h3c3579f0),
	.w8(32'h3d133fcc),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5537b8),
	.w1(32'hbc5eec7f),
	.w2(32'hbb866d0e),
	.w3(32'hbb3a782c),
	.w4(32'h3ac7661b),
	.w5(32'h3c03e485),
	.w6(32'h3c2569d0),
	.w7(32'hbb8347d3),
	.w8(32'h3bed7632),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07d802),
	.w1(32'hbc0a2e37),
	.w2(32'h3c1ef606),
	.w3(32'h3b84975c),
	.w4(32'hbb083bc9),
	.w5(32'h398f73b3),
	.w6(32'h3b6b2f4e),
	.w7(32'hbc261de0),
	.w8(32'h3c7494b8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ffa04),
	.w1(32'h3c302ec4),
	.w2(32'h3c45ec56),
	.w3(32'hbbc98817),
	.w4(32'hbc039cac),
	.w5(32'hbbfd2fef),
	.w6(32'h3b83a402),
	.w7(32'hbbe3c188),
	.w8(32'h3b4b1cb3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b946119),
	.w1(32'hbb2f86d1),
	.w2(32'h3b8ad7f0),
	.w3(32'hbbf210b4),
	.w4(32'h3a840b78),
	.w5(32'hbbe8c798),
	.w6(32'h3cb152f7),
	.w7(32'h3c31f92a),
	.w8(32'h3c3bbf74),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50486d),
	.w1(32'hb9dcedf6),
	.w2(32'h3c6a0ffb),
	.w3(32'hbc1ed996),
	.w4(32'hbc541a47),
	.w5(32'hbb69f679),
	.w6(32'h3bcf1951),
	.w7(32'h3c29ba37),
	.w8(32'h3c54bb39),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aaec4),
	.w1(32'h3b62bdbc),
	.w2(32'hba846622),
	.w3(32'hbbc57acf),
	.w4(32'h3b800060),
	.w5(32'h3c15c814),
	.w6(32'hbca34db5),
	.w7(32'hbc59500d),
	.w8(32'hba0eea24),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule