module layer_10_featuremap_256(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199f16),
	.w1(32'h3cb0e1b7),
	.w2(32'h3c0107c7),
	.w3(32'hbcdac919),
	.w4(32'hbca93ee3),
	.w5(32'hbc2587a8),
	.w6(32'h3be09928),
	.w7(32'hbb2564ec),
	.w8(32'hbaba44f6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65c7b0),
	.w1(32'h3bd38851),
	.w2(32'h3b18a89d),
	.w3(32'hbc3ca86b),
	.w4(32'h3b8fd08a),
	.w5(32'h3c03880f),
	.w6(32'h3b68ee1d),
	.w7(32'hbb33a29b),
	.w8(32'hba686d9a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33cd3e),
	.w1(32'h3ba960c4),
	.w2(32'hbb9e9712),
	.w3(32'h3be6eef8),
	.w4(32'hbb6ff77f),
	.w5(32'h3c2fd214),
	.w6(32'hbb243dee),
	.w7(32'hbc2f293e),
	.w8(32'h3ae83e7e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba811eb),
	.w1(32'hbb92b768),
	.w2(32'hba5b017b),
	.w3(32'h3ca6e13a),
	.w4(32'h3c89dabb),
	.w5(32'h3ac8b145),
	.w6(32'h3b384d85),
	.w7(32'h3bc65004),
	.w8(32'hbb440931),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23d090),
	.w1(32'h3c51392c),
	.w2(32'h3b37873e),
	.w3(32'h3ba9a3aa),
	.w4(32'h3ba73f77),
	.w5(32'h3bcee880),
	.w6(32'h3b8f85c9),
	.w7(32'hbb0dce52),
	.w8(32'h3bd83b20),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4bb68),
	.w1(32'h3b104fe2),
	.w2(32'h3b4ce6bd),
	.w3(32'h3c3f32c3),
	.w4(32'h3ba9dde0),
	.w5(32'hba128480),
	.w6(32'h3c7cc368),
	.w7(32'h3c17506a),
	.w8(32'hbb2dae72),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72adb5),
	.w1(32'hbb4faf34),
	.w2(32'hbbcef34c),
	.w3(32'h3c2c0677),
	.w4(32'h3b4346a2),
	.w5(32'h3c37b142),
	.w6(32'h3c4ba006),
	.w7(32'h3ad5b0da),
	.w8(32'h3c0d58d1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc103714),
	.w1(32'hbc23d45c),
	.w2(32'hbb2fab78),
	.w3(32'h3c4dd307),
	.w4(32'h3ba27de9),
	.w5(32'h3b172906),
	.w6(32'h3b9a9e3e),
	.w7(32'hbb30b9d0),
	.w8(32'h3a3225be),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6baa6),
	.w1(32'h3c51067b),
	.w2(32'h3bbbfe9a),
	.w3(32'h3c153acb),
	.w4(32'h3bceb02b),
	.w5(32'h3b908d12),
	.w6(32'h3c4bad9b),
	.w7(32'h3bfd4f18),
	.w8(32'h3b5f8db9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c6c5),
	.w1(32'h3a9fd8e7),
	.w2(32'h3befa0e9),
	.w3(32'h3be5e6db),
	.w4(32'h3bd5e1a9),
	.w5(32'h3c440a02),
	.w6(32'h3c52d831),
	.w7(32'h3c07484b),
	.w8(32'h3bb15ff2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85895c),
	.w1(32'h3af5acd3),
	.w2(32'h3b2aa0a1),
	.w3(32'h3c8db434),
	.w4(32'h3bcd0aca),
	.w5(32'h3b388018),
	.w6(32'h3c3e28e7),
	.w7(32'h3a8d5bf5),
	.w8(32'h3bf477ad),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb54b09),
	.w1(32'h3ab7a21c),
	.w2(32'hbbd0fd3f),
	.w3(32'h3beda099),
	.w4(32'hbc0a9623),
	.w5(32'hbc0c620f),
	.w6(32'hbb41e12e),
	.w7(32'hbc39419a),
	.w8(32'h3b9ab1cf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6839d9),
	.w1(32'h3c779e27),
	.w2(32'h3be9d214),
	.w3(32'hbcee7975),
	.w4(32'hbd0a10e4),
	.w5(32'hbb9f3ab0),
	.w6(32'hbb132b5a),
	.w7(32'hbb66f646),
	.w8(32'h3a6566c0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b855ef4),
	.w1(32'h3c1f25e6),
	.w2(32'h3b2727fa),
	.w3(32'hbc471432),
	.w4(32'h394cc6b7),
	.w5(32'h3b0bf744),
	.w6(32'hbab8f01a),
	.w7(32'h399f4666),
	.w8(32'hbb532cd0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c64a37),
	.w1(32'hbb5fe2ea),
	.w2(32'hbb1b9862),
	.w3(32'h3c010596),
	.w4(32'h3990d1e7),
	.w5(32'hbb7b418c),
	.w6(32'h3a39620c),
	.w7(32'hbb6a6b04),
	.w8(32'hbc09dc51),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f271ac),
	.w1(32'h3bf86a54),
	.w2(32'hbb483f17),
	.w3(32'hbc4fc641),
	.w4(32'hbb44646a),
	.w5(32'hbb84eca1),
	.w6(32'hbbb04ea7),
	.w7(32'hbafbc6b4),
	.w8(32'h3bc99f00),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8938339),
	.w1(32'h3af9558b),
	.w2(32'hba9eecc5),
	.w3(32'hbc056c6a),
	.w4(32'hbba251da),
	.w5(32'hbb05f8cc),
	.w6(32'h3c0cd07a),
	.w7(32'h3baadd23),
	.w8(32'h39f1e8c4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bc883),
	.w1(32'hbaeaac67),
	.w2(32'h3a67860b),
	.w3(32'hbc30e29f),
	.w4(32'hbc249fd5),
	.w5(32'h3bceb958),
	.w6(32'hbbad3afb),
	.w7(32'hbbb3da60),
	.w8(32'hbac316d4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70195a),
	.w1(32'hbbf4e1c5),
	.w2(32'h3a43df9e),
	.w3(32'h3ab8cf7d),
	.w4(32'hbbee9e48),
	.w5(32'h3b15bf2a),
	.w6(32'hbc056923),
	.w7(32'hbc61d665),
	.w8(32'h3a5b32b9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc024213),
	.w1(32'hbb46b348),
	.w2(32'h3b3599ad),
	.w3(32'hbbe5d6d1),
	.w4(32'h3b21b3aa),
	.w5(32'hbae54c8d),
	.w6(32'h3aad74f2),
	.w7(32'hbb222ae1),
	.w8(32'hbba93f29),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ff5bb),
	.w1(32'h3c9e4923),
	.w2(32'h3b91aec4),
	.w3(32'hbc921763),
	.w4(32'hbba8b4d4),
	.w5(32'h3c322740),
	.w6(32'h3919dbeb),
	.w7(32'h3adf05ce),
	.w8(32'h3a0eb8a8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b8abb),
	.w1(32'hbc552b45),
	.w2(32'hbb8f9eff),
	.w3(32'h3cccd779),
	.w4(32'h3cc059a3),
	.w5(32'h3b1620dc),
	.w6(32'h3baadf02),
	.w7(32'h3c67e251),
	.w8(32'h3addbb46),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd63fde),
	.w1(32'h37412407),
	.w2(32'hbbb02203),
	.w3(32'h3b1855bf),
	.w4(32'hbb831940),
	.w5(32'hbc6a0fc2),
	.w6(32'hbb1150db),
	.w7(32'hbbbeb0f5),
	.w8(32'hbbeba992),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5832b2),
	.w1(32'h3be5be87),
	.w2(32'hbb870bc2),
	.w3(32'hbc842310),
	.w4(32'hbc524f06),
	.w5(32'hba8fbc5a),
	.w6(32'hba91f1f0),
	.w7(32'hbc2e313d),
	.w8(32'h3b436c0b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8668a0),
	.w1(32'hba77cd5e),
	.w2(32'hbbd68dcb),
	.w3(32'hbb0c4619),
	.w4(32'hbb5daa68),
	.w5(32'h3b970e3f),
	.w6(32'hb976185d),
	.w7(32'hbaf670e8),
	.w8(32'h3a47ee84),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fbe8c),
	.w1(32'hbb7a7bfe),
	.w2(32'h3ab5036d),
	.w3(32'h3b094045),
	.w4(32'hbbe31f37),
	.w5(32'h3c98828d),
	.w6(32'h3a801e63),
	.w7(32'hbb04ff5d),
	.w8(32'h3a4fdac2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc245259),
	.w1(32'hbc06fb09),
	.w2(32'hbc82503d),
	.w3(32'h3cc0d4de),
	.w4(32'h3bead397),
	.w5(32'hbc3bd8b4),
	.w6(32'h3a8ac9ae),
	.w7(32'hbb6c7b1f),
	.w8(32'hbb2e988f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc72954),
	.w1(32'h3ca0ea5d),
	.w2(32'h3c8376eb),
	.w3(32'hbc9ccab3),
	.w4(32'hbc1bd7cc),
	.w5(32'hb7b41699),
	.w6(32'hb7d3c366),
	.w7(32'h3b5902d8),
	.w8(32'hbb5a1844),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bb12f),
	.w1(32'hb836fb2f),
	.w2(32'h3c0c0390),
	.w3(32'hbac3b725),
	.w4(32'h3bd05d92),
	.w5(32'h3aeb9e48),
	.w6(32'h3baa6f6e),
	.w7(32'h3b725db2),
	.w8(32'hba8b5a0b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45308b),
	.w1(32'h39a84027),
	.w2(32'hbbde9466),
	.w3(32'hbc38d7c3),
	.w4(32'hbbec457c),
	.w5(32'hbbda103e),
	.w6(32'h3992d78d),
	.w7(32'hbc1c4ac1),
	.w8(32'hbc3fd527),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b845339),
	.w1(32'h3bb61a9a),
	.w2(32'h3b0975a1),
	.w3(32'hbba80b57),
	.w4(32'hbc0e3254),
	.w5(32'hbc0a4530),
	.w6(32'hbca8690d),
	.w7(32'hbce7236d),
	.w8(32'hbb389b69),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cea1c),
	.w1(32'hbc88998b),
	.w2(32'hbc1cd99b),
	.w3(32'hbbee8e62),
	.w4(32'hb83a70d6),
	.w5(32'hbca2ee8a),
	.w6(32'hbaaa15b4),
	.w7(32'h3abd1d62),
	.w8(32'hbb76c7f8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19c1de),
	.w1(32'hbc3d22dd),
	.w2(32'hb7aa6864),
	.w3(32'hbc4ae725),
	.w4(32'hbb61c985),
	.w5(32'hbb846688),
	.w6(32'h3b8c0a14),
	.w7(32'h3b1c5b7e),
	.w8(32'hbba8bca2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19e6b2),
	.w1(32'h3bcd88e6),
	.w2(32'h3b1daf72),
	.w3(32'hbc4273c0),
	.w4(32'hbbbb4304),
	.w5(32'h3bda9d37),
	.w6(32'hbb8d2717),
	.w7(32'hbbae3c5d),
	.w8(32'h3bcbe9f6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f68052),
	.w1(32'hbb284ed8),
	.w2(32'hba964891),
	.w3(32'h3ac27795),
	.w4(32'h39f9329f),
	.w5(32'hbb00da58),
	.w6(32'h3c1cfb12),
	.w7(32'h3a577838),
	.w8(32'hbc32efd2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fb5be),
	.w1(32'h3bdca611),
	.w2(32'hbbbff471),
	.w3(32'hbc2f1297),
	.w4(32'hbc23d7c0),
	.w5(32'hbc7254b1),
	.w6(32'hbbade9c7),
	.w7(32'hbc12c4e0),
	.w8(32'hbbff2cd8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8049e),
	.w1(32'hbbd4f2b0),
	.w2(32'h3bd44ad4),
	.w3(32'hbc7e27f1),
	.w4(32'hbc49fb79),
	.w5(32'h3c019b18),
	.w6(32'hbc172164),
	.w7(32'hbc93240c),
	.w8(32'h3b4d4ce9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84a6db),
	.w1(32'hbc0d44b3),
	.w2(32'hbc5e2b73),
	.w3(32'h3cbd6ef9),
	.w4(32'h3c3b5acd),
	.w5(32'h3b56b3cc),
	.w6(32'h3c45b1ed),
	.w7(32'hbaa3c670),
	.w8(32'h3bfabd66),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf4242),
	.w1(32'h3bf6af2e),
	.w2(32'h3c0e1f27),
	.w3(32'hbbf0641f),
	.w4(32'hbabb6c37),
	.w5(32'h3c538d96),
	.w6(32'h3c6a909d),
	.w7(32'hbb2a1efe),
	.w8(32'h3bf44c3c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb397f5),
	.w1(32'hbc748d99),
	.w2(32'hbb9f6612),
	.w3(32'h3c757915),
	.w4(32'h3b136bf0),
	.w5(32'hbb40c5f1),
	.w6(32'h3c4eb6bc),
	.w7(32'h3c445457),
	.w8(32'h3b2cc46e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48d15c),
	.w1(32'h3afcf037),
	.w2(32'h3b8dfbf0),
	.w3(32'hbbf4f2bf),
	.w4(32'hbbf377b2),
	.w5(32'hbb380881),
	.w6(32'hbb7e50a9),
	.w7(32'hbae2bc03),
	.w8(32'hbb428249),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a0b28),
	.w1(32'hbc3c5fbb),
	.w2(32'hbbc19f5a),
	.w3(32'h3c1db711),
	.w4(32'hb9d42baf),
	.w5(32'hbc2daa2c),
	.w6(32'h3bad82a2),
	.w7(32'h3b097efe),
	.w8(32'hbaf6192f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870375),
	.w1(32'hbb82770b),
	.w2(32'hbc1e09e0),
	.w3(32'h3af0647a),
	.w4(32'hbc31fd8d),
	.w5(32'hbba903bd),
	.w6(32'h3a74a2a1),
	.w7(32'hbc48e45b),
	.w8(32'hbc208df7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6544af),
	.w1(32'hbc33be9b),
	.w2(32'hbc6202f5),
	.w3(32'hbbff2a91),
	.w4(32'hbc48859d),
	.w5(32'hba86e6c1),
	.w6(32'hbbe7e238),
	.w7(32'hbc7592fb),
	.w8(32'hbb5b011c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7131d9),
	.w1(32'hbc3709b1),
	.w2(32'h3b8fe83b),
	.w3(32'h3c4f1509),
	.w4(32'h3c1e9290),
	.w5(32'hbc020057),
	.w6(32'h3c00214a),
	.w7(32'h3c27d855),
	.w8(32'hba1f0455),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88ff30),
	.w1(32'h3cb04893),
	.w2(32'h3c2190c9),
	.w3(32'hbc9ef6b4),
	.w4(32'hbc88ebc9),
	.w5(32'h3c57fd3a),
	.w6(32'hbc10af77),
	.w7(32'hbb98b6c5),
	.w8(32'h3ace39fc),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c8e20),
	.w1(32'hbbc8f994),
	.w2(32'hbc05a358),
	.w3(32'h3b2d5c87),
	.w4(32'hbb6aa2af),
	.w5(32'h3b789bb5),
	.w6(32'hbba3148d),
	.w7(32'hbc1842c8),
	.w8(32'h3b8dd354),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9898a9),
	.w1(32'hb876493d),
	.w2(32'hbaf59a4b),
	.w3(32'h3ba4150b),
	.w4(32'h3b0088d0),
	.w5(32'hbc8e34f9),
	.w6(32'h3b11cb25),
	.w7(32'h3a5fb6a3),
	.w8(32'hbc0ce998),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02c68e),
	.w1(32'h3be04021),
	.w2(32'hba95fe0b),
	.w3(32'hbcba0b4d),
	.w4(32'hbcddd32b),
	.w5(32'h3c256a35),
	.w6(32'hbbd92e4b),
	.w7(32'hbc74d398),
	.w8(32'h3b4a079d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80b9f2),
	.w1(32'hbc248cac),
	.w2(32'hbbdd2d5c),
	.w3(32'h3ccf46b3),
	.w4(32'h3cabf0a3),
	.w5(32'h3b111126),
	.w6(32'h3c79624c),
	.w7(32'h3c0903d1),
	.w8(32'hbb3d9ac1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27c1c9),
	.w1(32'h3a9625a5),
	.w2(32'hbbd282e2),
	.w3(32'hbbaf36fa),
	.w4(32'hbbe13c59),
	.w5(32'hbc03c580),
	.w6(32'hb9a28ffd),
	.w7(32'hbac3de21),
	.w8(32'hbafe8f94),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d9da9),
	.w1(32'hbb5813ea),
	.w2(32'hbb5507c9),
	.w3(32'hbbb040f3),
	.w4(32'hbaf12b81),
	.w5(32'h3ac8fb3e),
	.w6(32'hbc15b24b),
	.w7(32'hbbdc6113),
	.w8(32'hbc029ad0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393eb4ed),
	.w1(32'h3a66eee3),
	.w2(32'hbb233768),
	.w3(32'hb811fcfa),
	.w4(32'hbb574a09),
	.w5(32'h3ada4fd2),
	.w6(32'hbbfe378e),
	.w7(32'hbb9684ce),
	.w8(32'h3b658111),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d7aa2),
	.w1(32'hbb8c769f),
	.w2(32'h3b9ca7e5),
	.w3(32'hbc0a9a91),
	.w4(32'hbccb0560),
	.w5(32'hbba66b5a),
	.w6(32'hba79b006),
	.w7(32'hbc187428),
	.w8(32'hbb1a78da),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1a33b),
	.w1(32'h3a4e9954),
	.w2(32'h3a7e7e31),
	.w3(32'hbc04b602),
	.w4(32'h3a53924c),
	.w5(32'hbbbd0e42),
	.w6(32'hbb289876),
	.w7(32'hbb84caaf),
	.w8(32'h3b6c9365),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81b7ed),
	.w1(32'h3b809851),
	.w2(32'h3b42cd5d),
	.w3(32'hbba05f2d),
	.w4(32'h3bc0476b),
	.w5(32'h3a4ddef2),
	.w6(32'h3b10933a),
	.w7(32'h3b1f992a),
	.w8(32'h3b1cf78a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7efdd),
	.w1(32'hba735f89),
	.w2(32'h3adb64ad),
	.w3(32'hbad8abb5),
	.w4(32'h3aee42e6),
	.w5(32'h3a51e447),
	.w6(32'hbbdcc538),
	.w7(32'h3ac04839),
	.w8(32'hbb0e68a4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf573cb),
	.w1(32'hbb39de7f),
	.w2(32'hbba75afd),
	.w3(32'hbc1ae5ba),
	.w4(32'hbb8d50d6),
	.w5(32'h3be7a6b4),
	.w6(32'hb9db7bf3),
	.w7(32'hba3a123a),
	.w8(32'h394ce317),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaac571),
	.w1(32'hbc1af8ed),
	.w2(32'hbbdab0b3),
	.w3(32'h3c9e04c6),
	.w4(32'h3c593012),
	.w5(32'h3c6b2bb5),
	.w6(32'h3c7fae12),
	.w7(32'h3bad00ae),
	.w8(32'h3bd31356),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b0cad),
	.w1(32'hbcb973cc),
	.w2(32'h3c5386bd),
	.w3(32'h3cc397e6),
	.w4(32'h3c820cb7),
	.w5(32'h39771047),
	.w6(32'hbc072303),
	.w7(32'h3c265c61),
	.w8(32'h3b22bea0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee3f54),
	.w1(32'h3ad31469),
	.w2(32'hba13c469),
	.w3(32'hbbec04c4),
	.w4(32'hbbb1ab15),
	.w5(32'h3b4b6f04),
	.w6(32'h3c26d460),
	.w7(32'hbb918596),
	.w8(32'h39102e5e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadead0),
	.w1(32'hba4dd199),
	.w2(32'h3b8717eb),
	.w3(32'hbc02a0f1),
	.w4(32'hbbd5d1e8),
	.w5(32'hbbc41130),
	.w6(32'h3adfa733),
	.w7(32'hba0f0199),
	.w8(32'hbb2d50e2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c314c),
	.w1(32'hbabf5d23),
	.w2(32'hbb4fe8c1),
	.w3(32'hbc0b2ab8),
	.w4(32'hbc18d571),
	.w5(32'hba80c63e),
	.w6(32'h3aaf85fc),
	.w7(32'hbba397a5),
	.w8(32'h3a465562),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3dd0de),
	.w1(32'h3b258087),
	.w2(32'h39baa8db),
	.w3(32'hbba8d979),
	.w4(32'hbb8e6a13),
	.w5(32'h3b1ce025),
	.w6(32'hbaa908e9),
	.w7(32'hbb4b357d),
	.w8(32'h3925f773),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2bc34),
	.w1(32'h39909992),
	.w2(32'h39a29b69),
	.w3(32'hbb833562),
	.w4(32'hbb067be4),
	.w5(32'hbb453c7d),
	.w6(32'h3b5ddd2b),
	.w7(32'hbbdbf4fa),
	.w8(32'hbae6b014),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38a3e3),
	.w1(32'h3b91bb30),
	.w2(32'h3b5d10ad),
	.w3(32'hbba1ad31),
	.w4(32'hb9932b25),
	.w5(32'h3b5ae4d4),
	.w6(32'hbae12ddb),
	.w7(32'hbb55ce3c),
	.w8(32'h3a2017e3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba582f8),
	.w1(32'h3c79fb93),
	.w2(32'h3ae160ca),
	.w3(32'h3afd09b0),
	.w4(32'hbc02798c),
	.w5(32'hbc16e1fb),
	.w6(32'hbb0402f8),
	.w7(32'hbb90bc1d),
	.w8(32'hbbe64cb3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b351c),
	.w1(32'h3c02de02),
	.w2(32'hbbfb3036),
	.w3(32'hbc1de051),
	.w4(32'hbc035919),
	.w5(32'hbbea2d50),
	.w6(32'hbb962813),
	.w7(32'hbb9cf497),
	.w8(32'h3b14cf40),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d902a),
	.w1(32'hbb51458d),
	.w2(32'hbc353001),
	.w3(32'hbc8ce90b),
	.w4(32'h3a927bd8),
	.w5(32'h3c28b385),
	.w6(32'hbb8735c1),
	.w7(32'hba4d3ae2),
	.w8(32'hbae3628b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcb2c4),
	.w1(32'hbb9d2678),
	.w2(32'hbbaedbf1),
	.w3(32'h3b88f826),
	.w4(32'hbb18ed34),
	.w5(32'h3ba7ddcf),
	.w6(32'hbb6556cb),
	.w7(32'hbb38c363),
	.w8(32'h3a7fd04e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8607ed),
	.w1(32'hbc5a3abd),
	.w2(32'hbc03e4af),
	.w3(32'h3c1b19f7),
	.w4(32'h3afb062f),
	.w5(32'h3b200ca1),
	.w6(32'h3b6cfa75),
	.w7(32'hbb91098b),
	.w8(32'h3bc34777),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6be51),
	.w1(32'h3ca891bb),
	.w2(32'hbbd79752),
	.w3(32'hbc57bfa2),
	.w4(32'hbc086f2a),
	.w5(32'hba24ca39),
	.w6(32'h3a197f34),
	.w7(32'hbb393a4c),
	.w8(32'h3bd03a5c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b673aea),
	.w1(32'h3ba11f33),
	.w2(32'hbb0a45ec),
	.w3(32'hbbaa5142),
	.w4(32'hbbfd8693),
	.w5(32'hbc137a63),
	.w6(32'hb9b5744b),
	.w7(32'h3ac17634),
	.w8(32'hbba5be10),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb692c74),
	.w1(32'hba5ae0c9),
	.w2(32'h3b15ace7),
	.w3(32'hbca7785a),
	.w4(32'hbc788cb6),
	.w5(32'h3b2175bc),
	.w6(32'hbbc48d87),
	.w7(32'hbc27840a),
	.w8(32'h392dfa07),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcba97),
	.w1(32'h3c5b7648),
	.w2(32'h3b77b8dc),
	.w3(32'hba844010),
	.w4(32'hbc1179d2),
	.w5(32'hbbe73d5d),
	.w6(32'hb9d63f71),
	.w7(32'hbbba10ce),
	.w8(32'h3c387fef),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d070b18),
	.w1(32'h3ccc77aa),
	.w2(32'h3c6fcdae),
	.w3(32'hbcc21ead),
	.w4(32'hbcf6009b),
	.w5(32'h3a8bf360),
	.w6(32'hbbc827d3),
	.w7(32'hbbd4ed98),
	.w8(32'h3adfbf76),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b856a71),
	.w1(32'hba1651b8),
	.w2(32'h3a548d75),
	.w3(32'hbb98d883),
	.w4(32'hbc0af79d),
	.w5(32'hbb6bcd2f),
	.w6(32'hbb738891),
	.w7(32'hbb0cd268),
	.w8(32'hbc21283c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0afdb4),
	.w1(32'hbbce3c9d),
	.w2(32'hbb7ba646),
	.w3(32'h3b389231),
	.w4(32'h3b2b60cb),
	.w5(32'h3bb14524),
	.w6(32'hbbb1b8c1),
	.w7(32'hbb756536),
	.w8(32'h3c184111),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8198f8),
	.w1(32'h3c21485d),
	.w2(32'h3b8b66c8),
	.w3(32'hbb1bee11),
	.w4(32'hbbd8c738),
	.w5(32'hbb486606),
	.w6(32'hb9dbd12a),
	.w7(32'h3a84af96),
	.w8(32'h3bc6f8b6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c461e33),
	.w1(32'h3c8ab696),
	.w2(32'h3c11341e),
	.w3(32'hbc3dc559),
	.w4(32'hbc2a4712),
	.w5(32'h3b5a216a),
	.w6(32'h3bbc2426),
	.w7(32'h3aa929a3),
	.w8(32'h3bd92e5f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4f766),
	.w1(32'h3b560652),
	.w2(32'h3aa1a409),
	.w3(32'h3c048140),
	.w4(32'h3a2c4ac1),
	.w5(32'hbb8c73ef),
	.w6(32'hba424f10),
	.w7(32'h3abd3c4b),
	.w8(32'h3b86cd3b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20836a),
	.w1(32'h3bb0c350),
	.w2(32'h3b0bce3d),
	.w3(32'hbc35ba5b),
	.w4(32'hbc8618d3),
	.w5(32'hbaea2380),
	.w6(32'hbb4f60de),
	.w7(32'hbc01e987),
	.w8(32'hbb0fa030),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e406a),
	.w1(32'h3b3fab94),
	.w2(32'hbbdddbf1),
	.w3(32'hbb145e96),
	.w4(32'hbbfb9ce4),
	.w5(32'h3c428333),
	.w6(32'hba1d6f34),
	.w7(32'hbbf2b23b),
	.w8(32'hbbc6db2f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05c1d9),
	.w1(32'h38ec77bf),
	.w2(32'hbc1793a8),
	.w3(32'h3bdce6af),
	.w4(32'h3b438634),
	.w5(32'hbb92ca0c),
	.w6(32'hbca72a91),
	.w7(32'hbc178692),
	.w8(32'hbb97ea73),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb430ca4),
	.w1(32'h3af77886),
	.w2(32'hbb930a72),
	.w3(32'h39f68053),
	.w4(32'hbb2a50e3),
	.w5(32'hbb26471f),
	.w6(32'hbb30e46a),
	.w7(32'hbbb262f9),
	.w8(32'h3c07ff79),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab529cc),
	.w1(32'h3b0447e6),
	.w2(32'h3c275169),
	.w3(32'hbc983eab),
	.w4(32'hbc58bd90),
	.w5(32'h3c2302e7),
	.w6(32'h3b76fabd),
	.w7(32'h39ae3f82),
	.w8(32'h3b4b8f8e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab1806),
	.w1(32'hbbb790e8),
	.w2(32'hbc51b670),
	.w3(32'h3c56b20a),
	.w4(32'hbc1d8390),
	.w5(32'hbad0fcc3),
	.w6(32'h3b26d192),
	.w7(32'hbc2f3e00),
	.w8(32'h3ba67aed),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac13014),
	.w1(32'hbb9a1216),
	.w2(32'hbaff85ee),
	.w3(32'hbc365ce7),
	.w4(32'hbc064e3f),
	.w5(32'hbb3dfa63),
	.w6(32'h3bd76b3b),
	.w7(32'hba9a7793),
	.w8(32'hbb480712),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34ba54),
	.w1(32'hbbead442),
	.w2(32'hbb634797),
	.w3(32'h3b95b546),
	.w4(32'h3abf290f),
	.w5(32'h3b352bd9),
	.w6(32'h3c0dd28c),
	.w7(32'h3b2f58b9),
	.w8(32'h3b5a9044),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fce6f),
	.w1(32'h3c8e2000),
	.w2(32'h3b1d9c2d),
	.w3(32'hbc73c7af),
	.w4(32'hbc123c1b),
	.w5(32'hbc0b8418),
	.w6(32'hbb9d821e),
	.w7(32'hbb069ad8),
	.w8(32'hbc3e930c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbafdc),
	.w1(32'h3c982f5f),
	.w2(32'h3c2704c1),
	.w3(32'hbbe2860c),
	.w4(32'hbc04766e),
	.w5(32'h3aabc2b6),
	.w6(32'hbb6a2842),
	.w7(32'hbb437f2d),
	.w8(32'hb96be4f0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36dd29),
	.w1(32'hbbb2b3cf),
	.w2(32'h3ae4245a),
	.w3(32'hbb346801),
	.w4(32'h3bc0d13e),
	.w5(32'hbc69896d),
	.w6(32'hbb081a5c),
	.w7(32'hbb736492),
	.w8(32'hbc095dfe),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca90d82),
	.w1(32'hbc03bea7),
	.w2(32'hbcae1285),
	.w3(32'h3ad21b1f),
	.w4(32'h3bc998db),
	.w5(32'h3c32a2bd),
	.w6(32'h3bb651a0),
	.w7(32'h36ceb3fe),
	.w8(32'h3a40aaea),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2993a),
	.w1(32'hbc00d464),
	.w2(32'h3aa07fa9),
	.w3(32'hba9b549d),
	.w4(32'h3b86dcd9),
	.w5(32'hbba61bf9),
	.w6(32'hbc3f71ec),
	.w7(32'hbb946a52),
	.w8(32'hbc0d923c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5dd7),
	.w1(32'h3c33926e),
	.w2(32'hbb934dd3),
	.w3(32'hbb9066f4),
	.w4(32'hbbf463a2),
	.w5(32'h3aed6424),
	.w6(32'h38f6b6d0),
	.w7(32'hbbf0e029),
	.w8(32'hbbf21c5a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c231f),
	.w1(32'h3a9a0856),
	.w2(32'hbc43d80c),
	.w3(32'h3c4e9369),
	.w4(32'h3a6cf3a3),
	.w5(32'hb88cb26f),
	.w6(32'hbb314a5d),
	.w7(32'hbca23462),
	.w8(32'h3c074aff),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c810a96),
	.w1(32'h3b8f7866),
	.w2(32'h3c1f2e2b),
	.w3(32'hbbaf81d3),
	.w4(32'hbb6027ba),
	.w5(32'hbc6fd1d6),
	.w6(32'hbb7fa7f5),
	.w7(32'h3b103033),
	.w8(32'hbbc3e270),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97182a),
	.w1(32'hbc266ed3),
	.w2(32'hbb32106e),
	.w3(32'hbc2e20e4),
	.w4(32'hba7fb959),
	.w5(32'hba077826),
	.w6(32'hbb6ca6a5),
	.w7(32'h3a5bf246),
	.w8(32'hbaf07eb0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9c8b9),
	.w1(32'hbadc2216),
	.w2(32'h3b65c459),
	.w3(32'hb9349821),
	.w4(32'h3aef3ba1),
	.w5(32'h3a9145d6),
	.w6(32'hba946438),
	.w7(32'h39aca1fb),
	.w8(32'hbb49281b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912f9b),
	.w1(32'hbc08d5aa),
	.w2(32'hbbb9f150),
	.w3(32'hbbe4e3a5),
	.w4(32'hbbb33fc3),
	.w5(32'hbb1d62c7),
	.w6(32'hbbb79eac),
	.w7(32'hbbb702fc),
	.w8(32'hbac8b4ce),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbade2a9),
	.w1(32'hbabf081e),
	.w2(32'hba64876d),
	.w3(32'h38a83b74),
	.w4(32'h3b4ec30c),
	.w5(32'h3b099e77),
	.w6(32'h3934044b),
	.w7(32'hbb13dfae),
	.w8(32'h3b32b667),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b08db),
	.w1(32'h3a9c2adb),
	.w2(32'h3b8f231f),
	.w3(32'hba4d45d5),
	.w4(32'hbaa8b1ba),
	.w5(32'h3b32e97b),
	.w6(32'hbb0ca6ec),
	.w7(32'hbaa8dad1),
	.w8(32'h39adb563),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fafbc),
	.w1(32'hbac4567d),
	.w2(32'h3a8e3d84),
	.w3(32'hbb41aa3d),
	.w4(32'hbae40285),
	.w5(32'hba1d83a0),
	.w6(32'hbb21a4dc),
	.w7(32'hbaa2c4a2),
	.w8(32'hbb1a852e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d3bcf),
	.w1(32'h3a5c3efb),
	.w2(32'hbb2ad88e),
	.w3(32'hb96b34d1),
	.w4(32'hba6babba),
	.w5(32'hbb155741),
	.w6(32'h39ce24af),
	.w7(32'hbabe1a85),
	.w8(32'h3b046739),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65018e),
	.w1(32'hbba55887),
	.w2(32'hbbb66b87),
	.w3(32'hbae91fbd),
	.w4(32'hbae64ff0),
	.w5(32'hbb85193a),
	.w6(32'hb99a9eea),
	.w7(32'hbb96a0ea),
	.w8(32'h3a131c4e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7dd36),
	.w1(32'h38ca2df4),
	.w2(32'h3a2589bb),
	.w3(32'h3b230060),
	.w4(32'hba109561),
	.w5(32'hbabc996e),
	.w6(32'h3ade0440),
	.w7(32'hbb08973c),
	.w8(32'hba15a6e7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e1aca),
	.w1(32'hb9a5ef00),
	.w2(32'h3a4ad8de),
	.w3(32'hbb26e93d),
	.w4(32'hbb0e1d5c),
	.w5(32'hb9a8ce7f),
	.w6(32'h3b0b2a20),
	.w7(32'hb898723a),
	.w8(32'hba8e4aea),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f92fa),
	.w1(32'hbab0554d),
	.w2(32'hbab7ad42),
	.w3(32'hbab7a5a4),
	.w4(32'h3a42f387),
	.w5(32'hbabcf1cb),
	.w6(32'hbad6931a),
	.w7(32'hba87e37f),
	.w8(32'hbae92038),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcdaac),
	.w1(32'h37cbafc4),
	.w2(32'h3b74f88f),
	.w3(32'hbb3ef3eb),
	.w4(32'hba15fc04),
	.w5(32'h3aad580e),
	.w6(32'hbb7b17c9),
	.w7(32'h39205237),
	.w8(32'hb8e08184),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926b7a6),
	.w1(32'h3ac45584),
	.w2(32'h3b6d0587),
	.w3(32'hb999af68),
	.w4(32'h3b2499c2),
	.w5(32'h3b89b124),
	.w6(32'h3a2b937c),
	.w7(32'h3b1f9a59),
	.w8(32'h3b94024e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43c10e),
	.w1(32'hba2adcc1),
	.w2(32'hba15e8ca),
	.w3(32'h398b8091),
	.w4(32'h398764c8),
	.w5(32'h392ea76e),
	.w6(32'h3b20813d),
	.w7(32'h3b5f4146),
	.w8(32'hbb2bc522),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34a8f8),
	.w1(32'hb93b9f91),
	.w2(32'h3a376779),
	.w3(32'hbaa28239),
	.w4(32'h3abbb158),
	.w5(32'h3b01b607),
	.w6(32'hbaa07c1e),
	.w7(32'h3a3f38c1),
	.w8(32'h386f465c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb790dd4e),
	.w1(32'hbac2e314),
	.w2(32'h3b01afb7),
	.w3(32'h39b05b0d),
	.w4(32'h3af0a417),
	.w5(32'h3b40036b),
	.w6(32'hbb41466a),
	.w7(32'h3a91d75a),
	.w8(32'h397d8b72),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d9abe),
	.w1(32'hbab2c92c),
	.w2(32'hba753c65),
	.w3(32'h38c9242f),
	.w4(32'hba5681f2),
	.w5(32'hba4f071d),
	.w6(32'hbb42b4df),
	.w7(32'hbae1e70d),
	.w8(32'hbb0a3ebf),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40ad9b),
	.w1(32'h39de1ece),
	.w2(32'hbb0dbe13),
	.w3(32'h3ab09014),
	.w4(32'hba6b928e),
	.w5(32'h3b0c041b),
	.w6(32'h3a93bb3e),
	.w7(32'hb92b9c30),
	.w8(32'hbaa67641),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba860e8c),
	.w1(32'hba062817),
	.w2(32'h39ab6a12),
	.w3(32'h39ba0f45),
	.w4(32'h38f2d1f6),
	.w5(32'hb92f846c),
	.w6(32'hbb202f8a),
	.w7(32'hb8784a02),
	.w8(32'hba7c3935),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b9a25),
	.w1(32'h39a91489),
	.w2(32'hb9d1076f),
	.w3(32'h3a0e739f),
	.w4(32'hba373c1a),
	.w5(32'hbbcf51bf),
	.w6(32'h395b6837),
	.w7(32'hba244838),
	.w8(32'hbb18f5de),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387cc1ed),
	.w1(32'h3a0bc410),
	.w2(32'h3ae80e03),
	.w3(32'hbb3619b0),
	.w4(32'hbb0d7aff),
	.w5(32'hba9d0b99),
	.w6(32'hba9f45e4),
	.w7(32'hbae66640),
	.w8(32'hbb1ce075),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb113453),
	.w1(32'hbb565cfa),
	.w2(32'h39ee5493),
	.w3(32'hbb6b8e01),
	.w4(32'hba9c1e6a),
	.w5(32'hbb15cc42),
	.w6(32'hbb7423eb),
	.w7(32'hbaea3c06),
	.w8(32'hbba423ff),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ded12),
	.w1(32'hbb228827),
	.w2(32'h39c1a59e),
	.w3(32'hbb728b2d),
	.w4(32'hbb5c7e3c),
	.w5(32'h3b6d05c0),
	.w6(32'hbc0c65d3),
	.w7(32'hbb489aa6),
	.w8(32'h39f96ba6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f38d13),
	.w1(32'h3a9db165),
	.w2(32'h3a0e53a8),
	.w3(32'h3a6fe3f4),
	.w4(32'h3a4a1338),
	.w5(32'hb9e67ab0),
	.w6(32'hbad7da29),
	.w7(32'h3a05e509),
	.w8(32'hba9b1fa8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba753205),
	.w1(32'hb9505875),
	.w2(32'hbabfae2d),
	.w3(32'hba31186a),
	.w4(32'hbab6537f),
	.w5(32'h3ab5602d),
	.w6(32'hbaa4ca7a),
	.w7(32'hbac8fc50),
	.w8(32'h3aff5c4a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945af8b),
	.w1(32'h3abf879f),
	.w2(32'h3b381a3b),
	.w3(32'h3acd0ca5),
	.w4(32'h3ad791c6),
	.w5(32'h3a439dfb),
	.w6(32'h3a77a244),
	.w7(32'h3b521f47),
	.w8(32'h3b0c6c45),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add22a6),
	.w1(32'h397921c0),
	.w2(32'h3b0be566),
	.w3(32'hb9ca69db),
	.w4(32'h39a2c1b4),
	.w5(32'h3a456ca0),
	.w6(32'hbac94d66),
	.w7(32'h3a969f1a),
	.w8(32'h3aa0a6ef),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06b0b9),
	.w1(32'h3a3e36a6),
	.w2(32'h3ac0ee4c),
	.w3(32'h3850db35),
	.w4(32'h39497e5e),
	.w5(32'hbb337126),
	.w6(32'hba1ad41b),
	.w7(32'h3a628420),
	.w8(32'hbae3e096),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b2f4f),
	.w1(32'h3a9e7b87),
	.w2(32'h3a47f08b),
	.w3(32'hb8674b49),
	.w4(32'hba133555),
	.w5(32'hb8fd7229),
	.w6(32'hba19512f),
	.w7(32'hbad73d8a),
	.w8(32'h3ac6814b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a021641),
	.w1(32'hb999bf33),
	.w2(32'hba4d764a),
	.w3(32'h389fb733),
	.w4(32'hba5b30ff),
	.w5(32'h3a0fd133),
	.w6(32'h3b1d3aa9),
	.w7(32'h38df2a46),
	.w8(32'hba032fd8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb303166),
	.w1(32'hba7b75c2),
	.w2(32'hbadd5ab9),
	.w3(32'h3996221e),
	.w4(32'hba5d9f63),
	.w5(32'h3b8c60c5),
	.w6(32'hb9d2fccc),
	.w7(32'hbacf9777),
	.w8(32'h3b242a0c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c145c4),
	.w1(32'hba362989),
	.w2(32'h3b3a644e),
	.w3(32'h3abe1052),
	.w4(32'h3ad35337),
	.w5(32'hba7434bb),
	.w6(32'hb8e034fa),
	.w7(32'h3a3ffdae),
	.w8(32'h3aa035f2),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b223a93),
	.w1(32'hb8e2b60d),
	.w2(32'h3acbee85),
	.w3(32'hba5cc2e3),
	.w4(32'hb9d12137),
	.w5(32'hba60aeaa),
	.w6(32'hba9e74d2),
	.w7(32'h39eb23a7),
	.w8(32'hbab5604b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae7df1),
	.w1(32'hb9429b04),
	.w2(32'hbafba7d4),
	.w3(32'hbb129325),
	.w4(32'hbb641446),
	.w5(32'hba8da6bb),
	.w6(32'hbb2bf500),
	.w7(32'hba2ded7e),
	.w8(32'hbad741fb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba038714),
	.w1(32'hba6fd573),
	.w2(32'hba338bcd),
	.w3(32'hba342f8b),
	.w4(32'hba84757f),
	.w5(32'hbb6d544d),
	.w6(32'hbb36fb44),
	.w7(32'hba938b4e),
	.w8(32'hbb04e55e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7a0c),
	.w1(32'hbb84e1ef),
	.w2(32'hbb308ff1),
	.w3(32'hbbcaec5a),
	.w4(32'hbadd6490),
	.w5(32'hb94d5b7b),
	.w6(32'hbbd1c48b),
	.w7(32'hbb64d69d),
	.w8(32'hba46da76),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26377d),
	.w1(32'h39dee833),
	.w2(32'hb9c74e6b),
	.w3(32'hba763ae3),
	.w4(32'hb99d4adb),
	.w5(32'hb9f5346b),
	.w6(32'h3a7c8040),
	.w7(32'h3ac4b60e),
	.w8(32'h3a290658),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb938ca1),
	.w1(32'hbb79b00b),
	.w2(32'hbb752cb8),
	.w3(32'hbb5d16f5),
	.w4(32'hbb879e16),
	.w5(32'hba867d6f),
	.w6(32'hbaff7962),
	.w7(32'hbb8155a4),
	.w8(32'hbb194adf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38ca65),
	.w1(32'h3a0db414),
	.w2(32'h3a836ecd),
	.w3(32'hbac5b353),
	.w4(32'hbb02d183),
	.w5(32'h3ab59b02),
	.w6(32'hba9a9ad8),
	.w7(32'hbab7d0de),
	.w8(32'hba0cdc03),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb663fc0),
	.w1(32'hbafd3b36),
	.w2(32'h38aa2eae),
	.w3(32'hba487ed3),
	.w4(32'h39ada105),
	.w5(32'h3a6bdc6c),
	.w6(32'hbab25fa5),
	.w7(32'hba4b1540),
	.w8(32'h3ac8eb78),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49f8d4),
	.w1(32'hbaccba8f),
	.w2(32'hbac6f201),
	.w3(32'hbb3d426b),
	.w4(32'hbb3786d8),
	.w5(32'hbb023c95),
	.w6(32'hbb0606ef),
	.w7(32'hba66467e),
	.w8(32'hba5fd6ce),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3e0d5),
	.w1(32'hba290e01),
	.w2(32'hba50a578),
	.w3(32'hbb01aaee),
	.w4(32'hbab5da79),
	.w5(32'h3a8817cf),
	.w6(32'hba104403),
	.w7(32'hba6e7d61),
	.w8(32'hba8998d1),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b8168),
	.w1(32'h3aa44a01),
	.w2(32'hbb43b77c),
	.w3(32'hba2d50c2),
	.w4(32'hbb2f018c),
	.w5(32'hba607c7a),
	.w6(32'hbab42dca),
	.w7(32'hbab19f87),
	.w8(32'hbab853c2),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f02e9),
	.w1(32'hba8e1335),
	.w2(32'h3a521fce),
	.w3(32'hba36d9b8),
	.w4(32'hb9c04ed5),
	.w5(32'hba3c9b49),
	.w6(32'hbae1402e),
	.w7(32'hb79636b2),
	.w8(32'hb9eb05b1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af5c7),
	.w1(32'hbb21a84e),
	.w2(32'h3a04ecea),
	.w3(32'hbb25d6ab),
	.w4(32'h3b0cd600),
	.w5(32'h3add286f),
	.w6(32'h3a7a18b6),
	.w7(32'h3a7696bf),
	.w8(32'h395ab5db),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb155c55),
	.w1(32'hbb0333ac),
	.w2(32'hbb35751c),
	.w3(32'hba94f438),
	.w4(32'hbb32867c),
	.w5(32'hbb0258c9),
	.w6(32'hbaf34b28),
	.w7(32'hba89c8d0),
	.w8(32'hba1dc827),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b040e76),
	.w1(32'hbaa08602),
	.w2(32'hba1e1a9a),
	.w3(32'hb9c62cd2),
	.w4(32'h3a1724c0),
	.w5(32'h38d2231d),
	.w6(32'hba713581),
	.w7(32'h396517e8),
	.w8(32'h3a16e9e9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafcfea),
	.w1(32'hba9f7099),
	.w2(32'h38e36635),
	.w3(32'hba085b6d),
	.w4(32'h39fa819b),
	.w5(32'hb9409f88),
	.w6(32'hb9ba5cbf),
	.w7(32'hb86fbf42),
	.w8(32'hb9fd37ad),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98280fa),
	.w1(32'hbab21a4e),
	.w2(32'hba14007d),
	.w3(32'hba838a45),
	.w4(32'hba8f6a6d),
	.w5(32'h3ac86eab),
	.w6(32'hbaef2c31),
	.w7(32'hbac357dc),
	.w8(32'h3ba2c7b8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20b191),
	.w1(32'hbae4d11a),
	.w2(32'hbb002b69),
	.w3(32'h39ea6fea),
	.w4(32'h3b2393fe),
	.w5(32'hbb017b1a),
	.w6(32'h3b31dc47),
	.w7(32'h3ac332e4),
	.w8(32'hba1ebf3f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8527e4),
	.w1(32'hb90bc639),
	.w2(32'h3aaa5103),
	.w3(32'hb9b9e1f2),
	.w4(32'hb99903f7),
	.w5(32'h3a593aa4),
	.w6(32'h3a17d3cc),
	.w7(32'hb978d40e),
	.w8(32'h3aa2bcc7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa48c98),
	.w1(32'h3a195069),
	.w2(32'h3a1c4dbf),
	.w3(32'h39f47c97),
	.w4(32'hba6cf8e4),
	.w5(32'h37f1d2b9),
	.w6(32'h39cdbe28),
	.w7(32'h3a9e0866),
	.w8(32'hb95858a0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba062132),
	.w1(32'hb884f7b6),
	.w2(32'hb9e4b2ce),
	.w3(32'hbaa9bb18),
	.w4(32'hbad7e0fb),
	.w5(32'h3a910c90),
	.w6(32'hb79fdc49),
	.w7(32'hba82e3a0),
	.w8(32'h3a6a4e10),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974898d),
	.w1(32'h3aa0b726),
	.w2(32'h3a3705e5),
	.w3(32'h3ad3d0c1),
	.w4(32'h3aad593d),
	.w5(32'h3ac25562),
	.w6(32'h3a9dcbfa),
	.w7(32'h3a078fdd),
	.w8(32'hba26d6fa),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51963f),
	.w1(32'hbaf9810a),
	.w2(32'hba9594d0),
	.w3(32'hbaf3f9ba),
	.w4(32'hbb1ffc6f),
	.w5(32'hba92c64b),
	.w6(32'hbb1eb8d5),
	.w7(32'hbb9bdfac),
	.w8(32'hbaec9cf9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72a1f7),
	.w1(32'hb9099b5b),
	.w2(32'h3a4db21a),
	.w3(32'hbaad2c2a),
	.w4(32'hbb1752d2),
	.w5(32'h3ab8d764),
	.w6(32'hbb2b18ca),
	.w7(32'h38f42d72),
	.w8(32'h3a133e4a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3ca75),
	.w1(32'hb9dd52ff),
	.w2(32'hba938527),
	.w3(32'h3a3862b5),
	.w4(32'h3a0bba04),
	.w5(32'hbb023971),
	.w6(32'h3abdd616),
	.w7(32'hba915569),
	.w8(32'hba629766),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a008014),
	.w1(32'h38120eac),
	.w2(32'hb941e70f),
	.w3(32'h392fa200),
	.w4(32'h3a9cc780),
	.w5(32'h3b996e81),
	.w6(32'h3a18dfca),
	.w7(32'h3a2ef43c),
	.w8(32'h3b5e538f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ac6fb),
	.w1(32'hba95f76e),
	.w2(32'h3b2b8ca9),
	.w3(32'hbaea97db),
	.w4(32'h3ae3f667),
	.w5(32'hbb6a297c),
	.w6(32'hbac13366),
	.w7(32'h3b0a79f2),
	.w8(32'hba7afad2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c039e7),
	.w1(32'h3a7854c9),
	.w2(32'h3a737abd),
	.w3(32'h3a26ccbd),
	.w4(32'h3a2a5617),
	.w5(32'h39dffeaa),
	.w6(32'h3b358ccb),
	.w7(32'h3aa080d5),
	.w8(32'h3a867200),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62525d),
	.w1(32'h39382831),
	.w2(32'h3a860212),
	.w3(32'h3a4caa3d),
	.w4(32'h3a7ef163),
	.w5(32'h3b050d62),
	.w6(32'h393fd608),
	.w7(32'h3a791c49),
	.w8(32'h3ad5ac58),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37337074),
	.w1(32'hba07efc8),
	.w2(32'hba2d3d28),
	.w3(32'hba3e97f2),
	.w4(32'hba44ab7e),
	.w5(32'h3b0dd191),
	.w6(32'hb9b13504),
	.w7(32'hbada3b1a),
	.w8(32'h3b0ddc34),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af477f7),
	.w1(32'h3b2cdb78),
	.w2(32'h3979e185),
	.w3(32'h3ae01847),
	.w4(32'hba0164b8),
	.w5(32'h39493b43),
	.w6(32'h398733f6),
	.w7(32'h3b03249f),
	.w8(32'hb9d215d1),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69ba4f),
	.w1(32'hbb170773),
	.w2(32'hb9cb4181),
	.w3(32'h3a53b37d),
	.w4(32'h39b3cece),
	.w5(32'hba9c0cd8),
	.w6(32'hbb9534b4),
	.w7(32'hbb545f1b),
	.w8(32'h394f448f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc177b),
	.w1(32'hba832817),
	.w2(32'hb9b8479f),
	.w3(32'hbac8858c),
	.w4(32'hba7cf09d),
	.w5(32'h39b6ae71),
	.w6(32'hbad59c86),
	.w7(32'hba06a9fc),
	.w8(32'h3a21b432),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ef11f),
	.w1(32'h3a9d9a5d),
	.w2(32'h39f0d7a1),
	.w3(32'hbae44868),
	.w4(32'hbaa9c7f2),
	.w5(32'h3b421e48),
	.w6(32'hb98da7ae),
	.w7(32'hbaa796d7),
	.w8(32'hb9b25190),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb045d56),
	.w1(32'hba0fcfc7),
	.w2(32'hba1ad7f7),
	.w3(32'hb904e034),
	.w4(32'h39fab755),
	.w5(32'hba21ad03),
	.w6(32'h3a357126),
	.w7(32'hba6e13a9),
	.w8(32'h3929fef0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b426967),
	.w1(32'h3adbfb47),
	.w2(32'h3b0a3ec7),
	.w3(32'h3b49aded),
	.w4(32'h3abd6cf0),
	.w5(32'h3adb3c7c),
	.w6(32'h38e61502),
	.w7(32'hba65dbbf),
	.w8(32'h3a15746a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936be69),
	.w1(32'h3a334c5f),
	.w2(32'h38a6ad7b),
	.w3(32'hba847f5d),
	.w4(32'hba9efa31),
	.w5(32'h3ab41dc4),
	.w6(32'h3a825f68),
	.w7(32'hb8c18322),
	.w8(32'h3a8e72de),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac83fae),
	.w1(32'h3accb971),
	.w2(32'h3b736e5f),
	.w3(32'h3aa47c12),
	.w4(32'h3adeb3e4),
	.w5(32'h399d8667),
	.w6(32'hbac84fae),
	.w7(32'h3a4f3afd),
	.w8(32'hba1cf42b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25bcb8),
	.w1(32'hbb1f3f95),
	.w2(32'hbb951bed),
	.w3(32'hbaafb716),
	.w4(32'hbb1d126f),
	.w5(32'hba963208),
	.w6(32'h3a411cd3),
	.w7(32'hbb69ce7f),
	.w8(32'hbaa18ee5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e3328),
	.w1(32'hbb0e7c75),
	.w2(32'hbb22fc90),
	.w3(32'hbb209b5e),
	.w4(32'hb6540655),
	.w5(32'hbac2d32a),
	.w6(32'hbb767cbc),
	.w7(32'hbb211167),
	.w8(32'hbb7bc951),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a124be),
	.w1(32'hba8dbca6),
	.w2(32'hbaa9af76),
	.w3(32'h39aa8aab),
	.w4(32'hba8112ed),
	.w5(32'h3b0bf484),
	.w6(32'h3a3d60ce),
	.w7(32'hbaa3f7ba),
	.w8(32'h3af22827),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4b281),
	.w1(32'hb94046a2),
	.w2(32'h3a43a773),
	.w3(32'h3a970118),
	.w4(32'h3b198729),
	.w5(32'h3abf79e0),
	.w6(32'hbad10387),
	.w7(32'hba2f3c8b),
	.w8(32'hb9754012),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed1ba),
	.w1(32'hbabd7d40),
	.w2(32'h39c5cad1),
	.w3(32'hba8d1ffa),
	.w4(32'h3a4d47a7),
	.w5(32'hbafa4b06),
	.w6(32'h3aae87ce),
	.w7(32'h39f9258e),
	.w8(32'hbb81dcf0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabd9ec),
	.w1(32'hbb99d9ac),
	.w2(32'hbb491eca),
	.w3(32'hbb78fecd),
	.w4(32'hbb84ca44),
	.w5(32'hbaac3985),
	.w6(32'hbb91ae0f),
	.w7(32'hbb9117e3),
	.w8(32'hb99ff9f4),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb354e),
	.w1(32'hbabb8f4c),
	.w2(32'hbb48efff),
	.w3(32'hbab51a9a),
	.w4(32'hb7cc7aa1),
	.w5(32'hbb034ff3),
	.w6(32'hb90b7066),
	.w7(32'hbb3de738),
	.w8(32'hbb05afe6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8984f4),
	.w1(32'hbadb093c),
	.w2(32'hbaf1a63a),
	.w3(32'hbb7feb2c),
	.w4(32'hbb5b5623),
	.w5(32'h3b08f02c),
	.w6(32'hbb184ca3),
	.w7(32'hbb821337),
	.w8(32'h3b02823a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b617711),
	.w1(32'h3b2d0006),
	.w2(32'h3b1b884f),
	.w3(32'h3a93f84e),
	.w4(32'h3a82f024),
	.w5(32'h3b17c5ef),
	.w6(32'h39980c0a),
	.w7(32'h3aab7c53),
	.w8(32'h39dfa184),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47530f),
	.w1(32'h3a62c0cc),
	.w2(32'h3acff5ac),
	.w3(32'hb91ecbeb),
	.w4(32'hba260397),
	.w5(32'hba757486),
	.w6(32'hb892deda),
	.w7(32'h3a1eb3f3),
	.w8(32'hbadade15),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d3a56b),
	.w1(32'h383515ea),
	.w2(32'hba69b2a4),
	.w3(32'hb9ad9af9),
	.w4(32'hbabc70a1),
	.w5(32'h3a923382),
	.w6(32'hba35c3de),
	.w7(32'hba985a8f),
	.w8(32'hba87af76),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b1329),
	.w1(32'hbb613d2c),
	.w2(32'hb9af8814),
	.w3(32'hbb5e7366),
	.w4(32'hba5ecbe2),
	.w5(32'hbb806e6b),
	.w6(32'hbb24f5cc),
	.w7(32'hba0cf80f),
	.w8(32'hbb6cad8c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36ada0),
	.w1(32'hba66204f),
	.w2(32'hbaf3591e),
	.w3(32'hbad542f3),
	.w4(32'hbac4666c),
	.w5(32'h3aa34a59),
	.w6(32'hb999d584),
	.w7(32'hbb2df7c8),
	.w8(32'hbac9de65),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dac3e),
	.w1(32'h398075cf),
	.w2(32'hbb059ab3),
	.w3(32'h3a16faee),
	.w4(32'hba3d4530),
	.w5(32'hba6a81db),
	.w6(32'h3a7de99c),
	.w7(32'hbae71ecf),
	.w8(32'h3a04e882),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd904f),
	.w1(32'hba34fb5d),
	.w2(32'hbb678789),
	.w3(32'h3a553fb3),
	.w4(32'hbab21b9b),
	.w5(32'hba01ea3a),
	.w6(32'hbaa2a602),
	.w7(32'hbb7b309a),
	.w8(32'h3a65d001),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39819800),
	.w1(32'h3aa733d6),
	.w2(32'hba512ff2),
	.w3(32'h3a41fbc7),
	.w4(32'hb6e9e303),
	.w5(32'h39ec46e8),
	.w6(32'h3adc890e),
	.w7(32'hba5d7512),
	.w8(32'h3adaf8c0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8f3ef),
	.w1(32'h392a48bd),
	.w2(32'hb9e11bc3),
	.w3(32'hb897777d),
	.w4(32'hb8fbddff),
	.w5(32'h38ff97ea),
	.w6(32'h3a407062),
	.w7(32'h3a999407),
	.w8(32'hb8cb9fbd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83f7a7),
	.w1(32'hba8e5bb3),
	.w2(32'h397c8c80),
	.w3(32'hb991af76),
	.w4(32'h39a46be1),
	.w5(32'h3ae7fc75),
	.w6(32'h3b04ce8a),
	.w7(32'h37976378),
	.w8(32'hb96af14f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa26d7c),
	.w1(32'hbaaed944),
	.w2(32'h3847dc10),
	.w3(32'h39851a2e),
	.w4(32'h3b0537c1),
	.w5(32'h3ac71c9f),
	.w6(32'hba386768),
	.w7(32'h3a466652),
	.w8(32'h3aacf271),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a48cb2),
	.w1(32'hb858c0c3),
	.w2(32'hbad7a34a),
	.w3(32'h37927396),
	.w4(32'hbaa0be0e),
	.w5(32'h396741e8),
	.w6(32'hba59c0c0),
	.w7(32'hbaa9888a),
	.w8(32'hba226e34),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada354d),
	.w1(32'h3b25cbf9),
	.w2(32'h3b704991),
	.w3(32'hba2059c9),
	.w4(32'h39ac10b1),
	.w5(32'hb8efb70e),
	.w6(32'hba7c1f90),
	.w7(32'hb93a48d6),
	.w8(32'h3a048510),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0980cf),
	.w1(32'h3ade007c),
	.w2(32'h3b30938e),
	.w3(32'hb97e4b30),
	.w4(32'h3ad338e8),
	.w5(32'hb99e724a),
	.w6(32'h3ac0d2d3),
	.w7(32'h3b2a5c2b),
	.w8(32'h3b27130a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38ffe7),
	.w1(32'hb8c05890),
	.w2(32'hb9ca8852),
	.w3(32'h39824f91),
	.w4(32'h3a63092a),
	.w5(32'hbafb6acf),
	.w6(32'h3ad9c976),
	.w7(32'hb9f131f2),
	.w8(32'hb96ca52e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae6ee8),
	.w1(32'h3a48a61f),
	.w2(32'hb9d4938a),
	.w3(32'hbb2a386d),
	.w4(32'hbadc9705),
	.w5(32'h39b156ef),
	.w6(32'hbb22f7c6),
	.w7(32'hbb34f0a3),
	.w8(32'h3aa290c5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc57a5),
	.w1(32'hba16775f),
	.w2(32'hb9a2ef37),
	.w3(32'hba55afcd),
	.w4(32'h39e4f2b2),
	.w5(32'h39ecfccd),
	.w6(32'h3a8b451a),
	.w7(32'h395cd9d1),
	.w8(32'h3b20aef4),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefa628),
	.w1(32'h3b05674e),
	.w2(32'h3a1b1d2d),
	.w3(32'hba2583ee),
	.w4(32'hba921019),
	.w5(32'hba5e2efe),
	.w6(32'h3a88dcbb),
	.w7(32'hba5fa069),
	.w8(32'h38f5c143),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4ebea),
	.w1(32'hba38a2a7),
	.w2(32'hb9ae7ca8),
	.w3(32'hb998ffbe),
	.w4(32'hb97bfb0f),
	.w5(32'h38fab33d),
	.w6(32'hbacd27aa),
	.w7(32'hbb05181e),
	.w8(32'h39bb25e1),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1de346),
	.w1(32'hba36c5d6),
	.w2(32'hbb188441),
	.w3(32'h3a7a0e16),
	.w4(32'hb99db5f0),
	.w5(32'hbb775ac0),
	.w6(32'h394636d5),
	.w7(32'hba9c06b6),
	.w8(32'hbb6fccf5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24293c),
	.w1(32'hbb4244c5),
	.w2(32'hba36e70d),
	.w3(32'hbbaa22ed),
	.w4(32'hbb529974),
	.w5(32'h3b23d135),
	.w6(32'hbb80cfda),
	.w7(32'hbb51eda7),
	.w8(32'h3a9bc7e2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba186f9d),
	.w1(32'hba505439),
	.w2(32'hb9db8be9),
	.w3(32'hbb203b37),
	.w4(32'hb982ee14),
	.w5(32'h3b2202f3),
	.w6(32'hb96f3564),
	.w7(32'hba1aad6c),
	.w8(32'h3a606b03),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab05148),
	.w1(32'hba981d0d),
	.w2(32'h39f335dd),
	.w3(32'hbaef24ee),
	.w4(32'hbae74125),
	.w5(32'h38fa7e75),
	.w6(32'h3a242ba5),
	.w7(32'hba4022ad),
	.w8(32'h3a708892),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21e240),
	.w1(32'hbad425b6),
	.w2(32'h386879e1),
	.w3(32'h3a890f83),
	.w4(32'hb9a2615c),
	.w5(32'h3aaa22fb),
	.w6(32'hbabbf1a4),
	.w7(32'hbaee641f),
	.w8(32'hba754e28),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7fc39),
	.w1(32'hb8f4f393),
	.w2(32'h39a1f0f0),
	.w3(32'h3a823d6e),
	.w4(32'hba370085),
	.w5(32'h3b431861),
	.w6(32'h3a854e14),
	.w7(32'h39e68c8d),
	.w8(32'h3b1a70b4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09120b),
	.w1(32'h38a30ab3),
	.w2(32'h3a351479),
	.w3(32'hb7a33ea9),
	.w4(32'h3a510a49),
	.w5(32'hbb16bda3),
	.w6(32'h3a9405af),
	.w7(32'h3af81550),
	.w8(32'hba210ee7),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f9dff),
	.w1(32'hba7d86b7),
	.w2(32'h3a89d186),
	.w3(32'hba207b1b),
	.w4(32'hba08597a),
	.w5(32'h3aad1359),
	.w6(32'hbb1aa223),
	.w7(32'h3936396f),
	.w8(32'h3a474d0a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1459f5),
	.w1(32'hb7875147),
	.w2(32'hb9f07bbf),
	.w3(32'h3adbee7a),
	.w4(32'h39ecde27),
	.w5(32'h3a653ebd),
	.w6(32'h3a1408d0),
	.w7(32'hb9a52cf1),
	.w8(32'h39b94b01),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58c5f1),
	.w1(32'h3aa357c7),
	.w2(32'h39d84257),
	.w3(32'h3b2e2506),
	.w4(32'h3b4a6d15),
	.w5(32'h3a25f718),
	.w6(32'h3b41b938),
	.w7(32'h3b37f36c),
	.w8(32'h3a0d0887),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff57d5),
	.w1(32'hba960de7),
	.w2(32'hb9ff9435),
	.w3(32'hba2a9e45),
	.w4(32'h3ab18b44),
	.w5(32'hbab12e7b),
	.w6(32'hbb0c38ed),
	.w7(32'hb8c1e869),
	.w8(32'hbb43d6ac),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad724cb),
	.w1(32'hba6db088),
	.w2(32'hbacb8a34),
	.w3(32'hba9e01a6),
	.w4(32'hba9b61b7),
	.w5(32'hbb091113),
	.w6(32'hb9faa02f),
	.w7(32'hbaf4861f),
	.w8(32'hba922623),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab02769),
	.w1(32'h380a5165),
	.w2(32'hba329853),
	.w3(32'hbafb9658),
	.w4(32'h39a55925),
	.w5(32'h38f37b21),
	.w6(32'h3a66c1fe),
	.w7(32'h3ae793d6),
	.w8(32'h3a088575),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb835ef2b),
	.w1(32'h39037168),
	.w2(32'h3a8d5d92),
	.w3(32'hbb2db37d),
	.w4(32'hb9621abb),
	.w5(32'h3b30a21f),
	.w6(32'hbac7c9f0),
	.w7(32'hb9873269),
	.w8(32'h3a804858),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb229a4b),
	.w1(32'h3a3c5944),
	.w2(32'h3b112fe3),
	.w3(32'h3a93fa7b),
	.w4(32'hbb1c666a),
	.w5(32'h3b3d47a9),
	.w6(32'h39abcb16),
	.w7(32'hba8a3802),
	.w8(32'h3ac40ca8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba371b40),
	.w1(32'hbafc920d),
	.w2(32'hba2717fb),
	.w3(32'h3a9d6727),
	.w4(32'h3a5a1493),
	.w5(32'h3a6877f5),
	.w6(32'hbaa51c7e),
	.w7(32'hb79338c3),
	.w8(32'h39095326),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f04bd),
	.w1(32'hb9cd2fd2),
	.w2(32'h3a7a53bf),
	.w3(32'hba1cea3d),
	.w4(32'hbaa1e8aa),
	.w5(32'hbb76be89),
	.w6(32'hba2b094e),
	.w7(32'hb9c4de3e),
	.w8(32'hbb00cbc0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d55f0),
	.w1(32'hb7e78326),
	.w2(32'h39f91470),
	.w3(32'hbb18051a),
	.w4(32'hbab9f22a),
	.w5(32'h3b017149),
	.w6(32'h398cf62e),
	.w7(32'hbae03dd1),
	.w8(32'h3ad1636e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb368acc),
	.w1(32'hbb1a7ef3),
	.w2(32'hba0a5e87),
	.w3(32'hbad5147b),
	.w4(32'hba9fba14),
	.w5(32'h3a64850f),
	.w6(32'hbb621732),
	.w7(32'hbb4a3706),
	.w8(32'hbab0c89c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fbf27),
	.w1(32'h3ab44581),
	.w2(32'h3955ffc2),
	.w3(32'hba9baf57),
	.w4(32'h3a41e0e7),
	.w5(32'h3a003db2),
	.w6(32'h3aef2009),
	.w7(32'h3a9c6c02),
	.w8(32'hbb17dea4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9566cc0),
	.w1(32'hbabaf18b),
	.w2(32'hbad53c83),
	.w3(32'hba941b93),
	.w4(32'hbb8fbc2d),
	.w5(32'hbb6c7dba),
	.w6(32'hbb2fec33),
	.w7(32'hbb1e043e),
	.w8(32'hbabbed0d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86906e),
	.w1(32'hb927badd),
	.w2(32'h3a0f097b),
	.w3(32'hba8200ea),
	.w4(32'hba2ab2a7),
	.w5(32'hba55d2e4),
	.w6(32'hbafa66b0),
	.w7(32'hbb05776b),
	.w8(32'hba98cc0f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab154b2),
	.w1(32'hbb14a295),
	.w2(32'hbaaa8efc),
	.w3(32'hba930c0a),
	.w4(32'hbaa1b2f7),
	.w5(32'h3a0df277),
	.w6(32'hba8bf9d2),
	.w7(32'hbab2663b),
	.w8(32'h3a11affd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39315225),
	.w1(32'h3afedb61),
	.w2(32'hb9c6b00d),
	.w3(32'h3b00911b),
	.w4(32'h398dafc8),
	.w5(32'hba30ec1f),
	.w6(32'h3adf9572),
	.w7(32'hbae5da8a),
	.w8(32'h3a80d3f1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560139),
	.w1(32'hbae3ca49),
	.w2(32'hbb4d7eb0),
	.w3(32'hbbe32c73),
	.w4(32'hbb449fa8),
	.w5(32'hbb0c48f9),
	.w6(32'hbbaf3f41),
	.w7(32'hbb03d1a1),
	.w8(32'hbac679b8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb062742),
	.w1(32'hbb396e19),
	.w2(32'hbb73905d),
	.w3(32'hbad72701),
	.w4(32'hb9b45243),
	.w5(32'hbb1aff73),
	.w6(32'hbaaf60a8),
	.w7(32'hbae576d3),
	.w8(32'h39213d15),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52dfe1),
	.w1(32'hbb637129),
	.w2(32'hbb3d4d88),
	.w3(32'hba0b32c5),
	.w4(32'h390bfbcb),
	.w5(32'h3aedf2c8),
	.w6(32'hbb2884c6),
	.w7(32'h3a889e19),
	.w8(32'h3a9e678c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0498dc),
	.w1(32'hbb1f5a70),
	.w2(32'h3a1bc9af),
	.w3(32'hbb8ad34f),
	.w4(32'hb8fe71f4),
	.w5(32'h3b20e0ba),
	.w6(32'hbb4ea7b0),
	.w7(32'hb98417fc),
	.w8(32'h3afb53cb),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ce0f6),
	.w1(32'h3a7f88e1),
	.w2(32'h3a644cec),
	.w3(32'h39928747),
	.w4(32'h381894dc),
	.w5(32'hb9a1005a),
	.w6(32'h3b11249e),
	.w7(32'h3a28aff9),
	.w8(32'hbb079f68),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8928bd),
	.w1(32'h3b33a289),
	.w2(32'h3a829850),
	.w3(32'h37b741e9),
	.w4(32'hba1150b5),
	.w5(32'hbb235cfd),
	.w6(32'h3856d0cd),
	.w7(32'h3aca02c7),
	.w8(32'hbace1745),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e0581),
	.w1(32'hba63cca9),
	.w2(32'hbaa1659e),
	.w3(32'hbab149df),
	.w4(32'h3a8320ce),
	.w5(32'hbabdd473),
	.w6(32'hba2725eb),
	.w7(32'h39aeea35),
	.w8(32'hbb369875),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e7e1),
	.w1(32'hbb02dae4),
	.w2(32'hba67e3c6),
	.w3(32'hbb03474d),
	.w4(32'hb90d71b9),
	.w5(32'hbafad05d),
	.w6(32'hbb2d845e),
	.w7(32'hbaaeb932),
	.w8(32'hbaeb5090),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc988d),
	.w1(32'hbbb4d64a),
	.w2(32'hb982aaea),
	.w3(32'hbb84cb0c),
	.w4(32'hba9c5452),
	.w5(32'hbaa3b115),
	.w6(32'hbbb68811),
	.w7(32'hba6fc23a),
	.w8(32'h3b472021),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f96f7),
	.w1(32'hbb00afff),
	.w2(32'h3bb4b0ba),
	.w3(32'hbc40a24f),
	.w4(32'h3a68694c),
	.w5(32'h3a3d6bd9),
	.w6(32'hbb867f12),
	.w7(32'h3b091abd),
	.w8(32'hb9d4fab0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae42c08),
	.w1(32'hbb68d7f8),
	.w2(32'h3a60989c),
	.w3(32'hbb40e821),
	.w4(32'hbb38dd73),
	.w5(32'hbb18e32b),
	.w6(32'hbbca5791),
	.w7(32'hbaa7c2e3),
	.w8(32'hbab752a0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f3c14),
	.w1(32'h3b0cf6d2),
	.w2(32'h3ae3c233),
	.w3(32'hbb14769f),
	.w4(32'h3b1c95ae),
	.w5(32'h381f0ada),
	.w6(32'hbaf45cc1),
	.w7(32'h38afb6d9),
	.w8(32'hbadaca27),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb800330),
	.w1(32'hbb8ee90a),
	.w2(32'hba84bb98),
	.w3(32'hbba52b5f),
	.w4(32'hbb3be9e7),
	.w5(32'h3a6de0e1),
	.w6(32'hbaab8388),
	.w7(32'hb9ae3bc2),
	.w8(32'h3b61534f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00f11c),
	.w1(32'h3ae5dd26),
	.w2(32'h3bf4af9a),
	.w3(32'h3b242000),
	.w4(32'h3b29b42c),
	.w5(32'hbae303e7),
	.w6(32'hba790e26),
	.w7(32'h3baa9989),
	.w8(32'hba8fbb65),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12e4eb),
	.w1(32'hbbbb6382),
	.w2(32'hbb7079c0),
	.w3(32'hbac35a7b),
	.w4(32'hbb571b81),
	.w5(32'hbb2bcc42),
	.w6(32'hbb38352b),
	.w7(32'hba9c6281),
	.w8(32'hb9f74f77),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb24a8),
	.w1(32'hbb7ae47a),
	.w2(32'h3b386e68),
	.w3(32'hbba6c9b5),
	.w4(32'h3b3160f1),
	.w5(32'hb92e35ec),
	.w6(32'hbb8bb751),
	.w7(32'hba1be229),
	.w8(32'h3a2e10ed),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee47e2),
	.w1(32'hbb4900c9),
	.w2(32'hbc122dbb),
	.w3(32'hbc457a93),
	.w4(32'hbbf0f237),
	.w5(32'h3b5d20b4),
	.w6(32'hbbdcbb45),
	.w7(32'hbbd22d44),
	.w8(32'h3ae32424),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c99bc),
	.w1(32'h3b20794a),
	.w2(32'h3960b131),
	.w3(32'h3b3c021b),
	.w4(32'hba999d97),
	.w5(32'hbb4cd91c),
	.w6(32'h3b513061),
	.w7(32'h39a63e77),
	.w8(32'hbb58f0fc),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb621a48),
	.w1(32'hbbb4730e),
	.w2(32'h3b05f615),
	.w3(32'hbbddb118),
	.w4(32'hba86318d),
	.w5(32'h3b10b9d8),
	.w6(32'hbbbafc5f),
	.w7(32'hb8f8809f),
	.w8(32'h3b110d02),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9138a7),
	.w1(32'h3b89c4cc),
	.w2(32'hba9a3c6c),
	.w3(32'h3b7f3c37),
	.w4(32'hb97ef370),
	.w5(32'hbb969c90),
	.w6(32'h3a87504a),
	.w7(32'hbaa13ac6),
	.w8(32'hbaf8326b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b9bea1),
	.w1(32'h3a001536),
	.w2(32'hbaee22f3),
	.w3(32'hbb2e8d97),
	.w4(32'h3a0fe438),
	.w5(32'h3b072ee0),
	.w6(32'h3b06a8cc),
	.w7(32'h3a815d00),
	.w8(32'h3b02cda1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3566b7),
	.w1(32'hbb60e48c),
	.w2(32'hbae97dde),
	.w3(32'hbbcdbc3e),
	.w4(32'h3adbed54),
	.w5(32'h3a9437d1),
	.w6(32'hbb2f85d3),
	.w7(32'hb9f6b4dd),
	.w8(32'hba1fd282),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab01ca8),
	.w1(32'h3a05e613),
	.w2(32'hbabe6a19),
	.w3(32'hbb081699),
	.w4(32'h3b143145),
	.w5(32'hb8d4a072),
	.w6(32'h3af0ec37),
	.w7(32'hbab65401),
	.w8(32'h38b95693),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73029a),
	.w1(32'hbb029990),
	.w2(32'hb982b9ad),
	.w3(32'hbb7ec137),
	.w4(32'hbbbbe3ac),
	.w5(32'hba56cef2),
	.w6(32'hbbb1397b),
	.w7(32'hbaa279a3),
	.w8(32'hbad5462c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49c11e),
	.w1(32'hbb52128c),
	.w2(32'h3a473694),
	.w3(32'h3b8755f7),
	.w4(32'h3b6d9b7f),
	.w5(32'hbaa333cd),
	.w6(32'h3a259711),
	.w7(32'h3bce1ac3),
	.w8(32'hb9fd566d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53088a),
	.w1(32'h3b2048f9),
	.w2(32'hb71f201b),
	.w3(32'hba52cb2c),
	.w4(32'h3b47dddd),
	.w5(32'h3ba65511),
	.w6(32'h3b190ba0),
	.w7(32'h3b85244b),
	.w8(32'h3acb722e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00c22d),
	.w1(32'hbacd891a),
	.w2(32'hba37b378),
	.w3(32'hba61d197),
	.w4(32'h3a4b9898),
	.w5(32'hbac713b7),
	.w6(32'hbb4814e0),
	.w7(32'hba796a3b),
	.w8(32'h3ab6a697),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fc7db),
	.w1(32'hbb4d110c),
	.w2(32'h3b560ab5),
	.w3(32'h38a8382a),
	.w4(32'h3ac25cd2),
	.w5(32'h3a5c2546),
	.w6(32'hbba1bfd0),
	.w7(32'h3a4daa11),
	.w8(32'h3962e210),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f41fd),
	.w1(32'hbc08a563),
	.w2(32'hbba0cb6d),
	.w3(32'hbbdbb6c9),
	.w4(32'hbb170ec9),
	.w5(32'hbab29802),
	.w6(32'hbbe8f7f1),
	.w7(32'hbaefe771),
	.w8(32'h3ad64b84),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6045bc),
	.w1(32'hbbba69b3),
	.w2(32'h39a6311f),
	.w3(32'hbb616c89),
	.w4(32'hbb245fac),
	.w5(32'hba6513a5),
	.w6(32'hbbddb996),
	.w7(32'h3a04f532),
	.w8(32'hb9994948),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954354e),
	.w1(32'hbadf566e),
	.w2(32'h3a759c90),
	.w3(32'h3a550a23),
	.w4(32'h3ab7b569),
	.w5(32'h3b31f0f5),
	.w6(32'h3acfed4c),
	.w7(32'h3b73b0fa),
	.w8(32'h3ac7ebe9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17f999),
	.w1(32'hba6570b8),
	.w2(32'hbb31d2f3),
	.w3(32'h396be282),
	.w4(32'hbb9743d1),
	.w5(32'hbb54cdc1),
	.w6(32'h3b670646),
	.w7(32'hbb5fca91),
	.w8(32'hbb8360a3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aefbc),
	.w1(32'hbb8c4966),
	.w2(32'h3aa0cc0e),
	.w3(32'h3b64f2d2),
	.w4(32'hba843a67),
	.w5(32'hbb34189b),
	.w6(32'hbbd6c7bb),
	.w7(32'hbb60cac6),
	.w8(32'h3a9c0eb3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3526e7),
	.w1(32'hbbb7a9da),
	.w2(32'hbb546ac0),
	.w3(32'hbbf56165),
	.w4(32'h3a05b140),
	.w5(32'hbbc4879e),
	.w6(32'hbb9e4085),
	.w7(32'h3b02c4c1),
	.w8(32'hbbcc3063),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cfabf),
	.w1(32'hbb43b8c8),
	.w2(32'h3b53f4c5),
	.w3(32'hb90443d7),
	.w4(32'h3a738f0f),
	.w5(32'hb8dd0664),
	.w6(32'hbb8fb4f5),
	.w7(32'hbb406783),
	.w8(32'h3a364a8b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc5edf),
	.w1(32'hba52b7c5),
	.w2(32'hbaffbeaf),
	.w3(32'hbb795ae1),
	.w4(32'hbb4277d1),
	.w5(32'hbb114526),
	.w6(32'hbbc2133f),
	.w7(32'hbb76a01a),
	.w8(32'hbae59781),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac681f3),
	.w1(32'h3acdf3b1),
	.w2(32'hbb762331),
	.w3(32'h3a9d473f),
	.w4(32'hbae4070a),
	.w5(32'hbb4b3928),
	.w6(32'h3b70a6c5),
	.w7(32'hbabfd47e),
	.w8(32'h399b6d2b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6429d8),
	.w1(32'h3b6fc62b),
	.w2(32'h3af94c5b),
	.w3(32'h3ad7b517),
	.w4(32'h3aa2019d),
	.w5(32'hb95735d8),
	.w6(32'hba4d33a8),
	.w7(32'h3b10973d),
	.w8(32'hbba406e0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule