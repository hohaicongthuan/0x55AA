module layer_10_featuremap_401(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cd132),
	.w1(32'h3c00b33d),
	.w2(32'h3a85beb7),
	.w3(32'h3bdae98e),
	.w4(32'h3c0bf066),
	.w5(32'h3a70aa0c),
	.w6(32'hbbf1b1a3),
	.w7(32'h3c555792),
	.w8(32'h3c978d11),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada4c48),
	.w1(32'hbc517815),
	.w2(32'hbb97e7e5),
	.w3(32'h3ae1a206),
	.w4(32'h3b46e870),
	.w5(32'h3b8bcb21),
	.w6(32'h3c51d191),
	.w7(32'h3b42120c),
	.w8(32'h3b9bf0cc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5df7d7),
	.w1(32'hbbe653c4),
	.w2(32'hbb7a987c),
	.w3(32'h3aaef1da),
	.w4(32'hbb136cbc),
	.w5(32'h3b95e525),
	.w6(32'hbb5030d3),
	.w7(32'hbb836ea3),
	.w8(32'hbaa9be98),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a54e8),
	.w1(32'hbbd457f6),
	.w2(32'hb9c41eee),
	.w3(32'h3b11424b),
	.w4(32'h39651227),
	.w5(32'h3a076a84),
	.w6(32'h3b0f8293),
	.w7(32'hbc278b4d),
	.w8(32'hbbd43146),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b574a4a),
	.w1(32'hba87f886),
	.w2(32'h3b1140e0),
	.w3(32'h3bc172ae),
	.w4(32'h3ba6a72b),
	.w5(32'hbb6306f5),
	.w6(32'h3b80e6e1),
	.w7(32'h3b270aa5),
	.w8(32'h3b38ead2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba593f0a),
	.w1(32'hbb802aed),
	.w2(32'hbbe99648),
	.w3(32'h3b88b5c1),
	.w4(32'hbbe394b2),
	.w5(32'hbb66daaa),
	.w6(32'hba3bd6b9),
	.w7(32'h3b5bb5da),
	.w8(32'hbc225049),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae08676),
	.w1(32'hbb723612),
	.w2(32'hba871f8b),
	.w3(32'h3b924347),
	.w4(32'hbb7f9a77),
	.w5(32'h3c615d42),
	.w6(32'hbc12b584),
	.w7(32'h3b7e2d04),
	.w8(32'h3b8603a4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07559b),
	.w1(32'h3ba78406),
	.w2(32'h3b798b0d),
	.w3(32'hbb2673ff),
	.w4(32'h3ac018f4),
	.w5(32'hbc36656b),
	.w6(32'h3b0a6c39),
	.w7(32'hbc0b2b73),
	.w8(32'hbbe2e5dc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b95e5),
	.w1(32'hbc1f878b),
	.w2(32'hbbd76f9e),
	.w3(32'h3ab4ed1f),
	.w4(32'hbba84b0d),
	.w5(32'hbc286a1c),
	.w6(32'hbc00eebc),
	.w7(32'hbae33733),
	.w8(32'hba0ac765),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8adf05),
	.w1(32'h399519ac),
	.w2(32'h3b451420),
	.w3(32'h3b1b9922),
	.w4(32'hb905c92e),
	.w5(32'h3bd486a9),
	.w6(32'h3be2625e),
	.w7(32'hbb0309d6),
	.w8(32'h39d10f1c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26f804),
	.w1(32'h3ac4dbde),
	.w2(32'h3ae907c6),
	.w3(32'h3a5c8fb4),
	.w4(32'h3c198f9e),
	.w5(32'h3cd26475),
	.w6(32'hba825d7a),
	.w7(32'hbb75def4),
	.w8(32'hbaec35bc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923700a),
	.w1(32'hbc7719e9),
	.w2(32'hbb285ae9),
	.w3(32'h3c8e65c9),
	.w4(32'hbc38ee42),
	.w5(32'h3aabdd38),
	.w6(32'h3be0e6bc),
	.w7(32'hbc20fe04),
	.w8(32'h3ab7bd60),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb655c0a),
	.w1(32'hbc08cc4e),
	.w2(32'h3b849643),
	.w3(32'h3b64337f),
	.w4(32'hbaf5b766),
	.w5(32'h3c0b2691),
	.w6(32'h3b41dd86),
	.w7(32'hbb8e6f43),
	.w8(32'h3ba648b4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40e5b6),
	.w1(32'hb9d7caaa),
	.w2(32'h3b826b20),
	.w3(32'h3aa48516),
	.w4(32'h3b5a3729),
	.w5(32'h3c2ec14d),
	.w6(32'h3c1c4878),
	.w7(32'h3b32b451),
	.w8(32'h3b35974c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b498024),
	.w1(32'hb9f329c5),
	.w2(32'h3aa4b126),
	.w3(32'h3b830416),
	.w4(32'hbbc2f981),
	.w5(32'h3ba93c7b),
	.w6(32'hba1e3266),
	.w7(32'h3b13ec81),
	.w8(32'h3b919c8a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb487450),
	.w1(32'h37427ec4),
	.w2(32'h3c5158b8),
	.w3(32'hbbf7c537),
	.w4(32'hbbfa3f43),
	.w5(32'h3b480099),
	.w6(32'h3b797325),
	.w7(32'h3b20d978),
	.w8(32'h3be298d8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7eaf43),
	.w1(32'hbc93b8db),
	.w2(32'hbc83956d),
	.w3(32'hbab5d4ea),
	.w4(32'hbc3b2525),
	.w5(32'hbbe6e066),
	.w6(32'hba69ac9e),
	.w7(32'hbb69d140),
	.w8(32'hbb4d9a9b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96560b),
	.w1(32'hba19aaee),
	.w2(32'h3a75f3cd),
	.w3(32'hbc3e3435),
	.w4(32'hbb35ed3e),
	.w5(32'h3bebb8b3),
	.w6(32'hbb724f67),
	.w7(32'hb90a948a),
	.w8(32'h3a9c791f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a2925),
	.w1(32'hbbc3f512),
	.w2(32'hb9af24cc),
	.w3(32'hbbef0a8d),
	.w4(32'hb981b518),
	.w5(32'h3c0d58f1),
	.w6(32'hbc14b794),
	.w7(32'h3b8e5aa2),
	.w8(32'h3c1e46d2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0decd3),
	.w1(32'h3a3f286e),
	.w2(32'hbbfd68b0),
	.w3(32'h3c5db849),
	.w4(32'hbbd56011),
	.w5(32'h3ad60300),
	.w6(32'h3c0b1359),
	.w7(32'hbb30e2c0),
	.w8(32'hbba08da1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba87c21),
	.w1(32'hbb9d42d1),
	.w2(32'hbbf8615f),
	.w3(32'hbbedd8ba),
	.w4(32'hbb823171),
	.w5(32'hbc4184a0),
	.w6(32'h3ac34058),
	.w7(32'hbc3ff2c8),
	.w8(32'hbc5809f3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e8bd1),
	.w1(32'h3aa2fab7),
	.w2(32'hb8793718),
	.w3(32'hbc15ff83),
	.w4(32'hbc0b5c4c),
	.w5(32'h3aa18dd8),
	.w6(32'hbc5168fa),
	.w7(32'hbc3da396),
	.w8(32'hbbead0d6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03ba59),
	.w1(32'hbc2d0664),
	.w2(32'h3bbc305b),
	.w3(32'hbc61a150),
	.w4(32'hbca347fc),
	.w5(32'hbac817ae),
	.w6(32'hbc0824e0),
	.w7(32'hbc83e75b),
	.w8(32'hbc227ba3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14173e),
	.w1(32'hbb8323f4),
	.w2(32'hbbfbd481),
	.w3(32'hbc05857f),
	.w4(32'h3b469e95),
	.w5(32'hbb3db935),
	.w6(32'h3a37afdd),
	.w7(32'h3b74ccd9),
	.w8(32'h3bcf70fc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b050add),
	.w1(32'h399ab932),
	.w2(32'hbb29ddd2),
	.w3(32'h3bff4cc4),
	.w4(32'hbb0634b8),
	.w5(32'hbbfaa0ce),
	.w6(32'h3cc55ef9),
	.w7(32'hbaf5edf3),
	.w8(32'hbc57f7ac),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b321bd5),
	.w1(32'h3afe0b84),
	.w2(32'h3a8c8120),
	.w3(32'hbbb2b442),
	.w4(32'hbbc5eb97),
	.w5(32'hbc834544),
	.w6(32'hbb58c5e0),
	.w7(32'hbc4bad3a),
	.w8(32'hbc0dddd7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c024824),
	.w1(32'hbb132b7c),
	.w2(32'h3b5e5035),
	.w3(32'hbaccf6ce),
	.w4(32'h3bdaf273),
	.w5(32'h3c477041),
	.w6(32'hbbc61ad3),
	.w7(32'h3c0c2ba6),
	.w8(32'h3c0645c6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c624fda),
	.w1(32'hbc1de0f5),
	.w2(32'hbbf414c3),
	.w3(32'h3c825572),
	.w4(32'hbbc91d9a),
	.w5(32'hbc02585f),
	.w6(32'h3c74190b),
	.w7(32'h39b9e228),
	.w8(32'hbc31d6c5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2cbee2),
	.w1(32'hbc581baf),
	.w2(32'hbcc6a698),
	.w3(32'hbb2e174a),
	.w4(32'hbc392549),
	.w5(32'hbbab4be0),
	.w6(32'hbbf525e6),
	.w7(32'hbb1bb678),
	.w8(32'hbbceb4ed),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8205),
	.w1(32'hbaf01682),
	.w2(32'hbb8633cd),
	.w3(32'h3bbc9c05),
	.w4(32'h3b82ff0d),
	.w5(32'hba6f211c),
	.w6(32'h3c1df34a),
	.w7(32'h3c010ea6),
	.w8(32'h39ef3ba3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f446d7),
	.w1(32'hbc39d2b9),
	.w2(32'hbc8a3ceb),
	.w3(32'hbaca35fa),
	.w4(32'hbc2615b4),
	.w5(32'hbba4b379),
	.w6(32'hbb5f28b5),
	.w7(32'h3c2110fd),
	.w8(32'h3b91f6ac),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a573b),
	.w1(32'h3b2d7398),
	.w2(32'h3b34cf2f),
	.w3(32'hbbc16b41),
	.w4(32'h3a309678),
	.w5(32'h3a7f3aee),
	.w6(32'h3bc70208),
	.w7(32'hbac41a0e),
	.w8(32'hbb046a60),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99f410),
	.w1(32'hbc004085),
	.w2(32'h3b29ac08),
	.w3(32'h3b031d92),
	.w4(32'hbb124f99),
	.w5(32'h3c2adf26),
	.w6(32'hbb72e0d9),
	.w7(32'hbc1931e6),
	.w8(32'h3bedafd6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64e770),
	.w1(32'hba6f034b),
	.w2(32'hbbd27875),
	.w3(32'h3bc949c4),
	.w4(32'hbb47407a),
	.w5(32'h3954b1c6),
	.w6(32'h3b2a7dea),
	.w7(32'hbbabff42),
	.w8(32'hbbe10279),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac77487),
	.w1(32'hbb783e60),
	.w2(32'hbc4c0125),
	.w3(32'h3bf49df6),
	.w4(32'hbbcffd12),
	.w5(32'hbc82ad66),
	.w6(32'hb7aadae4),
	.w7(32'hbbfdcade),
	.w8(32'hbc479c18),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40948f),
	.w1(32'h3b190e59),
	.w2(32'h3b918798),
	.w3(32'hbb982cc8),
	.w4(32'hbac3453d),
	.w5(32'hb81c993c),
	.w6(32'hbc8cb880),
	.w7(32'hbbe281bc),
	.w8(32'hb94471f6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8280a7),
	.w1(32'hbcc190dc),
	.w2(32'hbbc38866),
	.w3(32'h3c892c2a),
	.w4(32'hbcee04a3),
	.w5(32'h3cbf0be5),
	.w6(32'h3cb2e765),
	.w7(32'hbc8260f0),
	.w8(32'h3c1d155d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27995f),
	.w1(32'hbc34832b),
	.w2(32'hbc89420f),
	.w3(32'h3c13e572),
	.w4(32'hbc211efd),
	.w5(32'hbbde18fe),
	.w6(32'h3c826286),
	.w7(32'hbc3145ef),
	.w8(32'hbc685f0a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bfbd4),
	.w1(32'h3b4d2bac),
	.w2(32'hbc813197),
	.w3(32'h3c4efcdb),
	.w4(32'hbc28524c),
	.w5(32'hbc6df251),
	.w6(32'h3bf6e2dd),
	.w7(32'hbbfc695d),
	.w8(32'hbc6e0f5f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a5c9c),
	.w1(32'h3b7886d4),
	.w2(32'h3c17d9db),
	.w3(32'h3b274dfc),
	.w4(32'h3ba23b03),
	.w5(32'h3b79c010),
	.w6(32'h3c045a3e),
	.w7(32'hbae4b9b8),
	.w8(32'hb9b0a690),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd14f14),
	.w1(32'hbc2de69e),
	.w2(32'h3b0941f9),
	.w3(32'h3c2ad77d),
	.w4(32'h388129da),
	.w5(32'h3c257d03),
	.w6(32'hbb13110a),
	.w7(32'h3a91d61b),
	.w8(32'h3bc780aa),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad2d79),
	.w1(32'hbbad392b),
	.w2(32'hbb89633a),
	.w3(32'hba20fe1a),
	.w4(32'h3b6a9078),
	.w5(32'h3bd4ef1c),
	.w6(32'hbbae999d),
	.w7(32'h3b71ff2b),
	.w8(32'h3aa4069d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6a710),
	.w1(32'hbc02d425),
	.w2(32'hbb98974c),
	.w3(32'h37c4b709),
	.w4(32'hbaac0706),
	.w5(32'h3a792fec),
	.w6(32'hbb917339),
	.w7(32'hbc16a1b4),
	.w8(32'hbb5af9e1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9e932),
	.w1(32'h3ba5c324),
	.w2(32'h3bef7101),
	.w3(32'hb9e20c39),
	.w4(32'hbb8f3f2e),
	.w5(32'hbaa3c2b9),
	.w6(32'hbb8918c5),
	.w7(32'hbba694c3),
	.w8(32'hb9f37b0b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a65ec),
	.w1(32'hbb3b6232),
	.w2(32'hbb912f39),
	.w3(32'h39206bb5),
	.w4(32'h3a97696c),
	.w5(32'h3a86f954),
	.w6(32'hbadaecd1),
	.w7(32'hbb6e1b9c),
	.w8(32'hbb050377),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11c756),
	.w1(32'hbb8b613e),
	.w2(32'h3bd6c647),
	.w3(32'h3b818af0),
	.w4(32'hbc0f852f),
	.w5(32'hbc03ac69),
	.w6(32'hbb693475),
	.w7(32'hbb9ac074),
	.w8(32'hbb64ad14),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcf444),
	.w1(32'h3c9fe09c),
	.w2(32'h3ca75eef),
	.w3(32'hbbda6e09),
	.w4(32'h39d347af),
	.w5(32'hbb846278),
	.w6(32'hbae5a94b),
	.w7(32'hbc275181),
	.w8(32'hbc233eaa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8e5b5),
	.w1(32'h3b20b80d),
	.w2(32'h3be56635),
	.w3(32'h3a81f864),
	.w4(32'hbc0e1a15),
	.w5(32'h3c13c7c6),
	.w6(32'hbc41bb88),
	.w7(32'h3861498c),
	.w8(32'h3bb39b63),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96610a),
	.w1(32'h3c410445),
	.w2(32'h3bc05ff9),
	.w3(32'h3b016814),
	.w4(32'h3a8193df),
	.w5(32'hbc9d7e52),
	.w6(32'hb9cee8bc),
	.w7(32'hbb0f8c96),
	.w8(32'hbba4ca82),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21c3de),
	.w1(32'h3c265295),
	.w2(32'h3b916590),
	.w3(32'hbb6ad585),
	.w4(32'hbb48372b),
	.w5(32'hbc7168f6),
	.w6(32'hbb939f8e),
	.w7(32'h3b6fcf77),
	.w8(32'h3b357f16),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9f06f),
	.w1(32'hbbe1bfff),
	.w2(32'hbc095622),
	.w3(32'hba97a30c),
	.w4(32'h3b6d0367),
	.w5(32'hbbd144be),
	.w6(32'hbb681ea7),
	.w7(32'h3b7ab84a),
	.w8(32'h3b2be97f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a095ef4),
	.w1(32'hba19c305),
	.w2(32'hbb1aaa19),
	.w3(32'h3b12661e),
	.w4(32'h3a3fa5d4),
	.w5(32'h3c092a09),
	.w6(32'h3a42f6ab),
	.w7(32'hbbd96204),
	.w8(32'hbbb33c89),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b564ff3),
	.w1(32'hbb03ca81),
	.w2(32'hbbad7805),
	.w3(32'h3a277fa7),
	.w4(32'hbb96e91d),
	.w5(32'hbb8147c6),
	.w6(32'h3c129e6b),
	.w7(32'hbb5ea5e4),
	.w8(32'hbad0bfb9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29f5c8),
	.w1(32'hbb911734),
	.w2(32'hbace3c90),
	.w3(32'h3a82966c),
	.w4(32'h3c0a4cfd),
	.w5(32'h3ad87eef),
	.w6(32'hbc02fe29),
	.w7(32'h39d49233),
	.w8(32'h3a5bd412),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17843e),
	.w1(32'hbbfe47a4),
	.w2(32'hbbe63ba4),
	.w3(32'h3b0ffac2),
	.w4(32'hbb979ef1),
	.w5(32'hbb2c7fe4),
	.w6(32'hbbe7f2ed),
	.w7(32'hbc48b3fb),
	.w8(32'hbbdecde7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4abd56),
	.w1(32'hb8cf9040),
	.w2(32'hbb3bb9a8),
	.w3(32'h3baf65b8),
	.w4(32'h3b5288ba),
	.w5(32'h3aa6536a),
	.w6(32'h3b81b1a9),
	.w7(32'h39d830bc),
	.w8(32'h385bd911),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac47885),
	.w1(32'h3ac282d3),
	.w2(32'h3b83b44b),
	.w3(32'hba25c5f7),
	.w4(32'h3b6f0d6b),
	.w5(32'hba12d829),
	.w6(32'hbb977048),
	.w7(32'h3c1147d5),
	.w8(32'hba70b11e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a8823),
	.w1(32'hbb3a6eaf),
	.w2(32'h3ba9dafd),
	.w3(32'h3ba9acb3),
	.w4(32'hbbd0b6e2),
	.w5(32'hbc768f1e),
	.w6(32'hba502759),
	.w7(32'hbc81d14d),
	.w8(32'hbc987f06),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebd0ad),
	.w1(32'hbc4af348),
	.w2(32'hbc85f9bf),
	.w3(32'hbc107095),
	.w4(32'hbc564a22),
	.w5(32'hbc1ef48e),
	.w6(32'hbbfcfecc),
	.w7(32'hbc23f6e1),
	.w8(32'hbb517758),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc12d97),
	.w1(32'h3bf666d0),
	.w2(32'h3c90e832),
	.w3(32'hbc088435),
	.w4(32'h393d328b),
	.w5(32'h3bc3aa69),
	.w6(32'h3883736f),
	.w7(32'hbba8334e),
	.w8(32'hbbd1db43),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5eb2),
	.w1(32'h3a911dbf),
	.w2(32'h3c962c6d),
	.w3(32'h3be81a46),
	.w4(32'hbb87aae4),
	.w5(32'hbc6f9835),
	.w6(32'h3b35682e),
	.w7(32'hbc392b3d),
	.w8(32'hbbf26f13),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc82439),
	.w1(32'hbb44b48b),
	.w2(32'h3aa82db5),
	.w3(32'hbb4ff6ec),
	.w4(32'hbbc57054),
	.w5(32'h393ed95b),
	.w6(32'hbbe2ea71),
	.w7(32'hbb09e918),
	.w8(32'h3b201e8d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ab261),
	.w1(32'hbb13f379),
	.w2(32'hb9b8e650),
	.w3(32'h3c1851ee),
	.w4(32'h3bbeb821),
	.w5(32'h3ba5dac6),
	.w6(32'h3c0e1782),
	.w7(32'hbc4372b3),
	.w8(32'hbbeffe62),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd14539),
	.w1(32'hbab9b829),
	.w2(32'hbb82bfe6),
	.w3(32'hbaae2ac9),
	.w4(32'h3bfc48be),
	.w5(32'hbbc3c0ef),
	.w6(32'hbb197cd2),
	.w7(32'h3b8a0dab),
	.w8(32'h3c2be701),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb449e3b),
	.w1(32'h3cba2cbc),
	.w2(32'h3c5abff2),
	.w3(32'h3bbf6d5a),
	.w4(32'h3c67bff7),
	.w5(32'hbb1de352),
	.w6(32'h3c38c3d8),
	.w7(32'h3b8b0563),
	.w8(32'hb9cbc37c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a66d7),
	.w1(32'hbbca2619),
	.w2(32'hbc4a7986),
	.w3(32'h3b74ac48),
	.w4(32'hbb4cdba4),
	.w5(32'hbb8e610e),
	.w6(32'h39dd5f5c),
	.w7(32'hbc19cb4c),
	.w8(32'hbc082a2f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2133f8),
	.w1(32'hbaa6d5a2),
	.w2(32'h3bdc8557),
	.w3(32'hbc75ae7e),
	.w4(32'hbc204796),
	.w5(32'hbaf1f5a9),
	.w6(32'hbc236e36),
	.w7(32'h3b856d98),
	.w8(32'h3c96fb21),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86c964),
	.w1(32'h3ba79dc3),
	.w2(32'h3b573c83),
	.w3(32'hbc25314a),
	.w4(32'hba16774d),
	.w5(32'hbbfbd3b7),
	.w6(32'hbbeadc3a),
	.w7(32'hb9003f6d),
	.w8(32'h3b1df443),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e7b2),
	.w1(32'hbbaa48b3),
	.w2(32'hbbca5041),
	.w3(32'hbbeec25e),
	.w4(32'hbbb1e487),
	.w5(32'h3b21533b),
	.w6(32'hbc4c3890),
	.w7(32'hbbdc3c76),
	.w8(32'h3c132af7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cf38d),
	.w1(32'hbbbd8477),
	.w2(32'hbbfe120d),
	.w3(32'hbacf3cb6),
	.w4(32'hba2e9863),
	.w5(32'hbb1ff7a7),
	.w6(32'h3b3390a9),
	.w7(32'hba031755),
	.w8(32'h38a4f7c4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dd1aa),
	.w1(32'hbb8243c5),
	.w2(32'hbb66d7be),
	.w3(32'hbbec7031),
	.w4(32'h3936b36d),
	.w5(32'hbaf424a0),
	.w6(32'h3baea730),
	.w7(32'hbb3121cb),
	.w8(32'hbb4698c7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c68dd),
	.w1(32'h3c4bba0f),
	.w2(32'hbb4230ca),
	.w3(32'hbb1fb3a0),
	.w4(32'h3c09327e),
	.w5(32'h3bc35a27),
	.w6(32'hbb67c3b5),
	.w7(32'h3bf65e0c),
	.w8(32'h3b366a99),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68aa48),
	.w1(32'h3cb84962),
	.w2(32'h3cff9438),
	.w3(32'h3be5a06a),
	.w4(32'h3c5ccc49),
	.w5(32'h3cdf6097),
	.w6(32'hbbc22c5e),
	.w7(32'h3c6b1afc),
	.w8(32'h3c4fb8f5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac285e),
	.w1(32'hbaa20d6c),
	.w2(32'h3bd679db),
	.w3(32'h3c887e1f),
	.w4(32'h3986dedf),
	.w5(32'hbb9a6e2f),
	.w6(32'h3c0c5fbe),
	.w7(32'h3b74b808),
	.w8(32'hb8fe4dc9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e59a5d),
	.w1(32'hbb87e07f),
	.w2(32'hbb7425b1),
	.w3(32'hb99f6496),
	.w4(32'h3b564027),
	.w5(32'h3cd018e1),
	.w6(32'h3a4ec770),
	.w7(32'h3c2bcdcf),
	.w8(32'h3c5ad3b6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043d21),
	.w1(32'h3acb9c7a),
	.w2(32'h3be7986f),
	.w3(32'h3b9dd8ea),
	.w4(32'h3b20d13b),
	.w5(32'h3c02300f),
	.w6(32'h3b2fbf11),
	.w7(32'h3b6f43f4),
	.w8(32'h3c10dffd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a428441),
	.w1(32'h3be06054),
	.w2(32'h3c8a6c79),
	.w3(32'hb9c3cd40),
	.w4(32'h3b639688),
	.w5(32'h3ba9a5d7),
	.w6(32'hbb6aa2ac),
	.w7(32'hbc22188a),
	.w8(32'h3a200547),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59d0ec),
	.w1(32'hbb82ca62),
	.w2(32'hbafb2a90),
	.w3(32'h3c314343),
	.w4(32'h3be40bd1),
	.w5(32'h3bae1f1a),
	.w6(32'h3b91430d),
	.w7(32'h3c3e14fb),
	.w8(32'h3c5e62d5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3a0cb),
	.w1(32'hbb4a2be7),
	.w2(32'h3bc8e7e8),
	.w3(32'hbb35691d),
	.w4(32'hbad22bbb),
	.w5(32'h3b83ca3d),
	.w6(32'hbb5d4642),
	.w7(32'hbb1f8799),
	.w8(32'hb9cf8375),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e2287),
	.w1(32'h3b9542d2),
	.w2(32'h3b90e95c),
	.w3(32'h3c18abf7),
	.w4(32'h3b81a7f2),
	.w5(32'h3c0ce62e),
	.w6(32'h3b0b5571),
	.w7(32'h39a5bfff),
	.w8(32'h3c719d8d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad96e62),
	.w1(32'hba3f8591),
	.w2(32'h3c24a39d),
	.w3(32'hba80ecdf),
	.w4(32'h3a3504a9),
	.w5(32'hbb92fc70),
	.w6(32'h3b1a83ce),
	.w7(32'h3bbf925b),
	.w8(32'h3b4c53e4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06dfe2),
	.w1(32'h395675d1),
	.w2(32'h3b8af4c5),
	.w3(32'h3bf30cb1),
	.w4(32'hbb0ea242),
	.w5(32'hba37e3be),
	.w6(32'h3c0e288e),
	.w7(32'hb95c0bdd),
	.w8(32'h3b69a940),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b318dca),
	.w1(32'hbad8b86f),
	.w2(32'hbaad2683),
	.w3(32'h3b5a2a86),
	.w4(32'hbaf469c9),
	.w5(32'hbaa6e01e),
	.w6(32'h3b657920),
	.w7(32'hbb86d034),
	.w8(32'hb903f401),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9573d),
	.w1(32'h3b365a20),
	.w2(32'hb9adecfd),
	.w3(32'hbacfbbef),
	.w4(32'hbb268e4b),
	.w5(32'hbb13a552),
	.w6(32'hbb1c4d2e),
	.w7(32'hbc02786f),
	.w8(32'hbbcda5b2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa33f4d),
	.w1(32'h3bd8b1ca),
	.w2(32'h3c1dde88),
	.w3(32'hbafee537),
	.w4(32'hb99aee21),
	.w5(32'h3b474c71),
	.w6(32'hbb9e10f4),
	.w7(32'h3a126de9),
	.w8(32'hbb5706e9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b405d4f),
	.w1(32'hbb22e691),
	.w2(32'hbc445c01),
	.w3(32'h3ab28dc2),
	.w4(32'hbba4f9aa),
	.w5(32'hbbc9aaae),
	.w6(32'h3b1ae106),
	.w7(32'hbbe9acb3),
	.w8(32'hbb0e94ce),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384c13b9),
	.w1(32'hbb658eae),
	.w2(32'hbbcd018d),
	.w3(32'hbb5070ef),
	.w4(32'hbc075074),
	.w5(32'hbad1f568),
	.w6(32'hbb53ee66),
	.w7(32'hbc1c9782),
	.w8(32'hbbcb46c9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2f01f),
	.w1(32'hbb040c4f),
	.w2(32'h3ad7b26d),
	.w3(32'h3b7b0ffc),
	.w4(32'hbc165e32),
	.w5(32'hbb80c113),
	.w6(32'h396b09ab),
	.w7(32'hbc0a0348),
	.w8(32'hbbad6dca),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4399),
	.w1(32'hbaf4e7af),
	.w2(32'hbb54375c),
	.w3(32'h3b9d7477),
	.w4(32'h3bc08695),
	.w5(32'h3af2b8ec),
	.w6(32'hbb69f121),
	.w7(32'hbc23e09b),
	.w8(32'hbbbc40db),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe06ae),
	.w1(32'hbba5ac1b),
	.w2(32'h3b918902),
	.w3(32'hbbec6bc8),
	.w4(32'h3b29e6b0),
	.w5(32'hbb36c4c7),
	.w6(32'hbc76be16),
	.w7(32'h3b2a7270),
	.w8(32'hbb269c53),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf28e6),
	.w1(32'hbc0cf17d),
	.w2(32'hbb8c6d47),
	.w3(32'h3a80c945),
	.w4(32'hbc2b72d6),
	.w5(32'hbc365fe8),
	.w6(32'hb9fc8894),
	.w7(32'hbc424541),
	.w8(32'hbc42885a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd0aa5),
	.w1(32'hbb8592ff),
	.w2(32'h3c31dfa9),
	.w3(32'hbb8ff334),
	.w4(32'hbb6a62ed),
	.w5(32'h3c6daaa4),
	.w6(32'hbc05a68e),
	.w7(32'h3bd824ea),
	.w8(32'h3c9db12a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f06a6),
	.w1(32'hbaa4e27a),
	.w2(32'hbadbb701),
	.w3(32'h3a866899),
	.w4(32'hbb97a861),
	.w5(32'hbc55d70a),
	.w6(32'h3c05901a),
	.w7(32'hbc2209af),
	.w8(32'hbbd5d7e2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0c8c2),
	.w1(32'hbaa26668),
	.w2(32'h3bd1012e),
	.w3(32'hbb7b1be3),
	.w4(32'hba83cbe8),
	.w5(32'hbc2967f2),
	.w6(32'hbbb8b7e3),
	.w7(32'h3a0b459d),
	.w8(32'h3b43a4ed),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2558c9),
	.w1(32'h3bb6a70e),
	.w2(32'h3bd9700a),
	.w3(32'hbb89374e),
	.w4(32'h3ba7612a),
	.w5(32'h3c1e27a5),
	.w6(32'hba2dbc92),
	.w7(32'h3c3dac10),
	.w8(32'h3c89b72c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba75d66),
	.w1(32'hbb4744e4),
	.w2(32'hbc45bbf3),
	.w3(32'h3ba73699),
	.w4(32'hbab173eb),
	.w5(32'hbbdec786),
	.w6(32'h3c849c77),
	.w7(32'h3ba9427a),
	.w8(32'hbad19237),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6b1e4),
	.w1(32'hbb19c36d),
	.w2(32'hbb8187f2),
	.w3(32'hbc15722f),
	.w4(32'hbbac7683),
	.w5(32'hbbf68c3d),
	.w6(32'h3abcdc69),
	.w7(32'hbb7717ed),
	.w8(32'hbb82f79d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa4da1),
	.w1(32'h3c0ffe1b),
	.w2(32'h3c5dc5f4),
	.w3(32'hbbb65e3c),
	.w4(32'h3b0fe5d4),
	.w5(32'h3b972e11),
	.w6(32'hbb81e716),
	.w7(32'hbc50c59d),
	.w8(32'hbbdede17),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38e917),
	.w1(32'h3bd45a6a),
	.w2(32'h3d026957),
	.w3(32'hba3a00fd),
	.w4(32'h3b0971a6),
	.w5(32'h3bbc5f89),
	.w6(32'hbc109017),
	.w7(32'hbb0a805e),
	.w8(32'h3a5f21fa),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4f483),
	.w1(32'hbc78caae),
	.w2(32'hbaf290e2),
	.w3(32'h3cf21e64),
	.w4(32'hbac9c24e),
	.w5(32'h3c16de17),
	.w6(32'h3c32f673),
	.w7(32'hbb51a89d),
	.w8(32'h3c2b8ce6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b344553),
	.w1(32'hbc23d531),
	.w2(32'hbc310daf),
	.w3(32'h3ba6cc47),
	.w4(32'hbbf8affb),
	.w5(32'hbc2085a8),
	.w6(32'h3c2bcdc4),
	.w7(32'hbbdc586b),
	.w8(32'hbc069bbc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d469d),
	.w1(32'hbb911ed2),
	.w2(32'hbb96b668),
	.w3(32'h3b250d6b),
	.w4(32'hbbd42d56),
	.w5(32'hbb91148e),
	.w6(32'h3bb2f595),
	.w7(32'hbb82d93a),
	.w8(32'hbbd8e845),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b978f),
	.w1(32'hbaddfdff),
	.w2(32'h3bfb7331),
	.w3(32'hbb422619),
	.w4(32'hbbf4d94f),
	.w5(32'h3bfd12b1),
	.w6(32'hbbe5a4f3),
	.w7(32'hbb82bbdb),
	.w8(32'h3bb82118),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7b76d),
	.w1(32'hbb51db78),
	.w2(32'h3ab02507),
	.w3(32'hbb3df68e),
	.w4(32'hba8ee8d7),
	.w5(32'hbaf56b63),
	.w6(32'hbb0d3336),
	.w7(32'h3a9b7c78),
	.w8(32'hba5f9a82),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90aa54),
	.w1(32'hba220bad),
	.w2(32'hbadc88f4),
	.w3(32'h3c1bdc68),
	.w4(32'hbb642bf3),
	.w5(32'hb98c7840),
	.w6(32'h3c3a737f),
	.w7(32'h3b1685d3),
	.w8(32'h3a7b4775),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a583da3),
	.w1(32'h3a9305a5),
	.w2(32'h3bcb8eb9),
	.w3(32'h3bb16211),
	.w4(32'hbbc77f2f),
	.w5(32'hbb9348ee),
	.w6(32'hbafcbb13),
	.w7(32'hbbda537e),
	.w8(32'h3a63d521),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b562f60),
	.w1(32'hba5aafd9),
	.w2(32'hba43395e),
	.w3(32'h3b985ca8),
	.w4(32'h3a90467a),
	.w5(32'hb993431d),
	.w6(32'h3aa06647),
	.w7(32'h3b42cf13),
	.w8(32'h3b335fa8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfcfc9),
	.w1(32'h3bad8109),
	.w2(32'h3ca25db7),
	.w3(32'hbb2f5052),
	.w4(32'hbb85f70a),
	.w5(32'h3b9e7107),
	.w6(32'hba3965e7),
	.w7(32'hba73cfe5),
	.w8(32'hb99c966b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd23a83),
	.w1(32'hba785c54),
	.w2(32'h3b88fbac),
	.w3(32'h3c645405),
	.w4(32'hbac5a58d),
	.w5(32'h3ae2879e),
	.w6(32'h3bceca82),
	.w7(32'hba6efdc4),
	.w8(32'h3bc9fad6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06655b),
	.w1(32'hbadf6455),
	.w2(32'hbb650f23),
	.w3(32'hba65090c),
	.w4(32'hba2a3c01),
	.w5(32'hb99242d8),
	.w6(32'h3b202b87),
	.w7(32'h3afca59b),
	.w8(32'h3b7948b5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b892253),
	.w1(32'h3b43b10f),
	.w2(32'h3bf1568d),
	.w3(32'h3bc00f5f),
	.w4(32'h3bd239e3),
	.w5(32'h3b8beb53),
	.w6(32'h3bfd5093),
	.w7(32'h3b27d786),
	.w8(32'hbb8e9911),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28fcf6),
	.w1(32'h3a3b0092),
	.w2(32'hbaf6a707),
	.w3(32'h3c1c121b),
	.w4(32'h3be8e83c),
	.w5(32'h3b34679e),
	.w6(32'h3b144914),
	.w7(32'h3b883378),
	.w8(32'hbb7fe7c9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6bef3),
	.w1(32'h39d5fab2),
	.w2(32'h3bc99727),
	.w3(32'hbb4b53f1),
	.w4(32'hbab7b3af),
	.w5(32'h3a788727),
	.w6(32'hbbe108de),
	.w7(32'hbbd5c08f),
	.w8(32'h3a365e7e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40615f),
	.w1(32'h3a93bf43),
	.w2(32'h3c1f0e43),
	.w3(32'hbb4d408c),
	.w4(32'hba4d7376),
	.w5(32'h3a4aba48),
	.w6(32'h3a385ec4),
	.w7(32'h3bfbfd08),
	.w8(32'h3be39503),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0caeb3),
	.w1(32'hbb1484b6),
	.w2(32'h3b9a7ba5),
	.w3(32'h3b48ae61),
	.w4(32'hbbc0303b),
	.w5(32'hba47e0a1),
	.w6(32'h3b26ebea),
	.w7(32'hbc0871df),
	.w8(32'hbaa15f79),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e885d),
	.w1(32'h3c194ac5),
	.w2(32'h3c300186),
	.w3(32'h3adf87f5),
	.w4(32'hba17179d),
	.w5(32'h3ab15000),
	.w6(32'hbace4c11),
	.w7(32'h3b360790),
	.w8(32'h3bb82940),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb77462),
	.w1(32'h3b87174d),
	.w2(32'h3bd6b1e3),
	.w3(32'h3bebb539),
	.w4(32'hbac130dd),
	.w5(32'h3c21d2f9),
	.w6(32'h3bd3f797),
	.w7(32'hba9a69b4),
	.w8(32'h3ad4ab1e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa9ec8),
	.w1(32'hb9086ed3),
	.w2(32'hbb347c0e),
	.w3(32'h3bb9d269),
	.w4(32'hbb239552),
	.w5(32'hbc81ca7d),
	.w6(32'hbaa0a079),
	.w7(32'h38c57c05),
	.w8(32'hbb85d91f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2f909),
	.w1(32'hba537b09),
	.w2(32'hbb5e1d75),
	.w3(32'hb9a615b0),
	.w4(32'hba468123),
	.w5(32'hbb9f3589),
	.w6(32'hbadb4f87),
	.w7(32'h3b05dfb2),
	.w8(32'hbb93dfe9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb89313),
	.w1(32'hba224d24),
	.w2(32'h3b38d6ed),
	.w3(32'hbaf5c2fa),
	.w4(32'hba94b3cc),
	.w5(32'hb9f45136),
	.w6(32'hbc03a176),
	.w7(32'h3a4e59e6),
	.w8(32'hbb3a8cfe),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9719e),
	.w1(32'hbbbf32ac),
	.w2(32'hbae3f7c1),
	.w3(32'h3a42dfbd),
	.w4(32'hbb807a85),
	.w5(32'hbbb5cbe5),
	.w6(32'hb9c65f6e),
	.w7(32'hbbb430e1),
	.w8(32'hbb8a801b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91c42e),
	.w1(32'hbc621114),
	.w2(32'hbb5fd03b),
	.w3(32'hbbdd86bc),
	.w4(32'hbbd16628),
	.w5(32'hbc176c0b),
	.w6(32'hbbddf99c),
	.w7(32'hb982f01c),
	.w8(32'h3b39e113),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb6a67),
	.w1(32'hb9ff831a),
	.w2(32'hbbf06b57),
	.w3(32'hb9d689da),
	.w4(32'h3af7d3aa),
	.w5(32'hbb202718),
	.w6(32'h3bf51066),
	.w7(32'h3b0b2d42),
	.w8(32'h3a82e846),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc10fb5),
	.w1(32'hbb78cc8c),
	.w2(32'hba15459e),
	.w3(32'hbbc19209),
	.w4(32'h3a6dfa98),
	.w5(32'h38633e34),
	.w6(32'hbb86ef71),
	.w7(32'h3b56feea),
	.w8(32'h3b9c4878),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4bc13),
	.w1(32'h3bdcc324),
	.w2(32'hbb0771f1),
	.w3(32'hb922f66d),
	.w4(32'h3ac20756),
	.w5(32'hbb6da05f),
	.w6(32'h3ba28769),
	.w7(32'h3bcaecfa),
	.w8(32'h3b2764e8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ecc72),
	.w1(32'h3a7f28ff),
	.w2(32'hbb6bb521),
	.w3(32'hba8d8fe0),
	.w4(32'h393e4578),
	.w5(32'hbb4c1a14),
	.w6(32'hbb1f45e8),
	.w7(32'h381d4412),
	.w8(32'hba83ed27),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e4632),
	.w1(32'h391107cd),
	.w2(32'hbb273e7c),
	.w3(32'hbb220587),
	.w4(32'hbb9c116f),
	.w5(32'hbc35b6a0),
	.w6(32'hbb742c2b),
	.w7(32'h3b993734),
	.w8(32'hbaf06000),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93497f8),
	.w1(32'hbba453df),
	.w2(32'h3ac1e3d5),
	.w3(32'hbc0707a2),
	.w4(32'hbaffa02e),
	.w5(32'h3c8bd03d),
	.w6(32'hbc8e1e08),
	.w7(32'hbb3f857d),
	.w8(32'h3bb9048b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb338df6),
	.w1(32'hb9e1f8bc),
	.w2(32'h3c0cf94a),
	.w3(32'h390cfb87),
	.w4(32'h3b7bc9b8),
	.w5(32'h3b528674),
	.w6(32'hbb689168),
	.w7(32'h3b84c031),
	.w8(32'h3c12ff09),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5b812),
	.w1(32'hba5a93bf),
	.w2(32'h39d9a089),
	.w3(32'hb99b54b5),
	.w4(32'hbbbcfb22),
	.w5(32'hba5b9ba1),
	.w6(32'h3ab70a69),
	.w7(32'hbc04700a),
	.w8(32'hbc3e1dc8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b880960),
	.w1(32'h3b8a2cc6),
	.w2(32'h3ba0a642),
	.w3(32'hb98181cc),
	.w4(32'h3be71a1a),
	.w5(32'h3b3a36ca),
	.w6(32'hbc0d2623),
	.w7(32'h3b13e901),
	.w8(32'h3bc360db),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc96d1),
	.w1(32'h3abe6817),
	.w2(32'hbbd089b1),
	.w3(32'h3bab02dd),
	.w4(32'hbb927f17),
	.w5(32'hbbf160be),
	.w6(32'h3b570ffe),
	.w7(32'hbb17dfbf),
	.w8(32'hbb63f5f5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87a79d),
	.w1(32'hbb785af8),
	.w2(32'h3b2664ac),
	.w3(32'hbb9aa8b7),
	.w4(32'hbbbd3a02),
	.w5(32'hb9dba3b1),
	.w6(32'hbb86d3c2),
	.w7(32'h3a9aa6a2),
	.w8(32'hbb43d003),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b852850),
	.w1(32'h3b482820),
	.w2(32'hbb4cbd8d),
	.w3(32'hbbb828fe),
	.w4(32'h3bd04b30),
	.w5(32'h39f64726),
	.w6(32'hbba0d932),
	.w7(32'h3aefb7e4),
	.w8(32'h3b04fbe6),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a38c4),
	.w1(32'h3b0c6819),
	.w2(32'h3c3fbff5),
	.w3(32'hbbd81a43),
	.w4(32'h3b7b1af4),
	.w5(32'h3c1f9344),
	.w6(32'hbbacb497),
	.w7(32'h3bcc997f),
	.w8(32'h3bc398ab),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b351c1a),
	.w1(32'h3b6aeac2),
	.w2(32'h3b9e9063),
	.w3(32'h3ba82aae),
	.w4(32'h3b2ae2b9),
	.w5(32'hbc747bc2),
	.w6(32'h3a94ef06),
	.w7(32'hbb991174),
	.w8(32'hbb67b45e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43fcbb),
	.w1(32'hbb98306e),
	.w2(32'h3c1f5d6f),
	.w3(32'h3aa2b8bc),
	.w4(32'hbb87f702),
	.w5(32'h390c18b8),
	.w6(32'hbb6fbee2),
	.w7(32'hbab6d5b5),
	.w8(32'h3aafdb28),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe77e28),
	.w1(32'h3ba3d9d1),
	.w2(32'h3c542c83),
	.w3(32'hbbbcda51),
	.w4(32'h3a34c495),
	.w5(32'h3b5ad31a),
	.w6(32'hbac10a46),
	.w7(32'hbbb99b9e),
	.w8(32'hbab97c06),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1839bb),
	.w1(32'hba4aaa31),
	.w2(32'h3a7b91c2),
	.w3(32'hbc323b46),
	.w4(32'hbaceeb31),
	.w5(32'hb910aad0),
	.w6(32'hbc0cb920),
	.w7(32'h3830a40b),
	.w8(32'hbbbf02fc),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8a893),
	.w1(32'h3b5af325),
	.w2(32'h3c388a79),
	.w3(32'h3a8f7fdb),
	.w4(32'hbb9f6b37),
	.w5(32'h3b4936c5),
	.w6(32'hbb90484f),
	.w7(32'hbbeb4368),
	.w8(32'h3abe0ddf),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04e893),
	.w1(32'hba6bd321),
	.w2(32'hbbb379d4),
	.w3(32'h3ad78d10),
	.w4(32'hba4e1be3),
	.w5(32'hbb16b253),
	.w6(32'h3993803a),
	.w7(32'hba9733bd),
	.w8(32'h3baf43b8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaccfcc),
	.w1(32'h3afba2be),
	.w2(32'hbbab7d6b),
	.w3(32'h3bbc32c0),
	.w4(32'h3b5e49d9),
	.w5(32'hb9e16472),
	.w6(32'h3c262a6f),
	.w7(32'h3b8f2526),
	.w8(32'hbaae1ff7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ba9b5),
	.w1(32'h3abe8652),
	.w2(32'hbb6dafe9),
	.w3(32'h3b92d024),
	.w4(32'h3af01ec6),
	.w5(32'h3a34f706),
	.w6(32'hbb17a33c),
	.w7(32'h3b754a2b),
	.w8(32'h3b275c42),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a906535),
	.w1(32'h3a4f0d9e),
	.w2(32'h3b88e5ae),
	.w3(32'hbae3c388),
	.w4(32'hba97f4b3),
	.w5(32'hbb0b0e8d),
	.w6(32'hba5b5e76),
	.w7(32'hbb315cb1),
	.w8(32'hba29882b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb490235),
	.w1(32'h3be0485e),
	.w2(32'h3c68da2c),
	.w3(32'h3b99d5aa),
	.w4(32'h3bdedc33),
	.w5(32'h3c8a6cae),
	.w6(32'h3b291656),
	.w7(32'h3bca62e8),
	.w8(32'h3ae7c733),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba59919),
	.w1(32'hbb103a7b),
	.w2(32'h3ba18ff6),
	.w3(32'h3b942c83),
	.w4(32'hba6bb79b),
	.w5(32'hbc0c43ed),
	.w6(32'h3b335315),
	.w7(32'h3a8bf125),
	.w8(32'hb994eba2),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c616c65),
	.w1(32'hbaec67f8),
	.w2(32'hbb3eeed3),
	.w3(32'h3bc4741c),
	.w4(32'hbb200556),
	.w5(32'hbbafcad4),
	.w6(32'h3b515fdc),
	.w7(32'hbb47d73b),
	.w8(32'hbba07c77),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad278f8),
	.w1(32'h3c06b302),
	.w2(32'h3bcdab3a),
	.w3(32'hba4d2ebf),
	.w4(32'h3bc8d160),
	.w5(32'h3cc0f0db),
	.w6(32'hbb053846),
	.w7(32'h3af48720),
	.w8(32'hb9180f4d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09603e),
	.w1(32'hbb20d406),
	.w2(32'hb9d5bc66),
	.w3(32'h3aef0fef),
	.w4(32'h388f6612),
	.w5(32'h394c9620),
	.w6(32'h3b0ab08c),
	.w7(32'hbaee47b2),
	.w8(32'h3a4e4190),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d9c59),
	.w1(32'hbb9d3d9c),
	.w2(32'hb9f0b452),
	.w3(32'h3a94672c),
	.w4(32'hbba7acf9),
	.w5(32'h3b875a60),
	.w6(32'hb88c205c),
	.w7(32'hbc0826ab),
	.w8(32'h3bdf2972),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb995a98),
	.w1(32'hbb260676),
	.w2(32'hbb6bb00d),
	.w3(32'hbba4cf13),
	.w4(32'hbab60bc7),
	.w5(32'hbb231e70),
	.w6(32'hbb03e06e),
	.w7(32'hbb0f54e2),
	.w8(32'h3b513b07),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004717),
	.w1(32'h3bfe6a6a),
	.w2(32'h3bf57804),
	.w3(32'hbb374f27),
	.w4(32'h3be06e7e),
	.w5(32'h3b2227d7),
	.w6(32'hbb00e0e0),
	.w7(32'hbb051ec7),
	.w8(32'hb99d2649),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2960b),
	.w1(32'hbc452934),
	.w2(32'hbc7505fa),
	.w3(32'h3b077630),
	.w4(32'hbc455c20),
	.w5(32'hbbd07a0c),
	.w6(32'h3afb484c),
	.w7(32'hbb0a0b2e),
	.w8(32'hbbe2744c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b3b3b),
	.w1(32'h394629ce),
	.w2(32'h3bd010e9),
	.w3(32'hbb20bfe3),
	.w4(32'h3beaeeff),
	.w5(32'hbbc9981b),
	.w6(32'hbbe6af5b),
	.w7(32'h3be90030),
	.w8(32'h3beb82df),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e5edd),
	.w1(32'h3c5cdf6e),
	.w2(32'h3c9ac24d),
	.w3(32'hbbed913a),
	.w4(32'h3cbf4e50),
	.w5(32'h3cc1f58f),
	.w6(32'hbacf834d),
	.w7(32'h3c098033),
	.w8(32'h3b6502bf),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc3bee),
	.w1(32'hbbac6550),
	.w2(32'h3bb041d0),
	.w3(32'h3cbd8bce),
	.w4(32'hbba4c59d),
	.w5(32'hbaf4f6be),
	.w6(32'h3ba8b98b),
	.w7(32'hbba27fa4),
	.w8(32'hbbbcd017),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cb648),
	.w1(32'hbb4c99eb),
	.w2(32'hbb2c23f2),
	.w3(32'hbb88eb14),
	.w4(32'hbaaa824c),
	.w5(32'h3beae8b8),
	.w6(32'hbae66fdc),
	.w7(32'hbb87481e),
	.w8(32'hbb63d0de),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7495ad),
	.w1(32'hbb99f2f4),
	.w2(32'hbb6262e6),
	.w3(32'h3aa03dfa),
	.w4(32'h3a3fd529),
	.w5(32'hbbbaa17b),
	.w6(32'hbba74152),
	.w7(32'h3b49e7c0),
	.w8(32'hb8b062dd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1159a),
	.w1(32'h3b6999c5),
	.w2(32'h3bb224f2),
	.w3(32'h3ae7bb97),
	.w4(32'h3b23b682),
	.w5(32'h3c217156),
	.w6(32'hbafb53ca),
	.w7(32'hbbcc842b),
	.w8(32'hbbc29b60),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae61db5),
	.w1(32'hb894cf61),
	.w2(32'h3bc39a8f),
	.w3(32'h3a99e060),
	.w4(32'hba493d91),
	.w5(32'hba08da70),
	.w6(32'hbc0148b3),
	.w7(32'h3acdaaef),
	.w8(32'hbb91a970),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28e8eb),
	.w1(32'h3c151d97),
	.w2(32'h3c0155fa),
	.w3(32'h3af19e10),
	.w4(32'hbb08fa45),
	.w5(32'h3b5facbf),
	.w6(32'hba9a8c86),
	.w7(32'hbb16f968),
	.w8(32'hbb498af0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa202bc),
	.w1(32'hbaa5d1e0),
	.w2(32'h3b71eb30),
	.w3(32'hbb1d5805),
	.w4(32'hb97b92e1),
	.w5(32'hbba2faa6),
	.w6(32'h3aa92923),
	.w7(32'hb943fcc6),
	.w8(32'h39ec8f80),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd0f25),
	.w1(32'hbad54dce),
	.w2(32'h3a845566),
	.w3(32'hbc036a20),
	.w4(32'hbb58adb4),
	.w5(32'hbca23a49),
	.w6(32'h3b5443be),
	.w7(32'hbb80bd11),
	.w8(32'hbbac377d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00867e),
	.w1(32'hbba4d0ab),
	.w2(32'h3b4a3cf0),
	.w3(32'hbb8566cd),
	.w4(32'h3a841b3d),
	.w5(32'h3a595c24),
	.w6(32'hbacd6fca),
	.w7(32'hb737eaa7),
	.w8(32'h3b4662e6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39f38a),
	.w1(32'hbb8a8097),
	.w2(32'h3a89622f),
	.w3(32'h3bc13ea6),
	.w4(32'hbb64a5bf),
	.w5(32'h3c2c5da3),
	.w6(32'hbb116668),
	.w7(32'hbb46de91),
	.w8(32'h3aabbcb2),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa69372),
	.w1(32'h3a65daa0),
	.w2(32'h3b152777),
	.w3(32'h391aca04),
	.w4(32'hbb785033),
	.w5(32'h3b9e8401),
	.w6(32'hbacd64bf),
	.w7(32'hba379fd2),
	.w8(32'hbb2782bc),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60e929),
	.w1(32'hba0b8aca),
	.w2(32'h38fe7229),
	.w3(32'h3a2f0806),
	.w4(32'hbb1f5e57),
	.w5(32'hbb88cf75),
	.w6(32'hb84d0cb9),
	.w7(32'h3a26ec43),
	.w8(32'h3b8c4344),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3508ba),
	.w1(32'hba01e4b4),
	.w2(32'h3be990a2),
	.w3(32'h3af8d3fb),
	.w4(32'hbb8c55e0),
	.w5(32'hba9d8a73),
	.w6(32'h3bc7c8cd),
	.w7(32'hbb1f599f),
	.w8(32'h3a0eac79),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043329),
	.w1(32'hba86994f),
	.w2(32'hb9bb1ee7),
	.w3(32'h3be552ec),
	.w4(32'h3a28590a),
	.w5(32'h3c5804ee),
	.w6(32'hbb48d0e4),
	.w7(32'hbc42cba9),
	.w8(32'hbb979eb0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6659f9),
	.w1(32'hbbaaeb76),
	.w2(32'hbb2a8954),
	.w3(32'hbb2d0949),
	.w4(32'hbac2e676),
	.w5(32'h3b351308),
	.w6(32'hbba82336),
	.w7(32'hbb155d0e),
	.w8(32'hbb38471c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab9336),
	.w1(32'h3b8143ca),
	.w2(32'h3a9ef135),
	.w3(32'hbad717a9),
	.w4(32'h3b6cbef0),
	.w5(32'h3b1e2e4c),
	.w6(32'hbb833146),
	.w7(32'h3b00e5f3),
	.w8(32'h3a52acf0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f62c2),
	.w1(32'h3a31f21c),
	.w2(32'hbb3b5fe8),
	.w3(32'h3b8d7a1d),
	.w4(32'h391c6f4c),
	.w5(32'hb9f4ab77),
	.w6(32'h3b7dcddd),
	.w7(32'h3b994183),
	.w8(32'h3b512eb2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf2b04),
	.w1(32'h3bbbc1d8),
	.w2(32'h3c973167),
	.w3(32'h3a93a201),
	.w4(32'h3b645bb8),
	.w5(32'h3bb3cbdb),
	.w6(32'h3be7564d),
	.w7(32'h3c03c347),
	.w8(32'h3aed8c1b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b789f6c),
	.w1(32'hb9d05c60),
	.w2(32'h3bf62b01),
	.w3(32'hbbe6a5c8),
	.w4(32'hbb09642e),
	.w5(32'hbb47b94b),
	.w6(32'hbbd67340),
	.w7(32'hbc2b485b),
	.w8(32'hbbd8fb6c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37f6fb),
	.w1(32'h3ab17e22),
	.w2(32'hbad279fc),
	.w3(32'h3a8b8a39),
	.w4(32'hb9aa0c6e),
	.w5(32'hbb200d96),
	.w6(32'hbbae5ee8),
	.w7(32'hbad3fe85),
	.w8(32'hb9cea784),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb75b5),
	.w1(32'h393f450a),
	.w2(32'h3ab36d40),
	.w3(32'hba32caa3),
	.w4(32'h3a367871),
	.w5(32'hbab87658),
	.w6(32'hbb60e090),
	.w7(32'h3aa8f030),
	.w8(32'h3ab2fcf9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad2e1b),
	.w1(32'hbb7cb7b7),
	.w2(32'h3c45b23c),
	.w3(32'hbad01793),
	.w4(32'hb79276a6),
	.w5(32'h3b6e572b),
	.w6(32'h3a4e800f),
	.w7(32'h39b9832b),
	.w8(32'h3ba954b4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b830a07),
	.w1(32'hba8785db),
	.w2(32'h3c2b07b3),
	.w3(32'h3bf37120),
	.w4(32'h3b25577a),
	.w5(32'h3aadc28b),
	.w6(32'h3bd9d84a),
	.w7(32'hbba61528),
	.w8(32'hbb26b86d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2570a),
	.w1(32'h390ca6a1),
	.w2(32'hb94e53cc),
	.w3(32'h3bb05891),
	.w4(32'hba8448e1),
	.w5(32'h3b1e511a),
	.w6(32'hbb43369a),
	.w7(32'hbb84702f),
	.w8(32'hbaf127a6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e1abb),
	.w1(32'h3c1bf14a),
	.w2(32'h3a1c363d),
	.w3(32'hba030f00),
	.w4(32'hb91d8770),
	.w5(32'hbb385a6b),
	.w6(32'hbb70ff84),
	.w7(32'hbbcab36f),
	.w8(32'hbc8a19b1),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab31c67),
	.w1(32'h39d9f368),
	.w2(32'h3c2bd190),
	.w3(32'hba68ad77),
	.w4(32'hba52759c),
	.w5(32'hbc0e5652),
	.w6(32'hbac7636e),
	.w7(32'h3b993a64),
	.w8(32'h3b020569),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba122485),
	.w1(32'h354bbd60),
	.w2(32'h3b8e60b7),
	.w3(32'h3ab29b77),
	.w4(32'hbbb72b8e),
	.w5(32'hbc59a79b),
	.w6(32'h3a86fab5),
	.w7(32'hbbd549dd),
	.w8(32'hbbbfe484),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d2912),
	.w1(32'h3be8a1a1),
	.w2(32'h3ce2ac48),
	.w3(32'hba91a30c),
	.w4(32'hbb1de93a),
	.w5(32'h3c9fe203),
	.w6(32'hbac1d482),
	.w7(32'hba11830e),
	.w8(32'h3b8b6bed),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf1cfc),
	.w1(32'h3bad096e),
	.w2(32'h3c0d46bc),
	.w3(32'h3ca1f0ec),
	.w4(32'h3b36406b),
	.w5(32'h3beb0a7e),
	.w6(32'h3b864949),
	.w7(32'h39901f17),
	.w8(32'h3a8d7eb8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95da33),
	.w1(32'hba96b6a3),
	.w2(32'h3be1ad1e),
	.w3(32'h3c619b3f),
	.w4(32'h3bab4871),
	.w5(32'h3c1a0568),
	.w6(32'h3a461f71),
	.w7(32'h3b9ac318),
	.w8(32'h3c1c2612),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c425a50),
	.w1(32'hbbab70fb),
	.w2(32'hbbcc6bed),
	.w3(32'h3b9b5291),
	.w4(32'hbb3f0431),
	.w5(32'hbb1aeec5),
	.w6(32'h3bc86003),
	.w7(32'hba83cef9),
	.w8(32'h3c098b33),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37ce7a),
	.w1(32'h3bea7c36),
	.w2(32'h3ad35043),
	.w3(32'hbab3979a),
	.w4(32'h3bbda35c),
	.w5(32'h3c27540f),
	.w6(32'h3b2ad1a0),
	.w7(32'h3c18b399),
	.w8(32'h3ba5884f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b5212),
	.w1(32'h3c01bcbc),
	.w2(32'h3d03728a),
	.w3(32'h3b2ac847),
	.w4(32'hbb3c4a81),
	.w5(32'h3c925dbc),
	.w6(32'hbb43890c),
	.w7(32'h3b50fd26),
	.w8(32'h3bc3e89a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba88ff0),
	.w1(32'h3ca38dd0),
	.w2(32'h3d0e3b40),
	.w3(32'h3c478b11),
	.w4(32'h3c388b91),
	.w5(32'h3c2a2384),
	.w6(32'h3bbfb673),
	.w7(32'h3bbe231d),
	.w8(32'hbb3c4822),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e8ae3),
	.w1(32'h3bb3c819),
	.w2(32'h3c6decaf),
	.w3(32'h3ccd0447),
	.w4(32'hb968091d),
	.w5(32'h3baedb37),
	.w6(32'h39df0aca),
	.w7(32'hbb33b527),
	.w8(32'hbb58cbbd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3539e),
	.w1(32'h3b344a7a),
	.w2(32'hbb2401b9),
	.w3(32'h3bb23aa5),
	.w4(32'h3a09d514),
	.w5(32'hbba21556),
	.w6(32'hba64b8d7),
	.w7(32'hbab94108),
	.w8(32'hbb8a80d8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e8019),
	.w1(32'h3b812626),
	.w2(32'h3c0b1bb9),
	.w3(32'hbc098c07),
	.w4(32'h3aeb0a06),
	.w5(32'h3b50f995),
	.w6(32'hbc0dfffd),
	.w7(32'h3aa09925),
	.w8(32'h3bd3edf3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28a72d),
	.w1(32'hb7a152be),
	.w2(32'h3bb40635),
	.w3(32'h3b8dc012),
	.w4(32'h3b95734f),
	.w5(32'h3bafff2d),
	.w6(32'h3bf01f70),
	.w7(32'h3b5f8368),
	.w8(32'h3b8b1a4a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1727a),
	.w1(32'hbbd0efe4),
	.w2(32'h3aa1f26d),
	.w3(32'h3c13c872),
	.w4(32'hbbde0e21),
	.w5(32'hbba2399c),
	.w6(32'h3c1a39a0),
	.w7(32'hbbecd997),
	.w8(32'h3b7ee2bf),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b25e6),
	.w1(32'h3981927c),
	.w2(32'h3bc6cdec),
	.w3(32'h3aba39ad),
	.w4(32'hbb23fad2),
	.w5(32'hba117a87),
	.w6(32'h3b542d15),
	.w7(32'h3a3d6727),
	.w8(32'h3b8d1db4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7be484),
	.w1(32'h3bae2bbb),
	.w2(32'h3c73cb25),
	.w3(32'h3c148695),
	.w4(32'h3c1b1906),
	.w5(32'hbbac77d0),
	.w6(32'h3c130d27),
	.w7(32'h3b9ba310),
	.w8(32'h3bf1b3a1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15e117),
	.w1(32'h398f1315),
	.w2(32'hbb3766e4),
	.w3(32'h3bfe60a4),
	.w4(32'hb94f493c),
	.w5(32'hbb3ff6cb),
	.w6(32'hbb05e121),
	.w7(32'hbb0394e9),
	.w8(32'hbbd72151),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32de73),
	.w1(32'h39821454),
	.w2(32'h3c192db0),
	.w3(32'hbbc8e470),
	.w4(32'h3bb884f6),
	.w5(32'h3abff916),
	.w6(32'hbc30cc6b),
	.w7(32'h3944b0bc),
	.w8(32'h3b1d1ecb),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8531e),
	.w1(32'hbb462944),
	.w2(32'h3ae7786f),
	.w3(32'h3beedc69),
	.w4(32'hbc3db6b9),
	.w5(32'hbabfec5b),
	.w6(32'h3b8685f9),
	.w7(32'hbbcb65fa),
	.w8(32'hba8b9eda),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f9452),
	.w1(32'h3b360059),
	.w2(32'hbb9128cb),
	.w3(32'hbade27e0),
	.w4(32'h3beb35b1),
	.w5(32'hbc3dc675),
	.w6(32'hbb9c830c),
	.w7(32'h3ae1bce5),
	.w8(32'hbaf0b7bb),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7b502),
	.w1(32'hbb010631),
	.w2(32'h3b13451e),
	.w3(32'hba93f45a),
	.w4(32'hb9c0abd8),
	.w5(32'hbb6b41fe),
	.w6(32'h39832de0),
	.w7(32'h3b236484),
	.w8(32'hbb66ad5d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed2a0),
	.w1(32'hba70b520),
	.w2(32'hbb06e335),
	.w3(32'hbc3d845a),
	.w4(32'h39409215),
	.w5(32'h3b447964),
	.w6(32'hbc138975),
	.w7(32'hba8d0cd3),
	.w8(32'h3b2b1469),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb893187),
	.w1(32'h3c15820e),
	.w2(32'h3be71b7b),
	.w3(32'h3b00857a),
	.w4(32'hbc24665f),
	.w5(32'hbc49a418),
	.w6(32'hbb193429),
	.w7(32'h3b17a25b),
	.w8(32'h3a96e094),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2efc3c),
	.w1(32'h3b72586f),
	.w2(32'hbaa61c19),
	.w3(32'hbb00de26),
	.w4(32'h3abca15e),
	.w5(32'hbb5cd182),
	.w6(32'h3b796d2d),
	.w7(32'h3af11737),
	.w8(32'hbb4bdf92),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8a032),
	.w1(32'hbb6bc5ad),
	.w2(32'hba54cf1f),
	.w3(32'h398899fa),
	.w4(32'h3a3bcf54),
	.w5(32'h3b82efe7),
	.w6(32'hbaccdaed),
	.w7(32'hbbce09a6),
	.w8(32'hba2cc396),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb645d9),
	.w1(32'hbab1dbfd),
	.w2(32'h3b436976),
	.w3(32'h3c1b0cc6),
	.w4(32'hbc077124),
	.w5(32'hbadff0cf),
	.w6(32'h3b0ed408),
	.w7(32'hbb41ae2e),
	.w8(32'hba40bb7e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf969c2),
	.w1(32'h3bd2e7f8),
	.w2(32'h3c044b1b),
	.w3(32'hbb22032e),
	.w4(32'h35ca0954),
	.w5(32'h3c1a3fd8),
	.w6(32'h3b804dc8),
	.w7(32'h3b9b7053),
	.w8(32'h3c15c89e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe0495),
	.w1(32'h39d148c1),
	.w2(32'h3bb402ee),
	.w3(32'h3c056eed),
	.w4(32'hbbd35439),
	.w5(32'hbbc51fa2),
	.w6(32'h3c036c70),
	.w7(32'hbb292f6b),
	.w8(32'h399f37c5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c090c43),
	.w1(32'h39817977),
	.w2(32'h3aa81696),
	.w3(32'h3b7e3586),
	.w4(32'h3c5f9b2f),
	.w5(32'h3c6b5fd4),
	.w6(32'h3b45ea2a),
	.w7(32'h3b6cab22),
	.w8(32'h3aa8d41f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3c112),
	.w1(32'hbc0cfad8),
	.w2(32'hbb5b078e),
	.w3(32'h3c6c7b56),
	.w4(32'hbc7c9cbf),
	.w5(32'hbc8cd813),
	.w6(32'h3c00f073),
	.w7(32'hbc0bb60f),
	.w8(32'hbc00fd20),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b991f),
	.w1(32'hbba3cebf),
	.w2(32'hbbdf8bce),
	.w3(32'hbc6b0e5b),
	.w4(32'hbb8101d7),
	.w5(32'hbb5cb704),
	.w6(32'hbbdd045a),
	.w7(32'hbbed5ae0),
	.w8(32'hbb4ad308),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f870e),
	.w1(32'h3b2750f8),
	.w2(32'hbb57085a),
	.w3(32'h3aa3a6c9),
	.w4(32'hbb4af76f),
	.w5(32'hba23d7f7),
	.w6(32'hbb22838a),
	.w7(32'hbc09508b),
	.w8(32'hbb3d21bc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0578e6),
	.w1(32'hbbb789f3),
	.w2(32'h3bdf03d9),
	.w3(32'hbbf9aa2a),
	.w4(32'hbbe91df7),
	.w5(32'hbb217974),
	.w6(32'hbc3eab70),
	.w7(32'hbbda3ec9),
	.w8(32'hbaf3cd5e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fc747),
	.w1(32'hba8b0a35),
	.w2(32'hbaad3ae9),
	.w3(32'hba73a0e0),
	.w4(32'hbb0e9fa1),
	.w5(32'h3bd8a5df),
	.w6(32'h39ff70e2),
	.w7(32'hba0d2632),
	.w8(32'hba698c6b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f44f5),
	.w1(32'h3b3ed966),
	.w2(32'h3b88c81a),
	.w3(32'hbbd8cd47),
	.w4(32'h3ba15403),
	.w5(32'hba3e9824),
	.w6(32'hbad0e2aa),
	.w7(32'h3bfba632),
	.w8(32'h3b75c2b4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b519f96),
	.w1(32'h3bc3c9c4),
	.w2(32'h3ae60b0d),
	.w3(32'h3a94794b),
	.w4(32'h3c05c90e),
	.w5(32'h3a918483),
	.w6(32'hbbd6c741),
	.w7(32'h3ca47c84),
	.w8(32'hbaf2d8b3),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4f951),
	.w1(32'h3c07b2d6),
	.w2(32'h3a4b480e),
	.w3(32'hbbc862c0),
	.w4(32'h3bbd9927),
	.w5(32'h39da80be),
	.w6(32'hbc0ce0e8),
	.w7(32'hbb2c4171),
	.w8(32'hbacb34fd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8564ec),
	.w1(32'hbc9c164c),
	.w2(32'h3a5e4c79),
	.w3(32'h3c3e00a2),
	.w4(32'hbc808d09),
	.w5(32'h3b7fe031),
	.w6(32'h3b773d8b),
	.w7(32'hbc566c33),
	.w8(32'h3ac9a4b7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dbcdb),
	.w1(32'h3a8bd5b2),
	.w2(32'h3bd31334),
	.w3(32'hbb38e638),
	.w4(32'h3ae1dc7e),
	.w5(32'h3af49b40),
	.w6(32'hbc278521),
	.w7(32'hbbd6b136),
	.w8(32'h3763e852),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba451697),
	.w1(32'h3b90ad07),
	.w2(32'h3ba13cd0),
	.w3(32'hb96e91d2),
	.w4(32'hbb07ddfb),
	.w5(32'h3be9c896),
	.w6(32'hbb5fac84),
	.w7(32'hbaa081d5),
	.w8(32'h3c196a2f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a75a0),
	.w1(32'hbbbedb4e),
	.w2(32'hbbc66750),
	.w3(32'h3bbc94bb),
	.w4(32'h3b0d9fb8),
	.w5(32'hb99720b0),
	.w6(32'h3c59640d),
	.w7(32'h3b6a166f),
	.w8(32'hba624150),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3515bb),
	.w1(32'h3aff47a6),
	.w2(32'hba46dd73),
	.w3(32'h3c5ac1be),
	.w4(32'h3b934be9),
	.w5(32'h3bd63b06),
	.w6(32'h3bf27ebb),
	.w7(32'h3b541f49),
	.w8(32'hbbb61e55),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a256b0d),
	.w1(32'h3c4b9dde),
	.w2(32'hb9a28354),
	.w3(32'h3bcb2576),
	.w4(32'hbb2e9722),
	.w5(32'hbb86e1f1),
	.w6(32'hbb896768),
	.w7(32'h3aa2d4b7),
	.w8(32'h3bde47b2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a7964),
	.w1(32'h3b897914),
	.w2(32'hbbf0f24c),
	.w3(32'hbb10e6f7),
	.w4(32'h3ca189cd),
	.w5(32'h3b4f44c6),
	.w6(32'h3ba12c6c),
	.w7(32'h3a981461),
	.w8(32'hbc074c60),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8c057),
	.w1(32'hbaaaeaa3),
	.w2(32'h3b2ded5e),
	.w3(32'h3c02a14e),
	.w4(32'hbba66ad4),
	.w5(32'h3b27662c),
	.w6(32'hbb457978),
	.w7(32'h3ba2c913),
	.w8(32'h3bd5c954),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5fb4a),
	.w1(32'hbbe34366),
	.w2(32'hbbba4c4e),
	.w3(32'hbc5765c5),
	.w4(32'hbb828df8),
	.w5(32'hbb81e669),
	.w6(32'hbc033acd),
	.w7(32'hbc2b65cd),
	.w8(32'hbb39e37a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0942f4),
	.w1(32'hbc091642),
	.w2(32'h3b0e1b4a),
	.w3(32'h399192c4),
	.w4(32'hbab3c09e),
	.w5(32'h3be97bec),
	.w6(32'hba4dad14),
	.w7(32'hbbb42c33),
	.w8(32'h3b7a3142),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21d706),
	.w1(32'h3a6a4660),
	.w2(32'h3ca0c2f8),
	.w3(32'h3c106d68),
	.w4(32'h3c2df643),
	.w5(32'h3c976efc),
	.w6(32'hb9252d48),
	.w7(32'h3c12ee53),
	.w8(32'h3b34cf23),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90e2a4),
	.w1(32'h3b316e06),
	.w2(32'h3b871ab5),
	.w3(32'h3c8a4586),
	.w4(32'hbba75d6c),
	.w5(32'h3b6223c5),
	.w6(32'hbbcb49e6),
	.w7(32'hbb3e111c),
	.w8(32'h39d95c9a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79ec96),
	.w1(32'h3b002a43),
	.w2(32'h3ad29d0a),
	.w3(32'h3b2e72ee),
	.w4(32'hb951cd7a),
	.w5(32'h3bcd4b62),
	.w6(32'hb98e0980),
	.w7(32'h3997aaf6),
	.w8(32'h3aefda9d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc42a2b),
	.w1(32'hbb0c615e),
	.w2(32'h3bb3c13c),
	.w3(32'hbb776e2b),
	.w4(32'h3a187e6a),
	.w5(32'h3b60c3e1),
	.w6(32'hbbfa22e1),
	.w7(32'hbbb9d6c1),
	.w8(32'hbb7cfe1c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41be15),
	.w1(32'hbbb20d13),
	.w2(32'hbba22384),
	.w3(32'hbb260edf),
	.w4(32'hbbc94b53),
	.w5(32'hbc1374c4),
	.w6(32'hbb9c4c01),
	.w7(32'hbbc047f0),
	.w8(32'hbc07a320),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecfce7),
	.w1(32'h3bd97015),
	.w2(32'h3b19efde),
	.w3(32'hbc001747),
	.w4(32'hb4c6d902),
	.w5(32'hb7d6aa17),
	.w6(32'hbc156aae),
	.w7(32'hb82276c3),
	.w8(32'h3b850c6c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea82b2),
	.w1(32'hb820b2e4),
	.w2(32'h3ad9056f),
	.w3(32'h3aec53ed),
	.w4(32'hbafb3374),
	.w5(32'hbafd8d44),
	.w6(32'hbbbf894b),
	.w7(32'hbb60a06c),
	.w8(32'hba8858cd),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1429a),
	.w1(32'hbc1cdd74),
	.w2(32'hbb784374),
	.w3(32'hbc336542),
	.w4(32'hbc88262f),
	.w5(32'hbc04bc9b),
	.w6(32'hbb8e2bbb),
	.w7(32'hbbff3063),
	.w8(32'hbb541418),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8bba4),
	.w1(32'hbb1346dc),
	.w2(32'h39de5403),
	.w3(32'hbc2d8825),
	.w4(32'h3ab5358d),
	.w5(32'h3c0acaf8),
	.w6(32'hbc09ae14),
	.w7(32'h39ea88d5),
	.w8(32'h3bc61dd7),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba99d22),
	.w1(32'hbb18451c),
	.w2(32'h3aaac74d),
	.w3(32'hbbb6277e),
	.w4(32'h3b94841b),
	.w5(32'hbb74669d),
	.w6(32'h3b0cf3db),
	.w7(32'h3a8119a1),
	.w8(32'hba3f46ed),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09e46e),
	.w1(32'h3b7f9a6c),
	.w2(32'hbaafe592),
	.w3(32'hba3a1b72),
	.w4(32'h3b206037),
	.w5(32'hbbe9e9cc),
	.w6(32'hbb0fd492),
	.w7(32'h3b7ac0de),
	.w8(32'hbb5c4a74),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b909532),
	.w1(32'hbbd538d7),
	.w2(32'hbbb05012),
	.w3(32'h3c0865bb),
	.w4(32'hbb573510),
	.w5(32'hbb3ae365),
	.w6(32'hbaaf4ec1),
	.w7(32'h3a39930b),
	.w8(32'h3b84971d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9909e4),
	.w1(32'h3bf8f204),
	.w2(32'h3c36f5a1),
	.w3(32'hbb9ecc3e),
	.w4(32'hbb67229b),
	.w5(32'h3a1510eb),
	.w6(32'h3ae84493),
	.w7(32'h3ad5831d),
	.w8(32'h3bce7096),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31bae7),
	.w1(32'hbbac7be6),
	.w2(32'hba391589),
	.w3(32'hbc6f5367),
	.w4(32'hbbfedc34),
	.w5(32'h3a7b6631),
	.w6(32'hbc5cd3b7),
	.w7(32'hbc01e024),
	.w8(32'h393e05af),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51f9da),
	.w1(32'h3c0f0f85),
	.w2(32'h3c0209a6),
	.w3(32'hbb273e96),
	.w4(32'h3c18f939),
	.w5(32'h3bc323cf),
	.w6(32'h3b11a5f2),
	.w7(32'h3b52dc61),
	.w8(32'h3b565b77),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab225fc),
	.w1(32'h3b96662a),
	.w2(32'h3be26c58),
	.w3(32'h3b62dee8),
	.w4(32'h3b041966),
	.w5(32'h3c753b8b),
	.w6(32'h3abba72e),
	.w7(32'h3b20402d),
	.w8(32'h3c59a07c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed6bdf),
	.w1(32'hbbb61869),
	.w2(32'hbac20d6c),
	.w3(32'h3c9ef813),
	.w4(32'hbc0ab31e),
	.w5(32'hbbe38b49),
	.w6(32'h3c1e3034),
	.w7(32'hbb8e7dac),
	.w8(32'hbb18ba15),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb590444),
	.w1(32'hbb96d9b5),
	.w2(32'hbb9415ac),
	.w3(32'hbb902d71),
	.w4(32'hbba8cad7),
	.w5(32'hbc2b899b),
	.w6(32'hbb24980f),
	.w7(32'h39f9e6b2),
	.w8(32'hbbebe4f2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08b122),
	.w1(32'hbbc0684d),
	.w2(32'hbb1a4aa4),
	.w3(32'h3bdddc96),
	.w4(32'h3a9a5738),
	.w5(32'h3b9e7be1),
	.w6(32'h3b6266ae),
	.w7(32'hbbf7d466),
	.w8(32'hbba427bf),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae2d8),
	.w1(32'h3b8c3f46),
	.w2(32'h3bb362bc),
	.w3(32'hbba99cdd),
	.w4(32'h3b1f1127),
	.w5(32'h3bf17efc),
	.w6(32'hbc4bcf75),
	.w7(32'hbb344055),
	.w8(32'hbb19fba0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc054d),
	.w1(32'h3aabb08e),
	.w2(32'hbb944f96),
	.w3(32'h3bee7965),
	.w4(32'h3bf5cfe3),
	.w5(32'h3ab7cbfa),
	.w6(32'h3c15b35d),
	.w7(32'hbad52a64),
	.w8(32'hbb6c92ec),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bc54d),
	.w1(32'h3b478d45),
	.w2(32'hba1ad62c),
	.w3(32'h3adc38f6),
	.w4(32'h3b057d27),
	.w5(32'hba98aaa7),
	.w6(32'hb8ce41e0),
	.w7(32'hbb66dcba),
	.w8(32'hbb18f3db),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3182e),
	.w1(32'h3c092dd4),
	.w2(32'h3c01d80b),
	.w3(32'h3c42809e),
	.w4(32'h3c3b96a9),
	.w5(32'h3b845407),
	.w6(32'h3b85486b),
	.w7(32'h3bbc71bf),
	.w8(32'hb8a04dce),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c177428),
	.w1(32'hba8a31e3),
	.w2(32'hbb102f43),
	.w3(32'hbb4599a0),
	.w4(32'hbc282d79),
	.w5(32'hbbe62617),
	.w6(32'hbb955e07),
	.w7(32'hbb95dca5),
	.w8(32'hbb9e7b75),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc071e5),
	.w1(32'h3b8d1d8f),
	.w2(32'h3bb149c8),
	.w3(32'hbc4ceb8e),
	.w4(32'hbbbb6555),
	.w5(32'h3a2ff99c),
	.w6(32'hbc061077),
	.w7(32'h3a72496b),
	.w8(32'h3b4682ab),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba10739),
	.w1(32'h3bcdec76),
	.w2(32'h3b6165c6),
	.w3(32'hbc16c116),
	.w4(32'h3c05a9b4),
	.w5(32'hbbed9aa6),
	.w6(32'h3a9e0cfe),
	.w7(32'h3c20c949),
	.w8(32'hba0cd2f5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff7990),
	.w1(32'h3b49be9e),
	.w2(32'h3bc78319),
	.w3(32'hbc8f4dca),
	.w4(32'hbc14ca54),
	.w5(32'hbb8eeac7),
	.w6(32'hbb23971a),
	.w7(32'hbb602b3b),
	.w8(32'hb9bbc286),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba418d3c),
	.w1(32'h3bce22c1),
	.w2(32'h3ba30ad2),
	.w3(32'hba7fdb82),
	.w4(32'hbbf533a4),
	.w5(32'h3b09c411),
	.w6(32'hbba1fb29),
	.w7(32'hb89db71b),
	.w8(32'h3b6169ab),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb41a1d),
	.w1(32'h3b2526b4),
	.w2(32'hbae28d8c),
	.w3(32'h3b4ec7b3),
	.w4(32'hbbf47f05),
	.w5(32'hbbafb0b1),
	.w6(32'h3b207009),
	.w7(32'hbc3111a2),
	.w8(32'hbc161f6b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule