module layer_10_featuremap_272(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3fef3),
	.w1(32'h3bc85b2d),
	.w2(32'h3af35bd5),
	.w3(32'h3c16b4e4),
	.w4(32'h3b88e532),
	.w5(32'h3aa17043),
	.w6(32'h3c4cebbb),
	.w7(32'h3a91739b),
	.w8(32'h3a7d121e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9549238),
	.w1(32'hbbb17f2c),
	.w2(32'hbbf08763),
	.w3(32'h39849ad5),
	.w4(32'hbba71db2),
	.w5(32'h3a21e0c0),
	.w6(32'hba66c7e9),
	.w7(32'hbb926ea1),
	.w8(32'hbb383e61),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14c2b1),
	.w1(32'h3a0f7595),
	.w2(32'h3ad38d9c),
	.w3(32'hbb8ee7f0),
	.w4(32'h3baf10f6),
	.w5(32'hbb82a48f),
	.w6(32'hbb7a29b3),
	.w7(32'hbb521ef9),
	.w8(32'hbb739961),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb284064),
	.w1(32'hbb1a0058),
	.w2(32'hbb3d89e9),
	.w3(32'hbae71cb2),
	.w4(32'hbb6b5c60),
	.w5(32'h3a35c7bb),
	.w6(32'hbb4490f4),
	.w7(32'hbb6dc249),
	.w8(32'h3b8f664c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0675b6),
	.w1(32'hbc3f9540),
	.w2(32'hbb7154e6),
	.w3(32'hbb26192b),
	.w4(32'h3aba2baf),
	.w5(32'h3b63dc78),
	.w6(32'hbbaf1e69),
	.w7(32'hbb6791f4),
	.w8(32'h3b7a5e60),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920702),
	.w1(32'h3a8ac662),
	.w2(32'hbadefd77),
	.w3(32'h3b38da2e),
	.w4(32'h3b38f569),
	.w5(32'hbb01ec9e),
	.w6(32'h3a8c908b),
	.w7(32'hb9ae106f),
	.w8(32'hbb1b2c6d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d8f4),
	.w1(32'h3afc91d2),
	.w2(32'hbb35080c),
	.w3(32'h3aa0bdd4),
	.w4(32'hba8a5c09),
	.w5(32'h3aff3ce7),
	.w6(32'h3b906ff0),
	.w7(32'hbba2d929),
	.w8(32'hb933b316),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba908fcd),
	.w1(32'h3c096778),
	.w2(32'h3bff4a28),
	.w3(32'hba91964f),
	.w4(32'h3a76fe53),
	.w5(32'h3bccbc24),
	.w6(32'h3bbfc31e),
	.w7(32'h3c0455ba),
	.w8(32'h3b6916d3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48e660),
	.w1(32'h3b1e35eb),
	.w2(32'h3ae8bb54),
	.w3(32'h3b22beec),
	.w4(32'h3b520038),
	.w5(32'h3b440732),
	.w6(32'h3b885b33),
	.w7(32'h3b6baef7),
	.w8(32'h3b363726),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54dfb0),
	.w1(32'h39773400),
	.w2(32'hbb3f64a4),
	.w3(32'h3b544c5f),
	.w4(32'hbac855eb),
	.w5(32'hbb07145f),
	.w6(32'hb9853e27),
	.w7(32'hbb8a9dba),
	.w8(32'hbb4e9558),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39803c),
	.w1(32'h3a07d72c),
	.w2(32'hbb1142e2),
	.w3(32'h3ba1fdbe),
	.w4(32'h3a29eda0),
	.w5(32'hbb10b5e6),
	.w6(32'h3b8fdd85),
	.w7(32'hbb96da65),
	.w8(32'h3b545775),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19ad0c),
	.w1(32'h3b3ee536),
	.w2(32'h3b0f1cb7),
	.w3(32'hbb94a852),
	.w4(32'h3a584007),
	.w5(32'h3b9c1a3d),
	.w6(32'hba881d08),
	.w7(32'h3b4f1f99),
	.w8(32'h3b80d351),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b303220),
	.w1(32'h3b352970),
	.w2(32'hb86c26ed),
	.w3(32'h3bc0f4f6),
	.w4(32'h3af6aa0e),
	.w5(32'h391796e1),
	.w6(32'h3b247d82),
	.w7(32'h3b15b619),
	.w8(32'hba8146e1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a60c4d),
	.w1(32'hba2c0a92),
	.w2(32'h399bd6db),
	.w3(32'h3b9a0ab1),
	.w4(32'hb8d4e028),
	.w5(32'hbbaba35e),
	.w6(32'h3be35920),
	.w7(32'h398bd3ae),
	.w8(32'hbb8386db),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97a541),
	.w1(32'hbb4f5fbb),
	.w2(32'hbb923bb7),
	.w3(32'hbb16c9b3),
	.w4(32'hbbb8eceb),
	.w5(32'h3b0918bf),
	.w6(32'hba568dcc),
	.w7(32'hbbc6b651),
	.w8(32'h3b4ab256),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb705cde),
	.w1(32'hbb4d4e8c),
	.w2(32'hbb626657),
	.w3(32'h3b82ec3d),
	.w4(32'h3ad72f7b),
	.w5(32'h3b97ff8f),
	.w6(32'h3c22c64a),
	.w7(32'hbacc9850),
	.w8(32'h3bcc1e55),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aa58a),
	.w1(32'hbb49a7b5),
	.w2(32'hb9e6f80e),
	.w3(32'hb7dccfaf),
	.w4(32'h3a14168b),
	.w5(32'hb802ba9a),
	.w6(32'hbbc1c8f5),
	.w7(32'h3aca95f7),
	.w8(32'hba9d8a2f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2e833),
	.w1(32'hba9e6ac4),
	.w2(32'h3af34cd7),
	.w3(32'h3b3890be),
	.w4(32'h3b8b1764),
	.w5(32'h3a3150f9),
	.w6(32'h3b1a53e1),
	.w7(32'h3b5b3b72),
	.w8(32'h3b44806a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d88ed),
	.w1(32'hbaa8ea6b),
	.w2(32'hb9cd08d2),
	.w3(32'hbaa68499),
	.w4(32'hbb0286fd),
	.w5(32'hba6780b2),
	.w6(32'h3a370879),
	.w7(32'h39d419c6),
	.w8(32'h3b158e49),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b92da),
	.w1(32'hba7ab6c4),
	.w2(32'hbb5e1323),
	.w3(32'h3b427d38),
	.w4(32'hb8edf821),
	.w5(32'h3ae1a8a5),
	.w6(32'h3a899199),
	.w7(32'hbace0b27),
	.w8(32'h3a272180),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbd973),
	.w1(32'hb9991ec5),
	.w2(32'hbb5a2d6d),
	.w3(32'h3c29c903),
	.w4(32'h3bf38a34),
	.w5(32'h3af3393d),
	.w6(32'h3c4ae855),
	.w7(32'h3b249942),
	.w8(32'h3b002174),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd70c31),
	.w1(32'h3c07da6a),
	.w2(32'h3bb4be97),
	.w3(32'hbb4fed19),
	.w4(32'hbb4463b3),
	.w5(32'hbb738c20),
	.w6(32'hbb062237),
	.w7(32'h3b96c10a),
	.w8(32'h3a40d7ff),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7543e8),
	.w1(32'hba484da2),
	.w2(32'hba505719),
	.w3(32'h3b05c971),
	.w4(32'h3b9a824c),
	.w5(32'hbb908136),
	.w6(32'h3b5085b4),
	.w7(32'hbaa04442),
	.w8(32'hbc24e2dd),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43ded6),
	.w1(32'hbb337bed),
	.w2(32'hbb8b19b8),
	.w3(32'h3c063294),
	.w4(32'h3a93fa54),
	.w5(32'h3ae2f579),
	.w6(32'h3c0569e7),
	.w7(32'hbb471b92),
	.w8(32'hba933d6d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a849508),
	.w1(32'h396f9765),
	.w2(32'h3b6fdddd),
	.w3(32'hb965861a),
	.w4(32'hbafc09bb),
	.w5(32'hbb2d747e),
	.w6(32'hbb9a6c47),
	.w7(32'hbb64d27c),
	.w8(32'hba0d0b8c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb158f44),
	.w1(32'h3b7a4e94),
	.w2(32'hbaafd583),
	.w3(32'h3b98f71c),
	.w4(32'hbbcb8e0b),
	.w5(32'h3a8a7aed),
	.w6(32'h3bdac822),
	.w7(32'hbbd47241),
	.w8(32'h3abdef93),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b203984),
	.w1(32'h3bb11c3e),
	.w2(32'h3b1163bd),
	.w3(32'h3b23a24f),
	.w4(32'hba706cc9),
	.w5(32'h3c4ca528),
	.w6(32'h3bccc17c),
	.w7(32'hb76862d8),
	.w8(32'h3c2c348d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c340b0c),
	.w1(32'h3af5bbec),
	.w2(32'h3b332fb3),
	.w3(32'h3b3a04fb),
	.w4(32'h3bf67af8),
	.w5(32'hbb1eb9f5),
	.w6(32'h3bb076b5),
	.w7(32'h3b6854e6),
	.w8(32'hbb557bec),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a51c8),
	.w1(32'hbae387dd),
	.w2(32'hbb986826),
	.w3(32'h3a52a5ab),
	.w4(32'hbb761e1e),
	.w5(32'hbc164d40),
	.w6(32'h3af314f4),
	.w7(32'hbb5a3ad4),
	.w8(32'hbbed323d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafa6be),
	.w1(32'hbb2100e5),
	.w2(32'hbb22ada9),
	.w3(32'h3b81c7a1),
	.w4(32'hbb56be8c),
	.w5(32'hbb2f3198),
	.w6(32'h3c359d01),
	.w7(32'hbb5cc023),
	.w8(32'h3b1d4759),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc12dd7),
	.w1(32'hbb372739),
	.w2(32'hbacbc99f),
	.w3(32'hbbb2e2ad),
	.w4(32'hba61ec0d),
	.w5(32'h3aa0f543),
	.w6(32'hba730308),
	.w7(32'hbb022fb1),
	.w8(32'h3b043988),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b8011),
	.w1(32'h3b606a73),
	.w2(32'h3ba5d564),
	.w3(32'hbacf436a),
	.w4(32'h3b40e5c1),
	.w5(32'h3a8c29aa),
	.w6(32'hbb262224),
	.w7(32'h3b82ae89),
	.w8(32'h3b507d2d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf7996),
	.w1(32'hbafb4296),
	.w2(32'h3b790426),
	.w3(32'h3aa4727d),
	.w4(32'hbbb64c02),
	.w5(32'hbafeb457),
	.w6(32'h3b303119),
	.w7(32'hba4f28e2),
	.w8(32'hbae96555),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea269c),
	.w1(32'hbb406422),
	.w2(32'hbaff984a),
	.w3(32'h3b4a0d96),
	.w4(32'h3b5def20),
	.w5(32'hba97d9fd),
	.w6(32'hb90080ad),
	.w7(32'h3b9a8556),
	.w8(32'hbb330383),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f6665),
	.w1(32'hba0b9127),
	.w2(32'h348cc9d0),
	.w3(32'hb97066d2),
	.w4(32'hbac8c668),
	.w5(32'hbb20e9a4),
	.w6(32'h3ac6a8f7),
	.w7(32'h3b16b46a),
	.w8(32'hbbe0a92c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb59dad),
	.w1(32'hbad318b3),
	.w2(32'hbb19228f),
	.w3(32'h3accb956),
	.w4(32'h3b532c18),
	.w5(32'hba2ffe85),
	.w6(32'h3b4422ef),
	.w7(32'hbacb8cc6),
	.w8(32'h3ac6f021),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba926e3d),
	.w1(32'hb9363ef4),
	.w2(32'hb90e8cb0),
	.w3(32'hb9b390fa),
	.w4(32'hbb111de3),
	.w5(32'h3baf3022),
	.w6(32'h3ab5f129),
	.w7(32'hba966e78),
	.w8(32'h3bf8351a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc30ce),
	.w1(32'h3c2ad1e3),
	.w2(32'hbb6b13ed),
	.w3(32'h3c362c60),
	.w4(32'hbb2caa19),
	.w5(32'h3bb1075d),
	.w6(32'h3ca955e0),
	.w7(32'hbb28cfe9),
	.w8(32'h3be83bc2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46d09e),
	.w1(32'hbb7f6eec),
	.w2(32'hbb8b6d47),
	.w3(32'h3ab7ace4),
	.w4(32'hbc07ff3f),
	.w5(32'hbb33e941),
	.w6(32'hbbe8b00f),
	.w7(32'hbc239418),
	.w8(32'hb906d0c2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b510296),
	.w1(32'h3b394f77),
	.w2(32'h3c06047f),
	.w3(32'h3a7eb9ff),
	.w4(32'h3b16edfd),
	.w5(32'h3b1aab0e),
	.w6(32'hbb20d99f),
	.w7(32'h3c3340fc),
	.w8(32'h3bab1f5d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda1f18),
	.w1(32'h3b6c8868),
	.w2(32'h3aee89c1),
	.w3(32'h3b261750),
	.w4(32'h3b4f829f),
	.w5(32'hba04a559),
	.w6(32'h3baf6710),
	.w7(32'h3bd3f084),
	.w8(32'h3a2b0838),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989450a),
	.w1(32'h3b850e9d),
	.w2(32'hbaa646b7),
	.w3(32'h3b78da15),
	.w4(32'hbb30cc4e),
	.w5(32'h395b68e0),
	.w6(32'h3b2714e3),
	.w7(32'hbbb43470),
	.w8(32'hb9be0dfa),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba585885),
	.w1(32'hba1bf56b),
	.w2(32'hbae5ec79),
	.w3(32'hb9ecd6e6),
	.w4(32'h3adf5e59),
	.w5(32'hbb92ae0a),
	.w6(32'h3ba8448f),
	.w7(32'hbaa969b0),
	.w8(32'hbbb6dc1e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac8143),
	.w1(32'hbb64f93c),
	.w2(32'h3a80e653),
	.w3(32'hbb6571b1),
	.w4(32'h3bc73823),
	.w5(32'hbb3bd899),
	.w6(32'hbb06f277),
	.w7(32'hba184dfc),
	.w8(32'hbb3b9157),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaad422),
	.w1(32'h3b336cfb),
	.w2(32'hba36bd8b),
	.w3(32'hbac4d599),
	.w4(32'hbba1d42d),
	.w5(32'h3b6d208d),
	.w6(32'h3acded4f),
	.w7(32'hb92be919),
	.w8(32'h3b5afe62),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be81486),
	.w1(32'h3bee337d),
	.w2(32'h3b96e111),
	.w3(32'hbae1cb9f),
	.w4(32'h3bd277f3),
	.w5(32'h3a45eac9),
	.w6(32'hbc173d12),
	.w7(32'hba47f893),
	.w8(32'h3b0424d5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b6be),
	.w1(32'h3b69bef7),
	.w2(32'h3b9bf405),
	.w3(32'h3b161a99),
	.w4(32'h3b53c2c4),
	.w5(32'h3c0bd240),
	.w6(32'h3b45116f),
	.w7(32'h3b8c0f19),
	.w8(32'h3bfae94b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd68404),
	.w1(32'h3b5f3b9c),
	.w2(32'h3a724796),
	.w3(32'h3ac4d12d),
	.w4(32'hbb25eeaf),
	.w5(32'hbb14ccc9),
	.w6(32'h3aeba1fe),
	.w7(32'h3ae868d3),
	.w8(32'hbb6604d8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb711335),
	.w1(32'hbb75cab6),
	.w2(32'hbb819e8e),
	.w3(32'hbad5ad3a),
	.w4(32'hbae2f7f2),
	.w5(32'hb92ee441),
	.w6(32'h39b7165d),
	.w7(32'hbb8a52d1),
	.w8(32'h3b179083),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b701254),
	.w1(32'h3baa415c),
	.w2(32'h3b498379),
	.w3(32'hba2418df),
	.w4(32'hbba990fd),
	.w5(32'h3b1f1fc6),
	.w6(32'h3b82cf7f),
	.w7(32'h3acf9250),
	.w8(32'hb9c0952a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b253dcc),
	.w1(32'hbb4713ee),
	.w2(32'h3acc759f),
	.w3(32'hba0580fe),
	.w4(32'hba490e7c),
	.w5(32'h3a781aab),
	.w6(32'hbac9f49e),
	.w7(32'h3a0b8a99),
	.w8(32'h3b2ca044),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9f795),
	.w1(32'hbad10bee),
	.w2(32'h3a294a62),
	.w3(32'hbac04c23),
	.w4(32'h3b56d2f2),
	.w5(32'hbb89dc41),
	.w6(32'hbaa2e581),
	.w7(32'h387eed4d),
	.w8(32'hbb7aaf53),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba787ea3),
	.w1(32'hbad3aa59),
	.w2(32'hbb6da220),
	.w3(32'h3951f0e3),
	.w4(32'h3b1e097b),
	.w5(32'hbbbad0e9),
	.w6(32'h3b83b62e),
	.w7(32'hbb7a426a),
	.w8(32'h3a8c0563),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1342fb),
	.w1(32'h3b2529ed),
	.w2(32'h3b056e09),
	.w3(32'h3b012590),
	.w4(32'h3b7a5cdf),
	.w5(32'h3a4aa0f6),
	.w6(32'h3bc249fe),
	.w7(32'h3aeaa8b1),
	.w8(32'h3bbcb9c1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15a1c3),
	.w1(32'h39ffa426),
	.w2(32'hbb1c8425),
	.w3(32'h3a0f6c06),
	.w4(32'h3b2c0e34),
	.w5(32'h3a338c43),
	.w6(32'hba481727),
	.w7(32'hbb489606),
	.w8(32'hbaf4c993),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a6bfc),
	.w1(32'hbae59d32),
	.w2(32'hbb800ccd),
	.w3(32'h3b8522cb),
	.w4(32'h3a622dbe),
	.w5(32'h3b3408df),
	.w6(32'h3adb34cc),
	.w7(32'hbab4a03d),
	.w8(32'h3b226786),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcc8e6),
	.w1(32'hba1b7a10),
	.w2(32'h3a04f6d4),
	.w3(32'hba8306a9),
	.w4(32'h3aa3315e),
	.w5(32'hbb593ba1),
	.w6(32'hbb4ac5cf),
	.w7(32'h3b1e3b6d),
	.w8(32'h39c58a58),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab6ab2),
	.w1(32'hb9acca00),
	.w2(32'hba9caa50),
	.w3(32'h3aedf5ce),
	.w4(32'h3b0e0752),
	.w5(32'hbb1babc1),
	.w6(32'h3b2fa675),
	.w7(32'h3a6beb17),
	.w8(32'hbaaf8443),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70ad49),
	.w1(32'h3b722ded),
	.w2(32'h3b746dde),
	.w3(32'hb886f1b5),
	.w4(32'hbb96a463),
	.w5(32'h3ac8dfcd),
	.w6(32'h3bdb97d2),
	.w7(32'hba8b8e22),
	.w8(32'h3a09c50f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc87a38),
	.w1(32'h3a3c6368),
	.w2(32'hbb139174),
	.w3(32'hbc438b6d),
	.w4(32'hbc14bd01),
	.w5(32'h3b05a6f6),
	.w6(32'hbc70fec7),
	.w7(32'hbc251a11),
	.w8(32'h3bd65dda),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b201ac9),
	.w1(32'hb9fb0914),
	.w2(32'hba74e868),
	.w3(32'h3b289702),
	.w4(32'hbbac9294),
	.w5(32'hbaca443c),
	.w6(32'hba02efb8),
	.w7(32'hbb8cc855),
	.w8(32'h39d093e7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8467de),
	.w1(32'hbb52f25f),
	.w2(32'h3a273e7e),
	.w3(32'hba8eabd9),
	.w4(32'h3981b534),
	.w5(32'hbb1488e0),
	.w6(32'hbb2f8722),
	.w7(32'hbba88e8b),
	.w8(32'h3b8ec91d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7b1bb),
	.w1(32'hbb2483d1),
	.w2(32'h393e1e85),
	.w3(32'hbb3b0069),
	.w4(32'hbb548a82),
	.w5(32'h3aa84ed9),
	.w6(32'hbb3b5b8f),
	.w7(32'hbb942ef4),
	.w8(32'h3aa09ebf),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad7dd),
	.w1(32'h3ba4c349),
	.w2(32'h3a5d142c),
	.w3(32'h3c0404da),
	.w4(32'h3b02710c),
	.w5(32'h372d744c),
	.w6(32'h3c3d9943),
	.w7(32'h3b39ecdc),
	.w8(32'hba4a79e4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f634d),
	.w1(32'hb9471e55),
	.w2(32'hbb5b3310),
	.w3(32'h3b3c2653),
	.w4(32'h3b04b3b6),
	.w5(32'hbb418b90),
	.w6(32'h3b9a691f),
	.w7(32'hba2f4d22),
	.w8(32'h3bf9e28b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978a370),
	.w1(32'hbb727d92),
	.w2(32'hbbe4db74),
	.w3(32'hbb642a47),
	.w4(32'h3b3844d2),
	.w5(32'h3b110412),
	.w6(32'hbb522c8d),
	.w7(32'hbb8bfe0d),
	.w8(32'h3b184b2b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a425caa),
	.w1(32'h3b58ebcb),
	.w2(32'h3a627e3c),
	.w3(32'hb9be374d),
	.w4(32'h3b9b2e00),
	.w5(32'h3b80d496),
	.w6(32'h3b75e33f),
	.w7(32'h3b39e8c2),
	.w8(32'h38e26e9f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0754b6),
	.w1(32'hbb9ccf0c),
	.w2(32'h39dcb368),
	.w3(32'hbb52209c),
	.w4(32'hb9c2514f),
	.w5(32'h3b9c79ae),
	.w6(32'hbb10ec04),
	.w7(32'hbba00d0d),
	.w8(32'h3ba7a30e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f305e),
	.w1(32'h3a34db91),
	.w2(32'h3b28b772),
	.w3(32'h3b3ddc56),
	.w4(32'h3af64045),
	.w5(32'hbb95826a),
	.w6(32'h3bb4675c),
	.w7(32'h39492072),
	.w8(32'hbbb151c0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d0d16),
	.w1(32'h3995b92c),
	.w2(32'hba13bf75),
	.w3(32'hba52d5f5),
	.w4(32'h3b2e36f4),
	.w5(32'hb9bf3a54),
	.w6(32'hbae880ba),
	.w7(32'h3ae59829),
	.w8(32'hb998cbb3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b1876),
	.w1(32'h3ae0ca89),
	.w2(32'hbab8b0b3),
	.w3(32'h3a8da5d5),
	.w4(32'hbb7fff94),
	.w5(32'h3b1af788),
	.w6(32'h3b79ee12),
	.w7(32'hbac4a909),
	.w8(32'h3b6a8786),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb535a45),
	.w1(32'hba4c54ec),
	.w2(32'h3aa964c4),
	.w3(32'h3b79a33d),
	.w4(32'h3adc946f),
	.w5(32'h3bcfe0c1),
	.w6(32'h3b779b3c),
	.w7(32'h3b41bcad),
	.w8(32'h3b82b2d1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af07bb1),
	.w1(32'hbbb44b5f),
	.w2(32'hbb6fc6b7),
	.w3(32'hba838362),
	.w4(32'hbb80db0e),
	.w5(32'h3ae52328),
	.w6(32'hbaca76d6),
	.w7(32'hbc0aa4df),
	.w8(32'h3a5bacd5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd8a70),
	.w1(32'hba44b547),
	.w2(32'hbb1e5c3c),
	.w3(32'h3ba9735c),
	.w4(32'hba72c31a),
	.w5(32'h3bb5d22a),
	.w6(32'h3b325b02),
	.w7(32'hba7103a2),
	.w8(32'h3bec5af0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87bc25),
	.w1(32'h3b5589f9),
	.w2(32'hba8908e7),
	.w3(32'h3ad36c60),
	.w4(32'h3b558bc0),
	.w5(32'h3ba56e02),
	.w6(32'h3bc46fcd),
	.w7(32'h3b278726),
	.w8(32'h3aadf2e4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74d303),
	.w1(32'hbb870bea),
	.w2(32'hbb63adb6),
	.w3(32'h3b93640e),
	.w4(32'h3b691e6a),
	.w5(32'h3935da45),
	.w6(32'hba27d91c),
	.w7(32'hba9b8655),
	.w8(32'h3b96affa),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b319e19),
	.w1(32'hb90082e9),
	.w2(32'hbac51d9f),
	.w3(32'h3b5f16f3),
	.w4(32'h3b37d40f),
	.w5(32'hbb18ec01),
	.w6(32'h3b0336c1),
	.w7(32'hbaca1219),
	.w8(32'hb9ac0812),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9463c27),
	.w1(32'hbb320d11),
	.w2(32'h3b8aee14),
	.w3(32'hba35845e),
	.w4(32'h3bbccb0c),
	.w5(32'h3a6a5a04),
	.w6(32'hbaac94d8),
	.w7(32'h3bb9b5b0),
	.w8(32'h3a4c2a91),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac228d1),
	.w1(32'h3a2a48aa),
	.w2(32'hbac5d0b9),
	.w3(32'hbb1d919e),
	.w4(32'h3b49ed85),
	.w5(32'h3b457696),
	.w6(32'h38efd568),
	.w7(32'h3b09c771),
	.w8(32'h3b870771),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990697c),
	.w1(32'hbbc551ad),
	.w2(32'hbb2ced5a),
	.w3(32'hbb22cb13),
	.w4(32'h3aa6ac43),
	.w5(32'hbab7b073),
	.w6(32'hbbd4fa9c),
	.w7(32'hbaa1f673),
	.w8(32'hbb7c8749),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a7806),
	.w1(32'h3a9bc762),
	.w2(32'h3ae492ed),
	.w3(32'h391f06b0),
	.w4(32'h3ab6c13a),
	.w5(32'h3b569ca0),
	.w6(32'h3bda3eca),
	.w7(32'h3bccf645),
	.w8(32'h3b0061ed),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ff8b4),
	.w1(32'hb9bf9b41),
	.w2(32'hb9884ce3),
	.w3(32'h3b362189),
	.w4(32'h3ac80444),
	.w5(32'hba25fd4c),
	.w6(32'h3b76204a),
	.w7(32'hba0b9a03),
	.w8(32'hba4e2683),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac07961),
	.w1(32'h3a6cca1a),
	.w2(32'h3b4c7e85),
	.w3(32'h3b4100fe),
	.w4(32'h37a7e4ee),
	.w5(32'hba7105ba),
	.w6(32'h3b78b969),
	.w7(32'hba8b22f2),
	.w8(32'hba85b887),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48ce1d),
	.w1(32'hba953b5b),
	.w2(32'hbb397b96),
	.w3(32'h3a7f9131),
	.w4(32'hbb09c02b),
	.w5(32'hba95e9ea),
	.w6(32'h3b8cad8b),
	.w7(32'hba621024),
	.w8(32'hb8c43cad),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b380fc2),
	.w1(32'h3a2ae737),
	.w2(32'hb9a85f7f),
	.w3(32'h3ac36968),
	.w4(32'h3adda43c),
	.w5(32'hba012ecc),
	.w6(32'h3a40def0),
	.w7(32'hba71ce19),
	.w8(32'hbb13277f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e8d86),
	.w1(32'h3a2ee50e),
	.w2(32'h392a78da),
	.w3(32'hbb17aec1),
	.w4(32'h3ba5a7ff),
	.w5(32'hbb37769f),
	.w6(32'hbb9000f4),
	.w7(32'hbbf3d385),
	.w8(32'h3b0e8f13),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02a010),
	.w1(32'h3b87a09a),
	.w2(32'h3be5c81e),
	.w3(32'hbb0c6969),
	.w4(32'h3bb563af),
	.w5(32'hb88228af),
	.w6(32'h3b0370d6),
	.w7(32'h3b4903f8),
	.w8(32'h3ac7d0b7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8b3ba),
	.w1(32'hbb48d842),
	.w2(32'hbb813f31),
	.w3(32'h3b05a1c5),
	.w4(32'h3b3395fb),
	.w5(32'h3b4abc2f),
	.w6(32'hbb9057b1),
	.w7(32'hbb228d92),
	.w8(32'h3b88f266),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87395e),
	.w1(32'h3b15fcf8),
	.w2(32'h3b4d7349),
	.w3(32'h3aadccea),
	.w4(32'h3b0789f4),
	.w5(32'hbbca1ed7),
	.w6(32'h3b242cb2),
	.w7(32'h3b7dd2b0),
	.w8(32'hbbe44177),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4984bf),
	.w1(32'h38a89607),
	.w2(32'h3afa4f05),
	.w3(32'h3c821aa1),
	.w4(32'hbb9b1089),
	.w5(32'hbb13b08a),
	.w6(32'h3cb31441),
	.w7(32'h39d31532),
	.w8(32'h3ac0ad83),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb574d5),
	.w1(32'hbb3ee40e),
	.w2(32'hbb87a6e1),
	.w3(32'h3bf8232f),
	.w4(32'h3ba030f4),
	.w5(32'hbbda625d),
	.w6(32'hb9645f63),
	.w7(32'h3b4883ca),
	.w8(32'hbc240554),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13db36),
	.w1(32'hba9f97f9),
	.w2(32'h3a83828d),
	.w3(32'h3b3ad628),
	.w4(32'hba9fb4c8),
	.w5(32'hbaa2098d),
	.w6(32'h3bacf160),
	.w7(32'hbb2810e7),
	.w8(32'hbb64909a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba473f8),
	.w1(32'hba682a10),
	.w2(32'h3ba4802c),
	.w3(32'h3bc19e28),
	.w4(32'h3b501d6e),
	.w5(32'h3abdef81),
	.w6(32'h3bf01b9f),
	.w7(32'h3bbb6744),
	.w8(32'h3b599dc1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9cf42),
	.w1(32'h3b2ed3b3),
	.w2(32'h3be52732),
	.w3(32'hbb996a1a),
	.w4(32'h3bc515d1),
	.w5(32'h3b1fb48d),
	.w6(32'hbb48ab1b),
	.w7(32'h3bd04439),
	.w8(32'h3b8ad46d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14a83d),
	.w1(32'h3bae0f80),
	.w2(32'hbacff85e),
	.w3(32'h3c55d9c4),
	.w4(32'hbbc3e014),
	.w5(32'h3a333d61),
	.w6(32'h3c9a8c89),
	.w7(32'hbb6a9054),
	.w8(32'h3a4cea04),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25fb7d),
	.w1(32'h3bbd346d),
	.w2(32'h3aa8e61d),
	.w3(32'h3b06678e),
	.w4(32'h3b9c3546),
	.w5(32'h3a5d60d6),
	.w6(32'h3bb04290),
	.w7(32'hbb545f9b),
	.w8(32'h3a96b9b2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b590564),
	.w1(32'h3a4b9651),
	.w2(32'hba171f2a),
	.w3(32'h3a679af5),
	.w4(32'h3ae64395),
	.w5(32'h3b85ad3b),
	.w6(32'hbba97612),
	.w7(32'h3919fe1d),
	.w8(32'h3b4108d2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d0ffa),
	.w1(32'hba9d62b8),
	.w2(32'h3bd44694),
	.w3(32'h3b21c561),
	.w4(32'hbbb71c13),
	.w5(32'hbac7f6e8),
	.w6(32'h3b611b70),
	.w7(32'h3a4ddfc9),
	.w8(32'hbac5bc09),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefbe68),
	.w1(32'hba810c7a),
	.w2(32'hbb7599d3),
	.w3(32'h38fe57f6),
	.w4(32'hbb793b57),
	.w5(32'h3b853138),
	.w6(32'h390eba12),
	.w7(32'hbb48ae77),
	.w8(32'h3b3f6241),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48f5f4),
	.w1(32'hbb9b226d),
	.w2(32'hbb85f0fa),
	.w3(32'hba4aaf40),
	.w4(32'hbad28aef),
	.w5(32'hba7887da),
	.w6(32'hbb238625),
	.w7(32'hbbaeecde),
	.w8(32'h398dce39),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd1fdb),
	.w1(32'hb9076156),
	.w2(32'hbb1252af),
	.w3(32'h3a3a26f5),
	.w4(32'hbb000b72),
	.w5(32'h3aa6aa92),
	.w6(32'h3b6b0731),
	.w7(32'h39047041),
	.w8(32'h3b0d2b0d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc6d84),
	.w1(32'hbb1909fe),
	.w2(32'hbb219708),
	.w3(32'h3b509160),
	.w4(32'h3af529d4),
	.w5(32'hbb4b0569),
	.w6(32'hbadf2f9f),
	.w7(32'hbb94de7c),
	.w8(32'hbba06b14),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e57dc),
	.w1(32'h3b58534f),
	.w2(32'hbaa741ef),
	.w3(32'h3b3d16b1),
	.w4(32'hba8f1455),
	.w5(32'hbb19f7e5),
	.w6(32'h3b234f15),
	.w7(32'hbb059666),
	.w8(32'hba4f1746),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2088a9),
	.w1(32'h3a0c1402),
	.w2(32'hbaf737fe),
	.w3(32'hbb5ae7ab),
	.w4(32'hbb9c5329),
	.w5(32'hbb7fe582),
	.w6(32'h3b551d56),
	.w7(32'hbb0a6f91),
	.w8(32'hbb8620cf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bd74f),
	.w1(32'hbab3f440),
	.w2(32'hbafab964),
	.w3(32'h3b8637ac),
	.w4(32'h3ab4133d),
	.w5(32'h3afd6674),
	.w6(32'h3a9eddab),
	.w7(32'hbae0480b),
	.w8(32'h3b08eb71),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee7add),
	.w1(32'hba37a597),
	.w2(32'hb9bdb0a0),
	.w3(32'h3a6fd89b),
	.w4(32'h3a9e49d3),
	.w5(32'hba0da02c),
	.w6(32'h39bc17a0),
	.w7(32'h3a1d8f95),
	.w8(32'h3ad8e6bd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb886a5),
	.w1(32'h3bc1fc44),
	.w2(32'h3aa56c42),
	.w3(32'h3ae454fe),
	.w4(32'h3ac3762a),
	.w5(32'hbac82c31),
	.w6(32'h3bd928d3),
	.w7(32'h3b6e8aed),
	.w8(32'hb84efc46),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba146033),
	.w1(32'hbb45aeed),
	.w2(32'hbb6cc3f5),
	.w3(32'hbb347122),
	.w4(32'hbb714f96),
	.w5(32'hbb3cc6ee),
	.w6(32'hba9bd454),
	.w7(32'hbb5f4123),
	.w8(32'hbb69f9f3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60290e),
	.w1(32'hb99251ae),
	.w2(32'hbc5776ad),
	.w3(32'h37d5deee),
	.w4(32'hbc649b01),
	.w5(32'hbba667d0),
	.w6(32'hba00df44),
	.w7(32'hbc5d3972),
	.w8(32'hbb859ea1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4441),
	.w1(32'h3a901440),
	.w2(32'h3b4aa1fd),
	.w3(32'h3b118e9b),
	.w4(32'h3b169f7f),
	.w5(32'h3b2d4ab8),
	.w6(32'h3ac59022),
	.w7(32'h3b4fda5b),
	.w8(32'h3af3f9a7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace4e6f),
	.w1(32'hb9c6ff86),
	.w2(32'h3a19a348),
	.w3(32'h3b4025f9),
	.w4(32'h39dec9f0),
	.w5(32'h3b01903a),
	.w6(32'h3a71dd88),
	.w7(32'h38bc0e83),
	.w8(32'h3ae53f46),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d7fbe2),
	.w1(32'hbbe268ed),
	.w2(32'hbb621de2),
	.w3(32'hbb5fc0d6),
	.w4(32'hba2a149c),
	.w5(32'hbb583a6c),
	.w6(32'hbb3cef52),
	.w7(32'hbb4bef58),
	.w8(32'hbb8d11f9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb2bf),
	.w1(32'h3bc19c16),
	.w2(32'h3bfef021),
	.w3(32'h3b8cd316),
	.w4(32'h3bcc3b79),
	.w5(32'h3a60c552),
	.w6(32'h3b907fbc),
	.w7(32'h3c014332),
	.w8(32'hbaea21f7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03973b),
	.w1(32'h3aa11a2e),
	.w2(32'h3aa99189),
	.w3(32'h3b1fecc0),
	.w4(32'h3a7455ba),
	.w5(32'h3b5a0a22),
	.w6(32'hb8c18ab4),
	.w7(32'hba425123),
	.w8(32'h3babe708),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babd4a5),
	.w1(32'h3b015883),
	.w2(32'hbac3fd8c),
	.w3(32'hba1d62c4),
	.w4(32'hba9b70c7),
	.w5(32'h3ae8b0a0),
	.w6(32'h3b001e26),
	.w7(32'hbab9b74d),
	.w8(32'h3b9b9b1b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ca27f),
	.w1(32'hbb86e17c),
	.w2(32'hbb4566ea),
	.w3(32'hba1352e0),
	.w4(32'hba2cec88),
	.w5(32'h3bcfc2cd),
	.w6(32'h3a790f0b),
	.w7(32'hbb56f620),
	.w8(32'h3b7d07cf),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad010c),
	.w1(32'h3b87a834),
	.w2(32'h3c0a1e70),
	.w3(32'h3b9ea31b),
	.w4(32'h3c074a50),
	.w5(32'h3b4fefcb),
	.w6(32'h3b1b1c5c),
	.w7(32'h3bea997d),
	.w8(32'hba9579fa),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40ffd3),
	.w1(32'h3909ffcf),
	.w2(32'h3877525e),
	.w3(32'h3b3ecd51),
	.w4(32'h3afc0bbb),
	.w5(32'hbb3455cf),
	.w6(32'hbacca2d1),
	.w7(32'hbaa16df9),
	.w8(32'hbb83076e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ffa4f),
	.w1(32'hbbb3d871),
	.w2(32'hbaa12434),
	.w3(32'hbb0e4eb7),
	.w4(32'hb988fb9d),
	.w5(32'h3b8345eb),
	.w6(32'hbbb1be00),
	.w7(32'hbab27e4c),
	.w8(32'h3c0b497c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf0cbc),
	.w1(32'h3c04052f),
	.w2(32'h3b125d7b),
	.w3(32'h3b9c0ebb),
	.w4(32'hbb4553b7),
	.w5(32'h3bd9bf56),
	.w6(32'h3c1d087e),
	.w7(32'h3ac971f4),
	.w8(32'h3bd96d70),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b665fab),
	.w1(32'hbb289ea1),
	.w2(32'hbacf85a0),
	.w3(32'hba873136),
	.w4(32'h3b1c28e2),
	.w5(32'hbb77a53a),
	.w6(32'h3b1212ff),
	.w7(32'h3b3d6e7d),
	.w8(32'hbb2479bf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ebcad),
	.w1(32'h3814a8c6),
	.w2(32'hb74e0453),
	.w3(32'hbb46234a),
	.w4(32'h39c56d7a),
	.w5(32'hbb73b7e1),
	.w6(32'hbac0ad7f),
	.w7(32'hba8ed540),
	.w8(32'hbab38f3d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0f843),
	.w1(32'hbb0f09f1),
	.w2(32'hbae8b818),
	.w3(32'hbae20ab8),
	.w4(32'h39910b4a),
	.w5(32'hb80f4f0c),
	.w6(32'hba80ff4f),
	.w7(32'hba04f61b),
	.w8(32'hba8b6871),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc2115),
	.w1(32'h3ab52316),
	.w2(32'h3998b437),
	.w3(32'h3b0a1b1e),
	.w4(32'hbb3baed3),
	.w5(32'hbbde1712),
	.w6(32'hba432662),
	.w7(32'hba415e0d),
	.w8(32'hbb7c8a37),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67eaa3),
	.w1(32'hbaf24e06),
	.w2(32'hba2c0fbc),
	.w3(32'hbbc0e4c8),
	.w4(32'hbb1ba939),
	.w5(32'h3b423f13),
	.w6(32'hbb3d4c0a),
	.w7(32'hb9f933ee),
	.w8(32'h3b202e79),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b990de9),
	.w1(32'h3b71095c),
	.w2(32'h3b3f55e1),
	.w3(32'h3b260da8),
	.w4(32'h3bad37d5),
	.w5(32'h3b0e5211),
	.w6(32'h38ad0665),
	.w7(32'h3a4edf3f),
	.w8(32'h3b66269e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed3f5),
	.w1(32'h3b80d551),
	.w2(32'h3ade416c),
	.w3(32'h3b9dfe53),
	.w4(32'h3a5362d4),
	.w5(32'hb6f43760),
	.w6(32'h3ba53772),
	.w7(32'h3b045148),
	.w8(32'h3996f28b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfc5a2),
	.w1(32'hbb29c980),
	.w2(32'hb9b0e184),
	.w3(32'hba883a68),
	.w4(32'hba9fe826),
	.w5(32'hbc838eb3),
	.w6(32'hbb1d647e),
	.w7(32'hba29a131),
	.w8(32'hbc758aae),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc878283),
	.w1(32'h3b25aa84),
	.w2(32'hbb35b0f6),
	.w3(32'h3a9cab06),
	.w4(32'hbba148c8),
	.w5(32'h3b854f2c),
	.w6(32'h3b1ec4f8),
	.w7(32'hbb677cfa),
	.w8(32'h3b6b67a1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad6011),
	.w1(32'h3b69fe3a),
	.w2(32'h3b332993),
	.w3(32'h3b5bc18c),
	.w4(32'h3ab679a5),
	.w5(32'hbb2fedd5),
	.w6(32'h3b732242),
	.w7(32'h3b6ffa60),
	.w8(32'h3ab309c5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925dddb),
	.w1(32'hbb5e9346),
	.w2(32'hbb6a0c67),
	.w3(32'hbba57d15),
	.w4(32'hbb3a4998),
	.w5(32'h3c2ea7f0),
	.w6(32'hb99fa50a),
	.w7(32'hba88b7f0),
	.w8(32'h3c34f901),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c298827),
	.w1(32'h3bf32aee),
	.w2(32'h3b9f23b8),
	.w3(32'h3c11d1c6),
	.w4(32'h3bc9a996),
	.w5(32'hbbe52cc8),
	.w6(32'h3c0d0dea),
	.w7(32'h3bb476bd),
	.w8(32'h3a5923bc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb579d20),
	.w1(32'hbb4c4be7),
	.w2(32'hbb901677),
	.w3(32'hbb3c9ee9),
	.w4(32'hbbd3d496),
	.w5(32'h3bad71fa),
	.w6(32'hbb18be64),
	.w7(32'hbb01a8d4),
	.w8(32'h3bc22914),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98125b),
	.w1(32'h3bc3ea0e),
	.w2(32'h3ba9b63c),
	.w3(32'h3bd3cdff),
	.w4(32'h3bc0363b),
	.w5(32'h3b8b7b1a),
	.w6(32'h3bf16f3f),
	.w7(32'h3bd40b28),
	.w8(32'h3b9e9446),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b541caa),
	.w1(32'h3bc2a83d),
	.w2(32'h3bc88c38),
	.w3(32'h3b909df5),
	.w4(32'h3ba1dcdd),
	.w5(32'hbb4d339d),
	.w6(32'h3bb48927),
	.w7(32'h3bbd94f2),
	.w8(32'hbb1ab465),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e9449),
	.w1(32'hb9a2a65d),
	.w2(32'h3af285f7),
	.w3(32'h3aa72506),
	.w4(32'h3b97b21d),
	.w5(32'h3a420446),
	.w6(32'h3b03b633),
	.w7(32'h3b8345d7),
	.w8(32'h3a83fb17),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d9459),
	.w1(32'h3ba6363e),
	.w2(32'h3bb7a18f),
	.w3(32'h3b90f7cd),
	.w4(32'h3ba1ee77),
	.w5(32'h3bb19f0a),
	.w6(32'h3b8daa62),
	.w7(32'h3b9fb210),
	.w8(32'h3bbedee0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e040b),
	.w1(32'h3b5d7599),
	.w2(32'h3b82ec60),
	.w3(32'h3bca9d92),
	.w4(32'h3b9bf67f),
	.w5(32'h3bc999fc),
	.w6(32'h3ba9f9b6),
	.w7(32'h3baf1d00),
	.w8(32'h3c044b0a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8c698),
	.w1(32'h3b6681b0),
	.w2(32'h3b2a6410),
	.w3(32'h3b69f8d4),
	.w4(32'h3b935b66),
	.w5(32'hbb0a28f6),
	.w6(32'h3bcfe841),
	.w7(32'h3bad7ac2),
	.w8(32'hbae0bfe4),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a585a0e),
	.w1(32'h3b3791d2),
	.w2(32'hbafbb431),
	.w3(32'hbaa22592),
	.w4(32'h3a5da9ed),
	.w5(32'h3b7a9826),
	.w6(32'h3b625d69),
	.w7(32'h3b2b00c5),
	.w8(32'h3bdbcd7b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7c097),
	.w1(32'h3bf8e66e),
	.w2(32'h3be0a26a),
	.w3(32'h3bb0419b),
	.w4(32'h3b505791),
	.w5(32'hbb9a5a04),
	.w6(32'h3c098f08),
	.w7(32'h3c0bc34c),
	.w8(32'hbb20576b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb623bd0),
	.w1(32'hbb35542b),
	.w2(32'hbad08685),
	.w3(32'hbb6fbbc0),
	.w4(32'h3a911000),
	.w5(32'h3c18af6e),
	.w6(32'hbb1c6592),
	.w7(32'hba2df534),
	.w8(32'h3c1b6bcd),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9f012),
	.w1(32'h3b9fdfe8),
	.w2(32'h3ba0a2fe),
	.w3(32'h3be7c8de),
	.w4(32'h3b98d1f3),
	.w5(32'hbb47cbe5),
	.w6(32'h3bc3600a),
	.w7(32'h3b87a894),
	.w8(32'hbb371cd1),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac504b),
	.w1(32'hbba2a43e),
	.w2(32'hbb9f83c9),
	.w3(32'hbb6d893f),
	.w4(32'hbb609e0b),
	.w5(32'hbb58468f),
	.w6(32'hbb9b3fac),
	.w7(32'hbb8e0ff5),
	.w8(32'hbacd8af4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacad3e2),
	.w1(32'h3b04cce7),
	.w2(32'hba6f85d6),
	.w3(32'hb8be429e),
	.w4(32'hbb2c4742),
	.w5(32'h3a0f6b4b),
	.w6(32'h3b19cd00),
	.w7(32'hba1f61b4),
	.w8(32'h3b1b5bc0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b159209),
	.w1(32'hb89070cc),
	.w2(32'hbaa6ae44),
	.w3(32'hba84fd58),
	.w4(32'hba30a940),
	.w5(32'h3bb1dc68),
	.w6(32'h38103146),
	.w7(32'hb9819859),
	.w8(32'h3b7056bf),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ca04d),
	.w1(32'h3ac0422a),
	.w2(32'h3acfd2aa),
	.w3(32'h3b9a21c2),
	.w4(32'h3b5e96cb),
	.w5(32'hbaa63d24),
	.w6(32'h3b0da4a3),
	.w7(32'h3a72d8d4),
	.w8(32'hbacbcb6d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84750f),
	.w1(32'hbb8e152c),
	.w2(32'hbb2c17f6),
	.w3(32'hbbb47a78),
	.w4(32'hbb3467a0),
	.w5(32'h3a2ba9bc),
	.w6(32'hbbaeebd4),
	.w7(32'hbb93659f),
	.w8(32'hba666667),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a1e43),
	.w1(32'hbb9d36e8),
	.w2(32'hbb016540),
	.w3(32'hba93ca27),
	.w4(32'hba4ae5b5),
	.w5(32'h3b1b31a3),
	.w6(32'hbb42fdba),
	.w7(32'hbb207229),
	.w8(32'h39fbf9fa),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ef01a),
	.w1(32'h3b2c1e86),
	.w2(32'h3bb475cf),
	.w3(32'h3af416ec),
	.w4(32'h3b94086f),
	.w5(32'hba59117b),
	.w6(32'h39e7d152),
	.w7(32'h3b6415cf),
	.w8(32'hbb8fb50c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88c2e5),
	.w1(32'h3ade55f0),
	.w2(32'hba1d52d6),
	.w3(32'h38dd48a0),
	.w4(32'hbaaeffef),
	.w5(32'h3a2b48f6),
	.w6(32'hb8d16e6a),
	.w7(32'hba910cfb),
	.w8(32'h3b63bfcb),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00d513),
	.w1(32'hbb038a84),
	.w2(32'hbb09fc2c),
	.w3(32'hbab497ac),
	.w4(32'hbb63ee8a),
	.w5(32'hbb01af13),
	.w6(32'hbb08f3f9),
	.w7(32'hb96721e6),
	.w8(32'hb9db9054),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17e75e),
	.w1(32'hba68f465),
	.w2(32'hbb5e46cf),
	.w3(32'hba52e9e8),
	.w4(32'hbb0ab3ac),
	.w5(32'h3adc2ce0),
	.w6(32'hbafd3871),
	.w7(32'hbb6dae30),
	.w8(32'h3b40eb55),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b54ee),
	.w1(32'hbac16034),
	.w2(32'hbb0c28c5),
	.w3(32'h3b118f9b),
	.w4(32'hbae73e5c),
	.w5(32'hbb9c6ccc),
	.w6(32'h3adc563c),
	.w7(32'hbb2261f3),
	.w8(32'hbbbe550c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6293bc),
	.w1(32'h3b011644),
	.w2(32'hbc1a3485),
	.w3(32'h3a369f51),
	.w4(32'hbc1ceca5),
	.w5(32'hbc31794c),
	.w6(32'hba8888a9),
	.w7(32'hbc3a7421),
	.w8(32'hbc075231),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d4155),
	.w1(32'h3b38a3ba),
	.w2(32'h3b2a2a8a),
	.w3(32'h3b2ef43d),
	.w4(32'h3a9a68f5),
	.w5(32'h3b2f1f91),
	.w6(32'h3b47b0aa),
	.w7(32'h3b1c144b),
	.w8(32'h3b54fe96),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb42984),
	.w1(32'h3acf22a9),
	.w2(32'h3acf20f9),
	.w3(32'hbafb8d03),
	.w4(32'h3a062e4a),
	.w5(32'hbbb46903),
	.w6(32'hbb083e1e),
	.w7(32'hbae0cc4a),
	.w8(32'hbb9af233),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cf80f),
	.w1(32'hbad73ebf),
	.w2(32'hbaedb34d),
	.w3(32'hbad26d57),
	.w4(32'hbb631ffc),
	.w5(32'h3c06f6bd),
	.w6(32'hbacbfdd5),
	.w7(32'hbb4f8bf5),
	.w8(32'h3b4b934e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba298b69),
	.w1(32'hba849a22),
	.w2(32'hba173661),
	.w3(32'h3c0cf0c1),
	.w4(32'h3baebe61),
	.w5(32'hbaa70fbb),
	.w6(32'h3a0217e5),
	.w7(32'hbb81d5c6),
	.w8(32'hb9f93145),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842052e),
	.w1(32'hbb27a910),
	.w2(32'h3a206db3),
	.w3(32'hbb88e290),
	.w4(32'hbb2139df),
	.w5(32'h3a843312),
	.w6(32'hbb057f07),
	.w7(32'h3a9316a9),
	.w8(32'hb9a0af21),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1fa9c),
	.w1(32'hbbaed7a1),
	.w2(32'hb9b327c6),
	.w3(32'hba72813d),
	.w4(32'hbad6f202),
	.w5(32'hba04d1c1),
	.w6(32'hbb9857c2),
	.w7(32'hbbae0036),
	.w8(32'h3a9cf7be),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02144b),
	.w1(32'hbaa4b720),
	.w2(32'hbb1b8f78),
	.w3(32'hbaeaa229),
	.w4(32'hba7af357),
	.w5(32'hbb7b572b),
	.w6(32'hbb0970a7),
	.w7(32'hba889059),
	.w8(32'hbb5df372),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb403dd8),
	.w1(32'hbaf64746),
	.w2(32'hbb243acc),
	.w3(32'h39e8e66f),
	.w4(32'hba1ffdaf),
	.w5(32'h3bd4541b),
	.w6(32'hbafe218a),
	.w7(32'hba7ce9e4),
	.w8(32'h3b8fd004),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b124860),
	.w1(32'hbb57f9c3),
	.w2(32'hbaf251aa),
	.w3(32'h3ae6ebca),
	.w4(32'h3a2338f8),
	.w5(32'hbb2f74ba),
	.w6(32'hbb189f30),
	.w7(32'hbb134892),
	.w8(32'hbaaa6443),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fee96),
	.w1(32'hba9f137e),
	.w2(32'hba9ee238),
	.w3(32'h3a37f7cd),
	.w4(32'h3a5f36f9),
	.w5(32'hbb285d34),
	.w6(32'hbad8cb87),
	.w7(32'hbaec3c2a),
	.w8(32'hbb64024d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25bc5a),
	.w1(32'h39dce7de),
	.w2(32'hbaad873f),
	.w3(32'h3854e5e8),
	.w4(32'hba508fe3),
	.w5(32'hba678cd6),
	.w6(32'hba0623b8),
	.w7(32'hba1250e5),
	.w8(32'hbb8f11b3),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c988c),
	.w1(32'hbb424862),
	.w2(32'hbad55c8d),
	.w3(32'hba8e55ef),
	.w4(32'hbb0a7fd9),
	.w5(32'hb83ab32c),
	.w6(32'hbbc54d21),
	.w7(32'hbad284c8),
	.w8(32'h399bcb25),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b45da2),
	.w1(32'h3b929522),
	.w2(32'h3a4e2709),
	.w3(32'h3ae439d3),
	.w4(32'h3aab06fe),
	.w5(32'hba297e97),
	.w6(32'h3bbc8962),
	.w7(32'h3aaf4108),
	.w8(32'hbab3bf9e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b58a6),
	.w1(32'h3afd8791),
	.w2(32'hbb1b89d2),
	.w3(32'hb82ad3e5),
	.w4(32'hba28bcea),
	.w5(32'h3a94909d),
	.w6(32'h3a73d032),
	.w7(32'hbb1618ec),
	.w8(32'h3aee1c98),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977ada3),
	.w1(32'h396e4d1b),
	.w2(32'hbb067468),
	.w3(32'h3aaeb262),
	.w4(32'hbae31a5a),
	.w5(32'hba5e68ff),
	.w6(32'h3b526c08),
	.w7(32'h38600222),
	.w8(32'hbb4b49c4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d3841),
	.w1(32'hbb23fe62),
	.w2(32'hbb4fe12e),
	.w3(32'hb9303a35),
	.w4(32'hba4cdabb),
	.w5(32'h3c12746d),
	.w6(32'hbb4d31e7),
	.w7(32'hbb24183f),
	.w8(32'h3c10eb39),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb66ce3),
	.w1(32'h3bd13351),
	.w2(32'hbb317e92),
	.w3(32'h3c3882a1),
	.w4(32'h3b3f22e5),
	.w5(32'h3aa9bf8b),
	.w6(32'h3c1bba08),
	.w7(32'hba1ad1c5),
	.w8(32'h3b4e9cf9),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10bfee),
	.w1(32'h3b1cfa89),
	.w2(32'h39b38aa4),
	.w3(32'h3a5cf31f),
	.w4(32'hbb24d79d),
	.w5(32'hbbd1f5b3),
	.w6(32'h3bb16004),
	.w7(32'h3a195f41),
	.w8(32'hbbb37580),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb902682),
	.w1(32'hbb9bbde2),
	.w2(32'hbb3f0e6c),
	.w3(32'hbbaaff1c),
	.w4(32'hbb780543),
	.w5(32'h3a053d66),
	.w6(32'hbba6ea7d),
	.w7(32'hbb8cf697),
	.w8(32'h3aed71b4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7f66a),
	.w1(32'hbb0e7a7e),
	.w2(32'hbb9bc68d),
	.w3(32'hbb365efa),
	.w4(32'hbb8b1a19),
	.w5(32'h3bae8467),
	.w6(32'hb9bd2ee8),
	.w7(32'hbb91b145),
	.w8(32'h3b869acc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80b941),
	.w1(32'h3c194b07),
	.w2(32'h3c411684),
	.w3(32'h3c06e205),
	.w4(32'h3c221b2b),
	.w5(32'h3b9a5e42),
	.w6(32'h3be9cb72),
	.w7(32'h3c3de0c0),
	.w8(32'h3bc275f6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d0725),
	.w1(32'h3b8d565b),
	.w2(32'h3b80d485),
	.w3(32'h3bbd6d0c),
	.w4(32'h3b806637),
	.w5(32'hbb1a743d),
	.w6(32'h3bd7aa6a),
	.w7(32'h3bdc023d),
	.w8(32'hbb045eae),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e831e),
	.w1(32'h3ace67ab),
	.w2(32'h3a6f3f41),
	.w3(32'h3a65e2e4),
	.w4(32'h39d4dc57),
	.w5(32'hbbc10e9b),
	.w6(32'h3a1c04bf),
	.w7(32'h3a4012c8),
	.w8(32'hbb1044c1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d9fee),
	.w1(32'h3b956f3d),
	.w2(32'hbbaca648),
	.w3(32'h3b15a58a),
	.w4(32'hbaaea3e0),
	.w5(32'h3ba3ac16),
	.w6(32'h3c18d691),
	.w7(32'hbb63c5b8),
	.w8(32'h3b2199fb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b427845),
	.w1(32'h3b4ab450),
	.w2(32'h3b00d2ed),
	.w3(32'h3b515bbb),
	.w4(32'h3b10fcc5),
	.w5(32'h3bae47a0),
	.w6(32'h3b63153f),
	.w7(32'h3b36ecea),
	.w8(32'h3b616586),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b213bca),
	.w1(32'hba00538b),
	.w2(32'hba9c3f34),
	.w3(32'hba927941),
	.w4(32'h3b8e51c5),
	.w5(32'hbb08161e),
	.w6(32'h3b65f46b),
	.w7(32'h3b252091),
	.w8(32'hbb412269),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66b664),
	.w1(32'h3adcbb55),
	.w2(32'hba82c1d4),
	.w3(32'h3acdde96),
	.w4(32'h3a6fa2ea),
	.w5(32'h3b33d71e),
	.w6(32'h3a5e97cd),
	.w7(32'hbab2c9c4),
	.w8(32'h3a925a78),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ac4c8),
	.w1(32'hbaec8edd),
	.w2(32'hb84df8dc),
	.w3(32'hba003402),
	.w4(32'hba3fefa5),
	.w5(32'hbb81e95c),
	.w6(32'h3905e153),
	.w7(32'hba3d6424),
	.w8(32'hba1db8e2),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5abe79),
	.w1(32'h3b19130c),
	.w2(32'hba29975c),
	.w3(32'h39c96e26),
	.w4(32'hbb6b7b78),
	.w5(32'h3a180259),
	.w6(32'h3ad43027),
	.w7(32'hba1f4ffe),
	.w8(32'hb926533f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78426f),
	.w1(32'h3b0002ad),
	.w2(32'h3b12170c),
	.w3(32'h3b464dcd),
	.w4(32'h3afe0590),
	.w5(32'hbab12b05),
	.w6(32'h3a87abd6),
	.w7(32'h3adacbcf),
	.w8(32'hbb029a92),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03538f),
	.w1(32'hbb86f730),
	.w2(32'h3a9de964),
	.w3(32'hbb41b570),
	.w4(32'h3b9118cf),
	.w5(32'hbb2da0ad),
	.w6(32'hbb142fdb),
	.w7(32'h3b0010d9),
	.w8(32'hbad51df2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf6762),
	.w1(32'h3ace337b),
	.w2(32'h38913bf3),
	.w3(32'h3a76c47b),
	.w4(32'hb98e87fb),
	.w5(32'h3b04199b),
	.w6(32'h3a2b46f1),
	.w7(32'h398ff6da),
	.w8(32'h3b697fce),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94e449),
	.w1(32'h3bcdd594),
	.w2(32'h3c32f655),
	.w3(32'h3ba7c747),
	.w4(32'h3c3da3fe),
	.w5(32'hbb2db0d0),
	.w6(32'h3bf55963),
	.w7(32'h3c5fabab),
	.w8(32'hbb901eaa),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadf861),
	.w1(32'hbb45292d),
	.w2(32'hbaa77bdc),
	.w3(32'hba262ee2),
	.w4(32'hbaa56497),
	.w5(32'h3b14bef9),
	.w6(32'hbb89a107),
	.w7(32'hbb2faac1),
	.w8(32'h3b29d7e6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42105e),
	.w1(32'h3ada6c6c),
	.w2(32'hb98e896e),
	.w3(32'h3ba63fa3),
	.w4(32'hb998ff7e),
	.w5(32'hbad89f3a),
	.w6(32'h3bae75d6),
	.w7(32'h3a23c4e8),
	.w8(32'h3a6ad2aa),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8252788),
	.w1(32'hbb113efa),
	.w2(32'hbac8b1d1),
	.w3(32'h39ad61d5),
	.w4(32'hba6beb6d),
	.w5(32'hba0838ff),
	.w6(32'hb94e3314),
	.w7(32'h3a5bc0d0),
	.w8(32'h3a79a7ea),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a271552),
	.w1(32'h3bbb24ee),
	.w2(32'hba662f8a),
	.w3(32'h3b974fed),
	.w4(32'hbaa845d6),
	.w5(32'h3a655949),
	.w6(32'h3b998811),
	.w7(32'hba2f71a2),
	.w8(32'hbabb043a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71e2be),
	.w1(32'h3a9e68ac),
	.w2(32'h3ab22886),
	.w3(32'h3ba27b35),
	.w4(32'h3b0a986e),
	.w5(32'h39e161b5),
	.w6(32'h3b885f89),
	.w7(32'h3b99e632),
	.w8(32'hba5006bf),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a0a71),
	.w1(32'hba36ef66),
	.w2(32'hbaa4861e),
	.w3(32'hba700b01),
	.w4(32'h39965edd),
	.w5(32'hba1a1418),
	.w6(32'h3a9d9042),
	.w7(32'hb6aebaf3),
	.w8(32'hb936819e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac96f40),
	.w1(32'h3afa181e),
	.w2(32'h3aaaf952),
	.w3(32'h3b42650c),
	.w4(32'h3be2f5b1),
	.w5(32'h3cc564f2),
	.w6(32'h3b9242fc),
	.w7(32'h3b83b4d2),
	.w8(32'h3cd18aa1),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3d245),
	.w1(32'h3cd5f153),
	.w2(32'h3c93ca30),
	.w3(32'h3cd2caae),
	.w4(32'h3c63e721),
	.w5(32'hba60fae3),
	.w6(32'h3ccb28af),
	.w7(32'h3c75ddc4),
	.w8(32'h3aa5ad6d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5dafe),
	.w1(32'h3ad25a3d),
	.w2(32'hbb493744),
	.w3(32'h3b9257ee),
	.w4(32'hbb73a644),
	.w5(32'h3bdb39db),
	.w6(32'h3bb24c44),
	.w7(32'hbb83b968),
	.w8(32'h3b4d4468),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5af20d),
	.w1(32'h3b456ec8),
	.w2(32'h3a39a05c),
	.w3(32'h3c1f779a),
	.w4(32'h3b9e5175),
	.w5(32'h3aefb85d),
	.w6(32'h3b34f494),
	.w7(32'h3ab32c39),
	.w8(32'h3a549c44),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f76ca),
	.w1(32'h3a9a96d8),
	.w2(32'h393bdfd7),
	.w3(32'h3b460622),
	.w4(32'h3ab792e6),
	.w5(32'hba720c6a),
	.w6(32'h3aaec6ee),
	.w7(32'hba16093a),
	.w8(32'hb8208501),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb206192),
	.w1(32'hbaff94df),
	.w2(32'hbb3aa25d),
	.w3(32'hbad15b3c),
	.w4(32'hbb3b159f),
	.w5(32'hbafaedd8),
	.w6(32'hba99166b),
	.w7(32'hbb2582ca),
	.w8(32'hbb410dd2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba967e00),
	.w1(32'hb9cab391),
	.w2(32'h39de537d),
	.w3(32'hbb18b5cb),
	.w4(32'hbafc92b9),
	.w5(32'h3ac51d57),
	.w6(32'h385a451e),
	.w7(32'h3b6390fb),
	.w8(32'h39bfe223),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa70200),
	.w1(32'h3afe2eee),
	.w2(32'h3b0353ff),
	.w3(32'h3b112778),
	.w4(32'h3a881580),
	.w5(32'hbb603d20),
	.w6(32'h3b00ce64),
	.w7(32'h3ac8cba6),
	.w8(32'hbb522002),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13e636),
	.w1(32'h3b021e8f),
	.w2(32'h3a34ea2c),
	.w3(32'hbaa164ea),
	.w4(32'h3b6a99a5),
	.w5(32'hb94349ee),
	.w6(32'h3b1be8e4),
	.w7(32'h3b7de32f),
	.w8(32'h3a78c3dc),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927be9d),
	.w1(32'h3b0b1480),
	.w2(32'h3afc6a7f),
	.w3(32'h392f2ebf),
	.w4(32'hb95bfc61),
	.w5(32'hbb0d104f),
	.w6(32'h3b126985),
	.w7(32'h3b090179),
	.w8(32'hbb97c297),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6020),
	.w1(32'hb89bac07),
	.w2(32'hbb715416),
	.w3(32'h3ae483e0),
	.w4(32'hba8c7730),
	.w5(32'h3b3eab39),
	.w6(32'h3988ce67),
	.w7(32'hbb56ecc0),
	.w8(32'h3b586aba),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71da46),
	.w1(32'hbac2a33c),
	.w2(32'hbabcc3fb),
	.w3(32'hba8e2fa5),
	.w4(32'hbaa76049),
	.w5(32'hbb933c83),
	.w6(32'hb9d73d3d),
	.w7(32'hbad3e537),
	.w8(32'hbab4467b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cfdf6),
	.w1(32'h3a745f4a),
	.w2(32'hbb32d963),
	.w3(32'hba747a64),
	.w4(32'hbb17be62),
	.w5(32'h3a5f2974),
	.w6(32'h3b7cefc1),
	.w7(32'h369b65c3),
	.w8(32'h3ae79c30),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9583262),
	.w1(32'h3bb233c3),
	.w2(32'h3b9d3470),
	.w3(32'h3bef8785),
	.w4(32'h3bb99784),
	.w5(32'h3b1fcd53),
	.w6(32'h3bd9b67f),
	.w7(32'h3ba7ea72),
	.w8(32'h3aa40724),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4338ca),
	.w1(32'h3b8ec762),
	.w2(32'h3bff8223),
	.w3(32'h3b51f448),
	.w4(32'h3b9c501f),
	.w5(32'h3a4ad1de),
	.w6(32'h3b9d2640),
	.w7(32'h3bcbe8b0),
	.w8(32'hb9b442ad),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad79f01),
	.w1(32'hbafeebf8),
	.w2(32'hbb00aba8),
	.w3(32'h3a14dd90),
	.w4(32'hb9c18cea),
	.w5(32'h3aaa8cf0),
	.w6(32'hbac8294d),
	.w7(32'hbaca851d),
	.w8(32'h39b9f8cf),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38397e88),
	.w1(32'h3b4fb589),
	.w2(32'hba638c58),
	.w3(32'h3b2f336b),
	.w4(32'hb9e4c887),
	.w5(32'h3c501309),
	.w6(32'h3b2bddc3),
	.w7(32'hbb469019),
	.w8(32'h3c055a33),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e6f29),
	.w1(32'h3c616eba),
	.w2(32'h3bef0962),
	.w3(32'h3c53943f),
	.w4(32'h3bde6519),
	.w5(32'h3b29234e),
	.w6(32'h3c383971),
	.w7(32'h3beca02d),
	.w8(32'h36afc54d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25f59d),
	.w1(32'h3b0ccd81),
	.w2(32'h3a0820d2),
	.w3(32'h3b6c192d),
	.w4(32'h3b1c89c7),
	.w5(32'hba2a8053),
	.w6(32'h3aaf33b0),
	.w7(32'hba236269),
	.w8(32'hb926a0b4),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f3f89),
	.w1(32'hbab0cbd5),
	.w2(32'hbaf8a08a),
	.w3(32'hb7ede5f5),
	.w4(32'hb8f04686),
	.w5(32'hbbd5306e),
	.w6(32'h360648f2),
	.w7(32'hba860672),
	.w8(32'hbb6f7868),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99ceb8),
	.w1(32'hbb7780fa),
	.w2(32'hbbc27c5c),
	.w3(32'hbb9197c1),
	.w4(32'hbb937461),
	.w5(32'hba29dbeb),
	.w6(32'hbb108fc6),
	.w7(32'hbb8d87c8),
	.w8(32'hbab9ec3a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb0f03),
	.w1(32'hb76265e3),
	.w2(32'h3a0d0146),
	.w3(32'hb9073d1e),
	.w4(32'h3a92b713),
	.w5(32'h3a5c7213),
	.w6(32'hbb02ce2d),
	.w7(32'hba8f2a60),
	.w8(32'h3adccd35),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8996f61),
	.w1(32'h3b6579e0),
	.w2(32'h3b2a8451),
	.w3(32'h3b6e6cee),
	.w4(32'h3b3bd872),
	.w5(32'hbba6fe68),
	.w6(32'h3b6c6cb8),
	.w7(32'h3b1770e9),
	.w8(32'hba3d9780),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397fbdcf),
	.w1(32'hbb47c292),
	.w2(32'hbba46a9a),
	.w3(32'hbb0f08fc),
	.w4(32'hbbcb7434),
	.w5(32'hbafec9ab),
	.w6(32'hbae41bbf),
	.w7(32'hbbe4f227),
	.w8(32'hba680214),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86e351),
	.w1(32'hbb071b9f),
	.w2(32'hbb21a70f),
	.w3(32'hbb858a4a),
	.w4(32'hbb519efe),
	.w5(32'hb8c4e9b9),
	.w6(32'hbb4f802d),
	.w7(32'hbb10236c),
	.w8(32'h3a99a028),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4247a0),
	.w1(32'hbad0fad5),
	.w2(32'hbb30c53a),
	.w3(32'h3aa76900),
	.w4(32'hba845964),
	.w5(32'hbb71b882),
	.w6(32'h3a286158),
	.w7(32'hbb273f91),
	.w8(32'h3b67abe4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad28ab0),
	.w1(32'hbad819c1),
	.w2(32'hbb7b9e30),
	.w3(32'hbb25d852),
	.w4(32'hbb8dfe20),
	.w5(32'h3a8c5326),
	.w6(32'hbb2e47fe),
	.w7(32'hbb27291c),
	.w8(32'h3b0258af),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d560),
	.w1(32'hbb35bd65),
	.w2(32'h3b68178f),
	.w3(32'hbacf667e),
	.w4(32'h3bc34699),
	.w5(32'hbbd39768),
	.w6(32'hbac59f18),
	.w7(32'h3b973586),
	.w8(32'hbba8ed6b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4dfab),
	.w1(32'hbb9473a4),
	.w2(32'hbb86babd),
	.w3(32'hbb4e9021),
	.w4(32'hbb8e4b99),
	.w5(32'hbbbe8080),
	.w6(32'hbb86ef18),
	.w7(32'hbb8aa35b),
	.w8(32'hbbb3ba3d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecbd49),
	.w1(32'hbb13c7bc),
	.w2(32'hbb6a8538),
	.w3(32'hbbb74d9b),
	.w4(32'hbb953b5b),
	.w5(32'hbb740b7a),
	.w6(32'hbb658d20),
	.w7(32'hbb3c5541),
	.w8(32'hbb05d27b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2e4c8),
	.w1(32'h3b38da90),
	.w2(32'h3ad1b55f),
	.w3(32'hbae0d5d6),
	.w4(32'hba734676),
	.w5(32'hb998d697),
	.w6(32'h3b919272),
	.w7(32'h3b28e971),
	.w8(32'hbaeece09),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bf90b),
	.w1(32'hb97cde61),
	.w2(32'hbb255c49),
	.w3(32'h3b421199),
	.w4(32'hba89557f),
	.w5(32'h3b56ad78),
	.w6(32'h3a39e8fc),
	.w7(32'hbb8bcb97),
	.w8(32'hbaadf9a7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62ee70),
	.w1(32'hbb3dc583),
	.w2(32'h3b01342a),
	.w3(32'hbb87d59e),
	.w4(32'hb629a245),
	.w5(32'h3a3fd073),
	.w6(32'hbb72d36e),
	.w7(32'hba66d5fb),
	.w8(32'hba779544),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f944a),
	.w1(32'hbb92b959),
	.w2(32'hbb110e4d),
	.w3(32'hbbbe6b9b),
	.w4(32'hbbb0aa58),
	.w5(32'hba7a692c),
	.w6(32'h3c1d058a),
	.w7(32'hbc1721f4),
	.w8(32'h3b2681f5),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad340c8),
	.w1(32'h3a29c26b),
	.w2(32'h3b3661c9),
	.w3(32'h3982cc36),
	.w4(32'h3c3a8ea3),
	.w5(32'h3b456957),
	.w6(32'hbc365e62),
	.w7(32'h3be5af1c),
	.w8(32'hbbba06b9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc413c92),
	.w1(32'hba2afa01),
	.w2(32'h3c1b3d38),
	.w3(32'h3bb533df),
	.w4(32'hbb6fec4c),
	.w5(32'h3bd6a256),
	.w6(32'hbbd1c982),
	.w7(32'h3c54e038),
	.w8(32'h3b3b1a43),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebe751),
	.w1(32'h3b902fcc),
	.w2(32'hbbb9a805),
	.w3(32'h3c2d7b65),
	.w4(32'h3b826ec5),
	.w5(32'h3bc2b025),
	.w6(32'h3cb22c8e),
	.w7(32'h3b06c7bd),
	.w8(32'h3c2348ba),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e5895),
	.w1(32'hb86783af),
	.w2(32'hbb23b7dc),
	.w3(32'h3b09931d),
	.w4(32'hbb0d2847),
	.w5(32'h39cf68fa),
	.w6(32'h3b865222),
	.w7(32'hbb88f408),
	.w8(32'h3bda5fd9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad7470),
	.w1(32'hbae82084),
	.w2(32'hbbff95e1),
	.w3(32'h3a7a13a4),
	.w4(32'h3beb377b),
	.w5(32'hbb0b67cc),
	.w6(32'h371938ea),
	.w7(32'h3baea11b),
	.w8(32'hbac3578d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0b072),
	.w1(32'h3a1e4b86),
	.w2(32'hbbca0506),
	.w3(32'hbb8dfabd),
	.w4(32'h3a03cae1),
	.w5(32'h3b101db9),
	.w6(32'hbc67c690),
	.w7(32'hbbcb5cdc),
	.w8(32'h3bdd4536),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9be373),
	.w1(32'h3b16d609),
	.w2(32'hbb58ace8),
	.w3(32'h3b8f393d),
	.w4(32'h3b0f4317),
	.w5(32'hb99e11af),
	.w6(32'h3cd09269),
	.w7(32'hbbe4b6dc),
	.w8(32'hba071e99),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae56e4),
	.w1(32'h3c858f72),
	.w2(32'h3a0535cb),
	.w3(32'h3c5f602d),
	.w4(32'h3ab0bccb),
	.w5(32'h3b0208fa),
	.w6(32'h3c89f5d1),
	.w7(32'hbbdf8c9b),
	.w8(32'hbb911084),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b736b40),
	.w1(32'hbb52df21),
	.w2(32'h3798f4ad),
	.w3(32'h39aedf26),
	.w4(32'hbb9a4f3b),
	.w5(32'h3bab5c15),
	.w6(32'hba6e2800),
	.w7(32'hbba7dc28),
	.w8(32'h3b4195c9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97d57a),
	.w1(32'hb909e139),
	.w2(32'hbb79f3d8),
	.w3(32'h3b1ecdfa),
	.w4(32'hbadd55ba),
	.w5(32'hbc0d6d40),
	.w6(32'h39b0073e),
	.w7(32'hbb377c0f),
	.w8(32'hbb4f850c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb763842),
	.w1(32'hbb602b62),
	.w2(32'hbb0d6287),
	.w3(32'h3ab0c1fa),
	.w4(32'h3ba8545b),
	.w5(32'hbbdd040c),
	.w6(32'h3b5a387e),
	.w7(32'hbac57233),
	.w8(32'hbbc66e64),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc057950),
	.w1(32'hbc37b4ff),
	.w2(32'h3bcf9989),
	.w3(32'hbc3787d2),
	.w4(32'h3a9b0b11),
	.w5(32'hbb073f6b),
	.w6(32'h3b67b237),
	.w7(32'hba7db91d),
	.w8(32'hbb94e7f6),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83e1cff),
	.w1(32'hbafc72a6),
	.w2(32'h3b9e12cc),
	.w3(32'hb81c07d9),
	.w4(32'h3b8085b7),
	.w5(32'h3ab72bc1),
	.w6(32'h3af0938a),
	.w7(32'h3b992d49),
	.w8(32'h39a1af87),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6469f7),
	.w1(32'h3c6bc2b6),
	.w2(32'h3c0e2ce9),
	.w3(32'hbbb24557),
	.w4(32'h3c7ed758),
	.w5(32'hbc2da64e),
	.w6(32'hbb18f976),
	.w7(32'h3cf23584),
	.w8(32'hbc2fdf9e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6782c9),
	.w1(32'h3ab85300),
	.w2(32'hb9aebf66),
	.w3(32'hba1801f1),
	.w4(32'hbb85ae14),
	.w5(32'h3c776a27),
	.w6(32'hb9fa35d9),
	.w7(32'hbb5a217a),
	.w8(32'h3c09b61e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a970c),
	.w1(32'hbc1cc067),
	.w2(32'h3cc7e5d4),
	.w3(32'hbbaaa533),
	.w4(32'h3b0c9e8a),
	.w5(32'h3a60e45e),
	.w6(32'hbc3e26e6),
	.w7(32'h3c6f804a),
	.w8(32'h3b14195c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3fcf4),
	.w1(32'hbb93a2b2),
	.w2(32'hbb09d882),
	.w3(32'hbba3a988),
	.w4(32'hbb33f55d),
	.w5(32'h3c21276f),
	.w6(32'hbc118c7e),
	.w7(32'hbbbd4c29),
	.w8(32'h3b432c7f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5634b5),
	.w1(32'hbabb112b),
	.w2(32'h3b0f32bd),
	.w3(32'h3b44de81),
	.w4(32'hbb28a494),
	.w5(32'h3ab89bf2),
	.w6(32'h3c5de9b8),
	.w7(32'h3aa620df),
	.w8(32'hba97acf0),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9f6ab),
	.w1(32'h3b3e737b),
	.w2(32'hb9df6171),
	.w3(32'h39a9188e),
	.w4(32'h3b42be1b),
	.w5(32'h3b77382b),
	.w6(32'h3c0d74db),
	.w7(32'h3b96efaf),
	.w8(32'hbb997048),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdff55d),
	.w1(32'h3a6d27fc),
	.w2(32'h3abd62b8),
	.w3(32'h3ab5f42e),
	.w4(32'h3a3cf7ee),
	.w5(32'hbbb99129),
	.w6(32'hbb5faca8),
	.w7(32'h3b8e655a),
	.w8(32'hbb1cfe1a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc102a2c),
	.w1(32'h3b725ef7),
	.w2(32'h3bee4be1),
	.w3(32'hbbd8da1d),
	.w4(32'hbb23aad6),
	.w5(32'hbb359308),
	.w6(32'h3c633488),
	.w7(32'h3b2368b7),
	.w8(32'hba2e2ab0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef358f),
	.w1(32'hbb8f71be),
	.w2(32'hbb6eaba4),
	.w3(32'hbb24d851),
	.w4(32'h3a891d00),
	.w5(32'hbc0016a2),
	.w6(32'h3c13bb0e),
	.w7(32'hbbfba35a),
	.w8(32'hbb8bb1a0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6bfd3),
	.w1(32'hbbf071c3),
	.w2(32'hbc8b66bd),
	.w3(32'hb9a8bbe3),
	.w4(32'hbba62cb6),
	.w5(32'h3b60844b),
	.w6(32'hbc15ae5a),
	.w7(32'hbc310d4d),
	.w8(32'h3b233e3b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb893bff),
	.w1(32'h3c23eed0),
	.w2(32'hb9eef99e),
	.w3(32'hba7d04d3),
	.w4(32'hbbdc2bad),
	.w5(32'hbbb6870c),
	.w6(32'h3c2cbc71),
	.w7(32'hbc01529c),
	.w8(32'hbc08c75a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2127f6),
	.w1(32'hbc0cdda7),
	.w2(32'hbc7c06d0),
	.w3(32'hbba7e161),
	.w4(32'hbc183115),
	.w5(32'hbb5a9266),
	.w6(32'h39f47113),
	.w7(32'hbaa959ff),
	.w8(32'hbbb1ee77),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39a085),
	.w1(32'h3ba7ffba),
	.w2(32'hbbdf70d2),
	.w3(32'hbb93f46e),
	.w4(32'hba698250),
	.w5(32'h39bf4ad7),
	.w6(32'h3c2511e4),
	.w7(32'h3accf7fb),
	.w8(32'h3ad0ebc9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa79fcd),
	.w1(32'h3b2f3546),
	.w2(32'h3a5bb8db),
	.w3(32'h3a2a2a86),
	.w4(32'h3ab7a7df),
	.w5(32'h3b8436ff),
	.w6(32'hb99a8990),
	.w7(32'h3b0d569e),
	.w8(32'h3ac25610),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7a658),
	.w1(32'hbaea2447),
	.w2(32'h3bb60ea4),
	.w3(32'hbb75fce6),
	.w4(32'h3ba5ff28),
	.w5(32'hbb1b31d5),
	.w6(32'hba9d0e47),
	.w7(32'h3b9cd507),
	.w8(32'hbbaf4e18),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule