module layer_8_featuremap_201(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a11b0),
	.w1(32'hbb8a00f4),
	.w2(32'hbbab215a),
	.w3(32'hbc081665),
	.w4(32'hbb39f0f9),
	.w5(32'h3a3f2c5f),
	.w6(32'hbc2fa9fa),
	.w7(32'hbbcf8701),
	.w8(32'hbc23855b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59711e),
	.w1(32'hbb0f5a8e),
	.w2(32'hbb40287a),
	.w3(32'h3b203d1a),
	.w4(32'hbbf28b89),
	.w5(32'hbbeae8b8),
	.w6(32'hb9626422),
	.w7(32'h3992ba61),
	.w8(32'h3ad5cf0d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916a0a4),
	.w1(32'h3c689f7a),
	.w2(32'h3bf3dbfc),
	.w3(32'hbb1b7cf4),
	.w4(32'h3b0a366f),
	.w5(32'hbc074168),
	.w6(32'h3c115f76),
	.w7(32'h3c48d888),
	.w8(32'h3c3e59ed),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcffcc),
	.w1(32'hbc09f605),
	.w2(32'hbc4db379),
	.w3(32'hba7ba806),
	.w4(32'hba1fe9e7),
	.w5(32'hbc1abcdb),
	.w6(32'hbaa22e16),
	.w7(32'hbb68f61b),
	.w8(32'hbbc60a13),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2799fa),
	.w1(32'h3a79d7f8),
	.w2(32'h3bd0b4e3),
	.w3(32'hbbcc2a5f),
	.w4(32'h3a8105f8),
	.w5(32'h3bf1f2ac),
	.w6(32'hbb96731c),
	.w7(32'hbabfcb69),
	.w8(32'hbb1b66a1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c63e5),
	.w1(32'h396489d2),
	.w2(32'hbb09821c),
	.w3(32'h3be77545),
	.w4(32'h3a4c3405),
	.w5(32'h3b9f7a9b),
	.w6(32'hbab7de41),
	.w7(32'hbbdd5d63),
	.w8(32'hbae8479f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0044e),
	.w1(32'h3acb8565),
	.w2(32'h3bf06b15),
	.w3(32'h3c10946b),
	.w4(32'h3c15d42b),
	.w5(32'h3c6c0592),
	.w6(32'hbbc52ec7),
	.w7(32'hbb038070),
	.w8(32'hbb6d0c2a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a0536),
	.w1(32'hbbfb6c9e),
	.w2(32'hbbaa084e),
	.w3(32'h3c2f8435),
	.w4(32'hbbf49db0),
	.w5(32'h3a26ac5a),
	.w6(32'hbc6eae8c),
	.w7(32'hbbe17a84),
	.w8(32'hbbc4210b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d7fb6),
	.w1(32'hbc048497),
	.w2(32'hbc27035d),
	.w3(32'h3c698c79),
	.w4(32'hbc2b99f8),
	.w5(32'hbc41f511),
	.w6(32'hbb7ad2e5),
	.w7(32'hbb2be04b),
	.w8(32'hbbb0221e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd524e9),
	.w1(32'h3be20d24),
	.w2(32'h3c32d14f),
	.w3(32'hbbc3a456),
	.w4(32'hbba39d98),
	.w5(32'h3b93cf81),
	.w6(32'hbbc0e5c2),
	.w7(32'hb8876516),
	.w8(32'h3c0d8fd5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08264f),
	.w1(32'h3b847ab0),
	.w2(32'h3a75baeb),
	.w3(32'h3bfdda78),
	.w4(32'h3c53fa77),
	.w5(32'h3c203521),
	.w6(32'h3895c9a2),
	.w7(32'hbbe77f55),
	.w8(32'hbb57f0b1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6ac6c),
	.w1(32'h3c5ec51a),
	.w2(32'h3c982df1),
	.w3(32'hb9247569),
	.w4(32'h3c86a64a),
	.w5(32'h3cdc1613),
	.w6(32'h3b2c1355),
	.w7(32'h3b6d7619),
	.w8(32'h3b3369e2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c739e36),
	.w1(32'hbc0c5d81),
	.w2(32'hbc1e510d),
	.w3(32'h3ca5d0c7),
	.w4(32'hba409f1f),
	.w5(32'h3a12ea7e),
	.w6(32'hba8b70fa),
	.w7(32'hba0d2910),
	.w8(32'h3a9acd65),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb410fbe),
	.w1(32'h3b7e70e6),
	.w2(32'h3b40a975),
	.w3(32'h3987a7a8),
	.w4(32'h3c3735df),
	.w5(32'hbbe2147f),
	.w6(32'h3c09f1e8),
	.w7(32'h3c555180),
	.w8(32'hb8cce763),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa9a73),
	.w1(32'h38776741),
	.w2(32'hb882391b),
	.w3(32'h3b4e998d),
	.w4(32'h3b180282),
	.w5(32'h3ae5bc88),
	.w6(32'h39746646),
	.w7(32'h3b01bcc5),
	.w8(32'h3ad61a3b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0127ec),
	.w1(32'hbb76b99a),
	.w2(32'h3c2230a0),
	.w3(32'h3b775fe8),
	.w4(32'h3b23e3e0),
	.w5(32'hbb0a78ff),
	.w6(32'h3bfdcf66),
	.w7(32'h3b8e60d8),
	.w8(32'h3bb945f7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1382f3),
	.w1(32'hba11a884),
	.w2(32'h3ad5cc01),
	.w3(32'h3b9297cd),
	.w4(32'hbbd54196),
	.w5(32'h3b8ac390),
	.w6(32'hba5fcdb7),
	.w7(32'hbbd3195e),
	.w8(32'hbbbc178f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a3934),
	.w1(32'h3bbe2bce),
	.w2(32'hba82d376),
	.w3(32'h3b7431b2),
	.w4(32'h3c3b108d),
	.w5(32'hbc5522bb),
	.w6(32'h3c501865),
	.w7(32'h3c088128),
	.w8(32'h3c0db3e4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce2b66),
	.w1(32'h3bd7ebaf),
	.w2(32'h3b814b53),
	.w3(32'hbbb1d5db),
	.w4(32'h3a863227),
	.w5(32'h3c834720),
	.w6(32'hb9228bd9),
	.w7(32'hbc28e77a),
	.w8(32'h3abf1ca7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6c05e),
	.w1(32'hbbd00d4c),
	.w2(32'hbc19e03f),
	.w3(32'h3c36fe28),
	.w4(32'hbb3ed344),
	.w5(32'hbbf86016),
	.w6(32'hbbba15bb),
	.w7(32'hbbd904aa),
	.w8(32'hbbe083bd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef40ed),
	.w1(32'hbbc162f1),
	.w2(32'hbb72d78d),
	.w3(32'hbb91a9ba),
	.w4(32'h3bc553bf),
	.w5(32'hbb893729),
	.w6(32'hbc275774),
	.w7(32'hbc1c0fc3),
	.w8(32'h3b41db88),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c21764),
	.w1(32'h3c00fed1),
	.w2(32'hbbd66048),
	.w3(32'hbc0fe3c1),
	.w4(32'hbafd666b),
	.w5(32'hba694e92),
	.w6(32'h3b5adb9b),
	.w7(32'h3988e7f2),
	.w8(32'hbbdf3da0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb953c12),
	.w1(32'h3b6fea2e),
	.w2(32'h3bcaa970),
	.w3(32'h3970db03),
	.w4(32'h3aad4762),
	.w5(32'h3bc8820c),
	.w6(32'h3c20686a),
	.w7(32'h3bd461fb),
	.w8(32'h3ab96f3b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b762843),
	.w1(32'hbb59368a),
	.w2(32'hbbdef94a),
	.w3(32'hba6ebd77),
	.w4(32'h3b06056f),
	.w5(32'h3bce1d19),
	.w6(32'h3abad2c4),
	.w7(32'hbc0e47eb),
	.w8(32'hbb2dd7cc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e4f7),
	.w1(32'hbc027080),
	.w2(32'hbc160312),
	.w3(32'h3c114e98),
	.w4(32'h3a8feac6),
	.w5(32'h3a8d3a7d),
	.w6(32'hbb1c0f2b),
	.w7(32'hbbe835f6),
	.w8(32'hbb0dfefe),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9ca74),
	.w1(32'h3bc83ad4),
	.w2(32'h3be826ce),
	.w3(32'h3aee535d),
	.w4(32'h3bce0604),
	.w5(32'h3c0f2fa9),
	.w6(32'hbc1cde67),
	.w7(32'h3b9704a8),
	.w8(32'hbbbc8d38),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e6c41),
	.w1(32'hbc164fcd),
	.w2(32'hbb5164e0),
	.w3(32'h3bb4224c),
	.w4(32'h3b8beec4),
	.w5(32'h3c4aff6b),
	.w6(32'hbb963f4a),
	.w7(32'hbc04e4d1),
	.w8(32'hbb84f355),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7932d7),
	.w1(32'h3c0bc7dd),
	.w2(32'hba8305a2),
	.w3(32'h3c4585fb),
	.w4(32'h3c9774dc),
	.w5(32'hbb314c56),
	.w6(32'h3bc1ae83),
	.w7(32'h3c261adf),
	.w8(32'h39395b63),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40b847),
	.w1(32'hbba87f8e),
	.w2(32'hbb873f4b),
	.w3(32'hba42125e),
	.w4(32'hbc2988f8),
	.w5(32'hbbff4d7d),
	.w6(32'h3b70f575),
	.w7(32'hba68d94d),
	.w8(32'h3b645ad6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f48e3),
	.w1(32'h3ba6f57b),
	.w2(32'h3c29b428),
	.w3(32'hbb962242),
	.w4(32'h3cea1077),
	.w5(32'h3d0ed687),
	.w6(32'h3a7c51ab),
	.w7(32'h3b5af45e),
	.w8(32'h39e2e8ff),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd095a9),
	.w1(32'h39b62492),
	.w2(32'hb9aa0351),
	.w3(32'h3cfdc914),
	.w4(32'hba170897),
	.w5(32'hba8e985f),
	.w6(32'hba776653),
	.w7(32'hbb522634),
	.w8(32'hbbbae758),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affeb78),
	.w1(32'hbb910bb6),
	.w2(32'hbbf39679),
	.w3(32'hbb17b3ab),
	.w4(32'hbc6a8e31),
	.w5(32'hbc219fe6),
	.w6(32'h3bcf5f1b),
	.w7(32'hbadcce4d),
	.w8(32'h3a78c6c6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b575790),
	.w1(32'hbbabf538),
	.w2(32'hbc999fe7),
	.w3(32'hbc34e8cd),
	.w4(32'hba0934e1),
	.w5(32'hbc08d26f),
	.w6(32'h3b924e4a),
	.w7(32'h3b2ee675),
	.w8(32'h3b9f22ae),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f1755),
	.w1(32'h3a52ef19),
	.w2(32'h3c3c8e4b),
	.w3(32'hbc01f2dc),
	.w4(32'h3c2762c3),
	.w5(32'h3c610fe9),
	.w6(32'hbbb9f264),
	.w7(32'hba76f3cb),
	.w8(32'hbc44ddf3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ea4a1),
	.w1(32'hbb478b46),
	.w2(32'hbb9dd6df),
	.w3(32'hb9e395e3),
	.w4(32'hbbd151e1),
	.w5(32'hbc19e5de),
	.w6(32'h3b6874a0),
	.w7(32'h3ab849ff),
	.w8(32'hba57aec7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc77927),
	.w1(32'hbb60249e),
	.w2(32'h3c4f3a9a),
	.w3(32'hbbc7dba4),
	.w4(32'h3bce1616),
	.w5(32'h3c2ba1d4),
	.w6(32'hbc8459e7),
	.w7(32'hbc1d7091),
	.w8(32'hb9c3195a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f80d4),
	.w1(32'h3a647d43),
	.w2(32'hbb50e520),
	.w3(32'h3c35865e),
	.w4(32'h3b5e861e),
	.w5(32'h3ab211b1),
	.w6(32'h3a27c32e),
	.w7(32'hbaac697f),
	.w8(32'hbb8041ca),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8c5b3),
	.w1(32'hbc1f8ca9),
	.w2(32'hbc629d1e),
	.w3(32'hba8af880),
	.w4(32'hbc51654c),
	.w5(32'hbc973c96),
	.w6(32'h3991cbb9),
	.w7(32'h3880f7ba),
	.w8(32'h3b35cd92),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe21c93),
	.w1(32'hbb8658ea),
	.w2(32'hbb3a7f39),
	.w3(32'hbc35a52f),
	.w4(32'hbaba3912),
	.w5(32'hb99e5827),
	.w6(32'hbbf08e58),
	.w7(32'hbbe69add),
	.w8(32'hbbac7bac),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc1b0e),
	.w1(32'hbbc557b6),
	.w2(32'h3b8c7b1c),
	.w3(32'h3b217ac3),
	.w4(32'hb9420823),
	.w5(32'h3c5fa49c),
	.w6(32'hbc72da8e),
	.w7(32'hbbfe67f8),
	.w8(32'hbb3ae4e7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02fd7c),
	.w1(32'hbbe48736),
	.w2(32'hbc860a7b),
	.w3(32'h3c02f055),
	.w4(32'hbc441ab2),
	.w5(32'hbcbb229b),
	.w6(32'hba2bcd65),
	.w7(32'hbc169bed),
	.w8(32'hbaf0db3a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c9228),
	.w1(32'h3a300340),
	.w2(32'h3b4f6461),
	.w3(32'hbc849e3b),
	.w4(32'h3b0c0fae),
	.w5(32'h3b99d994),
	.w6(32'h3b7b4a56),
	.w7(32'h3b9c8afb),
	.w8(32'h3b37c0bf),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab92879),
	.w1(32'hbbcffd1e),
	.w2(32'hbb92ccd0),
	.w3(32'h3b6520a3),
	.w4(32'hbbb8ff08),
	.w5(32'h3a9968cc),
	.w6(32'hbada305f),
	.w7(32'hbb263f87),
	.w8(32'h3b15a494),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7bb96),
	.w1(32'h3b47dc57),
	.w2(32'h3b9f8898),
	.w3(32'hbab62322),
	.w4(32'h39f543e6),
	.w5(32'h3a2276bb),
	.w6(32'h3ad201e5),
	.w7(32'h3b313dcc),
	.w8(32'hbb159ae4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13af4b),
	.w1(32'h3bcd22fa),
	.w2(32'h3c0f0de0),
	.w3(32'hbbf72625),
	.w4(32'h3c43601b),
	.w5(32'h3bfe48d2),
	.w6(32'h3afe5604),
	.w7(32'hbb5031fc),
	.w8(32'hbbfeae34),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b020b),
	.w1(32'hba0a0a66),
	.w2(32'h3ac59c01),
	.w3(32'h3c0b9804),
	.w4(32'h3b3829c2),
	.w5(32'h3b62369b),
	.w6(32'hba8ae3e0),
	.w7(32'hbae67b7d),
	.w8(32'hbaec84d7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd4fd2),
	.w1(32'h3c4b9bb2),
	.w2(32'h3d09e0ac),
	.w3(32'h3b7563c1),
	.w4(32'h3cb881b6),
	.w5(32'h3d450e16),
	.w6(32'hbc4b84ee),
	.w7(32'hbbbab29b),
	.w8(32'hbc0f3a75),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2ef29),
	.w1(32'hba3b7285),
	.w2(32'h3a63f402),
	.w3(32'h3d0719a1),
	.w4(32'hbab4a1ad),
	.w5(32'h3c051154),
	.w6(32'hba5319f0),
	.w7(32'hbba0e955),
	.w8(32'hbb311ab1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c7252),
	.w1(32'h3ace0beb),
	.w2(32'hbbcd1039),
	.w3(32'hba2623e0),
	.w4(32'h3abfd08b),
	.w5(32'hbba159cc),
	.w6(32'h3aeb30b0),
	.w7(32'h3c505f0e),
	.w8(32'h3c20d9c6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb933385),
	.w1(32'h3b8b5b1e),
	.w2(32'hbb050011),
	.w3(32'hb841f77a),
	.w4(32'h39934b09),
	.w5(32'h39a044bb),
	.w6(32'h3c1b7206),
	.w7(32'hba739b41),
	.w8(32'h3c29c565),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9772bb),
	.w1(32'hbafa5322),
	.w2(32'hba748d2c),
	.w3(32'h3a9d5338),
	.w4(32'hbaa16d6f),
	.w5(32'hbb5e3e0a),
	.w6(32'hbaf9ee93),
	.w7(32'hbbac9e00),
	.w8(32'hba91a507),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4d5d1),
	.w1(32'hbb314678),
	.w2(32'hbbd3c43a),
	.w3(32'hbb2d3ad1),
	.w4(32'hbb5eef10),
	.w5(32'hbad423d1),
	.w6(32'hbba73329),
	.w7(32'hbc1f6445),
	.w8(32'hbbc070e1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4e78f),
	.w1(32'hbbf09979),
	.w2(32'hbb2f142a),
	.w3(32'h3aa684db),
	.w4(32'hbbf5f0da),
	.w5(32'hbb33b065),
	.w6(32'hbbb9e72e),
	.w7(32'hbb46aaa9),
	.w8(32'hba93e61e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d199a2),
	.w1(32'h3b5b792c),
	.w2(32'hbc110808),
	.w3(32'h39eca79a),
	.w4(32'h3a490256),
	.w5(32'hbc5d3cb2),
	.w6(32'hba1b7213),
	.w7(32'hbbac1295),
	.w8(32'hbbbd0368),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae03276),
	.w1(32'h3bd8b5b6),
	.w2(32'h3aafc322),
	.w3(32'hbbc7bf2f),
	.w4(32'hb90ca10b),
	.w5(32'h3c16532b),
	.w6(32'h3b8c58a5),
	.w7(32'hbb121f1e),
	.w8(32'h3c544093),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c186f93),
	.w1(32'h3a44fd7c),
	.w2(32'hbb82bbc9),
	.w3(32'h3bb40906),
	.w4(32'h3bbb615f),
	.w5(32'h39e10f6d),
	.w6(32'h3c046a92),
	.w7(32'h3bfcf91b),
	.w8(32'h3bd50ead),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7cc90),
	.w1(32'h3c244fbd),
	.w2(32'h3c134d2e),
	.w3(32'hbb074746),
	.w4(32'h3c5c31e0),
	.w5(32'h3b953224),
	.w6(32'h3c0c017e),
	.w7(32'h3a99867e),
	.w8(32'hbb8317ba),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb981e2b),
	.w1(32'h3b9a3df0),
	.w2(32'h3b92eb36),
	.w3(32'hbba58061),
	.w4(32'h3baba0ab),
	.w5(32'h3bf66e63),
	.w6(32'h3b910db7),
	.w7(32'h3b887439),
	.w8(32'hba3f43ee),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ac17),
	.w1(32'h3b27eb48),
	.w2(32'h3be972e6),
	.w3(32'hbb9b9783),
	.w4(32'h3b6958e1),
	.w5(32'h3beab3f5),
	.w6(32'hb9076674),
	.w7(32'h3adad478),
	.w8(32'h3b33c1c4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d8345),
	.w1(32'hbb7fb429),
	.w2(32'hbb1e87e8),
	.w3(32'h3c0382f5),
	.w4(32'h3b25cf7f),
	.w5(32'hba994895),
	.w6(32'h3b892725),
	.w7(32'hbbda8489),
	.w8(32'hbbacf4d8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0127f6),
	.w1(32'hbc029a3d),
	.w2(32'hbc733ae4),
	.w3(32'hbb673e07),
	.w4(32'hbbc79a1a),
	.w5(32'hbad6d38d),
	.w6(32'hbbe86985),
	.w7(32'hbafedd16),
	.w8(32'hb5f246e7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b889a21),
	.w1(32'hbc3b7b43),
	.w2(32'hbc1b9187),
	.w3(32'h3c20aef5),
	.w4(32'h3a6c0262),
	.w5(32'h3b451a02),
	.w6(32'hbc30019b),
	.w7(32'hbc7ca2de),
	.w8(32'hbc1f0f71),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda0531),
	.w1(32'hbc96db74),
	.w2(32'hbc7926ea),
	.w3(32'h3b352da3),
	.w4(32'hbcad921c),
	.w5(32'hbc8b84c5),
	.w6(32'hb8bca094),
	.w7(32'h3b9f1ac3),
	.w8(32'h3b80e826),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f2f19),
	.w1(32'h3c17d0fb),
	.w2(32'h3c00bc97),
	.w3(32'hbc44e7bc),
	.w4(32'h3c0d12e2),
	.w5(32'h3c22ecc6),
	.w6(32'h3bfc9aa6),
	.w7(32'h3be44026),
	.w8(32'h3c08c5f7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ac45d),
	.w1(32'h3b4d6c96),
	.w2(32'h3b3bea4d),
	.w3(32'h3bff2e35),
	.w4(32'h3ad76134),
	.w5(32'h3aab7281),
	.w6(32'h3bcbf44d),
	.w7(32'h3b9146f4),
	.w8(32'h3bc7dd1a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbf2c8),
	.w1(32'hbbc41831),
	.w2(32'h3b2e7018),
	.w3(32'h3b7e5464),
	.w4(32'h3bbb3b9c),
	.w5(32'h3c12e833),
	.w6(32'hbc4f0d20),
	.w7(32'hbb0f4fbf),
	.w8(32'hbbddac2e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b3d1),
	.w1(32'hbbe8787a),
	.w2(32'hba0bf27b),
	.w3(32'hba220c0b),
	.w4(32'hbbb32576),
	.w5(32'h3b8e4988),
	.w6(32'hbb3e40da),
	.w7(32'hbbe4997d),
	.w8(32'hbb650440),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f7410),
	.w1(32'h3c524c3c),
	.w2(32'h3ce55e8d),
	.w3(32'h3c365d52),
	.w4(32'h3cdd562d),
	.w5(32'h3d23b1ba),
	.w6(32'hbba473cd),
	.w7(32'h3b8bb77f),
	.w8(32'hbb3593ad),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42c3ae),
	.w1(32'hbb452eb4),
	.w2(32'hbbd87db7),
	.w3(32'h3ccfcef6),
	.w4(32'h3c721fdb),
	.w5(32'h3b802523),
	.w6(32'h39aa7f6f),
	.w7(32'h3966e6c2),
	.w8(32'hbc24b943),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33c9db),
	.w1(32'h3bf11077),
	.w2(32'hbc06230d),
	.w3(32'hbb13c919),
	.w4(32'hbbd3b3a7),
	.w5(32'hbc6645dd),
	.w6(32'h3c4c0365),
	.w7(32'h3c488580),
	.w8(32'h3c17ae30),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cfbfc),
	.w1(32'h3a6d7d76),
	.w2(32'h3bebdccb),
	.w3(32'hbbd05d0a),
	.w4(32'hbb7325bf),
	.w5(32'h3bf29b1b),
	.w6(32'h3b66d1d4),
	.w7(32'h3b5e683d),
	.w8(32'h3a4c5a6e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f9e3b),
	.w1(32'hbb2b794d),
	.w2(32'h3b9a7236),
	.w3(32'h3bd1f6c8),
	.w4(32'h3b783864),
	.w5(32'h3c128c05),
	.w6(32'hba3ab49d),
	.w7(32'hbbf0dbbf),
	.w8(32'hbb63436c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51c85a),
	.w1(32'hbac7897c),
	.w2(32'hba8506a3),
	.w3(32'h3bd2b723),
	.w4(32'hb882a550),
	.w5(32'h3acea6ae),
	.w6(32'hbc0f8c30),
	.w7(32'hbbad3d73),
	.w8(32'hbbc8ae54),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8433ec),
	.w1(32'hbb2ea720),
	.w2(32'hbb56905c),
	.w3(32'h3b31cf4a),
	.w4(32'hbbc2d596),
	.w5(32'hbb8c030d),
	.w6(32'h3a39f326),
	.w7(32'hba803c52),
	.w8(32'hbb94b979),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dca2d),
	.w1(32'hbb7393ed),
	.w2(32'hbb3b79f2),
	.w3(32'hbb20127b),
	.w4(32'hbaf088d4),
	.w5(32'h3b6dc6d5),
	.w6(32'hb97e10f0),
	.w7(32'hb90f740f),
	.w8(32'h399cd3fa),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57129c),
	.w1(32'h3c25adf8),
	.w2(32'hba076bc4),
	.w3(32'h3b200e42),
	.w4(32'h3b481071),
	.w5(32'hbc556ea5),
	.w6(32'h3c6b78c6),
	.w7(32'h3c198ffe),
	.w8(32'h3c450b65),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b265cf2),
	.w1(32'hbaef78ca),
	.w2(32'hbaeb55c4),
	.w3(32'hbb86d0db),
	.w4(32'hbb154205),
	.w5(32'hba8de8f7),
	.w6(32'h3a8235e5),
	.w7(32'hbb4dd536),
	.w8(32'h3af7cf51),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8de6ac),
	.w1(32'h3b88b416),
	.w2(32'hbae34622),
	.w3(32'hbb8a8915),
	.w4(32'h3b961990),
	.w5(32'h39d4915f),
	.w6(32'h3bdcba34),
	.w7(32'hba739313),
	.w8(32'h3a82689e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5916ff),
	.w1(32'h3b69ca0e),
	.w2(32'hba779dbd),
	.w3(32'hbb829c90),
	.w4(32'h3bbb6e88),
	.w5(32'h3b11eace),
	.w6(32'h39841149),
	.w7(32'hba253367),
	.w8(32'hbacc1721),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b70e21),
	.w1(32'hbb5a67a0),
	.w2(32'hbb82ff59),
	.w3(32'h3a5f4d67),
	.w4(32'h3bbbbe7b),
	.w5(32'h3bd63130),
	.w6(32'h3bd92d2b),
	.w7(32'h3c0b7632),
	.w8(32'hbb14ebdb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeae278),
	.w1(32'hbbc4a85d),
	.w2(32'hbb101f82),
	.w3(32'hbc11ad7e),
	.w4(32'h3ad77bce),
	.w5(32'hbc1087c7),
	.w6(32'h3c042290),
	.w7(32'h3c05292f),
	.w8(32'h3c1939bb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c68f7),
	.w1(32'hbb2d85f8),
	.w2(32'hbb8c3970),
	.w3(32'h3b20460f),
	.w4(32'h3b7790de),
	.w5(32'h3ba1da7d),
	.w6(32'hbb2b9e2a),
	.w7(32'h3b05921a),
	.w8(32'hbb9efa7e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb578259),
	.w1(32'h3bed2531),
	.w2(32'hbbbc4038),
	.w3(32'hbb6ffff3),
	.w4(32'h3c4500ce),
	.w5(32'hbc44c35b),
	.w6(32'h3c40cf50),
	.w7(32'h3c33f25e),
	.w8(32'h3bcf4373),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb28ada),
	.w1(32'hba9a31af),
	.w2(32'h3b1f3a9f),
	.w3(32'h3a1dc4ff),
	.w4(32'h3ba91f16),
	.w5(32'h3be36cec),
	.w6(32'h3ba63609),
	.w7(32'hbae9abf8),
	.w8(32'h3b603f19),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaf184),
	.w1(32'h3b9eb249),
	.w2(32'hbb1c1b8f),
	.w3(32'h3c8d3c69),
	.w4(32'h3b42f5b1),
	.w5(32'hbc0e2b96),
	.w6(32'h3bef7ec3),
	.w7(32'h3c28c392),
	.w8(32'h3c28cf16),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b317972),
	.w1(32'hbc00588e),
	.w2(32'hbbd3069b),
	.w3(32'hbc0289e0),
	.w4(32'h3c1808a6),
	.w5(32'h3c284617),
	.w6(32'h38d91fec),
	.w7(32'hbaed5f2c),
	.w8(32'hbb0a5dae),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c5724),
	.w1(32'h3b692c0a),
	.w2(32'h3b93935d),
	.w3(32'h3bad2acc),
	.w4(32'h3790df82),
	.w5(32'h3b8a53e9),
	.w6(32'h3b4ecbf0),
	.w7(32'h3b0a4919),
	.w8(32'h3a99f2c9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2124d9),
	.w1(32'h3a976228),
	.w2(32'h3b85d623),
	.w3(32'h3b4d5a64),
	.w4(32'h3b15a65b),
	.w5(32'h3b8f0afa),
	.w6(32'h3b614926),
	.w7(32'h3b89c59a),
	.w8(32'h3bffabd0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0dce9),
	.w1(32'h3b189c76),
	.w2(32'h3ba0d91a),
	.w3(32'h3b13d5a4),
	.w4(32'h3b996736),
	.w5(32'h3c15d41b),
	.w6(32'h3a50c73e),
	.w7(32'hbaa3e06d),
	.w8(32'h37d4f308),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81e071),
	.w1(32'h3c92d8d3),
	.w2(32'hbacee2e8),
	.w3(32'h3bf56ac8),
	.w4(32'h3b9752dd),
	.w5(32'hbb50424b),
	.w6(32'h3c5ca74a),
	.w7(32'h3be262f4),
	.w8(32'h3bc8189b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54d2b7),
	.w1(32'h3af0c89a),
	.w2(32'h3bc22788),
	.w3(32'hbb2950ac),
	.w4(32'hbaf3b927),
	.w5(32'h3be0d33c),
	.w6(32'hbbc84b72),
	.w7(32'h3991cfa4),
	.w8(32'hbc16ccd0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1e1f9),
	.w1(32'h3bc7cb1b),
	.w2(32'h3bb840c1),
	.w3(32'hbbac3226),
	.w4(32'h3c38d6de),
	.w5(32'h3caf45cf),
	.w6(32'hbbd95150),
	.w7(32'hbc1eea0d),
	.w8(32'hbc6ed9ea),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb1719),
	.w1(32'hb79e9c42),
	.w2(32'hba9af155),
	.w3(32'h3c248910),
	.w4(32'hbaa2d6ac),
	.w5(32'hbb301cfe),
	.w6(32'h3a71f348),
	.w7(32'hba9a5925),
	.w8(32'h3ae381d4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba179ec0),
	.w1(32'h3aaee4ae),
	.w2(32'h3bb9ec73),
	.w3(32'h39e48370),
	.w4(32'h3a3602ec),
	.w5(32'h3bf2a2f1),
	.w6(32'hbb4ecef3),
	.w7(32'hbade82e1),
	.w8(32'h383256f0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafaa11),
	.w1(32'h3bfdbff3),
	.w2(32'h3b16909c),
	.w3(32'h3be0ed25),
	.w4(32'hbafbbe47),
	.w5(32'h3c1e18db),
	.w6(32'h3b946a87),
	.w7(32'hbb25e233),
	.w8(32'h3b372351),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63daf8),
	.w1(32'h3b251d62),
	.w2(32'h39e89462),
	.w3(32'h3b324e83),
	.w4(32'h3ad0515a),
	.w5(32'hbab71337),
	.w6(32'h3ad35155),
	.w7(32'hbaa0c759),
	.w8(32'hbaaef4bb),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb300a19),
	.w1(32'hbb0943cd),
	.w2(32'hbbdbf34a),
	.w3(32'hbbd9e8cd),
	.w4(32'hbb537d25),
	.w5(32'hbb8cd495),
	.w6(32'h3bdfb5b1),
	.w7(32'hba1e4572),
	.w8(32'hbaa2091f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af788f9),
	.w1(32'h3b15cc25),
	.w2(32'hbb9d6ce7),
	.w3(32'hbb01be4c),
	.w4(32'hbb8dd969),
	.w5(32'hbc4dabd6),
	.w6(32'h3babbcde),
	.w7(32'hbbabb38c),
	.w8(32'h3b4183b9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20dfaf),
	.w1(32'hbb3a3c3f),
	.w2(32'hbaec0bf3),
	.w3(32'h3b889e75),
	.w4(32'hbb84ee78),
	.w5(32'hb8022878),
	.w6(32'h3ac76a0b),
	.w7(32'hbbe3cb8b),
	.w8(32'hbb56ba25),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00cb51),
	.w1(32'hb9e9eb1e),
	.w2(32'hbb9d7344),
	.w3(32'h3a68a1a1),
	.w4(32'h3bf7f3f5),
	.w5(32'h3c001035),
	.w6(32'hbbbcc2e3),
	.w7(32'hbc36ecd9),
	.w8(32'hbb664e73),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11cc2a),
	.w1(32'h3b698f56),
	.w2(32'hbbfcbd0e),
	.w3(32'hba4e65f6),
	.w4(32'h3ca18f2a),
	.w5(32'h3b81eeb5),
	.w6(32'h3b2c00ec),
	.w7(32'hbb9defe6),
	.w8(32'hba200a53),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2932ee),
	.w1(32'hbae36427),
	.w2(32'h3aeb32ba),
	.w3(32'hbba4f09d),
	.w4(32'hba9ad304),
	.w5(32'h3aac080e),
	.w6(32'hba208d19),
	.w7(32'hbbaa415c),
	.w8(32'h366a1ed8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb34ea2),
	.w1(32'hbbd33888),
	.w2(32'h3b306cae),
	.w3(32'h3c5e8d3a),
	.w4(32'h3bc63d90),
	.w5(32'h3bdca278),
	.w6(32'hbbd0ad0e),
	.w7(32'hbbd71fbf),
	.w8(32'hbc2c03a2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf53b94),
	.w1(32'h3a8b9864),
	.w2(32'h3bf7c5f8),
	.w3(32'h3b89fd34),
	.w4(32'hbc071c4c),
	.w5(32'h3a44ef00),
	.w6(32'h3c3192e2),
	.w7(32'h3c3e43b5),
	.w8(32'h39cfa3a5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8302f),
	.w1(32'h3bb80d3f),
	.w2(32'h3c99056c),
	.w3(32'h3aab6989),
	.w4(32'h3c3194f0),
	.w5(32'h3c91afab),
	.w6(32'h39fe661c),
	.w7(32'h3beb12b3),
	.w8(32'hba9c5516),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90fef58),
	.w1(32'h3b3eb5e2),
	.w2(32'h3bdd33ef),
	.w3(32'hbb211eff),
	.w4(32'h3b9c7510),
	.w5(32'h3bf66510),
	.w6(32'h3b3d880e),
	.w7(32'h3b8787ee),
	.w8(32'h3b24fd9b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0ddb2),
	.w1(32'h3ab8c511),
	.w2(32'h3ac53ccc),
	.w3(32'h3becabb5),
	.w4(32'h3b9324d8),
	.w5(32'h3bf431f4),
	.w6(32'h3aaf874a),
	.w7(32'hbab14c52),
	.w8(32'h39f35153),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bf2e4),
	.w1(32'hbb5d9a8e),
	.w2(32'hbc32dfa8),
	.w3(32'h3c1c8372),
	.w4(32'hba71df04),
	.w5(32'hbb83e373),
	.w6(32'hbb6253f6),
	.w7(32'hbb9a3e57),
	.w8(32'hbbc720aa),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc319b1b),
	.w1(32'h3c103d44),
	.w2(32'h3d0132e1),
	.w3(32'hbc0a21f7),
	.w4(32'h3c245adb),
	.w5(32'h3d1703b3),
	.w6(32'hbb087773),
	.w7(32'h3c447c53),
	.w8(32'h3c096ee8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f8862),
	.w1(32'hbacddb08),
	.w2(32'h3ae66354),
	.w3(32'h3cc92b48),
	.w4(32'hbb1b7978),
	.w5(32'hb95b6f33),
	.w6(32'hb985919d),
	.w7(32'h3ac9813a),
	.w8(32'h3a925c17),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac45105),
	.w1(32'hbbddf6ab),
	.w2(32'hbb07c530),
	.w3(32'hba0a3ccd),
	.w4(32'hbb87d16a),
	.w5(32'h3c1425e0),
	.w6(32'hba8e53eb),
	.w7(32'hbc6a4384),
	.w8(32'hbc42e6a9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977c5d),
	.w1(32'h3ba98aa8),
	.w2(32'h3b9570f7),
	.w3(32'h3aec96ac),
	.w4(32'h3c099820),
	.w5(32'h3c19908f),
	.w6(32'h3b1eca88),
	.w7(32'h3a9694a4),
	.w8(32'hba947159),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f6962),
	.w1(32'hbb38febc),
	.w2(32'h3aaba7df),
	.w3(32'h3bed4b18),
	.w4(32'h3c011bb9),
	.w5(32'h3c02cd53),
	.w6(32'h3be0d92a),
	.w7(32'hba3da7e2),
	.w8(32'h3ac1160b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadabfa1),
	.w1(32'h3b1b2b30),
	.w2(32'h3c13eb33),
	.w3(32'hb91f4393),
	.w4(32'h3bbb33c6),
	.w5(32'h3bdffd7c),
	.w6(32'h39209149),
	.w7(32'hbaa77ae4),
	.w8(32'h3a1e68ae),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb5f56),
	.w1(32'hbb1ca297),
	.w2(32'h39e7c9ec),
	.w3(32'h3ba52426),
	.w4(32'hbaedf9e3),
	.w5(32'h3aa6e3b2),
	.w6(32'hbb46a836),
	.w7(32'hbb953c2b),
	.w8(32'hbbb6f069),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0566e5),
	.w1(32'hbb25f0bd),
	.w2(32'hbb19b079),
	.w3(32'hbabb64ea),
	.w4(32'hbb846087),
	.w5(32'hbb956697),
	.w6(32'h3ae1f863),
	.w7(32'h3ab4e8a1),
	.w8(32'h3b37f422),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddfc3f),
	.w1(32'hbb6dd694),
	.w2(32'hbc33f450),
	.w3(32'hbb250987),
	.w4(32'h3b2fdcd6),
	.w5(32'hbbaa3cc8),
	.w6(32'hba654f7a),
	.w7(32'hbb7fbfdc),
	.w8(32'h3b71a076),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb848ef5),
	.w1(32'h3bc7d590),
	.w2(32'hbac4fb95),
	.w3(32'h3b370a61),
	.w4(32'h3c05561e),
	.w5(32'hbb1a2ef9),
	.w6(32'h3ba087d5),
	.w7(32'hbb9ae1eb),
	.w8(32'h3b923b73),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b338f),
	.w1(32'hbb4e9fb1),
	.w2(32'hbb8f95e2),
	.w3(32'h3b2362a9),
	.w4(32'h3c6c6a7c),
	.w5(32'h3c30d50d),
	.w6(32'hba976fab),
	.w7(32'hbb7c4532),
	.w8(32'h3bb83932),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc134222),
	.w1(32'hbbb3eda0),
	.w2(32'hbb84418b),
	.w3(32'h3981d2fc),
	.w4(32'hbaf9e785),
	.w5(32'h3b2cd7c8),
	.w6(32'hbb4b2e2f),
	.w7(32'hbb879b4d),
	.w8(32'hbb39e588),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba80104),
	.w1(32'hb6a3d80e),
	.w2(32'h3a8d2fc7),
	.w3(32'h3aa278ac),
	.w4(32'h3be4667e),
	.w5(32'h3aca26f9),
	.w6(32'hbbd55440),
	.w7(32'h3bc1cbda),
	.w8(32'hbb0764f0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc610eba),
	.w1(32'hbbe9c55b),
	.w2(32'hbc24277e),
	.w3(32'hbbf57f2c),
	.w4(32'hbbe4b30d),
	.w5(32'hbc26f499),
	.w6(32'hbc4ae312),
	.w7(32'hbc6a7404),
	.w8(32'hbb13461a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0dd18),
	.w1(32'h3bbc7705),
	.w2(32'h3c1beb57),
	.w3(32'hbc032106),
	.w4(32'h3bd64f37),
	.w5(32'h3c3540af),
	.w6(32'h3a87b568),
	.w7(32'h3a9f7ef0),
	.w8(32'h3aa98a8e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea5f71),
	.w1(32'h3b19d906),
	.w2(32'hbb3d3987),
	.w3(32'h3c1739df),
	.w4(32'h3bd8daab),
	.w5(32'hbb3c411c),
	.w6(32'h3b886e81),
	.w7(32'hbb919feb),
	.w8(32'h3c09536e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae131bd),
	.w1(32'h3be226c0),
	.w2(32'hbb7198ac),
	.w3(32'h3bdb2426),
	.w4(32'h3be065fe),
	.w5(32'h3990930c),
	.w6(32'hba7a0a6e),
	.w7(32'hba96915c),
	.w8(32'hbbb7c2b0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a349f),
	.w1(32'hbbcfdf09),
	.w2(32'hba595b28),
	.w3(32'hbc0c1867),
	.w4(32'hbba80670),
	.w5(32'h3b0129c3),
	.w6(32'hbb6b3003),
	.w7(32'hba7a9dab),
	.w8(32'hbbd78146),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f8d82),
	.w1(32'hbac01cec),
	.w2(32'hbb88d590),
	.w3(32'hba636f65),
	.w4(32'h39739246),
	.w5(32'hba4168a2),
	.w6(32'h39d4f6cf),
	.w7(32'hbb57641b),
	.w8(32'h3a9ae896),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b4cd0),
	.w1(32'hbc46020f),
	.w2(32'hbd0152b3),
	.w3(32'h3a5d8463),
	.w4(32'hbc56b8e6),
	.w5(32'hbced9a35),
	.w6(32'hbc82b1a6),
	.w7(32'hbd14a0b7),
	.w8(32'hbcfec7bf),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule