module layer_8_featuremap_87(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17c9c6),
	.w1(32'h3d0144a5),
	.w2(32'hbc3424e8),
	.w3(32'h3b379da7),
	.w4(32'h3cc6a97c),
	.w5(32'hbd3b94b3),
	.w6(32'h3ab83309),
	.w7(32'h3c27f78f),
	.w8(32'h3d2af6ad),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd52a46d),
	.w1(32'h3c4917fa),
	.w2(32'h3cb8cf03),
	.w3(32'h3bed70e1),
	.w4(32'h3c80b3f6),
	.w5(32'hbc036964),
	.w6(32'hbc0dd66f),
	.w7(32'h3c3f4466),
	.w8(32'h3c7d3a1d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3cabad),
	.w1(32'hbcb1de14),
	.w2(32'hbd000276),
	.w3(32'h3d0151fa),
	.w4(32'h3c946786),
	.w5(32'hbd143d33),
	.w6(32'hbbeeab70),
	.w7(32'hbc02da1f),
	.w8(32'h3cfdeca5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b928fd2),
	.w1(32'hbc423588),
	.w2(32'hbd890dcc),
	.w3(32'h3c2db42d),
	.w4(32'hba1190f0),
	.w5(32'hbd5a6656),
	.w6(32'h3d2da9d5),
	.w7(32'hbc4f21a9),
	.w8(32'h3ce0a41a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccea6c2),
	.w1(32'hbca054e0),
	.w2(32'hbd00a3eb),
	.w3(32'h3cc2f989),
	.w4(32'h3c901264),
	.w5(32'h3c720b60),
	.w6(32'h3b9a258f),
	.w7(32'h3d2a3bf5),
	.w8(32'hbc1d1479),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd897b5b),
	.w1(32'h3cc67aa5),
	.w2(32'hbcf217f0),
	.w3(32'h3d9191a5),
	.w4(32'h3aa36230),
	.w5(32'hbc86780a),
	.w6(32'hbbfe4482),
	.w7(32'h3b6240f8),
	.w8(32'hbc710406),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdaf642),
	.w1(32'h3ab7b19f),
	.w2(32'hbb684150),
	.w3(32'hbe3491ab),
	.w4(32'hbd275e29),
	.w5(32'h3c191ee9),
	.w6(32'h3c1ecf96),
	.w7(32'hbd49a269),
	.w8(32'hbc7395b3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e8733),
	.w1(32'hbc05f9ee),
	.w2(32'hbd09215c),
	.w3(32'h3c199ae5),
	.w4(32'h3bf6d47e),
	.w5(32'h3b9e92a7),
	.w6(32'h3d005c92),
	.w7(32'h3d3510a1),
	.w8(32'hbb33356a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e2f23),
	.w1(32'hbd0b3a64),
	.w2(32'h3897105f),
	.w3(32'hbb3582ec),
	.w4(32'hbd06c02a),
	.w5(32'hbcb26527),
	.w6(32'h3c4158b7),
	.w7(32'h3c8cfd5a),
	.w8(32'hbd8c5272),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80b18f),
	.w1(32'hbd1287d3),
	.w2(32'h3c3a4c83),
	.w3(32'hbc9f6bad),
	.w4(32'h3d0240f4),
	.w5(32'h3c4731c3),
	.w6(32'hbcb11f0d),
	.w7(32'hbcde9706),
	.w8(32'hbb846529),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c408c38),
	.w1(32'h3bd0c8af),
	.w2(32'hbb1ace2b),
	.w3(32'h3b7e6e99),
	.w4(32'h3c89f971),
	.w5(32'h3b9c389c),
	.w6(32'hbc657b54),
	.w7(32'h3bb0e1cf),
	.w8(32'h3c24ec0d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e9768),
	.w1(32'h3ca18ab3),
	.w2(32'h3a41a29c),
	.w3(32'h3c86e433),
	.w4(32'h3c484169),
	.w5(32'h3cf05716),
	.w6(32'h3c569ebd),
	.w7(32'hbb6c834b),
	.w8(32'hbc93dad6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f6e30),
	.w1(32'hbd37b27c),
	.w2(32'h3b511c9f),
	.w3(32'h3ba2e8df),
	.w4(32'h3c4b1c2f),
	.w5(32'hbbd7ecfa),
	.w6(32'h3c953be1),
	.w7(32'hbb9f4e50),
	.w8(32'h3c8b47ba),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f0efd),
	.w1(32'hbbfd6695),
	.w2(32'hbce74c52),
	.w3(32'h3b03977e),
	.w4(32'hbba1b384),
	.w5(32'hbd052e96),
	.w6(32'hbd0a0264),
	.w7(32'hbc0c3ad7),
	.w8(32'hbcba280c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd372d26),
	.w1(32'hbc9c45d6),
	.w2(32'h3bf09fd4),
	.w3(32'h3c5c480e),
	.w4(32'hbc9603a2),
	.w5(32'hbbd113c3),
	.w6(32'hbac31521),
	.w7(32'hbc988860),
	.w8(32'hbc793531),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ef501),
	.w1(32'h3c34fc95),
	.w2(32'h3cba5ea7),
	.w3(32'h3cabc593),
	.w4(32'h3da2ae9a),
	.w5(32'hbc067d8c),
	.w6(32'hba5f06fe),
	.w7(32'hbc8e63e8),
	.w8(32'h3c56bbb3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ee4cd),
	.w1(32'h3b7cadec),
	.w2(32'h3ad755d1),
	.w3(32'h3c4ac5a7),
	.w4(32'hbbdf5f6a),
	.w5(32'h3bb1dd6f),
	.w6(32'hbbd811d7),
	.w7(32'h3bc266ba),
	.w8(32'hbc6ff549),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8d0a4),
	.w1(32'hbba8fa76),
	.w2(32'hbbf2a209),
	.w3(32'hbba4ec75),
	.w4(32'hbc9f7216),
	.w5(32'h3bf5b8bc),
	.w6(32'h3b9f3f05),
	.w7(32'h3bd1623d),
	.w8(32'h3c87e6bd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1d20d),
	.w1(32'hbbda5c4d),
	.w2(32'hbb32b038),
	.w3(32'h3cc91c8b),
	.w4(32'hbc232f0e),
	.w5(32'hbb286290),
	.w6(32'h3cc5a57c),
	.w7(32'hbc4e5cdb),
	.w8(32'hbc890eca),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b176ff8),
	.w1(32'h3c8ed0ca),
	.w2(32'hbbd7fc18),
	.w3(32'hbc3c9e58),
	.w4(32'hbcb9a53e),
	.w5(32'hbb2b0dd1),
	.w6(32'hbc380359),
	.w7(32'h3933d9df),
	.w8(32'h3ab726ab),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd18e58e),
	.w1(32'h3bedefe0),
	.w2(32'hbc4ec553),
	.w3(32'h3d251332),
	.w4(32'hbc0d9571),
	.w5(32'h3b889f04),
	.w6(32'h3b90fa87),
	.w7(32'h3c14748c),
	.w8(32'hbb99e2e0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90ce70),
	.w1(32'hbbdf95eb),
	.w2(32'h3c06f770),
	.w3(32'hbba3bd04),
	.w4(32'hb9e3d65d),
	.w5(32'h3d04e50d),
	.w6(32'hbc07af0c),
	.w7(32'h3b9f6c50),
	.w8(32'hbc181094),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9063e6),
	.w1(32'h3b97a79f),
	.w2(32'hbb405577),
	.w3(32'hbc8ed7ac),
	.w4(32'hbba8233d),
	.w5(32'h3a1690eb),
	.w6(32'hbc26ec8b),
	.w7(32'h3c7b1b8d),
	.w8(32'hbc47c12a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92d583),
	.w1(32'h3c8a3eee),
	.w2(32'hbc315a6d),
	.w3(32'hbcf9963a),
	.w4(32'hbb0f5de4),
	.w5(32'hbb97897c),
	.w6(32'hbb72a8d2),
	.w7(32'hbcb21f3b),
	.w8(32'hbd56bf36),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8032e8),
	.w1(32'hbbbea9d0),
	.w2(32'h3ca42ea7),
	.w3(32'hb815aa1a),
	.w4(32'h3c566b0d),
	.w5(32'hba1688eb),
	.w6(32'hbbf090bd),
	.w7(32'hbc291f8b),
	.w8(32'hbb95d3cf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb468404),
	.w1(32'hbc0036a0),
	.w2(32'h3c456df3),
	.w3(32'h3c210e2e),
	.w4(32'hbba6d77f),
	.w5(32'hbb943264),
	.w6(32'h3c80b454),
	.w7(32'h3c0dd954),
	.w8(32'h3ce64916),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad78e8d),
	.w1(32'h3c042ea0),
	.w2(32'h3badcb93),
	.w3(32'hbc7d0809),
	.w4(32'hbd1aaa2b),
	.w5(32'hbc898ea1),
	.w6(32'h3b30278d),
	.w7(32'hbb4bff0f),
	.w8(32'h3c84b16e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90cf13),
	.w1(32'hbb26079d),
	.w2(32'hbc594e64),
	.w3(32'h3c55d095),
	.w4(32'hbc0579e0),
	.w5(32'h3c5aef8b),
	.w6(32'hbb04afd0),
	.w7(32'hbc05318b),
	.w8(32'hbdc8c279),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d28ebf7),
	.w1(32'h3c18c605),
	.w2(32'hbc77bb63),
	.w3(32'hbb96f073),
	.w4(32'h3b0175c0),
	.w5(32'h3c1584c0),
	.w6(32'hbd7fb5db),
	.w7(32'hbb813a15),
	.w8(32'hbc1f3924),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242e8c),
	.w1(32'h3c11ff63),
	.w2(32'hbcbcbc63),
	.w3(32'h3d1bd055),
	.w4(32'hbc5bb927),
	.w5(32'hbcbe0c0a),
	.w6(32'hbbf9a3db),
	.w7(32'hbb30f646),
	.w8(32'hbb2d4521),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b4fb9),
	.w1(32'h3cf29620),
	.w2(32'hbd487212),
	.w3(32'h3d2e2151),
	.w4(32'hbcef7f3f),
	.w5(32'h3a327968),
	.w6(32'hbdc2a81d),
	.w7(32'hbb9021b7),
	.w8(32'hbb39baee),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d9818),
	.w1(32'hbbc42430),
	.w2(32'hbc887f0d),
	.w3(32'h3b069f6f),
	.w4(32'h3b561613),
	.w5(32'h3bcb80b8),
	.w6(32'hbc8dfdff),
	.w7(32'hbca1fd10),
	.w8(32'h3b85ff31),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5568ab),
	.w1(32'hbc90fa66),
	.w2(32'hbb6873e8),
	.w3(32'h3b46db84),
	.w4(32'h3ccd7d82),
	.w5(32'h3bd11a46),
	.w6(32'hbc776670),
	.w7(32'hbd09862f),
	.w8(32'hbbca243b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc628f),
	.w1(32'hbc3c83e7),
	.w2(32'h3d41eb69),
	.w3(32'h3aaa8088),
	.w4(32'h3c053251),
	.w5(32'hbc02246e),
	.w6(32'h3c3339e8),
	.w7(32'h3d26b874),
	.w8(32'h3c86228d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46388d),
	.w1(32'h3c0f2c75),
	.w2(32'hbc417a72),
	.w3(32'hbc0faf58),
	.w4(32'hbbcb699f),
	.w5(32'hbc2fb683),
	.w6(32'h3cab0557),
	.w7(32'hbbff41f4),
	.w8(32'h3c30afc0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2753b0),
	.w1(32'hbd492a73),
	.w2(32'h3b67efcc),
	.w3(32'h3c41d53c),
	.w4(32'hbc63a5be),
	.w5(32'h3c8b1c7e),
	.w6(32'h3bd91ea4),
	.w7(32'hbd9cb09b),
	.w8(32'hbc346522),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77a8e2),
	.w1(32'h391a1b68),
	.w2(32'hbd852b70),
	.w3(32'hbc7230b4),
	.w4(32'hbd212f2b),
	.w5(32'hbc9a1b44),
	.w6(32'hbc883980),
	.w7(32'hbc4092de),
	.w8(32'h3bf8d842),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe24dc4),
	.w1(32'hbd1d5cb9),
	.w2(32'hbc0b9f6b),
	.w3(32'hbc0e7c2a),
	.w4(32'hbcc0ce30),
	.w5(32'hbb9ceec1),
	.w6(32'h3c377d73),
	.w7(32'hbd14ae97),
	.w8(32'hbc1730f4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce09735),
	.w1(32'h3cbbfa8f),
	.w2(32'hbdcab664),
	.w3(32'hbc030a16),
	.w4(32'hbbd97030),
	.w5(32'h3c665f6e),
	.w6(32'hbb2f5e4a),
	.w7(32'hb8f4b2d0),
	.w8(32'h3c164597),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae03d2f),
	.w1(32'h3a7c7ca6),
	.w2(32'hbba57926),
	.w3(32'h3b8869c4),
	.w4(32'hbb34ec2e),
	.w5(32'h3d8d777a),
	.w6(32'h3cc28472),
	.w7(32'hbd70c77a),
	.w8(32'hbaa44f2f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9294905),
	.w1(32'hbc6c5ad1),
	.w2(32'hbb849c3d),
	.w3(32'h3c43e7c6),
	.w4(32'h3c86d04e),
	.w5(32'hbc1bd865),
	.w6(32'hba6ad761),
	.w7(32'h3b16aa4e),
	.w8(32'hba700146),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc808a7),
	.w1(32'h3bb9479b),
	.w2(32'hbca2d511),
	.w3(32'h3d125a7b),
	.w4(32'hbd388806),
	.w5(32'hbbc93ec4),
	.w6(32'h3b6cde00),
	.w7(32'hbbaa70f0),
	.w8(32'hbba3296c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb732cec),
	.w1(32'hbc50c336),
	.w2(32'h3a0524c4),
	.w3(32'hbcda91ea),
	.w4(32'hbd2ad47f),
	.w5(32'hbcad0ab8),
	.w6(32'hbc06ffb5),
	.w7(32'h3d3fb50b),
	.w8(32'hbd19a2f6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f8fb2),
	.w1(32'h3cad1565),
	.w2(32'hbcfbaccf),
	.w3(32'h3b854c14),
	.w4(32'hbcd24929),
	.w5(32'h3c6f6e9c),
	.w6(32'hbc1ab6aa),
	.w7(32'hbcf3998a),
	.w8(32'h3c7cc9f2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab79e19),
	.w1(32'h3c160ae8),
	.w2(32'hbb8f4750),
	.w3(32'hbc285584),
	.w4(32'h3c4b4829),
	.w5(32'h3d43f633),
	.w6(32'h3a7a137e),
	.w7(32'hbc242c40),
	.w8(32'hbb54f526),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd213486),
	.w1(32'hbcae5580),
	.w2(32'hbc3ca1ce),
	.w3(32'hbc862baf),
	.w4(32'hbcfa56dd),
	.w5(32'h3c53f16e),
	.w6(32'hbc48326e),
	.w7(32'hbb788295),
	.w8(32'hbc2aa51e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb150352),
	.w1(32'hbd72537c),
	.w2(32'hbbc5c75e),
	.w3(32'hba79bdb8),
	.w4(32'hbd4641dd),
	.w5(32'h3b6c6b27),
	.w6(32'hbc860501),
	.w7(32'h3ca97286),
	.w8(32'h3b61ede4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7b292),
	.w1(32'hbacb9b29),
	.w2(32'hbd0d720f),
	.w3(32'h3d622a96),
	.w4(32'hbc86df13),
	.w5(32'hbcdd4df3),
	.w6(32'h3b0d341b),
	.w7(32'h3c043508),
	.w8(32'hbc7e2b8b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc921298),
	.w1(32'hbcbb042c),
	.w2(32'h3ca4cf4e),
	.w3(32'h3c33ec50),
	.w4(32'h3b9c97dd),
	.w5(32'hbc98815e),
	.w6(32'h3bf49cc4),
	.w7(32'hbcc59c17),
	.w8(32'hbca2c90c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2efbf),
	.w1(32'hbcb4a703),
	.w2(32'h3a899387),
	.w3(32'hbca1f498),
	.w4(32'hbc4e30a8),
	.w5(32'h3d0ddf3a),
	.w6(32'hbd331ed5),
	.w7(32'hbc403ea0),
	.w8(32'h39d41735),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e4009),
	.w1(32'hbc43c1b8),
	.w2(32'hbc8d7f4d),
	.w3(32'h3c04a80d),
	.w4(32'h3d7433cb),
	.w5(32'hbc230595),
	.w6(32'hbb8228ff),
	.w7(32'hba922276),
	.w8(32'hbbd0417b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08b81a),
	.w1(32'hbbb747c8),
	.w2(32'hbc023a9a),
	.w3(32'hbc09e1da),
	.w4(32'hb739fd15),
	.w5(32'hbc5e8535),
	.w6(32'h3d676a95),
	.w7(32'h3b469756),
	.w8(32'hbc616487),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc9f823),
	.w1(32'h3b79a2fb),
	.w2(32'hbc5a08a1),
	.w3(32'hbd3f9442),
	.w4(32'h3d03911a),
	.w5(32'h3a2e8ee5),
	.w6(32'hba88acc1),
	.w7(32'h3c159751),
	.w8(32'h3ccf6cc1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68b59a),
	.w1(32'h3c0e888d),
	.w2(32'h3b8d6781),
	.w3(32'h3b75dcf1),
	.w4(32'hb9bca2d8),
	.w5(32'hbaf5c033),
	.w6(32'hbbd2fc87),
	.w7(32'hbc3a9a25),
	.w8(32'h3a1bd914),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad97f29),
	.w1(32'hbd23ea47),
	.w2(32'h3baf41b9),
	.w3(32'h3b708a78),
	.w4(32'h3c82100f),
	.w5(32'hbc3b7cbb),
	.w6(32'h3c6e7cd5),
	.w7(32'h3d0bcacd),
	.w8(32'h3cae3465),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4a8d76),
	.w1(32'hbc97272f),
	.w2(32'hbc707b72),
	.w3(32'hba969ae3),
	.w4(32'h3b0ca02f),
	.w5(32'h3b49c2e0),
	.w6(32'h3cd51c55),
	.w7(32'hbd5dd96b),
	.w8(32'hbbe6cef2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d166721),
	.w1(32'h3d26a716),
	.w2(32'hbd805342),
	.w3(32'hbb8bea05),
	.w4(32'hbc57edb8),
	.w5(32'hbd375ef1),
	.w6(32'h3c161f23),
	.w7(32'h3c155726),
	.w8(32'h3c33f4d0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92a07c),
	.w1(32'hbcbb6c7f),
	.w2(32'hbbd9b551),
	.w3(32'h3c1258e1),
	.w4(32'hbc2f9144),
	.w5(32'hbd86ef9f),
	.w6(32'hbd3eb910),
	.w7(32'hbc343ff9),
	.w8(32'hbc856856),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95724a4),
	.w1(32'h3ca179cb),
	.w2(32'hbcd1a1d0),
	.w3(32'h3c79a35b),
	.w4(32'hbb38ea66),
	.w5(32'hbe005acc),
	.w6(32'h3c0921ad),
	.w7(32'h3cfbb56e),
	.w8(32'h3ca06bbb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b799c),
	.w1(32'h3cc3ccb7),
	.w2(32'h3b19e602),
	.w3(32'h3c10af0d),
	.w4(32'h3c96e407),
	.w5(32'hbbbced08),
	.w6(32'hbc0802f3),
	.w7(32'hbb6b1986),
	.w8(32'h3b11e267),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53ef25),
	.w1(32'h3bda8206),
	.w2(32'hbbed165e),
	.w3(32'hbc25a8b7),
	.w4(32'hbaf84617),
	.w5(32'hbbb568a3),
	.w6(32'hbcc153cb),
	.w7(32'hbc43e147),
	.w8(32'h3b89c247),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d261d55),
	.w1(32'h3c847e8a),
	.w2(32'h3cae828b),
	.w3(32'hba17eaf4),
	.w4(32'hbcdd934d),
	.w5(32'hbbb11130),
	.w6(32'hbbb34871),
	.w7(32'hba337a45),
	.w8(32'hbcc3abb4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d51054d),
	.w1(32'hbb1e7020),
	.w2(32'hbce4005a),
	.w3(32'h3d3160b2),
	.w4(32'hbb04a08f),
	.w5(32'hbcddda93),
	.w6(32'hb94e16e9),
	.w7(32'hbc2a73ed),
	.w8(32'h3bb4a624),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d92f44c),
	.w1(32'hbc0c6361),
	.w2(32'hbd3f53b8),
	.w3(32'h3cead10c),
	.w4(32'h3ab7d81d),
	.w5(32'h3c3a421e),
	.w6(32'hbc2fc2d7),
	.w7(32'h3c27329c),
	.w8(32'h3cbe78ec),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd16c6),
	.w1(32'hbc51b841),
	.w2(32'hbc03b513),
	.w3(32'hbc161276),
	.w4(32'h3d0c39a0),
	.w5(32'hbc8c6db3),
	.w6(32'h3cf0a66b),
	.w7(32'hbb1b61dd),
	.w8(32'h3cf859bd),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a32aa),
	.w1(32'hbc037c34),
	.w2(32'h3c72720e),
	.w3(32'h3c35a6a8),
	.w4(32'h3b5e8870),
	.w5(32'hbbc6a8d3),
	.w6(32'hbdde8938),
	.w7(32'h3c477021),
	.w8(32'h3c8d99b2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd004ae0),
	.w1(32'hbdb66b9f),
	.w2(32'hbc915568),
	.w3(32'hbbc0acf3),
	.w4(32'h3cb71199),
	.w5(32'h3be9bfbb),
	.w6(32'hbcdcec21),
	.w7(32'h3c84bcc2),
	.w8(32'hbca177f3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48e0b2),
	.w1(32'h3d0b3916),
	.w2(32'h3c927bf2),
	.w3(32'hbb403e7d),
	.w4(32'h3bbc0779),
	.w5(32'h3be08d28),
	.w6(32'hbc672744),
	.w7(32'hbc222171),
	.w8(32'hbd40f6be),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c864fca),
	.w1(32'h3a53dea3),
	.w2(32'hbcb40bfa),
	.w3(32'h3b5ec13c),
	.w4(32'hbc478a01),
	.w5(32'hbdcc78f4),
	.w6(32'hbc9159fc),
	.w7(32'h3d09bd71),
	.w8(32'h3c121f9c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2eb3a),
	.w1(32'h3bc18c25),
	.w2(32'hbb1b107c),
	.w3(32'hbc994dec),
	.w4(32'hbc28d76d),
	.w5(32'hbb2d632f),
	.w6(32'hbcd8be54),
	.w7(32'h3a81e075),
	.w8(32'h3950ce93),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4acd73),
	.w1(32'hbb5be53f),
	.w2(32'hbb0b80ca),
	.w3(32'h3aa4929d),
	.w4(32'hbc3735ab),
	.w5(32'h3cc3aa53),
	.w6(32'h3a792d77),
	.w7(32'h3bdaf5a7),
	.w8(32'hbc837f0b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6ad86),
	.w1(32'hba8dac73),
	.w2(32'hbbc98e9c),
	.w3(32'hbc212ad7),
	.w4(32'hba913501),
	.w5(32'h3a9ef817),
	.w6(32'hb8fe9228),
	.w7(32'hbc26d111),
	.w8(32'hbca10b68),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7d120),
	.w1(32'hbac3aaeb),
	.w2(32'h3b04cd09),
	.w3(32'hbca78bf4),
	.w4(32'h3b8f9a43),
	.w5(32'h3cc93b72),
	.w6(32'hbb396d61),
	.w7(32'h3acb0209),
	.w8(32'h3b030492),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0982),
	.w1(32'hbb04346a),
	.w2(32'hbcaaa5ba),
	.w3(32'h3bd6b110),
	.w4(32'hbbe606cf),
	.w5(32'hbbb852fc),
	.w6(32'hbc1a193b),
	.w7(32'hbae748b0),
	.w8(32'hbbad27b7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd14285),
	.w1(32'h3a2720fb),
	.w2(32'hbabd64e3),
	.w3(32'hbc3d000f),
	.w4(32'h3c59942c),
	.w5(32'hbc90cbec),
	.w6(32'hbaaab636),
	.w7(32'h3c23e221),
	.w8(32'hbc3cbc09),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4028c6),
	.w1(32'hbb00fbc2),
	.w2(32'hbc26f8a4),
	.w3(32'h3d3f2564),
	.w4(32'hbbd3c93d),
	.w5(32'h3c0a0a72),
	.w6(32'h3c4a4b44),
	.w7(32'h3b41c641),
	.w8(32'hb9df4b75),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9461c),
	.w1(32'hbb1309d0),
	.w2(32'h398e2589),
	.w3(32'hbc8ea2f7),
	.w4(32'h39a08df7),
	.w5(32'hbbddeea3),
	.w6(32'hb9567874),
	.w7(32'h3d81c812),
	.w8(32'h3b2ed3ea),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b9dbc),
	.w1(32'h3b639e1c),
	.w2(32'hbba21c9c),
	.w3(32'hbc9c1b6d),
	.w4(32'hbbea49ce),
	.w5(32'h3ba22218),
	.w6(32'h3b8dff89),
	.w7(32'hbc2bc5a9),
	.w8(32'hbb3528ff),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66fda2),
	.w1(32'hbbbdb4dd),
	.w2(32'h3c7b2a3b),
	.w3(32'hbb991d80),
	.w4(32'h3bed2913),
	.w5(32'h3c4a1851),
	.w6(32'hbbfbe3b7),
	.w7(32'hbccc83c9),
	.w8(32'h3bc3f163),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07b1c9),
	.w1(32'hbbe2bc56),
	.w2(32'hbbeb3f85),
	.w3(32'h3b8574d0),
	.w4(32'h3bce19c0),
	.w5(32'h3b5d1534),
	.w6(32'h3b3ef876),
	.w7(32'hbc31abc4),
	.w8(32'hba7dd826),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02fc96),
	.w1(32'hbb0bdd2d),
	.w2(32'hbb1d70f8),
	.w3(32'h383f20ea),
	.w4(32'hba95384f),
	.w5(32'hbcacd688),
	.w6(32'h3bd678c5),
	.w7(32'hbbf7952a),
	.w8(32'hbca95802),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b859f9e),
	.w1(32'h3b8c8ec4),
	.w2(32'hbba90088),
	.w3(32'h3ba1ee91),
	.w4(32'h39ffadf8),
	.w5(32'hbc0316f8),
	.w6(32'h3be1bc63),
	.w7(32'hbbfe6a98),
	.w8(32'h3bec6647),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2af8d0),
	.w1(32'hbaf23cd0),
	.w2(32'h3b339b21),
	.w3(32'h3c1f0de1),
	.w4(32'hbbf3677b),
	.w5(32'hbb886ca0),
	.w6(32'hbba8a2bb),
	.w7(32'hbcb458a5),
	.w8(32'hbcb3de83),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e4dd6),
	.w1(32'h3becb572),
	.w2(32'hbb578163),
	.w3(32'h3ab0adbf),
	.w4(32'hbcbb6643),
	.w5(32'h3b88f9ac),
	.w6(32'hbd11a33e),
	.w7(32'h3adf021d),
	.w8(32'h3ab1f1b8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3c42a1),
	.w1(32'h3b5df604),
	.w2(32'hbc78b716),
	.w3(32'h3bb5b8d8),
	.w4(32'h3caeecd8),
	.w5(32'h3d45db2b),
	.w6(32'h3c979e96),
	.w7(32'h3c7358db),
	.w8(32'h3d081ecd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94c564),
	.w1(32'h3bf2ad79),
	.w2(32'h3c5a6ba5),
	.w3(32'hbd69c4f8),
	.w4(32'hbc25a189),
	.w5(32'h3c22df4a),
	.w6(32'h3b5f87aa),
	.w7(32'h3adc11a4),
	.w8(32'hbc8ac918),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d831b),
	.w1(32'hbb46bc0b),
	.w2(32'hbc926c68),
	.w3(32'h3b807b0a),
	.w4(32'h3ba9dc57),
	.w5(32'h38f228e5),
	.w6(32'hbc880360),
	.w7(32'hbc5ac2c9),
	.w8(32'hbb389be4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1df8b1),
	.w1(32'hbd2aac5f),
	.w2(32'h3c98eb2d),
	.w3(32'h3cbe66b6),
	.w4(32'hbb841225),
	.w5(32'hbc101bcf),
	.w6(32'hbd7e2cfc),
	.w7(32'h3cde4633),
	.w8(32'h3bae977b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be899db),
	.w1(32'h3b8860e6),
	.w2(32'h3b8902d3),
	.w3(32'hbc03b094),
	.w4(32'hbc8481df),
	.w5(32'hbb9f9186),
	.w6(32'hbcb34e21),
	.w7(32'h3bb27cb7),
	.w8(32'h3d0966eb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2c676),
	.w1(32'hbb9249c2),
	.w2(32'hbccddc53),
	.w3(32'h3ba26984),
	.w4(32'hbcb8245f),
	.w5(32'hbc4321c6),
	.w6(32'h3b28ff5f),
	.w7(32'hbc8eee8c),
	.w8(32'h3bb35af1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08d077),
	.w1(32'h3b9a2ae8),
	.w2(32'hbd059044),
	.w3(32'h3bc97d22),
	.w4(32'hbdb668f3),
	.w5(32'hbc154e35),
	.w6(32'hbbf1948f),
	.w7(32'h3c130c40),
	.w8(32'h3b803196),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc272183),
	.w1(32'hb971f6c8),
	.w2(32'h3bfc931a),
	.w3(32'hbc43d228),
	.w4(32'h3d362516),
	.w5(32'h3d34692e),
	.w6(32'hbc6a6fb4),
	.w7(32'hbc539069),
	.w8(32'h3ccab8d7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a90ac),
	.w1(32'hbc188953),
	.w2(32'h3bb0c1b5),
	.w3(32'hbaf632a2),
	.w4(32'h39850b4b),
	.w5(32'hbb935f35),
	.w6(32'h3c20a2f8),
	.w7(32'h3bafe91c),
	.w8(32'hbd1a2928),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd3e1e),
	.w1(32'hbc3ffc8e),
	.w2(32'h3d29b716),
	.w3(32'h3d2584ad),
	.w4(32'h3b9b406c),
	.w5(32'h3d171427),
	.w6(32'h3c8da881),
	.w7(32'hbc8e6bb9),
	.w8(32'h3b0e8181),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc568480),
	.w1(32'hbc0c0498),
	.w2(32'h3c26a8f0),
	.w3(32'h3c9e9c09),
	.w4(32'h3c096cba),
	.w5(32'hbcdef6ca),
	.w6(32'h3c85ec89),
	.w7(32'h37db4fcc),
	.w8(32'h3ce3d9ee),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be444d5),
	.w1(32'h3ae1be4c),
	.w2(32'hbce3dcea),
	.w3(32'h3d0aab6f),
	.w4(32'h3bb03869),
	.w5(32'h3cedc147),
	.w6(32'hbb7bb4f4),
	.w7(32'h3c30aba3),
	.w8(32'h3baaa41d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30702d),
	.w1(32'hbd336363),
	.w2(32'hbcbea821),
	.w3(32'h3ce886af),
	.w4(32'hbb859064),
	.w5(32'h3cb9bd6a),
	.w6(32'h3cc54b63),
	.w7(32'hbc3084a7),
	.w8(32'hbbb46557),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78e574),
	.w1(32'h3c68546f),
	.w2(32'h3d06f3d3),
	.w3(32'hbb873ab8),
	.w4(32'h3ca99f89),
	.w5(32'h3c105ee3),
	.w6(32'hbc6bc8cc),
	.w7(32'hbc6f8c04),
	.w8(32'h3c38b079),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a8e36),
	.w1(32'hbcb6709c),
	.w2(32'hbbd1b4ba),
	.w3(32'h3bd30e1b),
	.w4(32'hbaa28551),
	.w5(32'hbcbff94e),
	.w6(32'hbd8e26d8),
	.w7(32'hbc5c3972),
	.w8(32'h3c9a0578),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82df02),
	.w1(32'hbcc52d30),
	.w2(32'h3c13b5a8),
	.w3(32'h3d789c42),
	.w4(32'hbd015cb7),
	.w5(32'hbbe98110),
	.w6(32'hbaf8666b),
	.w7(32'h3a226461),
	.w8(32'h3d0d9f50),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc88810),
	.w1(32'hbc623421),
	.w2(32'hbe015782),
	.w3(32'h3a3033d1),
	.w4(32'hbd69395b),
	.w5(32'hbce2a742),
	.w6(32'h3b6f4663),
	.w7(32'h3b69b19d),
	.w8(32'hbc8d8667),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9f57f),
	.w1(32'h3c651627),
	.w2(32'hbaf34410),
	.w3(32'h3bd1733d),
	.w4(32'h3c6f3c80),
	.w5(32'h3c716a6b),
	.w6(32'h3d34fa03),
	.w7(32'hbc07bffd),
	.w8(32'hbd04fc3e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce5817),
	.w1(32'hbb39ad56),
	.w2(32'hbd224aa1),
	.w3(32'hbb72455d),
	.w4(32'h3c9f0577),
	.w5(32'h3cbb8636),
	.w6(32'h3bbdae98),
	.w7(32'hbc9dece2),
	.w8(32'hbd04a33c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e08fd),
	.w1(32'hbc155b5e),
	.w2(32'hbccb6986),
	.w3(32'hbc7f12ae),
	.w4(32'h3b9bdca5),
	.w5(32'hbb9fb78b),
	.w6(32'hbc90dcf6),
	.w7(32'h3c47800c),
	.w8(32'h3b2b8109),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb12ecd),
	.w1(32'hbcb27293),
	.w2(32'hbd23a845),
	.w3(32'h3c8926a0),
	.w4(32'h3c192c00),
	.w5(32'hbd8f236c),
	.w6(32'hbc2e5996),
	.w7(32'hbd13b675),
	.w8(32'h3c09282f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5812d3),
	.w1(32'hbcc7b616),
	.w2(32'hbcb78a7e),
	.w3(32'h3baffe72),
	.w4(32'h3bc35d89),
	.w5(32'h3bee0529),
	.w6(32'hbc585135),
	.w7(32'hbbaf1501),
	.w8(32'hbcda95cd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd39d568),
	.w1(32'h3c3e1eba),
	.w2(32'hbcbbe48f),
	.w3(32'h3c72f267),
	.w4(32'hbc3c7e56),
	.w5(32'h3c6236af),
	.w6(32'hbda46015),
	.w7(32'hbc5f2733),
	.w8(32'hbc8c7139),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49f8e4),
	.w1(32'hbd0bb73d),
	.w2(32'hbd9378ca),
	.w3(32'h3b74c751),
	.w4(32'hbcff5690),
	.w5(32'hbc315199),
	.w6(32'hbc69da3c),
	.w7(32'h3cd68f07),
	.w8(32'hbde466c8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc981281),
	.w1(32'hbc04721f),
	.w2(32'hbb9c43d2),
	.w3(32'h3b151de8),
	.w4(32'h3b8d3d9e),
	.w5(32'hbc200ca5),
	.w6(32'h3caa9858),
	.w7(32'h3c8faf56),
	.w8(32'h3b4256ba),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19cda8),
	.w1(32'hbbde2dd4),
	.w2(32'h3be066ae),
	.w3(32'hbbc33d80),
	.w4(32'hbc10bfb3),
	.w5(32'hbb9210f4),
	.w6(32'h3b7082e0),
	.w7(32'hbbe1ddb9),
	.w8(32'hbdaee3ad),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fd9f4),
	.w1(32'h3cc886a6),
	.w2(32'h3c87eb22),
	.w3(32'hba97d714),
	.w4(32'hbaef0809),
	.w5(32'h3bec23a4),
	.w6(32'hba2458df),
	.w7(32'hbd12fb26),
	.w8(32'hbcc43b4e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a337038),
	.w1(32'h3babdcf3),
	.w2(32'hbbc62e78),
	.w3(32'hbcbe9cf1),
	.w4(32'hbd214fb1),
	.w5(32'hbc69a808),
	.w6(32'hbd711ab1),
	.w7(32'h3b224282),
	.w8(32'hbcdbd95d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd7d3),
	.w1(32'hbb1cead8),
	.w2(32'hbc1b629c),
	.w3(32'hbc809771),
	.w4(32'hbc2b026d),
	.w5(32'hbaa457f2),
	.w6(32'hbbc845ce),
	.w7(32'h3b5178f4),
	.w8(32'hbb3dda64),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc097b96),
	.w1(32'hbd6db8e1),
	.w2(32'hbc44e30e),
	.w3(32'h3c87f83c),
	.w4(32'hbb9100b8),
	.w5(32'h3c3ca838),
	.w6(32'hbcb90535),
	.w7(32'h3d4062dc),
	.w8(32'h3b7e013f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b12f2),
	.w1(32'h3b00aba9),
	.w2(32'h3cd152d4),
	.w3(32'hbd6304d2),
	.w4(32'h3b57bcfc),
	.w5(32'hbc2ec3e4),
	.w6(32'h3b802ba0),
	.w7(32'h3ce19f90),
	.w8(32'hbc83df4a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbe7ce),
	.w1(32'hbc938b36),
	.w2(32'hbbb753bf),
	.w3(32'hbbca2bfe),
	.w4(32'h3b716e78),
	.w5(32'hbc1fe742),
	.w6(32'hbcad2eec),
	.w7(32'hbc450220),
	.w8(32'hbcccff6b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef6518),
	.w1(32'h3c03aa5d),
	.w2(32'h3c070940),
	.w3(32'h3b8dac51),
	.w4(32'h3bbfb354),
	.w5(32'hbbc67d4e),
	.w6(32'h3aa1f196),
	.w7(32'hbbc28e08),
	.w8(32'hbcbef738),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c659c5b),
	.w1(32'h3b2b4ad4),
	.w2(32'hbc876b76),
	.w3(32'hbcaad521),
	.w4(32'hbc5b7dca),
	.w5(32'h3ca34f2d),
	.w6(32'hbc17ada7),
	.w7(32'hbc478f5b),
	.w8(32'h3d4fa696),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6385f3),
	.w1(32'hbcbfe202),
	.w2(32'hbb908f5b),
	.w3(32'h3cd93045),
	.w4(32'h3c543c3c),
	.w5(32'h3b0fe734),
	.w6(32'hbc257ffa),
	.w7(32'hbb8ccad1),
	.w8(32'hbbb53073),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bfc88),
	.w1(32'h3b3ffcf6),
	.w2(32'hbb8d3b03),
	.w3(32'hbc4b38be),
	.w4(32'hbc6f7b16),
	.w5(32'hbd178399),
	.w6(32'h3c9b9570),
	.w7(32'h3b1d1f89),
	.w8(32'hbd1961a1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02e010),
	.w1(32'hbd5f300b),
	.w2(32'hbcc5ff60),
	.w3(32'hbca7f592),
	.w4(32'h3cb54232),
	.w5(32'hbab0fd9a),
	.w6(32'hbc78c328),
	.w7(32'h3c793650),
	.w8(32'h3cb1e3ea),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0b725),
	.w1(32'h3d8bd77b),
	.w2(32'hbba908da),
	.w3(32'hbd7650a2),
	.w4(32'h3c6d6c56),
	.w5(32'h3b50ade6),
	.w6(32'hbcac5560),
	.w7(32'h3b43f7d8),
	.w8(32'hbb96601d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f455e),
	.w1(32'hbbd2267e),
	.w2(32'hbd48ff32),
	.w3(32'hbc19b4c9),
	.w4(32'h3aadcd1f),
	.w5(32'hbb573735),
	.w6(32'hbbb90c81),
	.w7(32'h3ae86f19),
	.w8(32'hbd1fff03),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1bfc75),
	.w1(32'h3c0b8413),
	.w2(32'h3c88d7b9),
	.w3(32'hbce844cd),
	.w4(32'hbd34cc20),
	.w5(32'hbc12ee4a),
	.w6(32'hbd96a402),
	.w7(32'hbc327a36),
	.w8(32'hbbaf9537),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2c02b),
	.w1(32'hbbc57e3e),
	.w2(32'hbb423ea2),
	.w3(32'hbd11eb74),
	.w4(32'hbbd437d0),
	.w5(32'hbbb72bed),
	.w6(32'h3ce497f6),
	.w7(32'h3c39cc3c),
	.w8(32'h3c057dc6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7f1d3),
	.w1(32'hbcb705b5),
	.w2(32'hbd3f7980),
	.w3(32'h3d274c86),
	.w4(32'h3cc8f50e),
	.w5(32'h3bc347a7),
	.w6(32'hbbd818ae),
	.w7(32'hbc90a532),
	.w8(32'h3ac95a50),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8000bf),
	.w1(32'hbb6adb5c),
	.w2(32'hbb779f8e),
	.w3(32'hbc433e17),
	.w4(32'hbbc368e9),
	.w5(32'h3c1814de),
	.w6(32'h3b3625ba),
	.w7(32'hbbb79c7f),
	.w8(32'hbc6d1398),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b61f4),
	.w1(32'hbccae021),
	.w2(32'hba286a41),
	.w3(32'hbb092f71),
	.w4(32'h3b55c647),
	.w5(32'hbc475801),
	.w6(32'hbb9bf0b0),
	.w7(32'h3b38e57d),
	.w8(32'hbc1fd6a6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule