module layer_10_featuremap_138(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35aeb88c),
	.w1(32'hb681abd0),
	.w2(32'h36343491),
	.w3(32'hb48a91b1),
	.w4(32'hb6928311),
	.w5(32'hb590c4b4),
	.w6(32'hb5500a36),
	.w7(32'hb6495455),
	.w8(32'hb49f73cd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3732dbd7),
	.w1(32'h370c2df7),
	.w2(32'h36e5ad38),
	.w3(32'h36d878f8),
	.w4(32'h36eb6296),
	.w5(32'h36d8dbaa),
	.w6(32'h36ad41f0),
	.w7(32'h361695e8),
	.w8(32'h353c519d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6911d4b),
	.w1(32'h3666bd22),
	.w2(32'h366bd05a),
	.w3(32'hb62912cc),
	.w4(32'h36494356),
	.w5(32'h366ef0c4),
	.w6(32'h34bf8183),
	.w7(32'h34e6240d),
	.w8(32'hb5d4caac),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e8815a),
	.w1(32'h3566a372),
	.w2(32'h367d1376),
	.w3(32'h35bdb180),
	.w4(32'hb6358211),
	.w5(32'hb57cc165),
	.w6(32'h35b305b3),
	.w7(32'h36e91032),
	.w8(32'h36bf09bd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h354b1ff1),
	.w1(32'hb5fb65d6),
	.w2(32'h35cee955),
	.w3(32'h36ba5e8a),
	.w4(32'hb5b5afd6),
	.w5(32'h3603eabc),
	.w6(32'hb4a971d5),
	.w7(32'h37002aba),
	.w8(32'h3576b785),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68799fc),
	.w1(32'h361b16c4),
	.w2(32'h34cdf933),
	.w3(32'hb5d96663),
	.w4(32'hb5a3452d),
	.w5(32'hb660d670),
	.w6(32'h3502b2ae),
	.w7(32'hb5e8879b),
	.w8(32'hb67f9535),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61dd9ec),
	.w1(32'hb617c91d),
	.w2(32'h365ad97c),
	.w3(32'hb7566446),
	.w4(32'hb6c44c9f),
	.w5(32'hb687804a),
	.w6(32'hb6123e9f),
	.w7(32'hb5e72b91),
	.w8(32'hb7403338),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a7659f),
	.w1(32'hb714e9fb),
	.w2(32'h38155c6d),
	.w3(32'hb875ec44),
	.w4(32'hb7bf2a25),
	.w5(32'h37a3e426),
	.w6(32'hb7ebcd87),
	.w7(32'hb69e3bc5),
	.w8(32'h3752e79a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8860011),
	.w1(32'h381810c1),
	.w2(32'h38c342e2),
	.w3(32'hb8c61be2),
	.w4(32'h36ab7cb3),
	.w5(32'h38939a7a),
	.w6(32'hb91781cf),
	.w7(32'h378b4523),
	.w8(32'h38b0426f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38330822),
	.w1(32'hb8e94207),
	.w2(32'hb8ad609e),
	.w3(32'h39078a9a),
	.w4(32'hb8d98147),
	.w5(32'hb8257e1f),
	.w6(32'h382d74f0),
	.w7(32'hb89b4a4c),
	.w8(32'h385a40cf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35215bba),
	.w1(32'h3898e51b),
	.w2(32'h380dfe93),
	.w3(32'hb69585d0),
	.w4(32'h381b6ab4),
	.w5(32'h38a37141),
	.w6(32'h3802a395),
	.w7(32'h37908217),
	.w8(32'hb80d87cc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ea1905),
	.w1(32'h370daf2f),
	.w2(32'hb80850c3),
	.w3(32'hb7a24171),
	.w4(32'h380c1f9e),
	.w5(32'hb801248d),
	.w6(32'h3677e3e8),
	.w7(32'h37a9fb16),
	.w8(32'hb7900f7d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb210d),
	.w1(32'hb8ab4e0f),
	.w2(32'hb82582d5),
	.w3(32'hb8b461b1),
	.w4(32'hb6b2a6bf),
	.w5(32'h376535fd),
	.w6(32'hb87d82c9),
	.w7(32'hb8411789),
	.w8(32'h3785df83),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ae4f3b),
	.w1(32'h37d5e492),
	.w2(32'hb8699278),
	.w3(32'h3758152e),
	.w4(32'h3736dbb2),
	.w5(32'hb8207183),
	.w6(32'hb4fec0e8),
	.w7(32'h37ff7ef8),
	.w8(32'hb7cb295a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87cf622),
	.w1(32'h37f6e020),
	.w2(32'hb7853158),
	.w3(32'h37e7c998),
	.w4(32'h37fcf453),
	.w5(32'h37a3a8f6),
	.w6(32'h368359a0),
	.w7(32'h388b8e3e),
	.w8(32'h3850326f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb871fa65),
	.w1(32'h382c776f),
	.w2(32'h383d7ea7),
	.w3(32'hb70b50ff),
	.w4(32'h3812aa59),
	.w5(32'h3890b232),
	.w6(32'hb889e6c2),
	.w7(32'h37eb9b4b),
	.w8(32'h37d87521),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3811c29b),
	.w1(32'h38b630d0),
	.w2(32'h383ca9b3),
	.w3(32'h37bfdbce),
	.w4(32'h379c4f11),
	.w5(32'h3787843b),
	.w6(32'h3856e078),
	.w7(32'h3887ca66),
	.w8(32'h37f47d91),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381944af),
	.w1(32'hb89c9ddb),
	.w2(32'hb90a3890),
	.w3(32'h381c7351),
	.w4(32'hb8122442),
	.w5(32'hb8faaad5),
	.w6(32'h3817c955),
	.w7(32'hb882cc05),
	.w8(32'hb8ff0b64),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83c40f3),
	.w1(32'hb7871811),
	.w2(32'hb81980ec),
	.w3(32'hb822ddcd),
	.w4(32'hb62384ae),
	.w5(32'hb7aed2da),
	.w6(32'hb710fa39),
	.w7(32'hb769c9a3),
	.w8(32'hb7c718e8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36039007),
	.w1(32'h36384cbc),
	.w2(32'h3606bd7f),
	.w3(32'h3687d3ee),
	.w4(32'h35d2852c),
	.w5(32'h35dcfc7d),
	.w6(32'h36572865),
	.w7(32'h3551aca7),
	.w8(32'h35a4500e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d41092),
	.w1(32'h36ef730c),
	.w2(32'h35d44b01),
	.w3(32'h35fd42b9),
	.w4(32'h3678cc69),
	.w5(32'hb61c4f5d),
	.w6(32'h36d16231),
	.w7(32'hb5ad924f),
	.w8(32'h35cdc217),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370c0df1),
	.w1(32'h378eb439),
	.w2(32'h376b8035),
	.w3(32'h371630e6),
	.w4(32'h369d4019),
	.w5(32'hb6c7ec51),
	.w6(32'hb6354a28),
	.w7(32'hb50b9eef),
	.w8(32'hb753a7af),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a65077),
	.w1(32'hb938f8fe),
	.w2(32'hb93b2d49),
	.w3(32'hb9775604),
	.w4(32'hb88cf712),
	.w5(32'hb938d316),
	.w6(32'hb8cd287c),
	.w7(32'hb93e08a2),
	.w8(32'h3768c5dd),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eec4f7),
	.w1(32'hb7d7237f),
	.w2(32'hb80eb9a9),
	.w3(32'hb8b845d7),
	.w4(32'hb8621e75),
	.w5(32'hb859bb77),
	.w6(32'hb8aa849e),
	.w7(32'hb8754bbb),
	.w8(32'hb84f208f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d73c3),
	.w1(32'hb6e269a2),
	.w2(32'hb948141e),
	.w3(32'hb888c650),
	.w4(32'h3900a0fe),
	.w5(32'hb928a202),
	.w6(32'hb84fbf38),
	.w7(32'h383ba6c3),
	.w8(32'hb8f1482a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d2707b),
	.w1(32'h3798dcd7),
	.w2(32'h37e5252d),
	.w3(32'hb8038e08),
	.w4(32'hb7697ca5),
	.w5(32'h37fbb50c),
	.w6(32'hb810dfdc),
	.w7(32'hb69ffc4e),
	.w8(32'h382b9929),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7262c62),
	.w1(32'h3685160b),
	.w2(32'hb6536067),
	.w3(32'hb5b5d670),
	.w4(32'h36d47817),
	.w5(32'hb5e66344),
	.w6(32'h36a9afd1),
	.w7(32'h368b1c25),
	.w8(32'h360efeb4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370ee993),
	.w1(32'h37f7288e),
	.w2(32'hb779bb67),
	.w3(32'h377c2298),
	.w4(32'h38273076),
	.w5(32'h376bac86),
	.w6(32'h37c65de4),
	.w7(32'h380040cd),
	.w8(32'h37061fc0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3825667d),
	.w1(32'h35a94239),
	.w2(32'hb70bb6b3),
	.w3(32'h380d393f),
	.w4(32'h38541590),
	.w5(32'hb8189820),
	.w6(32'hb6c785e9),
	.w7(32'h382faa17),
	.w8(32'hb83c7c31),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5f6a1),
	.w1(32'h370cef44),
	.w2(32'h3914db57),
	.w3(32'hb8004eb9),
	.w4(32'hb8c63d5e),
	.w5(32'h390f1036),
	.w6(32'hb84bf830),
	.w7(32'hb8994114),
	.w8(32'h39135e34),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb667a5ae),
	.w1(32'h37267979),
	.w2(32'hb60726bd),
	.w3(32'hb65a63e8),
	.w4(32'h37138e07),
	.w5(32'hb65d31ba),
	.w6(32'h36a924ba),
	.w7(32'h369c7037),
	.w8(32'hb672dfb1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bd8038),
	.w1(32'h37c4f556),
	.w2(32'hb7ba2484),
	.w3(32'h38707bce),
	.w4(32'h37e69e34),
	.w5(32'hb8396ba1),
	.w6(32'h382c84bf),
	.w7(32'h3544b269),
	.w8(32'hb816bacf),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3836e852),
	.w1(32'hb756b8f9),
	.w2(32'hb7dcbf89),
	.w3(32'h377d5957),
	.w4(32'hb835c325),
	.w5(32'hb8570818),
	.w6(32'hb82a8a86),
	.w7(32'hb86ad65d),
	.w8(32'hb8a7e264),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb863c46c),
	.w1(32'hb7f72afe),
	.w2(32'h376e4566),
	.w3(32'hb840a727),
	.w4(32'hb74a18de),
	.w5(32'h3750431d),
	.w6(32'hb7b96715),
	.w7(32'hb8366229),
	.w8(32'h384b170c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3632397d),
	.w1(32'hb6419696),
	.w2(32'hb6f63d04),
	.w3(32'h356680a1),
	.w4(32'hb5d1c19a),
	.w5(32'hb659eeaa),
	.w6(32'hb6afc3b1),
	.w7(32'hb6aaeeca),
	.w8(32'hb67adca8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f925bc),
	.w1(32'hb686a5c8),
	.w2(32'hb72f783f),
	.w3(32'hb5d9d187),
	.w4(32'hb66d2b4d),
	.w5(32'hb79d716b),
	.w6(32'hb686e71f),
	.w7(32'hb6775312),
	.w8(32'hb74732c3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39932c88),
	.w1(32'hb839cb60),
	.w2(32'hb94e477a),
	.w3(32'h39547978),
	.w4(32'hb927ad65),
	.w5(32'hb94d04eb),
	.w6(32'h3900803b),
	.w7(32'hb926aa12),
	.w8(32'hb77ca2b5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896fe1f),
	.w1(32'hb8575189),
	.w2(32'hb99d947a),
	.w3(32'h394fe7ce),
	.w4(32'h39287e23),
	.w5(32'hb92c2714),
	.w6(32'h39984a73),
	.w7(32'h392d1eb1),
	.w8(32'hb8c95a4d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb804b52b),
	.w1(32'h38036e4c),
	.w2(32'hb94d212d),
	.w3(32'h3933cadc),
	.w4(32'h392f4bd8),
	.w5(32'hb90ed0d3),
	.w6(32'h38db54a6),
	.w7(32'h389b73fd),
	.w8(32'hb96876b1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb722fd5a),
	.w1(32'hb75be4c4),
	.w2(32'hb7ad4e98),
	.w3(32'hb740314c),
	.w4(32'hb6a3fd74),
	.w5(32'hb792e8da),
	.w6(32'hb787521a),
	.w7(32'hb70dd168),
	.w8(32'hb7a8a9d4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807445d),
	.w1(32'hb7c03585),
	.w2(32'h388e894b),
	.w3(32'hb8ab9bc2),
	.w4(32'hb83e7b66),
	.w5(32'h38201875),
	.w6(32'hb7a7d14a),
	.w7(32'h3657c95a),
	.w8(32'h37efd320),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8274d29),
	.w1(32'hb7e7c7fa),
	.w2(32'hb73d3ebf),
	.w3(32'hb82d71ad),
	.w4(32'hb7c0c7df),
	.w5(32'hb7319be7),
	.w6(32'hb6626275),
	.w7(32'h37c5057e),
	.w8(32'h371784a1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37375b0f),
	.w1(32'h37c40157),
	.w2(32'hb8e1c77b),
	.w3(32'h381df991),
	.w4(32'h385a568e),
	.w5(32'hb883cad7),
	.w6(32'h37063a29),
	.w7(32'h37e5ba35),
	.w8(32'hb812daaa),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c6df0),
	.w1(32'hb9d7f34b),
	.w2(32'h38fa21db),
	.w3(32'hba092187),
	.w4(32'hb9df1c48),
	.w5(32'h399954a0),
	.w6(32'hb9d092d9),
	.w7(32'hb94b2608),
	.w8(32'h38891289),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aad795),
	.w1(32'hb7e81362),
	.w2(32'h35d3a6aa),
	.w3(32'hb80ec07d),
	.w4(32'hb8a84cf5),
	.w5(32'hb49c577c),
	.w6(32'hb83d89f6),
	.w7(32'hb852eab0),
	.w8(32'h370a541c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90253b8),
	.w1(32'hb9209917),
	.w2(32'h380845a0),
	.w3(32'hb92d0233),
	.w4(32'hb94f3aa8),
	.w5(32'hb67d0993),
	.w6(32'hb929345d),
	.w7(32'hb9219afc),
	.w8(32'h377f1584),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918705e),
	.w1(32'hb924046e),
	.w2(32'h39437748),
	.w3(32'hb965dcc7),
	.w4(32'hb986e4f7),
	.w5(32'h395ca74d),
	.w6(32'hb9425c9c),
	.w7(32'hb91e335e),
	.w8(32'h3976ffed),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9797413),
	.w1(32'hb904f33e),
	.w2(32'h3892ad30),
	.w3(32'hb9546182),
	.w4(32'hb8d727ee),
	.w5(32'h35e3b633),
	.w6(32'hb8fd9d25),
	.w7(32'hb7be4640),
	.w8(32'h3845d4c9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888993c),
	.w1(32'hb906c9ee),
	.w2(32'h35c95137),
	.w3(32'hb94ac703),
	.w4(32'hb92e54d0),
	.w5(32'h38f08df4),
	.w6(32'hb8bdf97c),
	.w7(32'hb81fcc4c),
	.w8(32'h37db7d86),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c07716),
	.w1(32'hb94a7d5b),
	.w2(32'h3901b1f6),
	.w3(32'hb9ba75b9),
	.w4(32'hb958a0f9),
	.w5(32'h37d3c79b),
	.w6(32'hb9a0ff9f),
	.w7(32'hb91cfa89),
	.w8(32'h38a3ab93),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b5de42),
	.w1(32'hb87ed3d3),
	.w2(32'hb8ea4bfe),
	.w3(32'hb8c4c713),
	.w4(32'h372317bc),
	.w5(32'hb874de77),
	.w6(32'h3604d64e),
	.w7(32'h37c8dd81),
	.w8(32'hb83ca756),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d0cb37),
	.w1(32'h35425b4d),
	.w2(32'hb606aeee),
	.w3(32'hb6963460),
	.w4(32'hb5bb8c45),
	.w5(32'hb684997c),
	.w6(32'h35c17835),
	.w7(32'h364540a6),
	.w8(32'h36bd3b8e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8201927),
	.w1(32'hb794a14a),
	.w2(32'hb73c5af6),
	.w3(32'hb7a22fa9),
	.w4(32'hb6a5310d),
	.w5(32'hb7767f43),
	.w6(32'hb72d9675),
	.w7(32'h35c23122),
	.w8(32'hb607f34a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883ac69),
	.w1(32'hb8843346),
	.w2(32'hb898a97d),
	.w3(32'hb850e3d0),
	.w4(32'hb826a376),
	.w5(32'hb873ac37),
	.w6(32'hb7c8fa40),
	.w7(32'hb7d8a88c),
	.w8(32'hb8586668),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74d061a),
	.w1(32'h374666b2),
	.w2(32'hb792c5dd),
	.w3(32'hb6f26f11),
	.w4(32'h37282742),
	.w5(32'hb7c8d41b),
	.w6(32'h374b37a6),
	.w7(32'h3750127b),
	.w8(32'hb7bc90c8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6328f0e),
	.w1(32'h36d58f9a),
	.w2(32'hb6999173),
	.w3(32'hb65333bf),
	.w4(32'h36038dd0),
	.w5(32'hb712308f),
	.w6(32'h370564bf),
	.w7(32'hb6a11551),
	.w8(32'hb6621a33),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb637d4a0),
	.w1(32'h35a56960),
	.w2(32'hb534e164),
	.w3(32'hb6f99a06),
	.w4(32'hb5aa9cd7),
	.w5(32'hb6231e46),
	.w6(32'hb698d301),
	.w7(32'hb6a96a58),
	.w8(32'hb6035865),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68ca1eb),
	.w1(32'hb72c4dd7),
	.w2(32'hb72ed057),
	.w3(32'hb649af96),
	.w4(32'hb688f3ba),
	.w5(32'h36203013),
	.w6(32'hb689a48a),
	.w7(32'h36946621),
	.w8(32'hb502bee9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3626a8dc),
	.w1(32'h36f82a3a),
	.w2(32'hb82f5fd1),
	.w3(32'h38057f6d),
	.w4(32'h37cf00c6),
	.w5(32'hb8426b03),
	.w6(32'h37cedbe4),
	.w7(32'h37a15197),
	.w8(32'hb83133a1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370542fe),
	.w1(32'h38663166),
	.w2(32'h385a4c9b),
	.w3(32'hb68b5d72),
	.w4(32'h37db29df),
	.w5(32'h38919459),
	.w6(32'hb7d6afdc),
	.w7(32'h3824091b),
	.w8(32'h335792e2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb821fc7c),
	.w1(32'hb6a03a6b),
	.w2(32'h3802db63),
	.w3(32'hb89405d4),
	.w4(32'hb75bee74),
	.w5(32'h37e501a0),
	.w6(32'hb860eb4a),
	.w7(32'h36bfa3b3),
	.w8(32'h36956171),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b66511),
	.w1(32'h379d326f),
	.w2(32'h377d3b16),
	.w3(32'hb76f8385),
	.w4(32'hb66d85e8),
	.w5(32'hb74723d4),
	.w6(32'hb607b108),
	.w7(32'hb7b4cb0d),
	.w8(32'h37144459),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e817f2),
	.w1(32'hb6711782),
	.w2(32'h36dcd32c),
	.w3(32'hb818abb7),
	.w4(32'h36c3babd),
	.w5(32'h377e79d2),
	.w6(32'hb78dc057),
	.w7(32'hb6437b7d),
	.w8(32'h37067ccd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b6250f),
	.w1(32'hb55a95a1),
	.w2(32'h34ad77c9),
	.w3(32'h369d3644),
	.w4(32'h3534475e),
	.w5(32'h3618e3d3),
	.w6(32'hb5bfafbd),
	.w7(32'hb646dde4),
	.w8(32'h352eec31),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3763714a),
	.w1(32'h3681de9e),
	.w2(32'hb6d17c89),
	.w3(32'h3767632b),
	.w4(32'h36aecd05),
	.w5(32'hb522fda5),
	.w6(32'hb68ec347),
	.w7(32'hb71db103),
	.w8(32'hb79e933e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36896ae2),
	.w1(32'hb5181d8b),
	.w2(32'h366abf17),
	.w3(32'h35f60648),
	.w4(32'h35aeff18),
	.w5(32'h36a3008c),
	.w6(32'hb68c987d),
	.w7(32'h360c94c4),
	.w8(32'h35a34f9f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ff4d61),
	.w1(32'hb78f1f7a),
	.w2(32'hb506ab32),
	.w3(32'hb74d6517),
	.w4(32'hb71d2821),
	.w5(32'h3718f1c2),
	.w6(32'hb717a8dd),
	.w7(32'hb77656ea),
	.w8(32'hb7529b07),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ed3a53),
	.w1(32'h374abafa),
	.w2(32'hb8a9bfcb),
	.w3(32'hb7ae7f99),
	.w4(32'h3758a9df),
	.w5(32'hb8aa8b1b),
	.w6(32'h375fd1c7),
	.w7(32'hb5f1ad9e),
	.w8(32'hb886e841),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df03f6),
	.w1(32'hb851509e),
	.w2(32'hb92179de),
	.w3(32'hb7b988bb),
	.w4(32'h374cff0f),
	.w5(32'hb9092df3),
	.w6(32'hb7cef3b2),
	.w7(32'hb7aabcbf),
	.w8(32'hb8bdd595),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb860c59f),
	.w1(32'hb76c01f3),
	.w2(32'hb911439b),
	.w3(32'hb806bc60),
	.w4(32'h38060452),
	.w5(32'hb8dae0c1),
	.w6(32'hb7f45f46),
	.w7(32'hb56a0ee8),
	.w8(32'hb8897c60),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70c8513),
	.w1(32'hb62b9104),
	.w2(32'hb452194a),
	.w3(32'hb63cf9ef),
	.w4(32'h349682cb),
	.w5(32'h352fc3a6),
	.w6(32'hb5f365b9),
	.w7(32'hb6356cfa),
	.w8(32'h35f3ea8d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64d80a0),
	.w1(32'hb4779868),
	.w2(32'h3679b93b),
	.w3(32'hb589202e),
	.w4(32'hb509be57),
	.w5(32'h36271e88),
	.w6(32'h3508b190),
	.w7(32'hb51872e9),
	.w8(32'h36968fb2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ff56d6),
	.w1(32'hb6492364),
	.w2(32'h34d85d50),
	.w3(32'hb60a2ca5),
	.w4(32'h34d68288),
	.w5(32'h369f1cac),
	.w6(32'h34686c0d),
	.w7(32'h35afaf59),
	.w8(32'h3637db79),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e66a79),
	.w1(32'h36e38983),
	.w2(32'hb747c32a),
	.w3(32'h376d0f1f),
	.w4(32'h36ee7dd7),
	.w5(32'hb75f3b3d),
	.w6(32'h36485412),
	.w7(32'h36b5a396),
	.w8(32'hb78adb57),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb860f221),
	.w1(32'hb78d81b4),
	.w2(32'h36b0b004),
	.w3(32'hb8696c5a),
	.w4(32'hb7b45806),
	.w5(32'h379a2647),
	.w6(32'hb81626a6),
	.w7(32'hb75f042c),
	.w8(32'h37165e8f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b09dd2),
	.w1(32'hb799289a),
	.w2(32'hb7294d13),
	.w3(32'hb7769382),
	.w4(32'hb5804f08),
	.w5(32'h361f995f),
	.w6(32'hb78c229c),
	.w7(32'hb6d61574),
	.w8(32'h35e63a62),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7abea32),
	.w1(32'hb612e607),
	.w2(32'hb811b66f),
	.w3(32'h34bd065b),
	.w4(32'hb6f797f5),
	.w5(32'hb7f39418),
	.w6(32'hb78b1c03),
	.w7(32'h36cf5eee),
	.w8(32'hb80b1fa2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d552af),
	.w1(32'h36b8213b),
	.w2(32'h36eba69b),
	.w3(32'hb7b15481),
	.w4(32'hb6495e2f),
	.w5(32'hb79b8bb6),
	.w6(32'hb7e424e0),
	.w7(32'h35b2647b),
	.w8(32'hb5eb6bb3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ada43f),
	.w1(32'hb766d1e2),
	.w2(32'hb86db85d),
	.w3(32'hb59dc990),
	.w4(32'hb69301c7),
	.w5(32'hb8653f62),
	.w6(32'h35e17ea5),
	.w7(32'hb63a0261),
	.w8(32'hb82f5386),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75ffc8e),
	.w1(32'hb6e9b15d),
	.w2(32'hb7bab0af),
	.w3(32'hb733734e),
	.w4(32'h368307d1),
	.w5(32'hb77de57e),
	.w6(32'h36c20030),
	.w7(32'h35c8d17e),
	.w8(32'hb78cc60f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379e8044),
	.w1(32'h38036911),
	.w2(32'hb81f6bea),
	.w3(32'h37874942),
	.w4(32'h376388c9),
	.w5(32'hb841c80a),
	.w6(32'h374d44ea),
	.w7(32'hb73bf9c3),
	.w8(32'hb7eb9c2f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb753f2cd),
	.w1(32'h376bddb1),
	.w2(32'hb799c263),
	.w3(32'hb78c3bf9),
	.w4(32'h375688fb),
	.w5(32'hb78ebcaf),
	.w6(32'h36a742ae),
	.w7(32'h369ed171),
	.w8(32'hb7cbb51b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3669a4ae),
	.w1(32'h36323d0b),
	.w2(32'h348feb79),
	.w3(32'h3698780a),
	.w4(32'h3639764c),
	.w5(32'h345d8c28),
	.w6(32'h364d9454),
	.w7(32'hb387a55e),
	.w8(32'h3615a269),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359fa9c7),
	.w1(32'h35e7c7fc),
	.w2(32'h35ad34e5),
	.w3(32'hb3a4dbed),
	.w4(32'hb5953b24),
	.w5(32'h33d54758),
	.w6(32'h359e8692),
	.w7(32'hb6867a29),
	.w8(32'hb6a94e97),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ba60a6),
	.w1(32'h37b04c1e),
	.w2(32'h371d76f0),
	.w3(32'h33ced1eb),
	.w4(32'h378ce98c),
	.w5(32'h35cd8d0b),
	.w6(32'h378c9a91),
	.w7(32'h36439703),
	.w8(32'hb4f8ef9e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36065f1a),
	.w1(32'h35fda09c),
	.w2(32'h36869f2b),
	.w3(32'hb6ca6db9),
	.w4(32'h361e52c1),
	.w5(32'h36372a4e),
	.w6(32'h361c3aec),
	.w7(32'h36029a93),
	.w8(32'h35282b29),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377db003),
	.w1(32'hb666e68c),
	.w2(32'hb7985ce2),
	.w3(32'hb69e2f10),
	.w4(32'h371c57da),
	.w5(32'h36566e03),
	.w6(32'h3608583f),
	.w7(32'h3735783c),
	.w8(32'h37493bc5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6868926),
	.w1(32'h3715c3f6),
	.w2(32'h376b267d),
	.w3(32'hb6c9220a),
	.w4(32'h3562ab1e),
	.w5(32'h3641b7e4),
	.w6(32'hb6a7ab6e),
	.w7(32'h35c5f563),
	.w8(32'h36878ffb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f26a09),
	.w1(32'h361d8400),
	.w2(32'hb6dd3f30),
	.w3(32'hb7520cc7),
	.w4(32'h3600ea94),
	.w5(32'hb7263d46),
	.w6(32'hb6b09dc7),
	.w7(32'h359bd54c),
	.w8(32'hb604c11a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dcb7b4),
	.w1(32'hb81c13a2),
	.w2(32'hb90fcfd4),
	.w3(32'hb85db46f),
	.w4(32'h372a1dc3),
	.w5(32'hb8803d15),
	.w6(32'h36c81eed),
	.w7(32'h35abcb68),
	.w8(32'hb7c977c4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37011d99),
	.w1(32'h38628a37),
	.w2(32'hb884fa0b),
	.w3(32'h3729658c),
	.w4(32'h38887ec0),
	.w5(32'hb835e93d),
	.w6(32'h3877f6de),
	.w7(32'h386c5c27),
	.w8(32'hb7fdb38d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8317072),
	.w1(32'hb79b836e),
	.w2(32'hb852580c),
	.w3(32'hb7d7cb5e),
	.w4(32'h370de5e2),
	.w5(32'hb78944c5),
	.w6(32'hb83ce9f3),
	.w7(32'hb79aa716),
	.w8(32'hb6c8f975),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b548f9),
	.w1(32'h373483be),
	.w2(32'hb930f2eb),
	.w3(32'h37aa7420),
	.w4(32'h388cf7c5),
	.w5(32'hb8d67c0c),
	.w6(32'h3829efff),
	.w7(32'h37f860dd),
	.w8(32'hb8be91a4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9405287),
	.w1(32'hb905db5e),
	.w2(32'hb89f00a0),
	.w3(32'hb92a5475),
	.w4(32'hb8dcc6f8),
	.w5(32'hb8cf6ede),
	.w6(32'hb8e59339),
	.w7(32'hb8d2d960),
	.w8(32'hb8a17c00),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bf60fc),
	.w1(32'hb680eafa),
	.w2(32'h385ecc84),
	.w3(32'hb8bd9814),
	.w4(32'h36924ef2),
	.w5(32'h36257ccb),
	.w6(32'hb77fff85),
	.w7(32'hb7a99299),
	.w8(32'h37e4f269),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a3bdd8),
	.w1(32'hb7313457),
	.w2(32'hb781aba0),
	.w3(32'hb78cc7b3),
	.w4(32'hb74a99db),
	.w5(32'hb7a2677a),
	.w6(32'hb7e3a997),
	.w7(32'hb66f8c7b),
	.w8(32'hb7caf40a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9810563),
	.w1(32'hb906af07),
	.w2(32'hb73dd775),
	.w3(32'hb9991c54),
	.w4(32'h37aa7e7b),
	.w5(32'hb746c258),
	.w6(32'hb96a359e),
	.w7(32'h3588dd5b),
	.w8(32'h38d9b3c4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0502cb),
	.w1(32'hb9e27c20),
	.w2(32'h36c885a0),
	.w3(32'hba00b52e),
	.w4(32'hb97e6d9c),
	.w5(32'h373cd84d),
	.w6(32'hb9a6322a),
	.w7(32'hb96a0c94),
	.w8(32'h390e1ec3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa006d),
	.w1(32'hb8a84e72),
	.w2(32'hb98c1163),
	.w3(32'hb8e5eff8),
	.w4(32'hb8b21e94),
	.w5(32'hb95d4eb1),
	.w6(32'hb90a587b),
	.w7(32'hb901bb65),
	.w8(32'hb84e1dd4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7752e1c),
	.w1(32'h363f360b),
	.w2(32'hb831b4da),
	.w3(32'hb697a69d),
	.w4(32'h37f959fc),
	.w5(32'hb819d0fd),
	.w6(32'h364486dc),
	.w7(32'h37d2b044),
	.w8(32'hb72fca3b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9301a14),
	.w1(32'hb9cae387),
	.w2(32'hb9c0057e),
	.w3(32'hb9ecf277),
	.w4(32'hb9b3aa6b),
	.w5(32'hb90d6dcb),
	.w6(32'hb99336b4),
	.w7(32'hb8d6f528),
	.w8(32'hb8df50e9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cffb69),
	.w1(32'hb921dc60),
	.w2(32'hb90856fc),
	.w3(32'hb9d5464e),
	.w4(32'hb838dce0),
	.w5(32'hb94e5589),
	.w6(32'hb932bcde),
	.w7(32'hb8a0b676),
	.w8(32'hb8a77371),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb717f2ac),
	.w1(32'hb981fb69),
	.w2(32'h38d5abe7),
	.w3(32'hb90a4af1),
	.w4(32'hb8a6f59b),
	.w5(32'h38b917da),
	.w6(32'hb91f57be),
	.w7(32'hb8b40807),
	.w8(32'h37de85be),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8feb8de),
	.w1(32'hb9c98145),
	.w2(32'hb92df834),
	.w3(32'hb9d4660a),
	.w4(32'hb90da1e2),
	.w5(32'hb91a9e11),
	.w6(32'hb99c7189),
	.w7(32'hb92989ec),
	.w8(32'hb927f9bc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7399ef4),
	.w1(32'hb7f502fd),
	.w2(32'h37ad919e),
	.w3(32'hb8f8ea64),
	.w4(32'h37d6df58),
	.w5(32'h37bdd474),
	.w6(32'hb8b3ceb1),
	.w7(32'h383c9424),
	.w8(32'h38197ac6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b8fea3),
	.w1(32'h375dc3ad),
	.w2(32'h37a85127),
	.w3(32'h3681e593),
	.w4(32'hb6c9f25d),
	.w5(32'h3687a968),
	.w6(32'hb8949164),
	.w7(32'h36c4b90d),
	.w8(32'h37476cf9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60c4e1b),
	.w1(32'h36eb2a17),
	.w2(32'hb69c141f),
	.w3(32'h368b111d),
	.w4(32'h3795f101),
	.w5(32'hb67e3f85),
	.w6(32'hb60e8b14),
	.w7(32'h36ae2714),
	.w8(32'hb782a1f5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb714e177),
	.w1(32'h3798c473),
	.w2(32'h36a323ec),
	.w3(32'hb7db70d7),
	.w4(32'h36d86c4a),
	.w5(32'hb73157c1),
	.w6(32'hb81d817f),
	.w7(32'h375b7b5c),
	.w8(32'hb62e3922),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b49e86),
	.w1(32'hb9abd93b),
	.w2(32'hb97e2cdc),
	.w3(32'hb93280e2),
	.w4(32'hb92f806b),
	.w5(32'hb82f2064),
	.w6(32'hb8f9d00c),
	.w7(32'hb96a2cf3),
	.w8(32'hb88843dc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99881e9),
	.w1(32'hb9dea166),
	.w2(32'h39578f48),
	.w3(32'hb9c93e71),
	.w4(32'hb9b19187),
	.w5(32'h3786d4e1),
	.w6(32'hb9a7c513),
	.w7(32'hb9b040df),
	.w8(32'h38ef9f20),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7be5850),
	.w1(32'hb8034912),
	.w2(32'h386d9eec),
	.w3(32'hb863ea04),
	.w4(32'hb832f2fa),
	.w5(32'hb78fc0e1),
	.w6(32'hb870e44c),
	.w7(32'hb7e6f9b7),
	.w8(32'h35979a30),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cdd24e),
	.w1(32'hb9346883),
	.w2(32'h374890a6),
	.w3(32'hb9096848),
	.w4(32'hb8d574a9),
	.w5(32'h389c9a1a),
	.w6(32'hb82e401f),
	.w7(32'hb7ecced3),
	.w8(32'h383a9a67),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ba7a61),
	.w1(32'h382d4ebd),
	.w2(32'hb87c9da3),
	.w3(32'h3825f4df),
	.w4(32'h383c18ed),
	.w5(32'hb84b602e),
	.w6(32'h38729b0e),
	.w7(32'h38465b11),
	.w8(32'hb811b185),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38288dc2),
	.w1(32'h35c16916),
	.w2(32'h3931ff0e),
	.w3(32'hb7684556),
	.w4(32'hb7f7dfe1),
	.w5(32'h389638dd),
	.w6(32'hb86119e7),
	.w7(32'h38b8100c),
	.w8(32'hb80eb875),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f5fdb),
	.w1(32'hb7cfaf95),
	.w2(32'hb79c2ff2),
	.w3(32'hb820f36f),
	.w4(32'hb7a4e257),
	.w5(32'hb7a0360d),
	.w6(32'hb7d974e6),
	.w7(32'hb6dba8e5),
	.w8(32'hb7668405),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d63e27),
	.w1(32'h35c39bb3),
	.w2(32'h36bee069),
	.w3(32'hb784b758),
	.w4(32'hb53147c8),
	.w5(32'h3657cddd),
	.w6(32'hb6ff72c0),
	.w7(32'h34d02238),
	.w8(32'hb5e208a2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36601ca8),
	.w1(32'h3623d10e),
	.w2(32'h361dd20d),
	.w3(32'h35be04a3),
	.w4(32'hb52e267a),
	.w5(32'hb4df9535),
	.w6(32'hb5e7ddc0),
	.w7(32'hb599676b),
	.w8(32'h352cc9e1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h354bed6f),
	.w1(32'h3582f772),
	.w2(32'h3523622c),
	.w3(32'hb5905358),
	.w4(32'hb5c54830),
	.w5(32'hb5da8018),
	.w6(32'hb5e019ba),
	.w7(32'hb639ee1f),
	.w8(32'hb5a51577),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d7b221),
	.w1(32'h369a89d1),
	.w2(32'h3731f9b7),
	.w3(32'h3698fc21),
	.w4(32'hb54fdf25),
	.w5(32'hb4f61aef),
	.w6(32'h3750c0f7),
	.w7(32'h35ab30cf),
	.w8(32'hb42d4502),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ea37a6),
	.w1(32'h38141fe8),
	.w2(32'hb7ed72e4),
	.w3(32'h37c2155d),
	.w4(32'h37c45961),
	.w5(32'hb8062f2a),
	.w6(32'h37c6bc19),
	.w7(32'h37bb5a73),
	.w8(32'hb8295264),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a9e1af),
	.w1(32'hb610451d),
	.w2(32'h37bc1dbb),
	.w3(32'hb69103ae),
	.w4(32'hb7f41220),
	.w5(32'h37ae1ca2),
	.w6(32'hb7f5c7da),
	.w7(32'hb7dd0536),
	.w8(32'h36a54f01),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb811c823),
	.w1(32'hb76857d2),
	.w2(32'h358f3dd8),
	.w3(32'hb7fa5743),
	.w4(32'h35a55005),
	.w5(32'hb70638cc),
	.w6(32'h3516034d),
	.w7(32'h36983d35),
	.w8(32'hb76cc931),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3745b9e0),
	.w1(32'h3797529f),
	.w2(32'h37a78efe),
	.w3(32'h371485c9),
	.w4(32'h378e22ff),
	.w5(32'h374ad746),
	.w6(32'h370e1d7d),
	.w7(32'h374a42a4),
	.w8(32'h369dd4c1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35fe447c),
	.w1(32'h35e27a46),
	.w2(32'h37388090),
	.w3(32'h34b9509a),
	.w4(32'hb65df87d),
	.w5(32'h3540e832),
	.w6(32'h349c1aa6),
	.w7(32'h33d42b7c),
	.w8(32'hb56f1e96),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361e711b),
	.w1(32'hb6d49d32),
	.w2(32'hb616383f),
	.w3(32'hb75a0bd7),
	.w4(32'hb70e394b),
	.w5(32'hb5b79b20),
	.w6(32'hb7350176),
	.w7(32'hb6dcbdb7),
	.w8(32'h35a7e603),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3643172c),
	.w1(32'h36c739ed),
	.w2(32'hb63a49be),
	.w3(32'h34085e4e),
	.w4(32'h36051556),
	.w5(32'hb78c4f3d),
	.w6(32'hb693e476),
	.w7(32'hb6f58ac5),
	.w8(32'hb77b01ba),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d54b9d),
	.w1(32'h3abfa70d),
	.w2(32'hbaa22155),
	.w3(32'hb6213beb),
	.w4(32'h3b372ed5),
	.w5(32'hbb5f23a9),
	.w6(32'h3b955114),
	.w7(32'hbafebc1b),
	.w8(32'hbb0dcadd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb829a3d),
	.w1(32'hbb91d31f),
	.w2(32'hbb75c6ce),
	.w3(32'hbb91118f),
	.w4(32'hbaf578e3),
	.w5(32'hbbc270a7),
	.w6(32'h39e4ddba),
	.w7(32'hbb9e106e),
	.w8(32'hbb97d495),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d4ba0),
	.w1(32'h3acfd5cf),
	.w2(32'hb97245a1),
	.w3(32'hbbf69cf6),
	.w4(32'hba844048),
	.w5(32'hbb5d2beb),
	.w6(32'h3b281839),
	.w7(32'hba1afd90),
	.w8(32'hba66e1c5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a4c08),
	.w1(32'h3bc26180),
	.w2(32'h3b98b0ce),
	.w3(32'hbbe6567f),
	.w4(32'h3ba86653),
	.w5(32'h3bc45e9f),
	.w6(32'h39594a06),
	.w7(32'h3b455f1e),
	.w8(32'h3a0cd48d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5c15a),
	.w1(32'h3b33e495),
	.w2(32'h398f7f35),
	.w3(32'h3b7afc4f),
	.w4(32'hb993500a),
	.w5(32'hba902ae3),
	.w6(32'hbb06b6dd),
	.w7(32'hbad913d4),
	.w8(32'hbb189c9d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a4d8b),
	.w1(32'h3c120c30),
	.w2(32'h3bb1fb9d),
	.w3(32'hbb8e3af0),
	.w4(32'h3ba36707),
	.w5(32'h3c097cd1),
	.w6(32'h3bae8846),
	.w7(32'hb89abcd9),
	.w8(32'hbb1add67),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b339ded),
	.w1(32'h3a2a4393),
	.w2(32'h3af46aad),
	.w3(32'h3b8ff8f6),
	.w4(32'h3a220d75),
	.w5(32'h3af2d712),
	.w6(32'h3b1c67f4),
	.w7(32'h3a664712),
	.w8(32'hbb87c67f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820b75),
	.w1(32'hbb92f9b1),
	.w2(32'hbb581543),
	.w3(32'hbba8348b),
	.w4(32'hba14178e),
	.w5(32'hbb9a0c5f),
	.w6(32'h3a94edb7),
	.w7(32'hbbaae428),
	.w8(32'hbb3bc93b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6d3f5),
	.w1(32'h3c1c844b),
	.w2(32'h3bf1ad0e),
	.w3(32'hbba4ce21),
	.w4(32'h3c18de51),
	.w5(32'h3c2b37e1),
	.w6(32'hba7c0086),
	.w7(32'h3b910a04),
	.w8(32'h3b07f23b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb2cc3),
	.w1(32'hbac2f63e),
	.w2(32'h3a55ad1a),
	.w3(32'h3bcfd462),
	.w4(32'h39a9bc22),
	.w5(32'hbb4b047b),
	.w6(32'h3bd3ee7d),
	.w7(32'h3b083fad),
	.w8(32'h3b01aa12),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba37a01),
	.w1(32'hbadfbc22),
	.w2(32'hbb22887b),
	.w3(32'hbb87f63a),
	.w4(32'hbb3b73b9),
	.w5(32'hbbba5c51),
	.w6(32'hba926251),
	.w7(32'hbbb703a4),
	.w8(32'hbb9488de),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1d1b0),
	.w1(32'h3c29c312),
	.w2(32'h39c0a799),
	.w3(32'hbbd680ad),
	.w4(32'h3c32dd90),
	.w5(32'h3c3a904e),
	.w6(32'hbaf5f492),
	.w7(32'hb989bcfa),
	.w8(32'h3afaca1b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56059f),
	.w1(32'h3b268285),
	.w2(32'h3b777d16),
	.w3(32'h3c667380),
	.w4(32'h3aeae278),
	.w5(32'h3ba88bfd),
	.w6(32'h3bc3ad9b),
	.w7(32'h3b93d7e3),
	.w8(32'h3b8bbed6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37220c6f),
	.w1(32'h39968e1d),
	.w2(32'h3ba899ea),
	.w3(32'h3b5eef20),
	.w4(32'h3bb6d7a6),
	.w5(32'h3bcf0697),
	.w6(32'h3adcd473),
	.w7(32'h3b8ecdc4),
	.w8(32'h3b0c6c3c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d014a),
	.w1(32'hbb37d189),
	.w2(32'hbb1761a7),
	.w3(32'h3b56f090),
	.w4(32'hbb307ce9),
	.w5(32'hbb8d3ef7),
	.w6(32'h39dd0547),
	.w7(32'hbb3a7143),
	.w8(32'hbb3294db),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c7ddd),
	.w1(32'hbb94378d),
	.w2(32'hba14d54b),
	.w3(32'hbb88d9ed),
	.w4(32'hbb6eb815),
	.w5(32'hbb96d946),
	.w6(32'h3c0d089f),
	.w7(32'h3b8fe495),
	.w8(32'h3be9af0f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb736e21),
	.w1(32'h3a871489),
	.w2(32'h3b97e49a),
	.w3(32'hbb129b38),
	.w4(32'h3b8096b3),
	.w5(32'h3bc8ac1c),
	.w6(32'hba0d557c),
	.w7(32'h3b2ae03b),
	.w8(32'hbaa42950),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb802de),
	.w1(32'hbb93d934),
	.w2(32'hbb7646ff),
	.w3(32'hb99d4de5),
	.w4(32'hbb982b92),
	.w5(32'hbbeedb27),
	.w6(32'hbb8a714f),
	.w7(32'hbc09e2ea),
	.w8(32'hbbf7dbcc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e8296),
	.w1(32'h3b12cc60),
	.w2(32'h3c0cd681),
	.w3(32'hbc09181b),
	.w4(32'hba15c8a6),
	.w5(32'h3b04e194),
	.w6(32'h3b94f4e3),
	.w7(32'h3c135e5d),
	.w8(32'h3b2f4d19),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b82705),
	.w1(32'h3b93d3b1),
	.w2(32'h3b39f9ea),
	.w3(32'hbb358ac0),
	.w4(32'h3b7aa600),
	.w5(32'h3c0be4b9),
	.w6(32'hbc1e166a),
	.w7(32'hbb0e118e),
	.w8(32'hbb97af2e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9cf75),
	.w1(32'hb9ef6028),
	.w2(32'h3a0c42a5),
	.w3(32'h3be11997),
	.w4(32'h3a945ebe),
	.w5(32'h3b424f26),
	.w6(32'hbb062d3e),
	.w7(32'h3aed2b48),
	.w8(32'hbb2decfb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f56c5),
	.w1(32'hb8c7c3cb),
	.w2(32'h3a125ffa),
	.w3(32'hbb1b849e),
	.w4(32'h392acc77),
	.w5(32'hbb1431c4),
	.w6(32'h3a41abe6),
	.w7(32'hbab8b49a),
	.w8(32'hb73452b5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb227925),
	.w1(32'hb9a71cb6),
	.w2(32'h3b305de9),
	.w3(32'hbaae367d),
	.w4(32'h3a822ad5),
	.w5(32'h3a15c4e8),
	.w6(32'h3b83d79f),
	.w7(32'h3a629960),
	.w8(32'hbae25856),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66bd30),
	.w1(32'h3ba8d298),
	.w2(32'h3c0c8048),
	.w3(32'hbb84f1ea),
	.w4(32'hbc13dc05),
	.w5(32'hbb76bb59),
	.w6(32'h3b234c4b),
	.w7(32'h3a8a2a99),
	.w8(32'hbbaeb907),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7bd43),
	.w1(32'h3b4af23a),
	.w2(32'hbb1e1f7d),
	.w3(32'hbbfb4899),
	.w4(32'hba355b4f),
	.w5(32'hbbbdb3e3),
	.w6(32'h3b93f7e7),
	.w7(32'hba590ce7),
	.w8(32'hba281d6b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb149f14),
	.w1(32'hbb2b5d1e),
	.w2(32'h3a20920e),
	.w3(32'hbb2a9294),
	.w4(32'hba8610af),
	.w5(32'hbb83a213),
	.w6(32'h3ba2574e),
	.w7(32'h3a31e149),
	.w8(32'h3a59c06c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8510d),
	.w1(32'h3b3d3f91),
	.w2(32'h3995e2b6),
	.w3(32'hbb946942),
	.w4(32'h3b1963af),
	.w5(32'hba92f87d),
	.w6(32'h3b528b2c),
	.w7(32'hba88a020),
	.w8(32'hbb1dcc43),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08a021),
	.w1(32'hbb5bff25),
	.w2(32'h3bc32ff2),
	.w3(32'hbad81fd6),
	.w4(32'hbc0de7bb),
	.w5(32'hbbf3746d),
	.w6(32'h3af61960),
	.w7(32'h3c0f7b9c),
	.w8(32'h3b2a5f22),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb943262),
	.w1(32'hbb3dadf6),
	.w2(32'hbaa71f37),
	.w3(32'hbbceef4e),
	.w4(32'hbaa54f55),
	.w5(32'hbb7a8181),
	.w6(32'hbaceb4af),
	.w7(32'hbb49377e),
	.w8(32'hbb0e8693),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83ae7e),
	.w1(32'h39ff4132),
	.w2(32'hbb6e5aa3),
	.w3(32'hbb3aae80),
	.w4(32'hb929cf00),
	.w5(32'hbaf54a48),
	.w6(32'hb9863ac8),
	.w7(32'hbbbc51de),
	.w8(32'hbb8fb506),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b531d),
	.w1(32'h3b3a3c3a),
	.w2(32'hbbc8a7fc),
	.w3(32'hbb5aeaac),
	.w4(32'h3bb6fdbc),
	.w5(32'hbb9242e7),
	.w6(32'h3c371b24),
	.w7(32'hba92e8eb),
	.w8(32'hb9ba7898),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf7310),
	.w1(32'h3b4d3297),
	.w2(32'h3bace84d),
	.w3(32'hbb5855e9),
	.w4(32'h38ce9a94),
	.w5(32'h3ab37e1c),
	.w6(32'h3bfc3a85),
	.w7(32'h3c0fa461),
	.w8(32'h3b77511c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad24b22),
	.w1(32'hbb30602e),
	.w2(32'hba0e770a),
	.w3(32'hb972a03c),
	.w4(32'hbb084274),
	.w5(32'hbb219095),
	.w6(32'hb89b3ee5),
	.w7(32'hbae0ede3),
	.w8(32'hbb2fdc47),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7072c0),
	.w1(32'hbb04b704),
	.w2(32'hb9b23e6f),
	.w3(32'hbb7d74c9),
	.w4(32'hba798d6c),
	.w5(32'hbb448236),
	.w6(32'h3ab9f27b),
	.w7(32'hba9303cf),
	.w8(32'hbaf6df19),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72bb14),
	.w1(32'h3c04d700),
	.w2(32'h3b617d39),
	.w3(32'hbb8d8146),
	.w4(32'h3ba70acb),
	.w5(32'h3ad74d85),
	.w6(32'h3bc9d9eb),
	.w7(32'h3b24f8bd),
	.w8(32'h3ae36d19),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae759ae),
	.w1(32'hbc01d99d),
	.w2(32'hba3a689d),
	.w3(32'hb9833613),
	.w4(32'hbaf99304),
	.w5(32'hbb87314d),
	.w6(32'hbbc55f0e),
	.w7(32'h3a730f18),
	.w8(32'h3be95d96),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16c1f3),
	.w1(32'hba5eb4a4),
	.w2(32'hbb18f1f4),
	.w3(32'h3b8b765c),
	.w4(32'h3a8cf35f),
	.w5(32'h3b966760),
	.w6(32'hbc335543),
	.w7(32'hbbc57f64),
	.w8(32'hbbb3bc5a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f0c71),
	.w1(32'hbaee3d67),
	.w2(32'hba60ea33),
	.w3(32'h3b80ef79),
	.w4(32'hba80650e),
	.w5(32'hbb2c24ac),
	.w6(32'h3afc5c93),
	.w7(32'hba37d74a),
	.w8(32'hbaecef11),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6b5a),
	.w1(32'h3bbf6f8e),
	.w2(32'h3b7e07ea),
	.w3(32'hba6354db),
	.w4(32'h3bf11cf9),
	.w5(32'h3c0e8c6a),
	.w6(32'hbb6ff704),
	.w7(32'h38a7de44),
	.w8(32'hbba198c2),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec5da0),
	.w1(32'h3bda5d55),
	.w2(32'h3bd4f73f),
	.w3(32'h3b595ce6),
	.w4(32'h3bad93fc),
	.w5(32'h3bf31056),
	.w6(32'hba5a344f),
	.w7(32'h3b82858e),
	.w8(32'h3aefef47),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb0ba4),
	.w1(32'hbba9b592),
	.w2(32'hbb0c0858),
	.w3(32'h3bb54ce7),
	.w4(32'hbb431cd9),
	.w5(32'hbbc45996),
	.w6(32'h3616da44),
	.w7(32'hbb756188),
	.w8(32'hbb5db892),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0108e3),
	.w1(32'h3b9d071b),
	.w2(32'h3b710f1e),
	.w3(32'hbbf02e73),
	.w4(32'h3b962074),
	.w5(32'h3bd4348c),
	.w6(32'h3a5e0d79),
	.w7(32'h3ba836f8),
	.w8(32'h3b03553f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fe316),
	.w1(32'h3adf6156),
	.w2(32'h3ab0ed52),
	.w3(32'h3b8d443b),
	.w4(32'hba109652),
	.w5(32'hb967918f),
	.w6(32'h3bee00fb),
	.w7(32'h3bd97401),
	.w8(32'h3b2ef278),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada6f3e),
	.w1(32'hba2a5d9a),
	.w2(32'hbabb0105),
	.w3(32'hba5df7c5),
	.w4(32'h3ab5ad74),
	.w5(32'h3b24204f),
	.w6(32'hbba4af99),
	.w7(32'hbb863685),
	.w8(32'hbbb91fa1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7abc6e),
	.w1(32'hb80d6d43),
	.w2(32'h3a69e6e9),
	.w3(32'hb8c40081),
	.w4(32'hb9b0e4fe),
	.w5(32'hbaafeca6),
	.w6(32'h3b47c23c),
	.w7(32'h388c74f7),
	.w8(32'hba1d9623),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359972),
	.w1(32'h3c6ecaba),
	.w2(32'h3a2d8c3c),
	.w3(32'hbb65b364),
	.w4(32'h3c7d0db8),
	.w5(32'h3c772491),
	.w6(32'hb98e7d91),
	.w7(32'h3ad73e0a),
	.w8(32'h3bf2a5a3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4dbf2),
	.w1(32'h3c4a7d49),
	.w2(32'h3abe9e5e),
	.w3(32'h3cbd7eca),
	.w4(32'h3c249696),
	.w5(32'h3baf5ccf),
	.w6(32'h3c276aa8),
	.w7(32'h3b5bb0c9),
	.w8(32'h3b9869ee),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c084fd2),
	.w1(32'h3ba19140),
	.w2(32'h3aed591b),
	.w3(32'h3c167248),
	.w4(32'h3bbfa770),
	.w5(32'h3b8bc21e),
	.w6(32'hba8ca730),
	.w7(32'h3a0e1f1d),
	.w8(32'h3a4d171d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4b406),
	.w1(32'h3b94c572),
	.w2(32'h3b98bf79),
	.w3(32'h3b350379),
	.w4(32'h3bf880d5),
	.w5(32'h3c20ea9f),
	.w6(32'hb9dc631d),
	.w7(32'h3b746a48),
	.w8(32'hb9ed4dfe),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb960807),
	.w1(32'h3a5de670),
	.w2(32'h3b315445),
	.w3(32'h3b8d0a98),
	.w4(32'h3a2ed852),
	.w5(32'h3a5aa2c7),
	.w6(32'h3bab9562),
	.w7(32'h3b9614c6),
	.w8(32'hba003e15),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c03c2),
	.w1(32'hba229dc0),
	.w2(32'h3acf4d9d),
	.w3(32'hbb409f62),
	.w4(32'h38bb74a9),
	.w5(32'hba249590),
	.w6(32'h3b5002db),
	.w7(32'h3ab5327d),
	.w8(32'h3ab1a074),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa518a),
	.w1(32'hbaa3ea82),
	.w2(32'h3a47298c),
	.w3(32'hbaed340f),
	.w4(32'hba293b45),
	.w5(32'hbb7d8165),
	.w6(32'h3bc5797e),
	.w7(32'h3b050b86),
	.w8(32'h3aa1c353),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafefbb),
	.w1(32'h3c015720),
	.w2(32'hbbaf4ded),
	.w3(32'hbba48228),
	.w4(32'h3c07c7a8),
	.w5(32'h3b042ba6),
	.w6(32'h3b5a3a07),
	.w7(32'h3a25e31b),
	.w8(32'h3b8fef36),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b558d99),
	.w1(32'h399af3de),
	.w2(32'hba6005c6),
	.w3(32'h3ba4184d),
	.w4(32'hba75b1bf),
	.w5(32'hbb1d8033),
	.w6(32'hb9cd6caa),
	.w7(32'hbb40d316),
	.w8(32'hbb9cfb5f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0891d),
	.w1(32'hbb9613bf),
	.w2(32'hbba23819),
	.w3(32'hbb1c47d7),
	.w4(32'hbb687cd2),
	.w5(32'hbc1e1c5e),
	.w6(32'hbb134f24),
	.w7(32'hbc1736df),
	.w8(32'hbbf9bd67),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e6572),
	.w1(32'hba3df6e6),
	.w2(32'hb9e12908),
	.w3(32'hbc215d92),
	.w4(32'h3b2ce96b),
	.w5(32'hba2ed691),
	.w6(32'hbb073b33),
	.w7(32'hba1dc93e),
	.w8(32'hbb887722),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c4c0e),
	.w1(32'hb9b96915),
	.w2(32'h3a177de9),
	.w3(32'hbbaa1440),
	.w4(32'hbb2aaa09),
	.w5(32'hba90c10e),
	.w6(32'hba18f3f6),
	.w7(32'h3ae60bd6),
	.w8(32'hbb84a542),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b4b85),
	.w1(32'hb988cc9e),
	.w2(32'hbb80e45d),
	.w3(32'hbb4930af),
	.w4(32'hba94d377),
	.w5(32'hbbc9152f),
	.w6(32'h3bce6cd3),
	.w7(32'h38ed3c2b),
	.w8(32'hb9ed4e00),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb908fe8),
	.w1(32'h3bc295d3),
	.w2(32'h399413b4),
	.w3(32'hba83e6ad),
	.w4(32'h3b8ba262),
	.w5(32'h3a92c1d7),
	.w6(32'h3bf1cf77),
	.w7(32'h3b7068e0),
	.w8(32'h39943490),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5ad8e),
	.w1(32'h3939a92c),
	.w2(32'hba829bba),
	.w3(32'h3ae353c3),
	.w4(32'h3b3534c5),
	.w5(32'hba1bc02b),
	.w6(32'h3b492719),
	.w7(32'h3b960c5f),
	.w8(32'hba226b4e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1416ec),
	.w1(32'h3c041535),
	.w2(32'h3bab81c1),
	.w3(32'hbb6c1efb),
	.w4(32'h3bc630df),
	.w5(32'h3be74dd4),
	.w6(32'h3b7ecd8d),
	.w7(32'h3b9d168f),
	.w8(32'h3ad55389),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0832a6),
	.w1(32'hbb9b3c71),
	.w2(32'hba8fee8c),
	.w3(32'h3bb63349),
	.w4(32'hbb4d8523),
	.w5(32'hbbaf09e4),
	.w6(32'h3ad4846a),
	.w7(32'hbaf63e17),
	.w8(32'hba9193cb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec9f15),
	.w1(32'h3b055517),
	.w2(32'h3a96fc58),
	.w3(32'hbbd74fb7),
	.w4(32'h3b93df67),
	.w5(32'h3b77b029),
	.w6(32'hbb20dd05),
	.w7(32'h3b1cc008),
	.w8(32'h39232abe),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50223d),
	.w1(32'hbb274f50),
	.w2(32'hb9e44cda),
	.w3(32'h3a0ec505),
	.w4(32'hbaf3471c),
	.w5(32'hbae9f6f3),
	.w6(32'h3b198a28),
	.w7(32'hba407328),
	.w8(32'hba5dfd54),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb16b3),
	.w1(32'h3bf71b23),
	.w2(32'hb89a3e0a),
	.w3(32'hbb8ea01f),
	.w4(32'h3b091e21),
	.w5(32'hba778934),
	.w6(32'h3be1b505),
	.w7(32'h3a9679ff),
	.w8(32'hbb002e24),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8d568),
	.w1(32'h3c0cce90),
	.w2(32'hba27f325),
	.w3(32'h3bac9700),
	.w4(32'h3c1f1db4),
	.w5(32'h3c1ef312),
	.w6(32'hbb05d634),
	.w7(32'hb9ca9c51),
	.w8(32'h3b4d039e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e3774),
	.w1(32'h3abd2b63),
	.w2(32'hbac273fc),
	.w3(32'h3c6e7557),
	.w4(32'h3b5b2039),
	.w5(32'h3b127d29),
	.w6(32'hbae20caa),
	.w7(32'hbb15c7f7),
	.w8(32'hbb4e8473),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fe76),
	.w1(32'hbaa6a32b),
	.w2(32'hbb09ac82),
	.w3(32'hb94d6904),
	.w4(32'h398ca92c),
	.w5(32'hba8e6e91),
	.w6(32'h3b830107),
	.w7(32'h3b08b286),
	.w8(32'h3a6ce01a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393360eb),
	.w1(32'hbb68dd11),
	.w2(32'h3b24e238),
	.w3(32'hbad2b2bc),
	.w4(32'hbb69d450),
	.w5(32'h39deff90),
	.w6(32'hbaadad9c),
	.w7(32'h3b26e232),
	.w8(32'hbacad040),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb080e00),
	.w1(32'h3aa15794),
	.w2(32'hbaeb3e35),
	.w3(32'hb913297b),
	.w4(32'hbb209c85),
	.w5(32'hbb7441a6),
	.w6(32'h3b9b675a),
	.w7(32'h3b5f14fd),
	.w8(32'hb80905d4),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb285ab6),
	.w1(32'hbc04feab),
	.w2(32'hbb1f7bec),
	.w3(32'hbb8404c0),
	.w4(32'hbbd7da81),
	.w5(32'hbc10aa70),
	.w6(32'hbbb8f447),
	.w7(32'hbc06fe98),
	.w8(32'hbc09b08c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2879a9),
	.w1(32'h3c82aaa3),
	.w2(32'h3a2a7e3d),
	.w3(32'hbc1353ab),
	.w4(32'h3c8921f1),
	.w5(32'h3be20fa3),
	.w6(32'h3c56ef0b),
	.w7(32'h3c098d6b),
	.w8(32'h3c26ff0e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc70374),
	.w1(32'h3b0952fa),
	.w2(32'h3b545285),
	.w3(32'h3c04a09b),
	.w4(32'h3ac0b1d0),
	.w5(32'h3ba91f67),
	.w6(32'hbbd97f1d),
	.w7(32'hba8cf719),
	.w8(32'hbb5f386e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0e0c4),
	.w1(32'hbb53136a),
	.w2(32'hba74cbe8),
	.w3(32'h3b9d3839),
	.w4(32'hbb038cc1),
	.w5(32'hbbafbfc4),
	.w6(32'h3aadf136),
	.w7(32'hbb1fb3ef),
	.w8(32'hbb61553a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb2157),
	.w1(32'hbb85ff3f),
	.w2(32'hba996a46),
	.w3(32'hbbbbb233),
	.w4(32'hbb235b6a),
	.w5(32'hbbae47a8),
	.w6(32'h39b62fb7),
	.w7(32'hbb364a58),
	.w8(32'hbb273e9f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe485db),
	.w1(32'hbb495972),
	.w2(32'hba1cf1ed),
	.w3(32'hbbbf6ac0),
	.w4(32'hba946327),
	.w5(32'hbb53dea9),
	.w6(32'h3adb62cc),
	.w7(32'hba55fabb),
	.w8(32'hbae08045),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5f14c),
	.w1(32'h3bce9454),
	.w2(32'h3baaf40c),
	.w3(32'hbb8662b4),
	.w4(32'h3bd16be5),
	.w5(32'h3be37ec1),
	.w6(32'h3b8e70e9),
	.w7(32'h3b9467ff),
	.w8(32'h3b22e312),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befca5a),
	.w1(32'h39e9490e),
	.w2(32'h3b7b2bd3),
	.w3(32'h3bd28b0e),
	.w4(32'h3b2ffab5),
	.w5(32'h3b9e97fc),
	.w6(32'hbaae3566),
	.w7(32'h3bbf0830),
	.w8(32'h3a4365d3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc071257),
	.w1(32'h3906cd25),
	.w2(32'h395d827e),
	.w3(32'h3b8c0f6f),
	.w4(32'h3aa0a274),
	.w5(32'hbb842c84),
	.w6(32'h3c2a3d75),
	.w7(32'h3b08437d),
	.w8(32'h3b942093),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a24ae),
	.w1(32'hb9e9d724),
	.w2(32'hbb233b90),
	.w3(32'hbb435085),
	.w4(32'h3a8482b0),
	.w5(32'h3ae1f38d),
	.w6(32'hb94ff67d),
	.w7(32'h3afda51d),
	.w8(32'hbaa1bc6f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b043e8f),
	.w1(32'h3c0312b2),
	.w2(32'h3bf6a35e),
	.w3(32'h3b299097),
	.w4(32'hba780c9d),
	.w5(32'hbb1165a4),
	.w6(32'h3beb6554),
	.w7(32'h3c0a06fb),
	.w8(32'hbbad1934),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08943b),
	.w1(32'hbb23bb3c),
	.w2(32'hba1608bd),
	.w3(32'hbc1d2cd7),
	.w4(32'hba95f4a0),
	.w5(32'hbb580c3e),
	.w6(32'h3aca24f1),
	.w7(32'hbb417393),
	.w8(32'hbb91e1cd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe12ebc),
	.w1(32'h392fa690),
	.w2(32'hbab60bc2),
	.w3(32'hbbdb4e49),
	.w4(32'h39d262ce),
	.w5(32'hbac31945),
	.w6(32'h3b5398ef),
	.w7(32'h3acca658),
	.w8(32'hb9fc764f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68a706),
	.w1(32'hba421e41),
	.w2(32'hb9936fd8),
	.w3(32'hbb18390f),
	.w4(32'h3aa8a7bd),
	.w5(32'h3b31ac67),
	.w6(32'hbb72195c),
	.w7(32'hb906aeb8),
	.w8(32'h38897100),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b105951),
	.w1(32'hb93cfdbe),
	.w2(32'hb8be5769),
	.w3(32'h3b299823),
	.w4(32'hba31a73a),
	.w5(32'hba9fe3b3),
	.w6(32'h3a361799),
	.w7(32'hbaba7978),
	.w8(32'hbb0fb0ea),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb373dbe),
	.w1(32'h3b9bf2ed),
	.w2(32'h3b33d99d),
	.w3(32'hb9d80799),
	.w4(32'h3bcabe08),
	.w5(32'h3bb5275d),
	.w6(32'h3b031b80),
	.w7(32'h3b868b7a),
	.w8(32'h3b4f3466),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1c531),
	.w1(32'hba8bf140),
	.w2(32'h3ba98f69),
	.w3(32'h3b841ea5),
	.w4(32'h3b982376),
	.w5(32'h3bb9f745),
	.w6(32'h3b641fbe),
	.w7(32'h3b6a2509),
	.w8(32'h3a125c50),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80cac4),
	.w1(32'h3be670a9),
	.w2(32'h3c12e717),
	.w3(32'h39e51b6a),
	.w4(32'h3bbdbcb6),
	.w5(32'h3bd9d812),
	.w6(32'h3bba4606),
	.w7(32'h3c083a1e),
	.w8(32'h3bc172b2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bcc5c),
	.w1(32'h3a7ce8bc),
	.w2(32'hba31ce25),
	.w3(32'h3bfbad79),
	.w4(32'h3b5fe91c),
	.w5(32'h3b648402),
	.w6(32'h3b203278),
	.w7(32'h3ba56ad8),
	.w8(32'h3bd19d53),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c155a51),
	.w1(32'hbb0cdf73),
	.w2(32'h36dd625d),
	.w3(32'h3bfe3d32),
	.w4(32'hbac34991),
	.w5(32'hbb1c62fe),
	.w6(32'h39c41c8b),
	.w7(32'hbabf1e9e),
	.w8(32'hbb179dea),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb664d82),
	.w1(32'h3857b12b),
	.w2(32'h371fc353),
	.w3(32'hbb8b79d7),
	.w4(32'hbac9aaba),
	.w5(32'hba83632a),
	.w6(32'hb8fff2f7),
	.w7(32'h3a4edb4a),
	.w8(32'hbb0dae6b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16c2d2),
	.w1(32'hbb273102),
	.w2(32'hba341611),
	.w3(32'hbb1a1eae),
	.w4(32'hbaa14d73),
	.w5(32'hbb66e0ad),
	.w6(32'h39c9e9c2),
	.w7(32'hbb4d4457),
	.w8(32'hbbaf6f70),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc68e5e),
	.w1(32'hbb1b4575),
	.w2(32'h394ee27c),
	.w3(32'hbbcaffce),
	.w4(32'hbac62fcc),
	.w5(32'hbabb47f4),
	.w6(32'h3b40dca2),
	.w7(32'h3ad6f918),
	.w8(32'h3ac5a56b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a3b5),
	.w1(32'h3bfa968c),
	.w2(32'h3baca8ea),
	.w3(32'hbb22e9ec),
	.w4(32'h3c05bb1a),
	.w5(32'h3c2aeda6),
	.w6(32'hbb02a4cc),
	.w7(32'h3b38347c),
	.w8(32'h3b5e4e80),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c443361),
	.w1(32'hbb25a020),
	.w2(32'hb983ad0f),
	.w3(32'h3c4d7385),
	.w4(32'hbb0f32ab),
	.w5(32'hbb17a5b2),
	.w6(32'hbb948db8),
	.w7(32'hbb08a517),
	.w8(32'hbb351e34),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32f6f8),
	.w1(32'hbb7bd6da),
	.w2(32'hbbf5913e),
	.w3(32'hbb0b4900),
	.w4(32'hbabb3c0f),
	.w5(32'hbbbc3970),
	.w6(32'h3b01a7b3),
	.w7(32'hbb8214a3),
	.w8(32'hbaff93df),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc65405),
	.w1(32'h3b3179a2),
	.w2(32'hb882ae7f),
	.w3(32'hbb5efbb6),
	.w4(32'hba8ff52b),
	.w5(32'hbb2605f9),
	.w6(32'hbb123b6d),
	.w7(32'hbb4520c5),
	.w8(32'hbb88070d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f89b01),
	.w1(32'hbb20b806),
	.w2(32'hbb315412),
	.w3(32'hbb730639),
	.w4(32'hba94f75d),
	.w5(32'hbb6d55ab),
	.w6(32'hb998905e),
	.w7(32'hba9b1825),
	.w8(32'hbb29d7c3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9deaa8),
	.w1(32'h3b64c305),
	.w2(32'h3b9ac277),
	.w3(32'hbbcf8981),
	.w4(32'hba682b07),
	.w5(32'h3aa64d99),
	.w6(32'h3ad36d7f),
	.w7(32'h3bd96223),
	.w8(32'hb9b1f3f8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968664c),
	.w1(32'h3c040973),
	.w2(32'hbb0dfbf7),
	.w3(32'hbae95190),
	.w4(32'h3c1199c0),
	.w5(32'hb9bc636e),
	.w6(32'h3c3f1563),
	.w7(32'h3aefb13e),
	.w8(32'hbaadada5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c84d16),
	.w1(32'hba6a2697),
	.w2(32'hba887126),
	.w3(32'hbac46c30),
	.w4(32'h3a76df5d),
	.w5(32'h3b87d20e),
	.w6(32'hbb744359),
	.w7(32'h39d758b9),
	.w8(32'hbb9df696),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6276db),
	.w1(32'hbbc44fc8),
	.w2(32'hbbd12d9b),
	.w3(32'h3977ebfe),
	.w4(32'hbbb32a66),
	.w5(32'hbc180949),
	.w6(32'hbb528efb),
	.w7(32'hbc10dcd6),
	.w8(32'hbc0a616c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f6222),
	.w1(32'h3aaf42f7),
	.w2(32'hbbf9b9fd),
	.w3(32'hbc1a3d94),
	.w4(32'h3b132660),
	.w5(32'hbbef9b28),
	.w6(32'h388d1c6f),
	.w7(32'h398ed2dc),
	.w8(32'hbc04174d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f63a5),
	.w1(32'h3bd05e92),
	.w2(32'h3beec08f),
	.w3(32'hbc425d03),
	.w4(32'h39e43dbb),
	.w5(32'hbace7fc8),
	.w6(32'h398ab9df),
	.w7(32'h3ab3ca15),
	.w8(32'hbc0eef61),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb95a2c),
	.w1(32'hb851ea20),
	.w2(32'h398af7d8),
	.w3(32'hbc028af3),
	.w4(32'h3acb076d),
	.w5(32'hbbc9df5a),
	.w6(32'h3c7feff9),
	.w7(32'h3b4eb539),
	.w8(32'h3be35a96),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeb581),
	.w1(32'hbb20830d),
	.w2(32'hba82a439),
	.w3(32'hbb9882db),
	.w4(32'h38482135),
	.w5(32'hbbb1cee1),
	.w6(32'h3aa567b2),
	.w7(32'hbb84386f),
	.w8(32'hbb7933c0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb150a6),
	.w1(32'h392608b8),
	.w2(32'h3964504f),
	.w3(32'hbbb4d7cf),
	.w4(32'h3a90e0cd),
	.w5(32'hbb402a7a),
	.w6(32'h3bff2f88),
	.w7(32'h3aaff016),
	.w8(32'h3b52c2a1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e1176),
	.w1(32'hb88637f9),
	.w2(32'h3a5cee89),
	.w3(32'hbb0cb61e),
	.w4(32'hb9d8d442),
	.w5(32'hbb0ce9af),
	.w6(32'h3a6cfea4),
	.w7(32'hbabf4229),
	.w8(32'hbac0a1ac),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dd0fe),
	.w1(32'h3aec7fad),
	.w2(32'hbac25964),
	.w3(32'hbaed6d56),
	.w4(32'hbac7c5a7),
	.w5(32'hbaf87733),
	.w6(32'hba0069d3),
	.w7(32'hbb84cf57),
	.w8(32'hbb9c2bc1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bd150),
	.w1(32'hbb37e8b7),
	.w2(32'h39d1eb85),
	.w3(32'h3774549b),
	.w4(32'hbae1dd75),
	.w5(32'hbaac8357),
	.w6(32'h3aed88c6),
	.w7(32'h3a344b2e),
	.w8(32'h38f6d77b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25db96),
	.w1(32'hb8aea451),
	.w2(32'h38bc96a0),
	.w3(32'hbb40ca44),
	.w4(32'h3a4a175e),
	.w5(32'hbb53c645),
	.w6(32'h3c08a9d2),
	.w7(32'h3af5b95c),
	.w8(32'h3b7433cb),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5161ca),
	.w1(32'h3c325f53),
	.w2(32'h39a407ad),
	.w3(32'hbb2b3ba9),
	.w4(32'h3c410afd),
	.w5(32'h3bd38a32),
	.w6(32'h3bc04cc1),
	.w7(32'h3827711f),
	.w8(32'h3ac89679),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cf7da),
	.w1(32'hbbeee6ff),
	.w2(32'hbb90c261),
	.w3(32'h3c1245e6),
	.w4(32'hbba5690d),
	.w5(32'hbc02b67d),
	.w6(32'hbb95daf4),
	.w7(32'hbbef9629),
	.w8(32'hbbdb9a70),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38be44),
	.w1(32'h3bb5f89c),
	.w2(32'hba72a255),
	.w3(32'hbc090ab3),
	.w4(32'h3b2f9251),
	.w5(32'hb8a73de7),
	.w6(32'h3bdeaabf),
	.w7(32'h3b15e23c),
	.w8(32'h3b7c8bc8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd7e5),
	.w1(32'hbbbb835b),
	.w2(32'hbb831770),
	.w3(32'h3ba47536),
	.w4(32'hbb91fa53),
	.w5(32'hbc1b811c),
	.w6(32'hbb8f45e1),
	.w7(32'hbc04e799),
	.w8(32'hbc080d07),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4460df),
	.w1(32'hba0c689d),
	.w2(32'hbb462585),
	.w3(32'hbc276ed3),
	.w4(32'hbb090fa3),
	.w5(32'hb8c2b70f),
	.w6(32'hbb49bb4d),
	.w7(32'hbb19c80b),
	.w8(32'hbb0cf13c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa555c),
	.w1(32'hba4efdad),
	.w2(32'h3ac45b15),
	.w3(32'h3a70ff9a),
	.w4(32'hba589572),
	.w5(32'hb9afa6e7),
	.w6(32'h3b5d433e),
	.w7(32'hba2b77b3),
	.w8(32'hbb5327d1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd7512),
	.w1(32'h38f68abc),
	.w2(32'h3991e0b3),
	.w3(32'hbbbffa22),
	.w4(32'h3ab0fe7d),
	.w5(32'hbb9470d4),
	.w6(32'h3c41080b),
	.w7(32'h3b1a30f1),
	.w8(32'h3ba8a411),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1aad),
	.w1(32'hba80c921),
	.w2(32'h3a9700c7),
	.w3(32'hbb5eb1df),
	.w4(32'h3a825362),
	.w5(32'hbb1b0ec0),
	.w6(32'h3ba4ff05),
	.w7(32'h3a52c027),
	.w8(32'h3aa3025a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb516bbd),
	.w1(32'hbae1b9de),
	.w2(32'h39e46a92),
	.w3(32'hbb33e2a8),
	.w4(32'h39162b8f),
	.w5(32'hbb419429),
	.w6(32'h3b9a0db1),
	.w7(32'hb9ea37f2),
	.w8(32'h3a8287ff),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f91bb),
	.w1(32'h3b772d7d),
	.w2(32'h3be42df6),
	.w3(32'hbb3aaf63),
	.w4(32'hbaa121dc),
	.w5(32'h3b53861d),
	.w6(32'h3b4543f7),
	.w7(32'h39c82520),
	.w8(32'h3b3acf50),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c2785),
	.w1(32'hba3b4975),
	.w2(32'hbb9d458d),
	.w3(32'h39f70659),
	.w4(32'h3b041666),
	.w5(32'hba4d3588),
	.w6(32'hbb829677),
	.w7(32'hb99163a5),
	.w8(32'hbbc31cc7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca27e),
	.w1(32'hbb950624),
	.w2(32'hbbcb21a1),
	.w3(32'hbbfbc2a0),
	.w4(32'hb9f82f91),
	.w5(32'hbb92a846),
	.w6(32'hba003282),
	.w7(32'hbbc47160),
	.w8(32'hbbc14459),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b75e2),
	.w1(32'hbb4ff6ab),
	.w2(32'hbbaac577),
	.w3(32'hbbab58d5),
	.w4(32'hbaa069f0),
	.w5(32'hbba10b60),
	.w6(32'hbae38ebe),
	.w7(32'hbb966f77),
	.w8(32'hbab26c0d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6b885),
	.w1(32'hbb60308d),
	.w2(32'h390f2973),
	.w3(32'hbb95a526),
	.w4(32'hbaec9f65),
	.w5(32'hbb98c315),
	.w6(32'h3b96d94f),
	.w7(32'h3946d75d),
	.w8(32'h39b6dc45),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb4d7f),
	.w1(32'h3ad4868f),
	.w2(32'h3b531626),
	.w3(32'hbbbf6066),
	.w4(32'hbab3b846),
	.w5(32'hba9df0d6),
	.w6(32'hbb487b01),
	.w7(32'hbb77d7e8),
	.w8(32'hbbd85d46),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba322f7),
	.w1(32'hbbbf2835),
	.w2(32'hbbbf6b33),
	.w3(32'hbb4b2e7f),
	.w4(32'hbb371f5d),
	.w5(32'hbc0cf15b),
	.w6(32'hbaa5d633),
	.w7(32'hbc2aff1e),
	.w8(32'hbc0f6c04),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc398560),
	.w1(32'hbb436b76),
	.w2(32'hbab2fdfd),
	.w3(32'hbc4c380c),
	.w4(32'hbb18689c),
	.w5(32'hbb7cbb10),
	.w6(32'h3ab73c5d),
	.w7(32'hbaeed452),
	.w8(32'hbb0fe2f8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4f62),
	.w1(32'h37659476),
	.w2(32'h364dd640),
	.w3(32'hbbb7e676),
	.w4(32'h3705a925),
	.w5(32'hb631458b),
	.w6(32'h37c1b0ac),
	.w7(32'hb68c2047),
	.w8(32'hb6e2f40a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b7c6c2),
	.w1(32'hb789dda0),
	.w2(32'hb7188f76),
	.w3(32'hb66d135e),
	.w4(32'hb7c2b52d),
	.w5(32'hb75b427c),
	.w6(32'h36ba0148),
	.w7(32'h3789692c),
	.w8(32'h36b90c87),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule