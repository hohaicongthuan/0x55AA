module layer_8_featuremap_189(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17fae0),
	.w1(32'hbb75849a),
	.w2(32'h3b85ba68),
	.w3(32'h3b761c40),
	.w4(32'hbb23b695),
	.w5(32'h3b795253),
	.w6(32'h3ade96d8),
	.w7(32'hbace137e),
	.w8(32'hbb200da0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b9cda),
	.w1(32'hba112f61),
	.w2(32'hbb2d3d38),
	.w3(32'h3ae1ce9c),
	.w4(32'h39e7dd9d),
	.w5(32'hba963848),
	.w6(32'hbae315bc),
	.w7(32'hbb21287b),
	.w8(32'hbba89bc4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d5aa6),
	.w1(32'hba33882b),
	.w2(32'hb974f953),
	.w3(32'hbae124c8),
	.w4(32'hbb1ad9a3),
	.w5(32'hbb0f2bd0),
	.w6(32'hbb68e461),
	.w7(32'hbb0057c3),
	.w8(32'hbb22093f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f1009),
	.w1(32'h3b871b5c),
	.w2(32'h3bbf9209),
	.w3(32'hbb8130af),
	.w4(32'h3b46b97a),
	.w5(32'h3bb1c712),
	.w6(32'h3c2a72e4),
	.w7(32'h3bb998ab),
	.w8(32'h3c0ff7a9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86b9b8),
	.w1(32'hb98edf5a),
	.w2(32'hbaac231f),
	.w3(32'h3b67e8d1),
	.w4(32'hbacab5fd),
	.w5(32'hbb882d68),
	.w6(32'h3aaf0f7b),
	.w7(32'h3a485713),
	.w8(32'h3af952fe),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b834524),
	.w1(32'h3b80896d),
	.w2(32'hbb048ace),
	.w3(32'hbad77198),
	.w4(32'hbbb9b889),
	.w5(32'hbb49fb24),
	.w6(32'h3bcc555a),
	.w7(32'h3afc1f82),
	.w8(32'h3a277b65),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc076b),
	.w1(32'hba55c304),
	.w2(32'hb91b3116),
	.w3(32'h3a3d10cf),
	.w4(32'hbaf6b58f),
	.w5(32'hbb04faf8),
	.w6(32'h3a8b1158),
	.w7(32'h394f3181),
	.w8(32'h3a51fd01),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4f775),
	.w1(32'hbaef7437),
	.w2(32'h3b3d94bf),
	.w3(32'hbb1c969e),
	.w4(32'hba878e00),
	.w5(32'h3aa77c5c),
	.w6(32'hbac26068),
	.w7(32'h3ae165eb),
	.w8(32'h3ac2ae4d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8728b5),
	.w1(32'hbb8a0378),
	.w2(32'hbbb48ad5),
	.w3(32'h3ade6924),
	.w4(32'hbb634e6e),
	.w5(32'hbbc6c276),
	.w6(32'hba8f8869),
	.w7(32'hbaac39f0),
	.w8(32'hba6b9a2e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc543efc),
	.w1(32'hbbc9f0c8),
	.w2(32'hb9824d01),
	.w3(32'hbbbd0b99),
	.w4(32'h3b8f2742),
	.w5(32'h3b9b9b62),
	.w6(32'hbc19c7f4),
	.w7(32'hbba21753),
	.w8(32'hbb99e7c2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9254a),
	.w1(32'hbb118817),
	.w2(32'h39a703a4),
	.w3(32'hba52b69a),
	.w4(32'h3a76f29b),
	.w5(32'h39fbe361),
	.w6(32'h3acc8898),
	.w7(32'h3b936b7a),
	.w8(32'hbad346e4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b36a3),
	.w1(32'hba780dc3),
	.w2(32'h399d1f2a),
	.w3(32'h3b245323),
	.w4(32'h3b318c25),
	.w5(32'hbadf1243),
	.w6(32'hb94a8c2b),
	.w7(32'h3a3f0bff),
	.w8(32'hbb416188),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c90031),
	.w1(32'hbaf0604c),
	.w2(32'h3b0214cd),
	.w3(32'hbb1d87e4),
	.w4(32'h3a453558),
	.w5(32'h3b4e078b),
	.w6(32'hbb290395),
	.w7(32'h3a097a43),
	.w8(32'hbafeacf1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae108ed),
	.w1(32'hbb70a5ee),
	.w2(32'hbbab1dd2),
	.w3(32'h3b466d53),
	.w4(32'hbac474ac),
	.w5(32'hbb242573),
	.w6(32'hbb311938),
	.w7(32'hbb3e4f79),
	.w8(32'hbafe0f4a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1a0ce),
	.w1(32'h3c39e84b),
	.w2(32'h3c2e0cbf),
	.w3(32'hba1f860c),
	.w4(32'h3c58913c),
	.w5(32'h3c74b210),
	.w6(32'h3c00e489),
	.w7(32'h3badac4b),
	.w8(32'h3baaaacb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c203210),
	.w1(32'hbb0c069c),
	.w2(32'hb9ce956f),
	.w3(32'h3c5244e3),
	.w4(32'h39d1e4d0),
	.w5(32'h3a87f377),
	.w6(32'hbaa6af74),
	.w7(32'h391d77c7),
	.w8(32'hbb8b8f12),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98b069),
	.w1(32'hbb4dd61b),
	.w2(32'h3a86dc07),
	.w3(32'hbbc7c7b6),
	.w4(32'hbb91b10c),
	.w5(32'h3953b61b),
	.w6(32'hbbb53b0c),
	.w7(32'hbb5edb8b),
	.w8(32'h3a68907b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94028f3),
	.w1(32'h3b6a52c0),
	.w2(32'h3aa9f719),
	.w3(32'h3bfc3fc9),
	.w4(32'h3c2fe3b7),
	.w5(32'hbaedc3ff),
	.w6(32'h3b9c2659),
	.w7(32'h3c05f62f),
	.w8(32'h3b0959f0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc812a5b),
	.w1(32'h3b42482e),
	.w2(32'h3ab74385),
	.w3(32'h3c1d4d48),
	.w4(32'h3b5a1fd5),
	.w5(32'h3b9a0a3e),
	.w6(32'h3aa64b1a),
	.w7(32'hbb91bc4c),
	.w8(32'hbc5a081d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b562339),
	.w1(32'h3b0d6517),
	.w2(32'h3b301ab8),
	.w3(32'hbbbbc286),
	.w4(32'hbb0faaed),
	.w5(32'hba14065d),
	.w6(32'hbb308346),
	.w7(32'hba246d46),
	.w8(32'h39eb6ff5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1c313),
	.w1(32'h3b9294d4),
	.w2(32'h3b8d951d),
	.w3(32'h3b380b8f),
	.w4(32'hbb953f7a),
	.w5(32'hbb2a1859),
	.w6(32'h3aa195b5),
	.w7(32'hbae23eea),
	.w8(32'hbb2b8a76),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d1fd6),
	.w1(32'h3a7504a2),
	.w2(32'h3b385122),
	.w3(32'hbb51d8d1),
	.w4(32'h3a4b88a2),
	.w5(32'h3ba95e4e),
	.w6(32'h3a0f3010),
	.w7(32'h3b5babae),
	.w8(32'h3b259d9c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc265b5e),
	.w1(32'hbbdba6c5),
	.w2(32'h3c00f4e3),
	.w3(32'h3aca80b1),
	.w4(32'h3a7724c6),
	.w5(32'h3be0adb9),
	.w6(32'hbbf18893),
	.w7(32'hbb95fa88),
	.w8(32'hbba099b3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ce251),
	.w1(32'hbab72dc5),
	.w2(32'h3ae96454),
	.w3(32'h3a43fcda),
	.w4(32'hbb88b354),
	.w5(32'hbb502ffd),
	.w6(32'hbacd9cb4),
	.w7(32'hbb0e05e4),
	.w8(32'hbb075fb0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5474cd),
	.w1(32'hbb516e13),
	.w2(32'hbaeed8fe),
	.w3(32'hbbcb6b53),
	.w4(32'hbbe81aeb),
	.w5(32'hbb90ea2d),
	.w6(32'h3b7f8e58),
	.w7(32'h3b511df0),
	.w8(32'h3b51675c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e6203),
	.w1(32'hbbdc8bea),
	.w2(32'hbb114d84),
	.w3(32'hba7d139d),
	.w4(32'h381b688e),
	.w5(32'hbb2bafc3),
	.w6(32'h3a3c917a),
	.w7(32'hb96ee2b0),
	.w8(32'hbab39768),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab96e2e),
	.w1(32'hbb1051d6),
	.w2(32'hbb406906),
	.w3(32'hbb3980aa),
	.w4(32'hbaffbb71),
	.w5(32'h39feb636),
	.w6(32'h3b64c561),
	.w7(32'h3ba9d2d2),
	.w8(32'h3bd1feed),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd138618),
	.w1(32'hbce7877a),
	.w2(32'h3c91c2c2),
	.w3(32'hbbd2a514),
	.w4(32'hbb73e8af),
	.w5(32'hbbc051c5),
	.w6(32'h3be1952b),
	.w7(32'h3bc2d8ca),
	.w8(32'hbba68fa6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64f75f),
	.w1(32'h3ac80014),
	.w2(32'h3aa0e94e),
	.w3(32'h3c015e14),
	.w4(32'h3adf4302),
	.w5(32'h3a8063e9),
	.w6(32'h3b91132a),
	.w7(32'h3afb2f82),
	.w8(32'hb5bb7e60),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b94d60),
	.w1(32'hbad873ab),
	.w2(32'hb8ee97f6),
	.w3(32'hbb2adb3d),
	.w4(32'h3c3f8c3d),
	.w5(32'h3c491578),
	.w6(32'hba8dccc5),
	.w7(32'hbac00a7b),
	.w8(32'hbb61a332),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb690178),
	.w1(32'hba06a65e),
	.w2(32'hbb67ef76),
	.w3(32'h3c1e2018),
	.w4(32'h3b0c674f),
	.w5(32'h3a5f6319),
	.w6(32'h3b585033),
	.w7(32'h3a59a47d),
	.w8(32'h3a84e540),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dc60e),
	.w1(32'hbb29d77b),
	.w2(32'hbb424473),
	.w3(32'hbb17a85c),
	.w4(32'hbb80c126),
	.w5(32'hbae26015),
	.w6(32'hbbe0d302),
	.w7(32'hbbd3ab96),
	.w8(32'hbbcd9f72),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49f765),
	.w1(32'h3b255d8f),
	.w2(32'h3b570c09),
	.w3(32'hbb15582d),
	.w4(32'h3b960469),
	.w5(32'hb994d987),
	.w6(32'h3c02dd79),
	.w7(32'h3b587be3),
	.w8(32'h3b9213eb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4ff94),
	.w1(32'hbacefc95),
	.w2(32'h3a92a236),
	.w3(32'h3a5f698b),
	.w4(32'hbb660783),
	.w5(32'hbacb2316),
	.w6(32'hbbcdfb25),
	.w7(32'hbb6f7446),
	.w8(32'hba61f8dd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7681d8),
	.w1(32'h3a7eb29d),
	.w2(32'h38826b89),
	.w3(32'hbacfcc73),
	.w4(32'h3a85c0d7),
	.w5(32'h389f2acb),
	.w6(32'hbb942679),
	.w7(32'hbaa21099),
	.w8(32'hbac74d54),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1651ca),
	.w1(32'hbbcdd13d),
	.w2(32'hbb81f138),
	.w3(32'hbafe5243),
	.w4(32'hbbb1d947),
	.w5(32'hbaa75e87),
	.w6(32'hb9b38d1a),
	.w7(32'hba03b16d),
	.w8(32'hbafa2568),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba982b13),
	.w1(32'h3aefbe2b),
	.w2(32'h3b2d1454),
	.w3(32'hbb175257),
	.w4(32'h39633139),
	.w5(32'h3ae955d5),
	.w6(32'h3b702d6e),
	.w7(32'h3b999635),
	.w8(32'h3bb9cb00),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e2e61),
	.w1(32'h3c1fd499),
	.w2(32'h3c0a7625),
	.w3(32'h3af6c014),
	.w4(32'h3c6a6835),
	.w5(32'h3c5ff980),
	.w6(32'h3c042123),
	.w7(32'h3ba6ba24),
	.w8(32'h3bb40ff8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be148bc),
	.w1(32'h3b6ef8eb),
	.w2(32'hbb66f283),
	.w3(32'h3c428a84),
	.w4(32'hb985ec32),
	.w5(32'h3a91f34f),
	.w6(32'h3a458b4e),
	.w7(32'h3994bab7),
	.w8(32'hb9f1638c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b991d6),
	.w1(32'hbb87f75f),
	.w2(32'hba93c75e),
	.w3(32'hbadc5cf1),
	.w4(32'hbb821615),
	.w5(32'hbb2f28f3),
	.w6(32'hba65906b),
	.w7(32'hbad75744),
	.w8(32'hb94b805e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23432b),
	.w1(32'h3bf2c5f2),
	.w2(32'h3bf3604c),
	.w3(32'h3c48d5e7),
	.w4(32'h3c5bc2c6),
	.w5(32'h3bd63ba2),
	.w6(32'h3c74d180),
	.w7(32'h3c08c67b),
	.w8(32'h3b725921),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56ffae),
	.w1(32'hba368a75),
	.w2(32'hba993f83),
	.w3(32'hbabfd5c0),
	.w4(32'hba80c08d),
	.w5(32'hbb5f7523),
	.w6(32'hbb55957c),
	.w7(32'hbb87cbfe),
	.w8(32'hbb0defbd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf49c4),
	.w1(32'hbabe5a04),
	.w2(32'hbb2d214f),
	.w3(32'hba927860),
	.w4(32'hbaf0030e),
	.w5(32'hbb84ad82),
	.w6(32'h3a394845),
	.w7(32'h3902ea9b),
	.w8(32'h3aec0f3a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e645ea),
	.w1(32'h3a20456b),
	.w2(32'hb94416f4),
	.w3(32'hb82f8fd4),
	.w4(32'h3b2e8297),
	.w5(32'h3b0af837),
	.w6(32'h3b22a9aa),
	.w7(32'hbb848007),
	.w8(32'hbb8462f0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3caa5b),
	.w1(32'hbb743ef4),
	.w2(32'h3b817857),
	.w3(32'hbb30374c),
	.w4(32'h3a061d26),
	.w5(32'h3b974db0),
	.w6(32'h3a70321e),
	.w7(32'hbb74d65d),
	.w8(32'hbb9efe35),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1879dd),
	.w1(32'hbba4194f),
	.w2(32'hbb0df0fa),
	.w3(32'hbaef129e),
	.w4(32'hbb571c68),
	.w5(32'hb96eacb0),
	.w6(32'hbbefa22b),
	.w7(32'hbc19bf0d),
	.w8(32'hbc3bc89a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5de14d),
	.w1(32'h3ad6e227),
	.w2(32'h3a93914b),
	.w3(32'hba4b8936),
	.w4(32'h3ab3b8ef),
	.w5(32'h3a2d1a08),
	.w6(32'h3b330cd9),
	.w7(32'h3a69683e),
	.w8(32'hb811de8e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b05dc),
	.w1(32'hbbf7913f),
	.w2(32'h3b6c6510),
	.w3(32'hbb89873c),
	.w4(32'hbb822331),
	.w5(32'hbb73ed5a),
	.w6(32'hbb95a00d),
	.w7(32'h3a6867c6),
	.w8(32'hbbf3bdbf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93bcb2),
	.w1(32'hbb561966),
	.w2(32'hbb700225),
	.w3(32'hbb8a933d),
	.w4(32'hbb4e3c27),
	.w5(32'h3a2a835e),
	.w6(32'hbb97500d),
	.w7(32'hbb07699c),
	.w8(32'hbac1cbaf),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4e1b3),
	.w1(32'h3b91d0ad),
	.w2(32'h3ab35e80),
	.w3(32'hbb425400),
	.w4(32'h3bf0d70a),
	.w5(32'h3b168ccb),
	.w6(32'h3b811c61),
	.w7(32'h3ba25ad8),
	.w8(32'h3b9042f1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2ffb3),
	.w1(32'h3af8efce),
	.w2(32'h39d06ad9),
	.w3(32'h3ba386ce),
	.w4(32'h3a8292d8),
	.w5(32'hba4ed937),
	.w6(32'h3955bca3),
	.w7(32'hbb1885d0),
	.w8(32'hbb56fbe4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26e8f1),
	.w1(32'hbb33d0ef),
	.w2(32'hbaafb3d3),
	.w3(32'h3a71b2fc),
	.w4(32'h3b17b5b9),
	.w5(32'h3b5f56c6),
	.w6(32'h3bc401bf),
	.w7(32'h39eb732f),
	.w8(32'hbab8dfcd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42a058),
	.w1(32'h3b93569d),
	.w2(32'h3b5ba134),
	.w3(32'hbadf031e),
	.w4(32'h3c370093),
	.w5(32'h3c329f16),
	.w6(32'hb7859902),
	.w7(32'hbb535af5),
	.w8(32'hbb971f63),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4248),
	.w1(32'hbb317b45),
	.w2(32'hb9cfbfd7),
	.w3(32'h3b9d5efc),
	.w4(32'h39c61252),
	.w5(32'hbab17a4a),
	.w6(32'hbbe7fdf7),
	.w7(32'hbb8188b6),
	.w8(32'hbbb436bc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a22de),
	.w1(32'h3afe63a9),
	.w2(32'h3a759034),
	.w3(32'hb96d0a35),
	.w4(32'h3bc2bff4),
	.w5(32'hb7d400ab),
	.w6(32'h3a7abf20),
	.w7(32'h39a970c4),
	.w8(32'h3b20538f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f70f4),
	.w1(32'hbbdb2afd),
	.w2(32'h3b3364c6),
	.w3(32'hbb81b890),
	.w4(32'h3b2a2335),
	.w5(32'hbadedd89),
	.w6(32'hbc497b9e),
	.w7(32'hbb8daf5b),
	.w8(32'hbbd371ef),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b490ce7),
	.w1(32'hbb351b24),
	.w2(32'hbb152cd4),
	.w3(32'h3b0fbe1c),
	.w4(32'hbb9efb08),
	.w5(32'hbbb71364),
	.w6(32'hbbd408d1),
	.w7(32'hbad79402),
	.w8(32'hba920aa3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb11f),
	.w1(32'hba66610c),
	.w2(32'h3b1803c5),
	.w3(32'hbb8c7a1d),
	.w4(32'hbafcc0dd),
	.w5(32'h3a25d43d),
	.w6(32'hb986ba33),
	.w7(32'h39b21261),
	.w8(32'hb7bde23d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277139),
	.w1(32'hbb509f45),
	.w2(32'h39e8e9b6),
	.w3(32'hbb8dbab6),
	.w4(32'hbade6e5b),
	.w5(32'h3ae10d9a),
	.w6(32'h383a1fd2),
	.w7(32'hbae1547d),
	.w8(32'hbb525196),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64ca66),
	.w1(32'hb7d7b2bc),
	.w2(32'h3b1db0b2),
	.w3(32'h3a8a6738),
	.w4(32'hba2fa799),
	.w5(32'h3bcaed6c),
	.w6(32'h39227c5b),
	.w7(32'h3bc040ff),
	.w8(32'h3b914225),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10d4ca),
	.w1(32'h3a2c199d),
	.w2(32'hbb5e479a),
	.w3(32'h3a82689f),
	.w4(32'hbb29f463),
	.w5(32'hba73c352),
	.w6(32'h3b875ed7),
	.w7(32'h3b530cc9),
	.w8(32'hb9892ff9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacad88d),
	.w1(32'h3b49fd29),
	.w2(32'h3b1641d5),
	.w3(32'hbacfd16b),
	.w4(32'h3b588258),
	.w5(32'h3b515bb0),
	.w6(32'h3c01a317),
	.w7(32'h3bc85be5),
	.w8(32'h3bb8c91b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8070c0),
	.w1(32'h398c5856),
	.w2(32'h3b4e4e0b),
	.w3(32'h3c11818a),
	.w4(32'h3c095272),
	.w5(32'h3b83edf2),
	.w6(32'h3bb85c94),
	.w7(32'h3b48755d),
	.w8(32'h3b672b03),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b719bed),
	.w1(32'h3934e099),
	.w2(32'hba2829d3),
	.w3(32'h3b878a84),
	.w4(32'hb96bb5e0),
	.w5(32'hba03043c),
	.w6(32'hb9dc7c26),
	.w7(32'hba880108),
	.w8(32'hbb0184d3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e438b),
	.w1(32'h3bc4c7aa),
	.w2(32'h3ba7c500),
	.w3(32'h392ba38c),
	.w4(32'h3c19e4a2),
	.w5(32'h3c20e412),
	.w6(32'h3ac5fad9),
	.w7(32'hbae9cba1),
	.w8(32'hbaeb472d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923fcd2),
	.w1(32'hbb211a0a),
	.w2(32'hbb9adc90),
	.w3(32'h3bd61204),
	.w4(32'hba210631),
	.w5(32'hba1fe8b0),
	.w6(32'hbb2de62f),
	.w7(32'hbb7b6921),
	.w8(32'hbb55e231),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7631462),
	.w1(32'h3a9e608f),
	.w2(32'h3afd33c3),
	.w3(32'hb99b94cb),
	.w4(32'hbb337913),
	.w5(32'h3aaaa86e),
	.w6(32'hbb950760),
	.w7(32'h3a8a8b4c),
	.w8(32'hbaa86089),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87cd3b),
	.w1(32'hbb11c283),
	.w2(32'hbb2fde6e),
	.w3(32'h3a7e03de),
	.w4(32'hbae7503d),
	.w5(32'hbb1cbee0),
	.w6(32'hbb110ff7),
	.w7(32'hbb831736),
	.w8(32'hbbe4b9eb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac8450),
	.w1(32'h3a22548c),
	.w2(32'hbb18a814),
	.w3(32'hbb639454),
	.w4(32'h3b3d7fb7),
	.w5(32'hb9cc526e),
	.w6(32'h3a188083),
	.w7(32'hbb081fbe),
	.w8(32'hbb0277e3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8a638),
	.w1(32'hbba0ccfa),
	.w2(32'h3bf6763a),
	.w3(32'hbafe01ac),
	.w4(32'hba43d666),
	.w5(32'h3be8ea08),
	.w6(32'h3b66c820),
	.w7(32'h3bda3e16),
	.w8(32'h3b252c9d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a887c1a),
	.w1(32'hb915e6c8),
	.w2(32'h385f2688),
	.w3(32'hbabdae8a),
	.w4(32'h3a89ed85),
	.w5(32'h3aafb369),
	.w6(32'h3a592c64),
	.w7(32'h3b1979a9),
	.w8(32'hba92f533),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72b4142),
	.w1(32'hbae9caca),
	.w2(32'hbad9422c),
	.w3(32'h3acd717e),
	.w4(32'hbb8b7c36),
	.w5(32'hbaebbd6e),
	.w6(32'hbaeb89af),
	.w7(32'h3aab077d),
	.w8(32'hbb0e045d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79d97b),
	.w1(32'h3a9c7811),
	.w2(32'hbb1a4c31),
	.w3(32'hbb96bc64),
	.w4(32'hbac7f7fa),
	.w5(32'hbb3fddbe),
	.w6(32'hbb5c2270),
	.w7(32'hbba8cb5b),
	.w8(32'hbbb24faf),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff9ac9),
	.w1(32'hbb9f4cd3),
	.w2(32'h3a097135),
	.w3(32'hbbba109c),
	.w4(32'hbadc70de),
	.w5(32'hbb0451c7),
	.w6(32'hbc1d0330),
	.w7(32'hbb15dc10),
	.w8(32'hbb70931a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4c78a),
	.w1(32'hba0ed047),
	.w2(32'hba2cf3fa),
	.w3(32'hbb930758),
	.w4(32'hbab79951),
	.w5(32'hbaf1512b),
	.w6(32'h3b5aa46b),
	.w7(32'h3b837617),
	.w8(32'h39c0216c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c49b25),
	.w1(32'hbbac82fb),
	.w2(32'hbb50ad22),
	.w3(32'hbb4b2759),
	.w4(32'hba903e7a),
	.w5(32'hba07e2f9),
	.w6(32'h3a9f1553),
	.w7(32'hbb4ec1ec),
	.w8(32'hbb4a3e2d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba931d6c),
	.w1(32'hb9a65343),
	.w2(32'hbacc0538),
	.w3(32'h3af252f6),
	.w4(32'hba7a204c),
	.w5(32'hbb234253),
	.w6(32'h3aa7cd62),
	.w7(32'h3aa6831f),
	.w8(32'h3a3d3d7e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82d338),
	.w1(32'h3b05a709),
	.w2(32'h3b7fe0fa),
	.w3(32'hba4d1c52),
	.w4(32'h3abecdc5),
	.w5(32'h3aa9403d),
	.w6(32'h3ba40b88),
	.w7(32'h3b6099ef),
	.w8(32'hba728a8a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc018ca8),
	.w1(32'hbc008ed2),
	.w2(32'h3a97c7f4),
	.w3(32'hbc042a67),
	.w4(32'hbb182a11),
	.w5(32'hba38f318),
	.w6(32'hbbcd6bc8),
	.w7(32'hbb0f4b5e),
	.w8(32'h3b1ef537),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5f760),
	.w1(32'h3a4a81e3),
	.w2(32'hba69b90b),
	.w3(32'hb994a907),
	.w4(32'h3bbc71fe),
	.w5(32'hba7eea49),
	.w6(32'hb9a7cd7a),
	.w7(32'h3affd912),
	.w8(32'hb8b5db1a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8692),
	.w1(32'h39f55b49),
	.w2(32'h3a9d7932),
	.w3(32'h3b3274ac),
	.w4(32'hbba20a3c),
	.w5(32'hbb4cc4fb),
	.w6(32'h3b92daa3),
	.w7(32'h3b11cc41),
	.w8(32'h39e03ec2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93df8f9),
	.w1(32'h3a90e998),
	.w2(32'h3a475a14),
	.w3(32'hbbfd236d),
	.w4(32'hbbb7238f),
	.w5(32'h3ac0ba4a),
	.w6(32'hbbba5961),
	.w7(32'hba04e3ce),
	.w8(32'h39b86c1e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63004f),
	.w1(32'hbac28d99),
	.w2(32'hbad7ef4f),
	.w3(32'hb699e1ba),
	.w4(32'hba877778),
	.w5(32'h3aad3d0a),
	.w6(32'h3bba688b),
	.w7(32'h39a9a67a),
	.w8(32'hbb2e9d66),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb341d6a),
	.w1(32'h3b4487a4),
	.w2(32'h3b3ef07c),
	.w3(32'h3c34cef0),
	.w4(32'h3c1bb068),
	.w5(32'h3c100f96),
	.w6(32'h3adbcd4c),
	.w7(32'h3be56e11),
	.w8(32'h3bce04f3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e834c),
	.w1(32'hbb957f20),
	.w2(32'h3bb1aae4),
	.w3(32'hbb0d6233),
	.w4(32'h3b011e9b),
	.w5(32'hba89f5cc),
	.w6(32'h3b9293d2),
	.w7(32'hbb41a655),
	.w8(32'hbb84342b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996ceda),
	.w1(32'h3952f6aa),
	.w2(32'h3b9756ae),
	.w3(32'hbae97c83),
	.w4(32'h3b482c2a),
	.w5(32'h3c3ad781),
	.w6(32'hbb13e876),
	.w7(32'h3a6f4a62),
	.w8(32'h3c1caeeb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af71d87),
	.w1(32'hba8ba0d7),
	.w2(32'hba84e627),
	.w3(32'h3b954b4d),
	.w4(32'h3b3657ae),
	.w5(32'h3b23059b),
	.w6(32'hbaa9eeaa),
	.w7(32'hba125d47),
	.w8(32'hba89e08b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04d8c2),
	.w1(32'h3b7f806d),
	.w2(32'h3baf90f7),
	.w3(32'h3b302a7d),
	.w4(32'hbb0cb59b),
	.w5(32'h39271bc7),
	.w6(32'h3c18a720),
	.w7(32'h3c146854),
	.w8(32'h3c29ed7f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbd902),
	.w1(32'hbb1916ad),
	.w2(32'hbb1e05f5),
	.w3(32'h3b047432),
	.w4(32'h3b3729bf),
	.w5(32'h3b27ef9b),
	.w6(32'hbac21c7b),
	.w7(32'hbada09de),
	.w8(32'hbada3942),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29ca31),
	.w1(32'hbae12169),
	.w2(32'h3a86059d),
	.w3(32'h3a3b2960),
	.w4(32'hbb544705),
	.w5(32'hbbac52b9),
	.w6(32'hba3d819a),
	.w7(32'hb88f91cd),
	.w8(32'hba01779c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ecb71),
	.w1(32'h3b0fd377),
	.w2(32'h3b7d65c1),
	.w3(32'hb9b7999a),
	.w4(32'hba513374),
	.w5(32'h3a060642),
	.w6(32'h399829cd),
	.w7(32'hbb75256a),
	.w8(32'h39efea3d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6145dc),
	.w1(32'hbaf2db98),
	.w2(32'hbb8a844e),
	.w3(32'h38f50e33),
	.w4(32'hba143f52),
	.w5(32'hbb3ac433),
	.w6(32'hbb20ecec),
	.w7(32'hba4a05ea),
	.w8(32'hbb2fd71e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd1ef5),
	.w1(32'h3acf2c67),
	.w2(32'hbaa5f7e7),
	.w3(32'hbb24f2ab),
	.w4(32'hba92ef6b),
	.w5(32'hbaebe7db),
	.w6(32'h3b2a151b),
	.w7(32'h3aed6ece),
	.w8(32'h3a9ee282),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7f129),
	.w1(32'hb9cb10a4),
	.w2(32'hba62f8e5),
	.w3(32'hbada60ac),
	.w4(32'hbacd6d35),
	.w5(32'hbb1081a0),
	.w6(32'hba5f3c97),
	.w7(32'hbb35ea7a),
	.w8(32'hbb74aabe),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1f451),
	.w1(32'hbaece49c),
	.w2(32'h3a09c226),
	.w3(32'hbb34158d),
	.w4(32'h3ba0bba1),
	.w5(32'hb9504f62),
	.w6(32'h3a92564c),
	.w7(32'h3a79dc8e),
	.w8(32'h3aecefab),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03871c),
	.w1(32'hbb5b401c),
	.w2(32'hbb4992a5),
	.w3(32'hbb92d491),
	.w4(32'hba5bfd45),
	.w5(32'hba74169f),
	.w6(32'hbb0c3e7b),
	.w7(32'hbb24839d),
	.w8(32'hbadd9889),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02cce0),
	.w1(32'h3b3db164),
	.w2(32'h3b0d0ae5),
	.w3(32'h369d35ae),
	.w4(32'h3babc846),
	.w5(32'h3aebac5b),
	.w6(32'h3b107561),
	.w7(32'h3b740546),
	.w8(32'h394e5e91),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3eaf2),
	.w1(32'h3a43ec55),
	.w2(32'hbafdc54e),
	.w3(32'h3a1d4001),
	.w4(32'h3967369d),
	.w5(32'h3a4eeefb),
	.w6(32'hba96b411),
	.w7(32'h39442249),
	.w8(32'hb7dd0f15),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1b5d9),
	.w1(32'hbb15388a),
	.w2(32'hbb1f7898),
	.w3(32'h3b89d6d0),
	.w4(32'hbad365ea),
	.w5(32'hbb1b8e3c),
	.w6(32'hbb90097a),
	.w7(32'hbb99d8ee),
	.w8(32'hbb9a76f7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc19774),
	.w1(32'hbb70b7b1),
	.w2(32'h389fc85b),
	.w3(32'hbaec8284),
	.w4(32'hbb88a548),
	.w5(32'hbb42cd65),
	.w6(32'hba31c3f8),
	.w7(32'h3b380b5e),
	.w8(32'h3bc8e111),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd425e),
	.w1(32'hba5f7324),
	.w2(32'hbaf6d095),
	.w3(32'h3b9782ad),
	.w4(32'hbb8f3af7),
	.w5(32'hbaf05995),
	.w6(32'hba90556e),
	.w7(32'hbb505347),
	.w8(32'hbba64d71),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba862fcb),
	.w1(32'hbb2f4713),
	.w2(32'hbadcf47c),
	.w3(32'hbacfcef8),
	.w4(32'h3a2410fb),
	.w5(32'hb9b9a6d0),
	.w6(32'hbaaf2e03),
	.w7(32'hbadea8ec),
	.w8(32'hb8038903),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc31d20),
	.w1(32'hbb48ed6b),
	.w2(32'hbad39bc7),
	.w3(32'hbb3c3314),
	.w4(32'hbab31ff8),
	.w5(32'hbb35f09e),
	.w6(32'hbb090e5e),
	.w7(32'hbbaea6b3),
	.w8(32'hbb504e3d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69fc9d),
	.w1(32'hbb691112),
	.w2(32'hbb70b648),
	.w3(32'hbbfcecf0),
	.w4(32'hbbc3e761),
	.w5(32'hbb088d3e),
	.w6(32'hbb083951),
	.w7(32'hbbea1922),
	.w8(32'hbba72423),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bd7ca),
	.w1(32'hbb1d633b),
	.w2(32'hba888862),
	.w3(32'hba4c4234),
	.w4(32'hb9d81151),
	.w5(32'hbaa7ad61),
	.w6(32'hbab2c829),
	.w7(32'hb978e466),
	.w8(32'hbb07fac9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d6b08),
	.w1(32'h3b82bb85),
	.w2(32'h3c41bc8d),
	.w3(32'hbb5aa14f),
	.w4(32'h3c228b4f),
	.w5(32'h3c9353dc),
	.w6(32'h39f47ba6),
	.w7(32'hbb0d6f10),
	.w8(32'hbba727c7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53e41f),
	.w1(32'hba8b907e),
	.w2(32'hbb8f025f),
	.w3(32'h3c427d02),
	.w4(32'h3a6e1714),
	.w5(32'h3988b4f4),
	.w6(32'h3b0c1d6a),
	.w7(32'hba686c69),
	.w8(32'hbaf5c1fa),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39114da0),
	.w1(32'hba87b755),
	.w2(32'hbac8d79b),
	.w3(32'hb89272e6),
	.w4(32'hbac0bc84),
	.w5(32'hbb54c8ef),
	.w6(32'h3b8afba4),
	.w7(32'h3b0f9b1a),
	.w8(32'h3b985f16),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b443712),
	.w1(32'h39e7f492),
	.w2(32'h3b25c7b1),
	.w3(32'h3a9ed14a),
	.w4(32'h3a0970bb),
	.w5(32'h3ac0239f),
	.w6(32'hbaf64fd9),
	.w7(32'hb8815a2e),
	.w8(32'h3a8ae1f8),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f5f63),
	.w1(32'h3a0df831),
	.w2(32'hba26318e),
	.w3(32'hb9ac6129),
	.w4(32'h3ab6491b),
	.w5(32'h3abd1f54),
	.w6(32'hb96152c8),
	.w7(32'hbad982a9),
	.w8(32'hbabf6451),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f95d5),
	.w1(32'hbb5c3592),
	.w2(32'h3a0ccdcd),
	.w3(32'h39eae6ed),
	.w4(32'hbbad400b),
	.w5(32'hbb49c39e),
	.w6(32'hbac81f42),
	.w7(32'h3a00f436),
	.w8(32'hbbc62000),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9973ebc),
	.w1(32'hba4820d0),
	.w2(32'hbb13974b),
	.w3(32'h38f51445),
	.w4(32'hbb2af52a),
	.w5(32'hbb2ab189),
	.w6(32'hbb4a1951),
	.w7(32'hbb8c73ff),
	.w8(32'hbb836a25),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe897d),
	.w1(32'hbaa29768),
	.w2(32'hbb6f2255),
	.w3(32'hbb67294a),
	.w4(32'hbb3f23ac),
	.w5(32'h3ae5ec90),
	.w6(32'hbaa99ac9),
	.w7(32'h3b2271af),
	.w8(32'hbb669ca5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b316821),
	.w1(32'hbb8a155f),
	.w2(32'hbb55e853),
	.w3(32'hba959aa3),
	.w4(32'hbb543c50),
	.w5(32'hbbaa4312),
	.w6(32'hbbb48930),
	.w7(32'hbb8ec9f5),
	.w8(32'hbb008397),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93bbd0),
	.w1(32'hbb582ed0),
	.w2(32'hbae801c5),
	.w3(32'hbb9d01f8),
	.w4(32'h3adda65f),
	.w5(32'h3b0d22bf),
	.w6(32'hbb2c4eef),
	.w7(32'hba31687e),
	.w8(32'h3ab54dd5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8539d),
	.w1(32'h3a70ff43),
	.w2(32'hb7466660),
	.w3(32'h39701039),
	.w4(32'h3b8d06a4),
	.w5(32'h3b6baa9e),
	.w6(32'hba945389),
	.w7(32'hbb54144b),
	.w8(32'hbb592778),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b5bad),
	.w1(32'hbb244a4e),
	.w2(32'hbb464f6f),
	.w3(32'h3b486afa),
	.w4(32'h3b43411c),
	.w5(32'h3b6434d7),
	.w6(32'h3a0158cf),
	.w7(32'h38307057),
	.w8(32'hbb80f91b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2c4ce),
	.w1(32'hbb2fe023),
	.w2(32'hba053617),
	.w3(32'h3b6c0afa),
	.w4(32'h3b0bf59e),
	.w5(32'hbb4f922f),
	.w6(32'h391819ae),
	.w7(32'hb9e74261),
	.w8(32'h3a00f669),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3019d),
	.w1(32'h399fc61f),
	.w2(32'hba9529a3),
	.w3(32'hbaf75373),
	.w4(32'h38a853a9),
	.w5(32'h398b0b56),
	.w6(32'h3a47d6cc),
	.w7(32'h3baa1ecf),
	.w8(32'hbac0be28),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac43ed4),
	.w1(32'hbb27d48e),
	.w2(32'hba0ca128),
	.w3(32'hbacbf1ee),
	.w4(32'hbac49df7),
	.w5(32'hba89fde8),
	.w6(32'hb977ff04),
	.w7(32'h3af7eeff),
	.w8(32'hba97cca7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a084b03),
	.w1(32'hbae56da7),
	.w2(32'hbb411a9f),
	.w3(32'hbb6a6bd5),
	.w4(32'h3b034c26),
	.w5(32'hb9e2280e),
	.w6(32'hbb827ad7),
	.w7(32'h3921119d),
	.w8(32'h3b33536b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb210e16),
	.w1(32'h3b1d4035),
	.w2(32'h3a8c0f2c),
	.w3(32'hba085fa1),
	.w4(32'h3a9b0f5e),
	.w5(32'hb9994072),
	.w6(32'hba78fd2b),
	.w7(32'hb93b74a9),
	.w8(32'hbb00b6fb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c7d74),
	.w1(32'hbb5c3219),
	.w2(32'hbb86ed2f),
	.w3(32'hbb1a59a0),
	.w4(32'hbb7ead64),
	.w5(32'hbbadfdbe),
	.w6(32'hbb3d7202),
	.w7(32'hbb473e5e),
	.w8(32'hbb6ffeaf),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb778904),
	.w1(32'h3af95a7f),
	.w2(32'h3a139f0e),
	.w3(32'hbb75ce19),
	.w4(32'h3ae0d59f),
	.w5(32'hbb68c292),
	.w6(32'hbac470a6),
	.w7(32'hbaa1508d),
	.w8(32'h3b7218d5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ac8c7),
	.w1(32'hbb58ba70),
	.w2(32'hbb83b6dc),
	.w3(32'h3a8b4c33),
	.w4(32'hbac5a602),
	.w5(32'hbb89e423),
	.w6(32'hbbb6f9d3),
	.w7(32'hbb934518),
	.w8(32'hbbc83ffc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3776d),
	.w1(32'hbc272413),
	.w2(32'hbb83d617),
	.w3(32'hbbf5eeb8),
	.w4(32'hbb41206b),
	.w5(32'hbb849afc),
	.w6(32'hbbc30285),
	.w7(32'hbb8c724a),
	.w8(32'hbb21c389),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f0778),
	.w1(32'hba44213b),
	.w2(32'h3b3ed267),
	.w3(32'hbba583a7),
	.w4(32'hbb01498c),
	.w5(32'h39653ea8),
	.w6(32'hbb257049),
	.w7(32'hba36b9dc),
	.w8(32'hba70ddd5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b46cb),
	.w1(32'hbbb7dbeb),
	.w2(32'hbbad76af),
	.w3(32'hbbaada90),
	.w4(32'hbc19e531),
	.w5(32'hb829a364),
	.w6(32'hbbd451b8),
	.w7(32'hbc036845),
	.w8(32'hbbf1d437),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule