module layer_8_featuremap_179(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc540fc7),
	.w1(32'hbc0ed50f),
	.w2(32'hbc3a45ad),
	.w3(32'h3b8e59d4),
	.w4(32'hbc0cb6e6),
	.w5(32'hbc171251),
	.w6(32'hbb84a337),
	.w7(32'h3c254514),
	.w8(32'h3c64f531),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a251d),
	.w1(32'hba34124d),
	.w2(32'h39b60b73),
	.w3(32'hbc777ed4),
	.w4(32'hbc143344),
	.w5(32'hbc3aa6ab),
	.w6(32'hbb817b2c),
	.w7(32'hbbb9fe44),
	.w8(32'hbbf1d5e3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb048db4),
	.w1(32'h3a8fc904),
	.w2(32'h3b5b93c8),
	.w3(32'hbc07fa5f),
	.w4(32'hbbc91975),
	.w5(32'hbbab247a),
	.w6(32'h3aeab21c),
	.w7(32'hbb80371b),
	.w8(32'hba271d20),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d8557),
	.w1(32'hbcd6dc41),
	.w2(32'hbcd68202),
	.w3(32'hb9bf435a),
	.w4(32'hbab50776),
	.w5(32'hbb901681),
	.w6(32'hbc455aff),
	.w7(32'hbb484906),
	.w8(32'h3c26f6e6),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58cc85),
	.w1(32'hba7c2277),
	.w2(32'hbba3d032),
	.w3(32'hbc3a792f),
	.w4(32'h3a5d6cb1),
	.w5(32'hbb0ec49d),
	.w6(32'h3b27b2cc),
	.w7(32'h3b87c631),
	.w8(32'h3ba99b21),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb764b8c),
	.w1(32'h3c21a107),
	.w2(32'h3c5e86e5),
	.w3(32'hbb77a7c1),
	.w4(32'hbc175379),
	.w5(32'hbbdda2d2),
	.w6(32'h3a1d9d71),
	.w7(32'h3bea302a),
	.w8(32'hb841c7e6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a820c4a),
	.w1(32'hbbd91727),
	.w2(32'hbc2de51a),
	.w3(32'hbc206107),
	.w4(32'hbac79e36),
	.w5(32'hba37d476),
	.w6(32'hbb23ae27),
	.w7(32'hbb4b3889),
	.w8(32'hba7247c5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5b23),
	.w1(32'h3b007801),
	.w2(32'hbc1d13f3),
	.w3(32'hbb94f996),
	.w4(32'hbacfcf8c),
	.w5(32'h3b19789a),
	.w6(32'h3be031b3),
	.w7(32'h3b248d7b),
	.w8(32'h3b0c8b88),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07cce1),
	.w1(32'h3b0e0fdd),
	.w2(32'hbc1cab33),
	.w3(32'hb8d7852b),
	.w4(32'h3c7f3ac7),
	.w5(32'h3c041d46),
	.w6(32'h3b3048ce),
	.w7(32'h3ab91236),
	.w8(32'h3c130eeb),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc69c80),
	.w1(32'hbca53a7c),
	.w2(32'hbd4e68a3),
	.w3(32'h3b72c5e1),
	.w4(32'hb9857382),
	.w5(32'hbc8cdd54),
	.w6(32'hbb937ab3),
	.w7(32'hb9b6910a),
	.w8(32'h3cbdc6b5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19c2e5),
	.w1(32'h3c41477e),
	.w2(32'h3d313b61),
	.w3(32'hbc9c6f67),
	.w4(32'hbccf914c),
	.w5(32'hbcbd9e7e),
	.w6(32'h3c074bbf),
	.w7(32'h3c71b0bd),
	.w8(32'hbbfdbb2a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d057976),
	.w1(32'hbb95ccff),
	.w2(32'hbac70cca),
	.w3(32'hbb512677),
	.w4(32'hbc0a8e95),
	.w5(32'hbbc21080),
	.w6(32'hbbbf2d61),
	.w7(32'hbb9912f6),
	.w8(32'hbc26730f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a9716),
	.w1(32'hbc37dce6),
	.w2(32'hbc28a54c),
	.w3(32'h3b4fc71d),
	.w4(32'hbc55efc3),
	.w5(32'hbd11db75),
	.w6(32'h3b9a834d),
	.w7(32'h3ca54a5e),
	.w8(32'h3cc25ec8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b604627),
	.w1(32'hbc58a369),
	.w2(32'hbb3b18c1),
	.w3(32'hbcdf45fc),
	.w4(32'hbc065519),
	.w5(32'hbc4f73cb),
	.w6(32'hb9122533),
	.w7(32'h3c64a667),
	.w8(32'h3c0f2e93),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb504e01),
	.w1(32'hbb6d7f16),
	.w2(32'hbc2f8f45),
	.w3(32'hbcb4af4d),
	.w4(32'h3b9e1930),
	.w5(32'h3bb21b75),
	.w6(32'hbb8bece9),
	.w7(32'hbb7f391d),
	.w8(32'hb8d80c71),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b0980),
	.w1(32'h3ae55e87),
	.w2(32'h3bc91a74),
	.w3(32'h39b7f267),
	.w4(32'h3c323a51),
	.w5(32'h3b7060cf),
	.w6(32'hbb354961),
	.w7(32'hbb2e21d8),
	.w8(32'hbb287782),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f5597),
	.w1(32'h3bcab922),
	.w2(32'h3bed69db),
	.w3(32'h3a7732f1),
	.w4(32'hba481150),
	.w5(32'hba93bbd4),
	.w6(32'hbb04fec1),
	.w7(32'hbb018f30),
	.w8(32'hbbd9d370),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a9ac2),
	.w1(32'hbad8af5d),
	.w2(32'h3b9a29a2),
	.w3(32'h3a870a9b),
	.w4(32'h3b224901),
	.w5(32'hbbb5eded),
	.w6(32'hbc0f219e),
	.w7(32'h3b175fa4),
	.w8(32'h3b4e818e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec686f),
	.w1(32'h3bb91142),
	.w2(32'h3bf0e450),
	.w3(32'hbb34d04a),
	.w4(32'h3b9a399b),
	.w5(32'hbbc63977),
	.w6(32'hba9fe5dd),
	.w7(32'h3c6b5e63),
	.w8(32'h3c90d9a2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49bd13),
	.w1(32'h3b97ea80),
	.w2(32'h3a114b98),
	.w3(32'hbc7fe6d6),
	.w4(32'h3bb68cd6),
	.w5(32'h3c03b895),
	.w6(32'h3ba8ec6f),
	.w7(32'h3b9f763b),
	.w8(32'h3c0c3210),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39739a02),
	.w1(32'hbb857eb2),
	.w2(32'h3b4c1f35),
	.w3(32'h3b371e56),
	.w4(32'hbc53d72a),
	.w5(32'hbcb7c248),
	.w6(32'h3c0c9f4e),
	.w7(32'hbb5e6ff8),
	.w8(32'hbb64b8d0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c235c60),
	.w1(32'hbb97b9d9),
	.w2(32'hb9727a3a),
	.w3(32'hbcc6a59c),
	.w4(32'hb9d3523a),
	.w5(32'hbb3d52a4),
	.w6(32'hba33fa1f),
	.w7(32'h3abd66f3),
	.w8(32'hbbf14c28),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a5435),
	.w1(32'hbc5b1205),
	.w2(32'hbba2f0fd),
	.w3(32'hbb9ec4d9),
	.w4(32'h3bb270c9),
	.w5(32'hba9c4065),
	.w6(32'hbc6182b4),
	.w7(32'hbc5e08d9),
	.w8(32'hbc17e71d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a855c),
	.w1(32'h3b9bdf90),
	.w2(32'h3b974d4e),
	.w3(32'hbba135b6),
	.w4(32'h3b8c941b),
	.w5(32'h3c108abb),
	.w6(32'hbc0d29a4),
	.w7(32'h3b4719b6),
	.w8(32'h3a958eaa),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59357a),
	.w1(32'h3b28534b),
	.w2(32'h3a9b92e9),
	.w3(32'h3a123e05),
	.w4(32'h3bf8b12c),
	.w5(32'h3c7e0fab),
	.w6(32'hbc3f03d6),
	.w7(32'hbcdc03c1),
	.w8(32'hbcd969b1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b9f5d),
	.w1(32'h3ad471e9),
	.w2(32'h3a96890b),
	.w3(32'h3c5d86c8),
	.w4(32'h3b901a50),
	.w5(32'h3bf636a3),
	.w6(32'h3ae4bba7),
	.w7(32'h3b37f0c8),
	.w8(32'hbae84ccb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe7d97),
	.w1(32'h3b01e523),
	.w2(32'h3ba4896d),
	.w3(32'h3c0fd10f),
	.w4(32'hbc0c3144),
	.w5(32'hbbe37df7),
	.w6(32'h3b532cc4),
	.w7(32'h3a5b672b),
	.w8(32'hbc05b2f2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca57ecb),
	.w1(32'hbc96287d),
	.w2(32'hbc9f7fe7),
	.w3(32'hbcc8fb06),
	.w4(32'hbbc16ff3),
	.w5(32'hbc7fbec9),
	.w6(32'hbcafe600),
	.w7(32'hbca65730),
	.w8(32'h3be25899),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4092f8),
	.w1(32'h3b2b6cb9),
	.w2(32'h3c12c527),
	.w3(32'hbb345f7e),
	.w4(32'hbbed461b),
	.w5(32'hbb4d1dfa),
	.w6(32'hbc452e80),
	.w7(32'hbc5977ae),
	.w8(32'hbc290619),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10cf44),
	.w1(32'hbaa8748c),
	.w2(32'hbb9ecf93),
	.w3(32'hbc050461),
	.w4(32'h3a745cf4),
	.w5(32'hba4c09fe),
	.w6(32'h3a35eea2),
	.w7(32'h3b061758),
	.w8(32'h3a191f48),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ec286f),
	.w1(32'h3bc8003e),
	.w2(32'h3c848a38),
	.w3(32'h3aa2ce59),
	.w4(32'hbc605a4b),
	.w5(32'hbd05537b),
	.w6(32'h3b91858e),
	.w7(32'h3c6fbd0b),
	.w8(32'h3c21ff35),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc909b4),
	.w1(32'h3c60265b),
	.w2(32'h3cae9caa),
	.w3(32'hbcb10b36),
	.w4(32'hbc7016ff),
	.w5(32'hbc8c10e9),
	.w6(32'h3b0ab433),
	.w7(32'h3b4011fe),
	.w8(32'hbb8f5a29),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c662112),
	.w1(32'hbc29225b),
	.w2(32'hbc67715e),
	.w3(32'hbbf9d196),
	.w4(32'hba86c9f8),
	.w5(32'hbbb89db4),
	.w6(32'hbbdb92e3),
	.w7(32'h3b6c0aad),
	.w8(32'h3be93cba),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabd704),
	.w1(32'h3b61854c),
	.w2(32'h3c33bdef),
	.w3(32'hbc184fc8),
	.w4(32'h3b6d4377),
	.w5(32'h3bbf5ed9),
	.w6(32'h3bae18e7),
	.w7(32'h3bfad777),
	.w8(32'h3bd5654e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65a0c8),
	.w1(32'h3bbb2ed0),
	.w2(32'h3ab76b6f),
	.w3(32'hbadf8ee9),
	.w4(32'h3a669321),
	.w5(32'hbc15a0a5),
	.w6(32'h3c9c61f5),
	.w7(32'h3cb34518),
	.w8(32'h3cd281b2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb12123),
	.w1(32'h3bf76abc),
	.w2(32'h3bfa88b4),
	.w3(32'hbc06c878),
	.w4(32'hbbd02ccb),
	.w5(32'hbb553b5c),
	.w6(32'hba3ab8ae),
	.w7(32'h38eec28a),
	.w8(32'h3b6bed71),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52c5d),
	.w1(32'h3c05fd9e),
	.w2(32'h3b8be72b),
	.w3(32'h3a080f63),
	.w4(32'h3c461cea),
	.w5(32'h3c988af9),
	.w6(32'hbc3250ef),
	.w7(32'hbc92ce7f),
	.w8(32'hbca23609),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee2e27),
	.w1(32'hb7253082),
	.w2(32'hbc17f3cb),
	.w3(32'h3c4c714a),
	.w4(32'h3c5b5e2a),
	.w5(32'h3c344529),
	.w6(32'hbb9bbd15),
	.w7(32'hbb9afb63),
	.w8(32'hbb0eabac),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3950c4),
	.w1(32'h3b9729b3),
	.w2(32'h3c083a66),
	.w3(32'h3b96a1ed),
	.w4(32'h3b525af2),
	.w5(32'h3c2bd636),
	.w6(32'hbada6a69),
	.w7(32'hbb230071),
	.w8(32'hba8832f8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cda55),
	.w1(32'hbb1bbf3f),
	.w2(32'h3bd3031a),
	.w3(32'h38e4d053),
	.w4(32'h3ad4f1b6),
	.w5(32'h3bacfda7),
	.w6(32'h3b26cddb),
	.w7(32'hbb0a4b21),
	.w8(32'h3b9be4f4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfaaa37),
	.w1(32'hba923b01),
	.w2(32'hb94b20d2),
	.w3(32'h3b75824a),
	.w4(32'hbb2fe508),
	.w5(32'hbb45b0ec),
	.w6(32'h3b0517dd),
	.w7(32'h3b6a5670),
	.w8(32'hb6d3879c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ddc72),
	.w1(32'h3b33ffda),
	.w2(32'h3c00a7fb),
	.w3(32'hbb13892f),
	.w4(32'hba172d02),
	.w5(32'hbc6187f5),
	.w6(32'h3be8130d),
	.w7(32'h3c13a89a),
	.w8(32'hba99c70c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c5b3d),
	.w1(32'h3c846850),
	.w2(32'h3c6a63fa),
	.w3(32'h3b58b160),
	.w4(32'h3c0e3fb1),
	.w5(32'h3c7a2fee),
	.w6(32'hbc077e6c),
	.w7(32'hbc8325f7),
	.w8(32'hbcb09fcc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a561d),
	.w1(32'h3ae911f1),
	.w2(32'h3b7136c6),
	.w3(32'h3c37d012),
	.w4(32'hbacf96f4),
	.w5(32'h3a6bf8fe),
	.w6(32'hbad09c4d),
	.w7(32'h39764d01),
	.w8(32'hbb22aea9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b6236),
	.w1(32'h3af50138),
	.w2(32'hbbf965af),
	.w3(32'h38571001),
	.w4(32'h3c1b788b),
	.w5(32'h39fcf15b),
	.w6(32'h3a1bb0b6),
	.w7(32'h3b69f013),
	.w8(32'h3c4e57be),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3343f3),
	.w1(32'h3b3d1779),
	.w2(32'h3ab13c4b),
	.w3(32'h3ab9df7a),
	.w4(32'hba4a1d66),
	.w5(32'hba362bc4),
	.w6(32'hb9ea2e69),
	.w7(32'hbb58c533),
	.w8(32'hbab593ef),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4dec1),
	.w1(32'hbc0b0cd5),
	.w2(32'hbbd381a2),
	.w3(32'hbb5da9fe),
	.w4(32'hbc58539d),
	.w5(32'hbc6ca31c),
	.w6(32'hbb3a1d4f),
	.w7(32'h3ba5ec7a),
	.w8(32'h3bd33478),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb837943),
	.w1(32'h3b86d874),
	.w2(32'hba2ddff4),
	.w3(32'hbc88e7e3),
	.w4(32'hbc022722),
	.w5(32'h3958b4f2),
	.w6(32'hbb85bd3b),
	.w7(32'h38592403),
	.w8(32'hba881ad6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4eb2c),
	.w1(32'hbbb986a3),
	.w2(32'hbb8c5468),
	.w3(32'h3b639d34),
	.w4(32'hbb9765b7),
	.w5(32'hbc957174),
	.w6(32'hbb86a382),
	.w7(32'h3b503aae),
	.w8(32'h3b9cb042),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e974c),
	.w1(32'hb85b775b),
	.w2(32'h3c24de52),
	.w3(32'h3b44a778),
	.w4(32'hbc0b5091),
	.w5(32'h3b883734),
	.w6(32'hbc36c455),
	.w7(32'hbc363dc1),
	.w8(32'hbba3e8d8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d6dc),
	.w1(32'hbba2e04b),
	.w2(32'hbb28c37b),
	.w3(32'hba66b708),
	.w4(32'h3b1421dd),
	.w5(32'hbabcc94a),
	.w6(32'h3b6a2628),
	.w7(32'h3aa8504e),
	.w8(32'h3b808840),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43fcc0),
	.w1(32'h3a550c46),
	.w2(32'h3b6d7a85),
	.w3(32'h3b058810),
	.w4(32'h3ab036f6),
	.w5(32'hbbcee6c9),
	.w6(32'h3c29fc29),
	.w7(32'h3c1d372b),
	.w8(32'h3c1f2931),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba916630),
	.w1(32'h3beae3e2),
	.w2(32'h3bbacb65),
	.w3(32'hbc0642fd),
	.w4(32'h3b19b64e),
	.w5(32'h3ab84205),
	.w6(32'h3ad5f5b4),
	.w7(32'h3a2fedde),
	.w8(32'h3a987b88),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca32bc),
	.w1(32'h3c564443),
	.w2(32'h3b6f08cc),
	.w3(32'hbb96eb47),
	.w4(32'h3bd94392),
	.w5(32'h3c2b13ac),
	.w6(32'h3b915450),
	.w7(32'hbc3bc2cf),
	.w8(32'hbbb31bbd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17079a),
	.w1(32'hbc19e1ab),
	.w2(32'hbc2926c2),
	.w3(32'h3bf88a6c),
	.w4(32'h3bc6ad7a),
	.w5(32'hbbf2ac8f),
	.w6(32'hb98ed69f),
	.w7(32'h3b381915),
	.w8(32'h3c2f649d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44c018),
	.w1(32'hbb8b4924),
	.w2(32'hba413dfc),
	.w3(32'hbb6570ff),
	.w4(32'hbb851152),
	.w5(32'h394a25ba),
	.w6(32'hbbc8dfba),
	.w7(32'h3ba5b613),
	.w8(32'h3b546ddb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b297150),
	.w1(32'h3c888b6b),
	.w2(32'h3cbdf820),
	.w3(32'hbb2ba0b3),
	.w4(32'hbb92f5d2),
	.w5(32'hbb54ebbb),
	.w6(32'h3bb6e385),
	.w7(32'h3c737694),
	.w8(32'h3c6248f7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f426f),
	.w1(32'hba9063a0),
	.w2(32'hbbd21dd8),
	.w3(32'hbc135c82),
	.w4(32'hba8d7f99),
	.w5(32'h3b28bb01),
	.w6(32'hbc388e1b),
	.w7(32'hbc84931d),
	.w8(32'hbbef004d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b761716),
	.w1(32'hbb85370f),
	.w2(32'h3ab98249),
	.w3(32'h3c10d74d),
	.w4(32'hbbac07f6),
	.w5(32'hbbc7a3a4),
	.w6(32'hbb13c4fb),
	.w7(32'h3a478a23),
	.w8(32'h3add6724),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49eb4d),
	.w1(32'hbab0b94c),
	.w2(32'hb98524eb),
	.w3(32'hbb61de73),
	.w4(32'hbc1555c5),
	.w5(32'h3bbfadce),
	.w6(32'h3ac10ca0),
	.w7(32'hbb827eff),
	.w8(32'h3884d485),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b850740),
	.w1(32'h3c479056),
	.w2(32'h3cd9b70a),
	.w3(32'h3ba80f55),
	.w4(32'hbc266309),
	.w5(32'hb9845193),
	.w6(32'hbc0463f2),
	.w7(32'hbb60341d),
	.w8(32'hbba62d79),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb53c01),
	.w1(32'h3c796893),
	.w2(32'h3b9c1181),
	.w3(32'hbb30b08a),
	.w4(32'h3cb9c007),
	.w5(32'h3d0ead6c),
	.w6(32'hbbe8a665),
	.w7(32'hbd031e97),
	.w8(32'hbd0876c5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa0b76),
	.w1(32'h3c6a7855),
	.w2(32'h3bcd4804),
	.w3(32'h3cd15781),
	.w4(32'h3bc857fe),
	.w5(32'h3bbb5e15),
	.w6(32'hbbbd5c55),
	.w7(32'hbca03172),
	.w8(32'hbcb92ae9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58f9e4),
	.w1(32'hbc7f4ee8),
	.w2(32'hbc9c29ac),
	.w3(32'h3ba527cb),
	.w4(32'hbc2c2c5e),
	.w5(32'hbc8e42fe),
	.w6(32'hbaaddc8f),
	.w7(32'h3ad3a0e5),
	.w8(32'h3b8a6518),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37266a),
	.w1(32'h3ba0aa61),
	.w2(32'h3bea2fab),
	.w3(32'hbc24d14e),
	.w4(32'hbac3530e),
	.w5(32'hbb787f6b),
	.w6(32'h3b5829a3),
	.w7(32'h3aebfe2a),
	.w8(32'hba408abb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc513a1),
	.w1(32'hbb16b89c),
	.w2(32'hbaf8e410),
	.w3(32'hb9e4bf2a),
	.w4(32'hba3281ed),
	.w5(32'h393803f6),
	.w6(32'h3b41231c),
	.w7(32'hbc17e5b6),
	.w8(32'hbc06fd24),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7285bb),
	.w1(32'hbc9a844f),
	.w2(32'hbca24c20),
	.w3(32'h3b649fec),
	.w4(32'hb93d7e9c),
	.w5(32'hbbce383d),
	.w6(32'hba875180),
	.w7(32'hbb182a06),
	.w8(32'hbb2099bd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86da13),
	.w1(32'hbb186686),
	.w2(32'hba83e15c),
	.w3(32'h372bdbb0),
	.w4(32'hbc305cca),
	.w5(32'hbbcc884f),
	.w6(32'hbb006973),
	.w7(32'hbbaaaa8b),
	.w8(32'hbc0c5cc3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb245f4),
	.w1(32'hbc3a7b45),
	.w2(32'hbb8598b5),
	.w3(32'hbc46cf01),
	.w4(32'hbacd9cd3),
	.w5(32'hbb9700ea),
	.w6(32'hbbcd84ed),
	.w7(32'h39e3d86e),
	.w8(32'hbb8f7c9e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbc4b3),
	.w1(32'hbc5d1c01),
	.w2(32'h3a49be21),
	.w3(32'hbc1dad71),
	.w4(32'hbbee09f3),
	.w5(32'hbb994854),
	.w6(32'hbc0680d7),
	.w7(32'h3b3f2a80),
	.w8(32'h3c05e90a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e6843),
	.w1(32'h38816f20),
	.w2(32'hbc6b7255),
	.w3(32'hbbe75d0f),
	.w4(32'h3c45b172),
	.w5(32'hbbfb5e1e),
	.w6(32'h3badf7e1),
	.w7(32'h3bfead75),
	.w8(32'h3be2bd6b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6e98a),
	.w1(32'hbb393558),
	.w2(32'hbba3e876),
	.w3(32'hbbf4a844),
	.w4(32'hbbce925e),
	.w5(32'hbb98936d),
	.w6(32'hbb67cede),
	.w7(32'h3ab207e0),
	.w8(32'hbabc5d97),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4beb4),
	.w1(32'h3b83f5b4),
	.w2(32'hb897c570),
	.w3(32'hbc4e17b7),
	.w4(32'hbc81aa53),
	.w5(32'hbc5d5612),
	.w6(32'hba3f7e7a),
	.w7(32'h3b1cbbfb),
	.w8(32'h3ba285e1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb489828),
	.w1(32'hbbe2b7cf),
	.w2(32'hbbfc1427),
	.w3(32'hbc3ce2f7),
	.w4(32'hbc19c04d),
	.w5(32'hbc8d8ad0),
	.w6(32'h3aa99a3f),
	.w7(32'h3c22f0f3),
	.w8(32'h3c717cb4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3fa4e),
	.w1(32'h3c36db6e),
	.w2(32'h3c4412b0),
	.w3(32'hbc3ef5fb),
	.w4(32'h3c649493),
	.w5(32'h3c6b624d),
	.w6(32'hbba0cb1e),
	.w7(32'hbc06a59b),
	.w8(32'hbc83d71b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6452fc),
	.w1(32'hbb0ac769),
	.w2(32'hbc542e86),
	.w3(32'h3c4626cb),
	.w4(32'h3bc3309f),
	.w5(32'h3ad9f703),
	.w6(32'hbaba0488),
	.w7(32'hba84781e),
	.w8(32'hbaffe7d7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d76de),
	.w1(32'hbbcc46ce),
	.w2(32'h3ab2ed5d),
	.w3(32'h3b187650),
	.w4(32'hbc0c9114),
	.w5(32'hbb258f5a),
	.w6(32'hbc1834d6),
	.w7(32'hbbad2e77),
	.w8(32'hbb35939e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8524c5),
	.w1(32'hb7d34ed9),
	.w2(32'h3c14e80f),
	.w3(32'hbaaae75b),
	.w4(32'hba348847),
	.w5(32'h3c2df68a),
	.w6(32'hbb925c82),
	.w7(32'hbaccedfe),
	.w8(32'h3ab5dea0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7b1e7),
	.w1(32'hbc9e26b2),
	.w2(32'hbc2228b3),
	.w3(32'h3bc4b77f),
	.w4(32'hbc8d723d),
	.w5(32'hbce691ec),
	.w6(32'hbbb02bd0),
	.w7(32'h3c40182e),
	.w8(32'h3c9d3e09),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcd3e9),
	.w1(32'hbc45e836),
	.w2(32'hbc513af5),
	.w3(32'hbc6871a9),
	.w4(32'h38e7a02f),
	.w5(32'hbc0665c5),
	.w6(32'hbb1634c7),
	.w7(32'h3c55f872),
	.w8(32'hbb1759bb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3ea9b),
	.w1(32'hbc20ba3a),
	.w2(32'hbb542980),
	.w3(32'hbbba3022),
	.w4(32'hbba0d909),
	.w5(32'hb85dd3a1),
	.w6(32'hbaeeaf3a),
	.w7(32'hbaf41342),
	.w8(32'h3c27987f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0a550),
	.w1(32'hbb58e530),
	.w2(32'hbba2ecc0),
	.w3(32'hbbc64cd8),
	.w4(32'h3a01bea6),
	.w5(32'hbb8993c0),
	.w6(32'hbb8fa3fd),
	.w7(32'h3b0accad),
	.w8(32'h3b8a436c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1e890),
	.w1(32'hba4de4d4),
	.w2(32'h3ab259f5),
	.w3(32'hbb78abd4),
	.w4(32'h3bebc906),
	.w5(32'h39799b54),
	.w6(32'hbb0b425f),
	.w7(32'hb9c11f84),
	.w8(32'h3b92e176),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf1fa6),
	.w1(32'hbc0d72ba),
	.w2(32'hbbedd8b5),
	.w3(32'hbc151740),
	.w4(32'hbbb43dcf),
	.w5(32'hba262024),
	.w6(32'hbab93014),
	.w7(32'h390f14b1),
	.w8(32'hbbaa285a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c2edd),
	.w1(32'hbbde2402),
	.w2(32'h3c177956),
	.w3(32'hbb5e59c0),
	.w4(32'hbc219cd2),
	.w5(32'hbc8bcb62),
	.w6(32'h3bf234b0),
	.w7(32'h3cbc7b8e),
	.w8(32'h3cafd81c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bc35f),
	.w1(32'hbbb4e237),
	.w2(32'h3ca6b7b5),
	.w3(32'hbc93ba20),
	.w4(32'hbbd9f3d8),
	.w5(32'hbc9a7fce),
	.w6(32'h3bb27bf3),
	.w7(32'h3cc8b8a6),
	.w8(32'h3cdf2c93),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05a1cc),
	.w1(32'hbc469771),
	.w2(32'hbc5b0785),
	.w3(32'hbc5d7903),
	.w4(32'hbc05275e),
	.w5(32'hbc8c6d50),
	.w6(32'hba839f8d),
	.w7(32'h3c43fc7c),
	.w8(32'h3c3a4879),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6855f8),
	.w1(32'h3c1d4d68),
	.w2(32'h3b1877ee),
	.w3(32'hbc04f722),
	.w4(32'h3b33d089),
	.w5(32'h3c6be808),
	.w6(32'hbcb9466a),
	.w7(32'hbd394a89),
	.w8(32'hbd396025),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc198f13),
	.w1(32'hbaa12cfe),
	.w2(32'h39acb75a),
	.w3(32'h3c7225ff),
	.w4(32'hbc7f7a7c),
	.w5(32'hbcc4eaa9),
	.w6(32'h3ba89d32),
	.w7(32'h3c85be7f),
	.w8(32'h3ca7c79e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8c28f),
	.w1(32'h3b899945),
	.w2(32'hbb56bb13),
	.w3(32'hbcbf372c),
	.w4(32'hbbac1f2b),
	.w5(32'hbc2b076b),
	.w6(32'hbb87c16d),
	.w7(32'h3c5cf735),
	.w8(32'h3c6635dc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd208b),
	.w1(32'hbc2c9930),
	.w2(32'hbc2d348f),
	.w3(32'hbc5b3d41),
	.w4(32'hbabd9328),
	.w5(32'hbc21c8e3),
	.w6(32'hbba560ec),
	.w7(32'hbb0e3ca3),
	.w8(32'hb93c0c70),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa430a),
	.w1(32'hba807e12),
	.w2(32'hbabb9f4e),
	.w3(32'hbc992aa3),
	.w4(32'h3b101606),
	.w5(32'h3a5414c2),
	.w6(32'hbb90d6fa),
	.w7(32'hbb370b3a),
	.w8(32'hbac61ea9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befbca7),
	.w1(32'hbb010f2b),
	.w2(32'hbb02fece),
	.w3(32'h3b2e2392),
	.w4(32'hbbd56a0e),
	.w5(32'hbc04beb7),
	.w6(32'h3b530d41),
	.w7(32'h3a7211c9),
	.w8(32'h3a4b07c5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb935ee2),
	.w1(32'h3a786421),
	.w2(32'h3b62a530),
	.w3(32'hbc1572b1),
	.w4(32'hbb803d88),
	.w5(32'hbbc268ad),
	.w6(32'hbadd1950),
	.w7(32'hbb77d32a),
	.w8(32'hbb9a9c37),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b222402),
	.w1(32'hb978fa58),
	.w2(32'hbbd0f4e2),
	.w3(32'hbb2a9aad),
	.w4(32'h3c0a72e3),
	.w5(32'h3c5b5fad),
	.w6(32'hbc45f308),
	.w7(32'hbc3a62ae),
	.w8(32'h3b476e45),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3df66d),
	.w1(32'hbb71455d),
	.w2(32'h3b8785dc),
	.w3(32'h3c8c0033),
	.w4(32'hbbbb993c),
	.w5(32'hbb552fe5),
	.w6(32'h3b479f5e),
	.w7(32'h3c2896ec),
	.w8(32'h3c7bbf8b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2da67f),
	.w1(32'h3b4fc41a),
	.w2(32'hbbb4f9e3),
	.w3(32'hbaa6da0c),
	.w4(32'hbc35aa31),
	.w5(32'hbb083a1e),
	.w6(32'h3bd1180a),
	.w7(32'hba302add),
	.w8(32'hbbc32f4a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb765d5),
	.w1(32'hbafc2427),
	.w2(32'hbac42b8f),
	.w3(32'hba5859ea),
	.w4(32'h3a01ce56),
	.w5(32'h3a9b7939),
	.w6(32'hbb55fae7),
	.w7(32'hbc028cfe),
	.w8(32'hbb878f38),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd59c8e),
	.w1(32'hbaccf8dd),
	.w2(32'h3b141232),
	.w3(32'h3bd6877e),
	.w4(32'h3bb31f9e),
	.w5(32'h3c15869e),
	.w6(32'hbb1874a6),
	.w7(32'hbbe13175),
	.w8(32'hbb30b3b8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f0d6e),
	.w1(32'hbb276bec),
	.w2(32'h3c3e2c70),
	.w3(32'hbb215a42),
	.w4(32'h3a6d51ce),
	.w5(32'h3b442d40),
	.w6(32'hbbdc4bea),
	.w7(32'hbbdade44),
	.w8(32'hbc294a35),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b8ff9),
	.w1(32'hbb251de9),
	.w2(32'hb993b72c),
	.w3(32'h3ad68358),
	.w4(32'hb8f6fef6),
	.w5(32'hbc833e20),
	.w6(32'h3c06ddd5),
	.w7(32'h3b891155),
	.w8(32'h3ba06810),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06210d),
	.w1(32'hbc016bc4),
	.w2(32'hbb3ac455),
	.w3(32'hbc52c988),
	.w4(32'hbba0f73d),
	.w5(32'hbba0cf2d),
	.w6(32'h38aba2c8),
	.w7(32'hbbba47a9),
	.w8(32'hbaa1f18b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba710170),
	.w1(32'hbbd8d8b4),
	.w2(32'hbc2186a1),
	.w3(32'h3b78c5cb),
	.w4(32'h3bf6c34c),
	.w5(32'h3ace70d1),
	.w6(32'hbc345e10),
	.w7(32'hbbc3cc3e),
	.w8(32'hbbb74015),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bd56d),
	.w1(32'hbc96f8a0),
	.w2(32'hbca18d44),
	.w3(32'hbc2c2458),
	.w4(32'hbc04913e),
	.w5(32'hba9f621a),
	.w6(32'h3c8638d3),
	.w7(32'h3d025a85),
	.w8(32'h3c7392ec),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82ebb8),
	.w1(32'hbb1fe01e),
	.w2(32'h3b9e0e13),
	.w3(32'hbc16c5ee),
	.w4(32'hba96a123),
	.w5(32'hbba26f47),
	.w6(32'hbbbae1bf),
	.w7(32'h3b1eb15d),
	.w8(32'h3ac114f5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0daf48),
	.w1(32'h3bd63c41),
	.w2(32'h3b50721c),
	.w3(32'hbace0a37),
	.w4(32'h3b89a42c),
	.w5(32'h3b79b54b),
	.w6(32'hba16cd55),
	.w7(32'hbb36499d),
	.w8(32'h39cf83f7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b680dc7),
	.w1(32'hbc5d1089),
	.w2(32'hbc43e02c),
	.w3(32'h3b0f3f80),
	.w4(32'hbc0be010),
	.w5(32'hbcbdf485),
	.w6(32'h3b98d166),
	.w7(32'h3c6fe00b),
	.w8(32'h3c47da07),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c595dd),
	.w1(32'h3c4e9deb),
	.w2(32'hbb62dbb7),
	.w3(32'hbcb4744e),
	.w4(32'h3c362811),
	.w5(32'h3c8c7acd),
	.w6(32'hbc7a0cd6),
	.w7(32'hbd2238a4),
	.w8(32'hbcdebb1a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc652128),
	.w1(32'h3a9ca3c5),
	.w2(32'hbb2b1a07),
	.w3(32'h3bfd714b),
	.w4(32'h3c06732c),
	.w5(32'h3c4f767e),
	.w6(32'hba3795fc),
	.w7(32'hbc19c15d),
	.w8(32'hbc5904fe),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c57ad),
	.w1(32'h3aa09ed9),
	.w2(32'h3b6a1c53),
	.w3(32'h3b7660c2),
	.w4(32'hbabb7ea8),
	.w5(32'hbb81e931),
	.w6(32'hbb78d5a0),
	.w7(32'hbb9bb968),
	.w8(32'hbc076191),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a872a98),
	.w1(32'hbc0dd0bc),
	.w2(32'hbb8a4ef7),
	.w3(32'hba98a6c2),
	.w4(32'hbaf8741c),
	.w5(32'hbc0a61ef),
	.w6(32'h3ac558f6),
	.w7(32'h3afe45cd),
	.w8(32'h3a99e078),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a3d81),
	.w1(32'h39c59fc9),
	.w2(32'h3b39c234),
	.w3(32'hbc119ce1),
	.w4(32'hbbbbec2c),
	.w5(32'hbbf137c8),
	.w6(32'h39bd1e1b),
	.w7(32'hba5b2162),
	.w8(32'h3a41024c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8e7d1),
	.w1(32'h3ada0f8b),
	.w2(32'hbbc60408),
	.w3(32'hbaf568d2),
	.w4(32'h3b8e2d39),
	.w5(32'hbb4b5dd5),
	.w6(32'hbaddd050),
	.w7(32'hbbef3ddc),
	.w8(32'hba5d1565),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3285a),
	.w1(32'h3b6110cf),
	.w2(32'h3c47dc62),
	.w3(32'hbc1784b9),
	.w4(32'h3c0d7697),
	.w5(32'h3c557711),
	.w6(32'hbc0da6f7),
	.w7(32'hbc7f9ccb),
	.w8(32'hbc880147),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c0486),
	.w1(32'h3b1fd1e6),
	.w2(32'h3be4bf5d),
	.w3(32'h3c85cdf5),
	.w4(32'hbc6d8d1c),
	.w5(32'hbcf3cec5),
	.w6(32'h3bcca944),
	.w7(32'h3c84ff07),
	.w8(32'h3c62118c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1b443),
	.w1(32'h3ba509e7),
	.w2(32'h3bf427ee),
	.w3(32'hbc57a806),
	.w4(32'hb9ceb51a),
	.w5(32'hbb1d0edd),
	.w6(32'hb92900ff),
	.w7(32'hba59d11d),
	.w8(32'hbb638933),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95bbf4),
	.w1(32'h3c3ea0f5),
	.w2(32'h3c242161),
	.w3(32'hbb09cfa8),
	.w4(32'h3c5eb7cd),
	.w5(32'h3ccbbb09),
	.w6(32'h3b16aedc),
	.w7(32'hbc291816),
	.w8(32'hbc88ea1c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43513c),
	.w1(32'hbb45fcaf),
	.w2(32'hbc4808fc),
	.w3(32'h3c961e56),
	.w4(32'hbbd03658),
	.w5(32'h39f2814a),
	.w6(32'hbbd7c09f),
	.w7(32'hbb3627bc),
	.w8(32'hbbfe6db9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44e44),
	.w1(32'hbbea15f4),
	.w2(32'hbc923cbe),
	.w3(32'hbb50990f),
	.w4(32'h3a0c2a5f),
	.w5(32'h3b0601e8),
	.w6(32'hbc202177),
	.w7(32'hbc9fbca8),
	.w8(32'h3abb38dc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a52de),
	.w1(32'hbb850c1a),
	.w2(32'hb8eabf6a),
	.w3(32'h39605844),
	.w4(32'h3bc7d5e3),
	.w5(32'h3c329cac),
	.w6(32'hbc037b5a),
	.w7(32'hbc0033de),
	.w8(32'hbc4f4f84),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00462a),
	.w1(32'h3ad23d54),
	.w2(32'hbb4b462f),
	.w3(32'h3be51db1),
	.w4(32'h3b911a75),
	.w5(32'h3a72e0c9),
	.w6(32'hbb98c9e4),
	.w7(32'h3bb17896),
	.w8(32'h3c0e4b22),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf16208),
	.w1(32'hbc15c61e),
	.w2(32'h3a415f3a),
	.w3(32'hbb9183b0),
	.w4(32'hbc42a424),
	.w5(32'hbc88cdd6),
	.w6(32'h3be5cdd8),
	.w7(32'h3cb2f355),
	.w8(32'h3c84c466),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c17fde),
	.w1(32'h3a609770),
	.w2(32'hba1b6158),
	.w3(32'hbc4edc3f),
	.w4(32'hbb74eb7e),
	.w5(32'hbc020204),
	.w6(32'h3b4ea7d5),
	.w7(32'h3b86a8d2),
	.w8(32'h3b900f61),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3628bf),
	.w1(32'h3bc466ce),
	.w2(32'hbb9cedca),
	.w3(32'hbb84f134),
	.w4(32'hbac24a5e),
	.w5(32'h3b11fb37),
	.w6(32'hbb16e238),
	.w7(32'h3ac939a8),
	.w8(32'hbb023acb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa9f03),
	.w1(32'h3875b0c1),
	.w2(32'hbc6cfd12),
	.w3(32'h374c2cfc),
	.w4(32'h3c5ffb7c),
	.w5(32'h3c5d9c0f),
	.w6(32'hbbff7140),
	.w7(32'h3b1a5e9b),
	.w8(32'h3c9ebeee),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1a9b3),
	.w1(32'hbb9ffa95),
	.w2(32'hbc01c24f),
	.w3(32'h3c547009),
	.w4(32'hba3b4930),
	.w5(32'h3af96c44),
	.w6(32'hbc01fa25),
	.w7(32'hbc3f840f),
	.w8(32'hbb2535e8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39842afb),
	.w1(32'h3ae76f13),
	.w2(32'h3ab4aeab),
	.w3(32'h3c2fdfe5),
	.w4(32'h39f61209),
	.w5(32'h3af03b05),
	.w6(32'h39811e07),
	.w7(32'h3b89f44a),
	.w8(32'hba462510),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2166c),
	.w1(32'h3c0efacc),
	.w2(32'h3b0038f2),
	.w3(32'hb89e1442),
	.w4(32'hbb001d82),
	.w5(32'hbc85ac20),
	.w6(32'h3b1ead27),
	.w7(32'h3c8b4660),
	.w8(32'hbb4ff987),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule