module layer_10_featuremap_354(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e57d6),
	.w1(32'hbaae549d),
	.w2(32'hb904a455),
	.w3(32'h39f67758),
	.w4(32'hb8c3b208),
	.w5(32'hbb0bb861),
	.w6(32'hb99e3269),
	.w7(32'hb97bdeef),
	.w8(32'hbaf41f06),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa29226),
	.w1(32'hbab9f161),
	.w2(32'hba569921),
	.w3(32'hbaf02c9e),
	.w4(32'hbababeae),
	.w5(32'h399162b0),
	.w6(32'h39b60bbc),
	.w7(32'hba1b32d5),
	.w8(32'h3a06d15d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8154ecb),
	.w1(32'hba12e8f1),
	.w2(32'h3a76784f),
	.w3(32'h3a72129b),
	.w4(32'h38b6d987),
	.w5(32'hb8c540a9),
	.w6(32'h3aa987ec),
	.w7(32'hb8de913c),
	.w8(32'hb9833350),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392cfc5c),
	.w1(32'hb7917893),
	.w2(32'h39b695e3),
	.w3(32'hb8f4575b),
	.w4(32'h38cfcf01),
	.w5(32'hbabdcfb0),
	.w6(32'hb79ae800),
	.w7(32'h3a1933b5),
	.w8(32'hba975eb5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1235ad),
	.w1(32'hbb42f368),
	.w2(32'hbae6ce50),
	.w3(32'hbb3fd225),
	.w4(32'hbb94d384),
	.w5(32'h3902e211),
	.w6(32'hbac448e3),
	.w7(32'hbb42474e),
	.w8(32'h38e99998),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc277b),
	.w1(32'hb9ba26a6),
	.w2(32'h37b2b50b),
	.w3(32'h39de7876),
	.w4(32'hb8b05e0a),
	.w5(32'hba834819),
	.w6(32'hb9d2b41e),
	.w7(32'hb9be941d),
	.w8(32'h38e065d9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cac4b),
	.w1(32'hba7fa9b2),
	.w2(32'hbacbe3e0),
	.w3(32'hba427334),
	.w4(32'hba66e26f),
	.w5(32'h39b8a986),
	.w6(32'hb92250a8),
	.w7(32'hba3ad400),
	.w8(32'hba30197a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba4264),
	.w1(32'hbadede09),
	.w2(32'hba92ffb6),
	.w3(32'hba0c647a),
	.w4(32'hbab24df8),
	.w5(32'hb99eee44),
	.w6(32'hbb2366c4),
	.w7(32'hbb015a13),
	.w8(32'h393104c3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0127a8),
	.w1(32'hb7c59bac),
	.w2(32'hba192d91),
	.w3(32'hba174e40),
	.w4(32'hba22d6ac),
	.w5(32'hb961f6e6),
	.w6(32'hb9ce63f1),
	.w7(32'hba001060),
	.w8(32'h39918ad2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a8677),
	.w1(32'hb96a862a),
	.w2(32'hb8f7ca24),
	.w3(32'hb943c243),
	.w4(32'hb88c9234),
	.w5(32'hb9a81bd8),
	.w6(32'hb862af69),
	.w7(32'hb93caab9),
	.w8(32'hb7f19e96),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997e00e),
	.w1(32'hba03247d),
	.w2(32'hb999d8b8),
	.w3(32'h3a6f15fc),
	.w4(32'hb98b8f04),
	.w5(32'h3ad04a60),
	.w6(32'h39916fdc),
	.w7(32'hba1ca03c),
	.w8(32'hb8eb2a7f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39842ada),
	.w1(32'h3a818f6c),
	.w2(32'h3a7e74d3),
	.w3(32'h3a3cbaa8),
	.w4(32'hba4408c3),
	.w5(32'hba0c3d42),
	.w6(32'h3a237698),
	.w7(32'hba774e0b),
	.w8(32'hb9d0b49c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ce19b),
	.w1(32'h3a42d8d8),
	.w2(32'h3a3eae93),
	.w3(32'h3a284c5e),
	.w4(32'h3a2d4d6a),
	.w5(32'h39903451),
	.w6(32'hba184d7f),
	.w7(32'hba260e40),
	.w8(32'h38ed44bf),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c1826a),
	.w1(32'hb8604da0),
	.w2(32'h3a8579ee),
	.w3(32'hba8b964c),
	.w4(32'hb78d0c30),
	.w5(32'h3a106cc3),
	.w6(32'h392fbaa2),
	.w7(32'h39a7a980),
	.w8(32'h39005061),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1bc34),
	.w1(32'h3a3d1f74),
	.w2(32'h3a9d3def),
	.w3(32'h39295ff9),
	.w4(32'h3a07685d),
	.w5(32'hbad1d53e),
	.w6(32'hba4e6b0f),
	.w7(32'h39b66327),
	.w8(32'hbafec560),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0093),
	.w1(32'hba5ac03b),
	.w2(32'hba160afd),
	.w3(32'hba2ba96a),
	.w4(32'h390ecc6a),
	.w5(32'hba8ca03c),
	.w6(32'hb977d597),
	.w7(32'hb99b6bb0),
	.w8(32'hba9e6486),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab604c4),
	.w1(32'hba45a921),
	.w2(32'h39a60442),
	.w3(32'hb93a3e7d),
	.w4(32'hb89acfb5),
	.w5(32'h391a6251),
	.w6(32'hb94999a2),
	.w7(32'hb98660b2),
	.w8(32'h3a344a7c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949235d),
	.w1(32'hbab8c6a6),
	.w2(32'hbaa6ac78),
	.w3(32'hba443982),
	.w4(32'hb981654b),
	.w5(32'hb9060224),
	.w6(32'hbab2224e),
	.w7(32'hba5e71ac),
	.w8(32'hb7866430),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b209d2),
	.w1(32'hb9a98568),
	.w2(32'hb9d45b64),
	.w3(32'hb9f0e06c),
	.w4(32'hb9ab0f6a),
	.w5(32'h399e9a9c),
	.w6(32'hbaae72b7),
	.w7(32'hb8d5a8d6),
	.w8(32'h39eb123e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c09fcb),
	.w1(32'hb9f706c6),
	.w2(32'h3a08d99a),
	.w3(32'h39acd542),
	.w4(32'h39cfc896),
	.w5(32'hba645edb),
	.w6(32'h3a290e86),
	.w7(32'h39217f1c),
	.w8(32'hbaca6c46),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60dcb7),
	.w1(32'h3a851356),
	.w2(32'h3a83716d),
	.w3(32'h3ae3091f),
	.w4(32'hb984b812),
	.w5(32'hb9df6ce3),
	.w6(32'h3a859b49),
	.w7(32'hba21a7dd),
	.w8(32'hb9ddb5d7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f2445),
	.w1(32'hb922f40c),
	.w2(32'hb8cd6291),
	.w3(32'hb9946f0f),
	.w4(32'h397ca417),
	.w5(32'h3aaa505e),
	.w6(32'hba631df1),
	.w7(32'hb8bdbd28),
	.w8(32'h3a55b26c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb887a421),
	.w1(32'h3ae0c164),
	.w2(32'h3a93b4a1),
	.w3(32'h3ad73e70),
	.w4(32'h3a35a929),
	.w5(32'hb97ae854),
	.w6(32'h3ad4c7d1),
	.w7(32'h3ae78db2),
	.w8(32'h3ac4d024),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26a1ad),
	.w1(32'h3aed8db7),
	.w2(32'hba923690),
	.w3(32'h3b548a7e),
	.w4(32'h39adcf74),
	.w5(32'hb86698a7),
	.w6(32'h3b0edcc4),
	.w7(32'hbae854c5),
	.w8(32'h391aee9a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9337d1e),
	.w1(32'hb9ec15c8),
	.w2(32'hba086474),
	.w3(32'h399b0c3d),
	.w4(32'hb9fdd866),
	.w5(32'hbad0a93a),
	.w6(32'h39814280),
	.w7(32'hba87287b),
	.w8(32'hba7de283),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c92107),
	.w1(32'h39be3a92),
	.w2(32'h3b01e45c),
	.w3(32'hb9d6be94),
	.w4(32'h3aa8004d),
	.w5(32'hb9f66a2e),
	.w6(32'hb894f81a),
	.w7(32'h3af16266),
	.w8(32'hb9bdff46),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16ccd3),
	.w1(32'hb9c11f3f),
	.w2(32'h39864238),
	.w3(32'hbaca95af),
	.w4(32'h39954811),
	.w5(32'hb9e51e60),
	.w6(32'hb8ee726e),
	.w7(32'h3a92ceac),
	.w8(32'hb87a7d42),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ab549),
	.w1(32'hba2fa8c6),
	.w2(32'h37cc23d0),
	.w3(32'hba9f1bdb),
	.w4(32'hba7b9df1),
	.w5(32'hb9542c4b),
	.w6(32'hba536847),
	.w7(32'hba09fdc6),
	.w8(32'h3905272a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882b1f1),
	.w1(32'hbb0ea5ca),
	.w2(32'h39864966),
	.w3(32'hbaa047b9),
	.w4(32'h38f0f078),
	.w5(32'hb9fcb05c),
	.w6(32'h39b56393),
	.w7(32'h3a172041),
	.w8(32'h39ad76ef),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dcdc1),
	.w1(32'hbb87d2f1),
	.w2(32'hba91158a),
	.w3(32'hbb1fec22),
	.w4(32'h39ab0acf),
	.w5(32'h3a9d74f8),
	.w6(32'hba33d1f2),
	.w7(32'h3a2e39ca),
	.w8(32'h3ab40bf8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c7067e),
	.w1(32'h3a5d75f4),
	.w2(32'hba8c486f),
	.w3(32'hb9559457),
	.w4(32'hbb0641ae),
	.w5(32'h3aa186d2),
	.w6(32'h3b1e2859),
	.w7(32'h39427dd7),
	.w8(32'h38ffe7e7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e1355),
	.w1(32'h38d2c566),
	.w2(32'hb99028cc),
	.w3(32'h3aca282b),
	.w4(32'hb9a86886),
	.w5(32'hb8d6a65f),
	.w6(32'h3a028115),
	.w7(32'hbad3f11b),
	.w8(32'h389e9950),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ede883),
	.w1(32'h3a938f60),
	.w2(32'h3a185c19),
	.w3(32'h397fa4c8),
	.w4(32'h3add1b9b),
	.w5(32'hb9c9b1af),
	.w6(32'h3b18cf69),
	.w7(32'h3b24b961),
	.w8(32'h39bfde56),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38917271),
	.w1(32'hbacd90a1),
	.w2(32'hbadc8cc9),
	.w3(32'hb9d31a86),
	.w4(32'hb9028a88),
	.w5(32'h3ae96550),
	.w6(32'hbaa832b2),
	.w7(32'hbac10658),
	.w8(32'h3a27f43f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78bd885),
	.w1(32'hba3ae37c),
	.w2(32'hba8b31b8),
	.w3(32'h3af230ff),
	.w4(32'h3aaa3a6f),
	.w5(32'h39b01193),
	.w6(32'h3a1541d3),
	.w7(32'hba72ae54),
	.w8(32'h3b2c290b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09b8af),
	.w1(32'h39c38feb),
	.w2(32'h3921c37f),
	.w3(32'h3ad58bb1),
	.w4(32'hba67e464),
	.w5(32'hba995b23),
	.w6(32'h3b2f4f16),
	.w7(32'h3a0ab3c3),
	.w8(32'h3a2e3abe),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa308a6),
	.w1(32'hbab305f9),
	.w2(32'hbb6ee041),
	.w3(32'hba615d87),
	.w4(32'hbad41108),
	.w5(32'hba54bf7e),
	.w6(32'h3a1d22c2),
	.w7(32'h3a2128d1),
	.w8(32'hba970ffe),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a415a),
	.w1(32'hb98b9abc),
	.w2(32'hba07f38a),
	.w3(32'h3986c5d9),
	.w4(32'h3a91e1d8),
	.w5(32'hbb048706),
	.w6(32'h39333386),
	.w7(32'h3a51792b),
	.w8(32'h3a7fdeed),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4767c),
	.w1(32'hbb2acabc),
	.w2(32'hbb087dda),
	.w3(32'hbae12abc),
	.w4(32'hba6e6861),
	.w5(32'h3a776fcc),
	.w6(32'h3a3c21a4),
	.w7(32'h3a82b4c3),
	.w8(32'h3ad2afb7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f33be),
	.w1(32'h3a4eb1f8),
	.w2(32'hbadb176d),
	.w3(32'h3a5dec0d),
	.w4(32'h3a96f0c1),
	.w5(32'h3aaf239a),
	.w6(32'h3ab35563),
	.w7(32'hb79f65c8),
	.w8(32'h39a8aa7e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93651ab),
	.w1(32'hba39dd05),
	.w2(32'h3af10ace),
	.w3(32'hbac7dcd8),
	.w4(32'hba5dde33),
	.w5(32'hbadd1861),
	.w6(32'hbaca8516),
	.w7(32'h3a474493),
	.w8(32'hba3a3a8d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab46408),
	.w1(32'hba12c70f),
	.w2(32'h399e0020),
	.w3(32'hb9e82708),
	.w4(32'h399f6807),
	.w5(32'h39efb07c),
	.w6(32'hba24e39c),
	.w7(32'h3a765256),
	.w8(32'h37f7c557),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d543d),
	.w1(32'h3a3c73df),
	.w2(32'h39f5520a),
	.w3(32'hba285ab2),
	.w4(32'hb9fa353a),
	.w5(32'hba545fe4),
	.w6(32'hba7d7998),
	.w7(32'hba2f56a2),
	.w8(32'hbb0276d5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a40de),
	.w1(32'hbad0061b),
	.w2(32'hba22f0f6),
	.w3(32'hbaf402b7),
	.w4(32'hbaea2ec4),
	.w5(32'h39dd268b),
	.w6(32'hba906756),
	.w7(32'hbaadcfb9),
	.w8(32'h3a9e041f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba238366),
	.w1(32'hbab33b6c),
	.w2(32'hba09b0ac),
	.w3(32'h39d89576),
	.w4(32'hba9f849f),
	.w5(32'hb8f2d5d6),
	.w6(32'hba19b520),
	.w7(32'hb9c3f14c),
	.w8(32'hba75de19),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40302b),
	.w1(32'hb9a2dfa3),
	.w2(32'hb9dc8273),
	.w3(32'hb9d34c1e),
	.w4(32'h3a2a9dd7),
	.w5(32'hbabc4579),
	.w6(32'hba7f6a46),
	.w7(32'hb8f013c7),
	.w8(32'hbaa97ddb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc4edf),
	.w1(32'hba96d147),
	.w2(32'hb99bd66b),
	.w3(32'hbad61bb8),
	.w4(32'hb9985e5b),
	.w5(32'h3990b140),
	.w6(32'hb9bc051f),
	.w7(32'h391ea96d),
	.w8(32'h397aa502),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861766f),
	.w1(32'hba035280),
	.w2(32'hb947e499),
	.w3(32'hb9dadf72),
	.w4(32'hb931ee9d),
	.w5(32'hb99ad14a),
	.w6(32'hba274c12),
	.w7(32'hb944a621),
	.w8(32'h394e6224),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62aadc),
	.w1(32'h3a8970d3),
	.w2(32'h3a93d24c),
	.w3(32'h3a10ed3a),
	.w4(32'hb7a97087),
	.w5(32'hb9a2a8dd),
	.w6(32'h38b8bd77),
	.w7(32'h396de0cd),
	.w8(32'hb94413af),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eaf63b),
	.w1(32'hb9be7111),
	.w2(32'hba3900a7),
	.w3(32'hb9fca60a),
	.w4(32'h3a167e7e),
	.w5(32'hba256846),
	.w6(32'hb9901060),
	.w7(32'h391e004c),
	.w8(32'hba935214),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba762eaf),
	.w1(32'hbb4df2fb),
	.w2(32'hbb27b934),
	.w3(32'hbb52dc23),
	.w4(32'hbaae8063),
	.w5(32'h3a2ed524),
	.w6(32'hbab2872b),
	.w7(32'hbabf5f36),
	.w8(32'h3975aa49),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54b65a),
	.w1(32'hba8e334a),
	.w2(32'hb9aa25bc),
	.w3(32'h3a0bf0fa),
	.w4(32'hba013da3),
	.w5(32'h3b5fc8cb),
	.w6(32'h38a86cf1),
	.w7(32'hba17d86c),
	.w8(32'h3a086c27),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c457ed),
	.w1(32'h3af5f784),
	.w2(32'h3ac69afc),
	.w3(32'h3a0f084d),
	.w4(32'hb9fed432),
	.w5(32'hb9275144),
	.w6(32'hb8176c17),
	.w7(32'h3a1b1cd0),
	.w8(32'h389533ca),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7487a6),
	.w1(32'hbb68f516),
	.w2(32'hbb3ab9ab),
	.w3(32'hbae13962),
	.w4(32'hbad6ea52),
	.w5(32'hb998df6e),
	.w6(32'hba951c6c),
	.w7(32'hbab379b0),
	.w8(32'hb93a6b53),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985597f),
	.w1(32'h39e02064),
	.w2(32'h3aa5bf1f),
	.w3(32'h3992dd66),
	.w4(32'h37a895db),
	.w5(32'hba9cbaec),
	.w6(32'hba07e3a7),
	.w7(32'hb988bedd),
	.w8(32'hbab04cf7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85a7e3),
	.w1(32'hbb0affdc),
	.w2(32'hba4c327e),
	.w3(32'hba9a7d83),
	.w4(32'hb9015af9),
	.w5(32'hb9a1de86),
	.w6(32'hba25853d),
	.w7(32'hbb03943d),
	.w8(32'hb9eaf067),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d5eab),
	.w1(32'hba1cb9f4),
	.w2(32'h3a65ac65),
	.w3(32'hb9eba398),
	.w4(32'h3931de57),
	.w5(32'h3aa42fa6),
	.w6(32'hb9d0003e),
	.w7(32'h39dc763a),
	.w8(32'h3aeecec2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad33f9e),
	.w1(32'h37e9c91a),
	.w2(32'h3a524078),
	.w3(32'hb953f4e8),
	.w4(32'h39a89635),
	.w5(32'hba8e85cf),
	.w6(32'h3a1fa283),
	.w7(32'h3a8d33ed),
	.w8(32'hb9267e52),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15bb1d),
	.w1(32'hb9f96c36),
	.w2(32'hbab9a80a),
	.w3(32'hba29824d),
	.w4(32'hb9ea42ca),
	.w5(32'hbab856c5),
	.w6(32'hba5526b1),
	.w7(32'hba1c1e05),
	.w8(32'hbb136b51),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd0421),
	.w1(32'hba646219),
	.w2(32'h39028255),
	.w3(32'hbb0b7bbf),
	.w4(32'hbab845a5),
	.w5(32'hba63e15d),
	.w6(32'hba4b79a5),
	.w7(32'hb9be09a2),
	.w8(32'h3a51f36f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd03ed),
	.w1(32'hbaccdb67),
	.w2(32'hba67304c),
	.w3(32'hbb1234c8),
	.w4(32'h38187962),
	.w5(32'hbad9b1a3),
	.w6(32'hba005525),
	.w7(32'h39b6873a),
	.w8(32'hbb26f37b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab82687),
	.w1(32'hba9cc257),
	.w2(32'h39dfb9c8),
	.w3(32'hbb03e5d0),
	.w4(32'hba471831),
	.w5(32'h3a772527),
	.w6(32'hbab71a8f),
	.w7(32'h392889f6),
	.w8(32'hb9b9f5c9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba518087),
	.w1(32'hb86b87ab),
	.w2(32'h39e04065),
	.w3(32'hba89f13c),
	.w4(32'hbaf7d246),
	.w5(32'hb98308c7),
	.w6(32'hba7ef1f8),
	.w7(32'hba9d6c11),
	.w8(32'hb8c8189b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a2fd5),
	.w1(32'hbaf1001e),
	.w2(32'hba284e4a),
	.w3(32'hb8754816),
	.w4(32'h376c82bb),
	.w5(32'h3a2e0963),
	.w6(32'hb90c2c8d),
	.w7(32'h38a2e0e9),
	.w8(32'h398ff34e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb8e9e),
	.w1(32'hba643510),
	.w2(32'h39d57d00),
	.w3(32'h3a0cce21),
	.w4(32'h3a812ed3),
	.w5(32'h391ac8f7),
	.w6(32'h39bd09ad),
	.w7(32'h395e71e9),
	.w8(32'hb99f5d4d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7d14c),
	.w1(32'h3b13341f),
	.w2(32'h3b0234b2),
	.w3(32'hb8f44f42),
	.w4(32'hbad54e8a),
	.w5(32'h3ad3b330),
	.w6(32'hba66684c),
	.w7(32'hbab4b7bc),
	.w8(32'h3a4aee20),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99133bc),
	.w1(32'hba955f74),
	.w2(32'hba11cb74),
	.w3(32'h3a34fc88),
	.w4(32'hba1360f6),
	.w5(32'hbaab9d65),
	.w6(32'hbaf5e8a0),
	.w7(32'hbac50b7e),
	.w8(32'hbb202413),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bb4bc),
	.w1(32'hbaa36cde),
	.w2(32'h39785678),
	.w3(32'hbb0ca679),
	.w4(32'hba98244a),
	.w5(32'h3a12f0b2),
	.w6(32'hbb049ce6),
	.w7(32'hba7b52c8),
	.w8(32'h3aabd89e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947da54),
	.w1(32'hb9f38535),
	.w2(32'h3a72dc7e),
	.w3(32'h3a8cc35f),
	.w4(32'h3ad8c327),
	.w5(32'h3a548ccd),
	.w6(32'h3aef07bb),
	.w7(32'h3ac78ffd),
	.w8(32'h3a4d3391),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7df99),
	.w1(32'h3a4b3c38),
	.w2(32'h3aa4b38f),
	.w3(32'h3a116ec2),
	.w4(32'hb96a16fa),
	.w5(32'hba0d6222),
	.w6(32'hbabb6fb4),
	.w7(32'h38ce4dfd),
	.w8(32'h392c547a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39179888),
	.w1(32'h3a4bcb22),
	.w2(32'h3a5b3844),
	.w3(32'hba358fd7),
	.w4(32'hba6f8e63),
	.w5(32'hbb6b2027),
	.w6(32'h3816e2a9),
	.w7(32'h3a1853b0),
	.w8(32'hbb82b952),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ba06f),
	.w1(32'h3b144673),
	.w2(32'hb9ece5cd),
	.w3(32'h39d78ffb),
	.w4(32'h3a43b35a),
	.w5(32'hbb59e9d7),
	.w6(32'h3b5bbb2c),
	.w7(32'h3a413840),
	.w8(32'h3a7314ac),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01bb08),
	.w1(32'hb919067e),
	.w2(32'hb9456482),
	.w3(32'hbba6b3ff),
	.w4(32'hbb36194b),
	.w5(32'hbb03fc97),
	.w6(32'h3b032c6d),
	.w7(32'h3b20eb17),
	.w8(32'hba89c89c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac535b3),
	.w1(32'hbac01740),
	.w2(32'hba88b3a1),
	.w3(32'hb9c27382),
	.w4(32'hba9b1575),
	.w5(32'h3acaf5dc),
	.w6(32'hb8a8f985),
	.w7(32'hba3f2cd8),
	.w8(32'h3a92bb78),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9c6d7),
	.w1(32'hba246412),
	.w2(32'h394777dd),
	.w3(32'h3accb819),
	.w4(32'h398442e0),
	.w5(32'hb5de0351),
	.w6(32'hba7a5fd6),
	.w7(32'hba9d9976),
	.w8(32'hb94e6270),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0deea3),
	.w1(32'h38ecd1a2),
	.w2(32'h38d423ce),
	.w3(32'h3905c46d),
	.w4(32'hb9a23b97),
	.w5(32'h3a791a93),
	.w6(32'hba13cd31),
	.w7(32'hba8960ff),
	.w8(32'h3a813a24),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd5e0c),
	.w1(32'h3acbb17b),
	.w2(32'h3b01c541),
	.w3(32'h3a8c11d2),
	.w4(32'hba34e523),
	.w5(32'h3ab666d8),
	.w6(32'h3af7c1f4),
	.w7(32'h3af058cd),
	.w8(32'h3a618520),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53d22b),
	.w1(32'hb9c43846),
	.w2(32'hbaaab512),
	.w3(32'h3a071f89),
	.w4(32'hba2ef029),
	.w5(32'h3a6d7e9f),
	.w6(32'hb9a06645),
	.w7(32'hba77794f),
	.w8(32'h39205434),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92ae79a),
	.w1(32'hba4e09ea),
	.w2(32'h38e2e858),
	.w3(32'h38e86b41),
	.w4(32'h3a410718),
	.w5(32'hba319fe4),
	.w6(32'hb87ae125),
	.w7(32'h3888cd57),
	.w8(32'hba209742),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c725d),
	.w1(32'hbaad888a),
	.w2(32'hba2d0dd2),
	.w3(32'hba77c62c),
	.w4(32'hba271372),
	.w5(32'h3a9d8665),
	.w6(32'hbabbc259),
	.w7(32'hb98aec12),
	.w8(32'hba5746a6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895957e),
	.w1(32'h39c1f26f),
	.w2(32'h3a3e1413),
	.w3(32'h392de015),
	.w4(32'hba52c55f),
	.w5(32'hba8bbcc3),
	.w6(32'hba5f634d),
	.w7(32'hba90373a),
	.w8(32'h39c56989),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7304579),
	.w1(32'h398c9c36),
	.w2(32'hb9df2693),
	.w3(32'hb97d1d32),
	.w4(32'hba3f5922),
	.w5(32'h3a04b26a),
	.w6(32'hb969494d),
	.w7(32'hb9b4fa65),
	.w8(32'h3a80f65f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93c8d5),
	.w1(32'h3abbe09c),
	.w2(32'h3ab00875),
	.w3(32'h3a3fe855),
	.w4(32'h3ab121d5),
	.w5(32'h3ab06bc7),
	.w6(32'h3b5cf6e6),
	.w7(32'h3b2c398d),
	.w8(32'h3a0cc005),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abc6d6),
	.w1(32'h3a0459f2),
	.w2(32'hb990f406),
	.w3(32'h3a971ddc),
	.w4(32'h3a939c77),
	.w5(32'h3a7dfa29),
	.w6(32'h3a69ad58),
	.w7(32'hba20f216),
	.w8(32'h3a15702f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a9eb6),
	.w1(32'h3aac4f09),
	.w2(32'h3a617404),
	.w3(32'h3ab02d2f),
	.w4(32'h3a3c2365),
	.w5(32'hb9e5aaa4),
	.w6(32'h3b1efa43),
	.w7(32'h3a4a1c79),
	.w8(32'hba253a2c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb08db),
	.w1(32'hbaa39029),
	.w2(32'h3aa298b6),
	.w3(32'hba221110),
	.w4(32'hba4d16b4),
	.w5(32'h3a0a0228),
	.w6(32'hbad05b38),
	.w7(32'h385455f4),
	.w8(32'hb94dfa4e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913e657),
	.w1(32'hbabc49df),
	.w2(32'hbaa5b6f1),
	.w3(32'h398b7d86),
	.w4(32'hb8b1dae4),
	.w5(32'hb9883155),
	.w6(32'h3914f285),
	.w7(32'hba15f9f3),
	.w8(32'h3a478bbf),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4baac),
	.w1(32'h3ae9a2dd),
	.w2(32'h3aafb155),
	.w3(32'h38eae0d8),
	.w4(32'hb9b84e8a),
	.w5(32'hba798e8d),
	.w6(32'h3aac35f1),
	.w7(32'h39f5c0a7),
	.w8(32'hba1d311b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba833c99),
	.w1(32'hb9d7629c),
	.w2(32'hba115f79),
	.w3(32'hb9f3bc98),
	.w4(32'h36fe5b7d),
	.w5(32'h3ac61e69),
	.w6(32'hb9f118c7),
	.w7(32'hb8647e05),
	.w8(32'h3ad94d28),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3f91b),
	.w1(32'hbb549c83),
	.w2(32'h3a2d3cb4),
	.w3(32'hbb4b3fff),
	.w4(32'h3ab4f3b2),
	.w5(32'h3a6e7f60),
	.w6(32'hba2d9d48),
	.w7(32'h3af6650e),
	.w8(32'h3a098e96),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a496c3a),
	.w1(32'h39bf92a7),
	.w2(32'hbac6ae35),
	.w3(32'h3a87fc27),
	.w4(32'hbaad59eb),
	.w5(32'hbb28503d),
	.w6(32'hb9af5933),
	.w7(32'hbaf05cbc),
	.w8(32'hbb5a61c3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b0243),
	.w1(32'hbb691321),
	.w2(32'hbb5f1554),
	.w3(32'hbb833aea),
	.w4(32'h39564381),
	.w5(32'hbace2810),
	.w6(32'hba10b06c),
	.w7(32'hba23453a),
	.w8(32'hba7ee6ed),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268f87),
	.w1(32'hbb33ecf2),
	.w2(32'hbb8827fd),
	.w3(32'hb9c4dcaf),
	.w4(32'hbacfcc3f),
	.w5(32'h3ab366d1),
	.w6(32'h39cd6abd),
	.w7(32'hbb0c1dd6),
	.w8(32'h3a567863),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba282e31),
	.w1(32'hbadfd6d3),
	.w2(32'hbaebc839),
	.w3(32'h3a16bc67),
	.w4(32'hb997bae6),
	.w5(32'hb9c8158a),
	.w6(32'hb959d2f8),
	.w7(32'hba11fd4a),
	.w8(32'hbaa5fef2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f8499),
	.w1(32'h39698dbb),
	.w2(32'h385734da),
	.w3(32'h396d0004),
	.w4(32'h3a4c5668),
	.w5(32'h3aaf3d94),
	.w6(32'h3aa04469),
	.w7(32'h3ab21d2d),
	.w8(32'hba6b21e7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f99eaa),
	.w1(32'hb9ddfc5f),
	.w2(32'hb9b41502),
	.w3(32'h3a99e3d9),
	.w4(32'h39b2185c),
	.w5(32'h3a8010e0),
	.w6(32'h3a892d0e),
	.w7(32'hbaa02dcc),
	.w8(32'h3a2fd9d0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cddfc6),
	.w1(32'hba04e55c),
	.w2(32'hb8222e40),
	.w3(32'h39e1acbb),
	.w4(32'h3a2223e7),
	.w5(32'hba461092),
	.w6(32'h3948a978),
	.w7(32'h3960f669),
	.w8(32'hba94f518),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10a65f),
	.w1(32'h3993d3da),
	.w2(32'h3949307f),
	.w3(32'hb90dec7e),
	.w4(32'hbad0208c),
	.w5(32'h3971739e),
	.w6(32'h3a9c9384),
	.w7(32'hb75081b2),
	.w8(32'h3aaff366),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0231c8),
	.w1(32'hbb00ad9a),
	.w2(32'hbb2430c2),
	.w3(32'hba465026),
	.w4(32'hbb17459f),
	.w5(32'hbb491a2f),
	.w6(32'h389c3f08),
	.w7(32'hbb34ab74),
	.w8(32'hbaccd55c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a850c53),
	.w1(32'h3ae8dad9),
	.w2(32'h3c0cce23),
	.w3(32'h3b83264b),
	.w4(32'hbae6c250),
	.w5(32'h3b8093d3),
	.w6(32'h3c0f133b),
	.w7(32'h3aef64c7),
	.w8(32'h3bacfd63),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84f9e7),
	.w1(32'h3c0db999),
	.w2(32'h39ce6d05),
	.w3(32'hbbbb0558),
	.w4(32'hbb17e08f),
	.w5(32'hbbd188f4),
	.w6(32'h3b5caa16),
	.w7(32'h3a979f9e),
	.w8(32'h3b108a7d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43a216),
	.w1(32'h3c4976c2),
	.w2(32'h3c025b68),
	.w3(32'hbbf49377),
	.w4(32'hbba053e0),
	.w5(32'hbb11bd92),
	.w6(32'hbb183e61),
	.w7(32'h3b1a9052),
	.w8(32'h36b18b4c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a25bc),
	.w1(32'h3a028f4a),
	.w2(32'h399fd367),
	.w3(32'h382231d2),
	.w4(32'hbac43955),
	.w5(32'hbb34b9cd),
	.w6(32'h39c15691),
	.w7(32'hbb1c788a),
	.w8(32'h3ac01948),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7876ca),
	.w1(32'h3b8be7af),
	.w2(32'h3b3a0b05),
	.w3(32'h3b62dfbb),
	.w4(32'hbbd913f4),
	.w5(32'h3b370c93),
	.w6(32'h3aa16a9f),
	.w7(32'hbbd33c6c),
	.w8(32'hbc04bc31),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b075703),
	.w1(32'hba80e71b),
	.w2(32'hbb848bf2),
	.w3(32'hbc074c4a),
	.w4(32'hbaa3d670),
	.w5(32'hb8ce203e),
	.w6(32'h3c2e036b),
	.w7(32'hbb6c0e94),
	.w8(32'hba8b9dad),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e319e),
	.w1(32'hba10b4be),
	.w2(32'h3b5fb41f),
	.w3(32'h3b5a0d3d),
	.w4(32'h3b4589ab),
	.w5(32'hbbe2d87e),
	.w6(32'h3b215417),
	.w7(32'h3b676184),
	.w8(32'hbc2c376a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a8142),
	.w1(32'h3a159628),
	.w2(32'h3b4921e4),
	.w3(32'hbc19df3e),
	.w4(32'hbbaccb16),
	.w5(32'hba2eac7f),
	.w6(32'h3a55c559),
	.w7(32'hbb480a2f),
	.w8(32'h3b0ac3ce),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6632ca),
	.w1(32'h3bb3ec8b),
	.w2(32'h3bce79aa),
	.w3(32'h3bb46885),
	.w4(32'h3b119c0d),
	.w5(32'hba1926d1),
	.w6(32'h3c34c190),
	.w7(32'h3b4ef47c),
	.w8(32'h3b4afa71),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ec185),
	.w1(32'h3a3a02c3),
	.w2(32'h3aaf232d),
	.w3(32'h3acf1478),
	.w4(32'hba3731e5),
	.w5(32'hbb1f44ca),
	.w6(32'h3a36bf09),
	.w7(32'hb98ea6d4),
	.w8(32'hbb19935a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4841b),
	.w1(32'hba533476),
	.w2(32'hbbad0644),
	.w3(32'hba886012),
	.w4(32'hbb519d8c),
	.w5(32'hbb790078),
	.w6(32'h39d0f81e),
	.w7(32'hbb42dce5),
	.w8(32'hbb88d737),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc13c87),
	.w1(32'h3b1082b3),
	.w2(32'hb9b65f14),
	.w3(32'hbbde3cc1),
	.w4(32'hbb9eece7),
	.w5(32'hbb68b08c),
	.w6(32'h3a8d3179),
	.w7(32'hbb9c818a),
	.w8(32'hbb961e5c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb506e94),
	.w1(32'h3a620895),
	.w2(32'h3b11270d),
	.w3(32'h3829b3c1),
	.w4(32'h3b00572a),
	.w5(32'hbb5d4b61),
	.w6(32'h3b8d107e),
	.w7(32'h3ba0a644),
	.w8(32'hbb699b8e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a68fb),
	.w1(32'h3b1a1223),
	.w2(32'hbc0445c8),
	.w3(32'hbbc0cb7b),
	.w4(32'hbbe12f0a),
	.w5(32'h38865ae8),
	.w6(32'h3b8b997a),
	.w7(32'hbbcf901c),
	.w8(32'h399ed647),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb244bc2),
	.w1(32'h39b2648c),
	.w2(32'h3b5dbccf),
	.w3(32'hba4f5ee9),
	.w4(32'h39fa512b),
	.w5(32'h3c0a7ed1),
	.w6(32'hbb00f1f1),
	.w7(32'hba03d824),
	.w8(32'h3bb78abb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b974bf4),
	.w1(32'hbc10f27a),
	.w2(32'h3c0b1163),
	.w3(32'h3b885475),
	.w4(32'h3bfdf1e2),
	.w5(32'hbb461cfa),
	.w6(32'hbc1b24b1),
	.w7(32'h3c32d2ff),
	.w8(32'hbb20aa2d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3cf92),
	.w1(32'h3b8d6e2e),
	.w2(32'h3b864f77),
	.w3(32'hbb8713c6),
	.w4(32'h3b0d2677),
	.w5(32'h398cc447),
	.w6(32'h388e5ab6),
	.w7(32'h3bdb09a3),
	.w8(32'hb9972666),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d30f5),
	.w1(32'hba7de830),
	.w2(32'hbb612795),
	.w3(32'hbb30e28c),
	.w4(32'hbb135319),
	.w5(32'h3c08db1f),
	.w6(32'hbb4dbf2c),
	.w7(32'hbab5893c),
	.w8(32'h39c34784),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf226ad),
	.w1(32'hbaf7c5fa),
	.w2(32'hbb934849),
	.w3(32'h3ba82611),
	.w4(32'h3c29a588),
	.w5(32'h3add1a4d),
	.w6(32'h3c429160),
	.w7(32'hbaa07def),
	.w8(32'h3b586906),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ebeb4),
	.w1(32'h3982b5ed),
	.w2(32'h397020fe),
	.w3(32'h391d40f0),
	.w4(32'h3bb0a7df),
	.w5(32'hbbb4737a),
	.w6(32'h3bdcf7d3),
	.w7(32'h3b946a16),
	.w8(32'hbb2c04a0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce556),
	.w1(32'hbc050178),
	.w2(32'hbbc3980c),
	.w3(32'hbb2f55ef),
	.w4(32'hbb943303),
	.w5(32'hbb3d9a0a),
	.w6(32'hbbbb90f9),
	.w7(32'hbbbef92c),
	.w8(32'hbb193d6d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f0b1b),
	.w1(32'h3bac1805),
	.w2(32'h3b2e8abd),
	.w3(32'hba364a7c),
	.w4(32'h3bc25bc4),
	.w5(32'h390a503f),
	.w6(32'hbb86023b),
	.w7(32'h3ba94142),
	.w8(32'hbb596c8a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae52fd),
	.w1(32'hbb712920),
	.w2(32'h3b7644e2),
	.w3(32'h3b2cea46),
	.w4(32'h3a975e0a),
	.w5(32'hbb5a2205),
	.w6(32'hb980eaba),
	.w7(32'h397bafbf),
	.w8(32'hbb64999e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a095771),
	.w1(32'h3be4157d),
	.w2(32'h3afbe583),
	.w3(32'hbad9cdda),
	.w4(32'hbb9293f5),
	.w5(32'hbbe74496),
	.w6(32'h3b19a8f5),
	.w7(32'hb899ff0e),
	.w8(32'hbb416564),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac27056),
	.w1(32'hbb6f797f),
	.w2(32'h3b395b0f),
	.w3(32'hb8e9782a),
	.w4(32'hba91e6c9),
	.w5(32'hba4d25c9),
	.w6(32'h3b5df900),
	.w7(32'h3b3f7bdb),
	.w8(32'hbac6287b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4fb97),
	.w1(32'hba8b3080),
	.w2(32'h3b386962),
	.w3(32'h3a70c153),
	.w4(32'hbb356d93),
	.w5(32'h3ab4f1ed),
	.w6(32'hb95e4294),
	.w7(32'hbb3aa634),
	.w8(32'hbabc3ced),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3b1e4),
	.w1(32'hbb20e7da),
	.w2(32'h3aa91168),
	.w3(32'h3abcad94),
	.w4(32'hbadb88c7),
	.w5(32'hb904739b),
	.w6(32'h3bc07a81),
	.w7(32'h3b39c749),
	.w8(32'hba885ba3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad53fe7),
	.w1(32'hbb3b652c),
	.w2(32'hbba69e22),
	.w3(32'h3adb7188),
	.w4(32'h3b0ba500),
	.w5(32'hba0e6ee3),
	.w6(32'h3a590f99),
	.w7(32'h3a53e637),
	.w8(32'h3bbbc500),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19f42c),
	.w1(32'hbbb4f81e),
	.w2(32'h3b16541d),
	.w3(32'hbb5992cc),
	.w4(32'hbbe06bcc),
	.w5(32'hbab38e41),
	.w6(32'hbbbe0010),
	.w7(32'hbb25815b),
	.w8(32'hbaad5f52),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8a86d),
	.w1(32'hbb5dab52),
	.w2(32'hbbd8d731),
	.w3(32'hbb5676be),
	.w4(32'hbb2779f7),
	.w5(32'hb96a1dc4),
	.w6(32'hbadef7ae),
	.w7(32'hbb7ff1e6),
	.w8(32'hbb7b6469),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba160de4),
	.w1(32'h3a6d13cc),
	.w2(32'hbc0048c6),
	.w3(32'h3b9088fd),
	.w4(32'h3be499fe),
	.w5(32'hbb69d716),
	.w6(32'h3c155548),
	.w7(32'hba0ed879),
	.w8(32'hbabb3705),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba852aa0),
	.w1(32'h3bf27d33),
	.w2(32'h3bea0bf7),
	.w3(32'hbb81ac73),
	.w4(32'h39abdfcb),
	.w5(32'hb99339d3),
	.w6(32'hbb415fba),
	.w7(32'hbac3ee06),
	.w8(32'hb9d1bcb2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15a1f9),
	.w1(32'h3afac13a),
	.w2(32'hbb24a7de),
	.w3(32'h3856d4e9),
	.w4(32'hb9b6a588),
	.w5(32'hbb9097aa),
	.w6(32'h3a8980e5),
	.w7(32'hbaf2a4a1),
	.w8(32'hbb92b3f8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb66d8),
	.w1(32'h3c88c243),
	.w2(32'h3baa5664),
	.w3(32'h38f2a636),
	.w4(32'hbc0ee6e6),
	.w5(32'hba26ec37),
	.w6(32'h3bed0234),
	.w7(32'hbba91939),
	.w8(32'hba9025df),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d80d3),
	.w1(32'h3b030927),
	.w2(32'hbb40f650),
	.w3(32'h390b2aa4),
	.w4(32'hbab7d4b8),
	.w5(32'h3a76f059),
	.w6(32'h3b771bfb),
	.w7(32'hbb0401e2),
	.w8(32'hba9e11e7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea7b12),
	.w1(32'hbb00160a),
	.w2(32'hbb9aaa2f),
	.w3(32'hba7f7e61),
	.w4(32'h3a446ae9),
	.w5(32'h390e614b),
	.w6(32'h39f7bef5),
	.w7(32'hbae6633c),
	.w8(32'hbb82517a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3d897),
	.w1(32'h3b9a2d07),
	.w2(32'hbb9e5a79),
	.w3(32'hba4ab278),
	.w4(32'hbb2d0dd8),
	.w5(32'hbb2e1f74),
	.w6(32'h3b136473),
	.w7(32'hbb5471b6),
	.w8(32'hbb460bc9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87666c),
	.w1(32'hbb1e8051),
	.w2(32'hbbd0716b),
	.w3(32'hbb51ef1e),
	.w4(32'hbbbd8626),
	.w5(32'hbaa92027),
	.w6(32'hbb1b24f1),
	.w7(32'hbbc87235),
	.w8(32'hba630db6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5365c3),
	.w1(32'h39d9ac16),
	.w2(32'hbb828471),
	.w3(32'hbab3f5ac),
	.w4(32'hbabaf97b),
	.w5(32'hba39ba22),
	.w6(32'h3b055ede),
	.w7(32'hbaa3b7fe),
	.w8(32'h3aaeb927),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e6eda),
	.w1(32'h3b37a669),
	.w2(32'hbb0bae63),
	.w3(32'hba8e50c2),
	.w4(32'hbad6f8dc),
	.w5(32'hba1cd23b),
	.w6(32'h3bc53b5d),
	.w7(32'hbad420ef),
	.w8(32'hbb3d09b3),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a38377),
	.w1(32'h3a01079c),
	.w2(32'h3b059b42),
	.w3(32'hbb075e65),
	.w4(32'hbb549c76),
	.w5(32'hba3915fe),
	.w6(32'hba93a2c7),
	.w7(32'hbbb0a902),
	.w8(32'hbb9ef56e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d8c34),
	.w1(32'h3c3dae65),
	.w2(32'h3b94d4a7),
	.w3(32'h3c08a898),
	.w4(32'hb883932f),
	.w5(32'hbb8b90e1),
	.w6(32'h3c2c2cb9),
	.w7(32'hb9fa4c3c),
	.w8(32'hbbe88bbd),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87c983),
	.w1(32'hba0e379d),
	.w2(32'hbb2b463e),
	.w3(32'h3b807084),
	.w4(32'hbb743978),
	.w5(32'hb995818f),
	.w6(32'hbb2bd0de),
	.w7(32'hbb05dcd0),
	.w8(32'h3a5dbaec),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e1594),
	.w1(32'h3b135c88),
	.w2(32'h3b30a851),
	.w3(32'hba9ea6de),
	.w4(32'hb9e048e5),
	.w5(32'hbb0426a9),
	.w6(32'h3b88fd20),
	.w7(32'hb8df8f43),
	.w8(32'hbbde1ff7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b00f6),
	.w1(32'h3be850bb),
	.w2(32'hbb178420),
	.w3(32'hba59efce),
	.w4(32'hbb381977),
	.w5(32'hb9bdf3a8),
	.w6(32'h3bc86fa4),
	.w7(32'hbb93e284),
	.w8(32'hbb5c17be),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b745039),
	.w1(32'h3baf6888),
	.w2(32'h3a598559),
	.w3(32'h3b584b1e),
	.w4(32'h3bea6bf0),
	.w5(32'hbaefe261),
	.w6(32'h3bda89a6),
	.w7(32'h3b1fae62),
	.w8(32'hb9354018),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a802bc5),
	.w1(32'h3a7cfe2a),
	.w2(32'h3a2cf912),
	.w3(32'hba61168d),
	.w4(32'hbb14c285),
	.w5(32'hbc20ce94),
	.w6(32'h3a624f83),
	.w7(32'hbb3f5ab7),
	.w8(32'hbbc854c8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ccbf),
	.w1(32'h3bd7c6fb),
	.w2(32'h3afa713c),
	.w3(32'hbc282993),
	.w4(32'hbb971861),
	.w5(32'hb9e45c36),
	.w6(32'hbb6233c2),
	.w7(32'hbb83d85e),
	.w8(32'hbaf38f5a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0460d2),
	.w1(32'hbbc94c40),
	.w2(32'h3b375253),
	.w3(32'h3b8e8db5),
	.w4(32'h3999965a),
	.w5(32'hbaa3654e),
	.w6(32'h3b8074ac),
	.w7(32'h3bfdfb35),
	.w8(32'hbbb19a00),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1918fd),
	.w1(32'h39284196),
	.w2(32'hbaa53343),
	.w3(32'h3a8603c7),
	.w4(32'h3a9554bf),
	.w5(32'h3b1af59e),
	.w6(32'hbb2428cc),
	.w7(32'h3aff5480),
	.w8(32'hba045af0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebfa28),
	.w1(32'h3ab1635c),
	.w2(32'hbb6c671b),
	.w3(32'hba19d2b6),
	.w4(32'hbae731b9),
	.w5(32'hbb61bfff),
	.w6(32'hbb01918b),
	.w7(32'hbac4621f),
	.w8(32'hbafb9ad9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba943341),
	.w1(32'hb9f58536),
	.w2(32'hbaea58a5),
	.w3(32'hbb85659e),
	.w4(32'hb9e830f6),
	.w5(32'hbb7556b7),
	.w6(32'hbb80fef0),
	.w7(32'hbb070615),
	.w8(32'hbb31bb57),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f0726),
	.w1(32'hbb0b71bf),
	.w2(32'hbb952de1),
	.w3(32'hb9a5d69a),
	.w4(32'hbaeb4e72),
	.w5(32'hbb532727),
	.w6(32'h38ac35fb),
	.w7(32'hbb74b275),
	.w8(32'hba6f2178),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cdcdf),
	.w1(32'h3aada78d),
	.w2(32'hb9884af5),
	.w3(32'hbb37cadb),
	.w4(32'hba866803),
	.w5(32'hbb25780d),
	.w6(32'hbbada2fa),
	.w7(32'h3b1f7625),
	.w8(32'h3b59fdfb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0cb45),
	.w1(32'h3bbfeef6),
	.w2(32'h3b05bf93),
	.w3(32'hbb38441b),
	.w4(32'hbb25814c),
	.w5(32'hba2a732c),
	.w6(32'h3b770028),
	.w7(32'hb9f34171),
	.w8(32'hb90153e9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad66f4a),
	.w1(32'h3bb06e90),
	.w2(32'h3a943a40),
	.w3(32'hbb878721),
	.w4(32'h3ac12169),
	.w5(32'hbb7f26c3),
	.w6(32'hbb51fb2a),
	.w7(32'hbb17487e),
	.w8(32'hbb92f806),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4a2ef),
	.w1(32'hbb3e8489),
	.w2(32'hbbf3680b),
	.w3(32'hbb793779),
	.w4(32'hbbb5ae23),
	.w5(32'h39d5a4a8),
	.w6(32'hbb30983a),
	.w7(32'hbbc5409d),
	.w8(32'hba49d1f7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66def4),
	.w1(32'hbb4b70a5),
	.w2(32'hbb8c1842),
	.w3(32'h3a4d8f8c),
	.w4(32'hb9fa4833),
	.w5(32'hbb785554),
	.w6(32'hba98536f),
	.w7(32'hbb8a1483),
	.w8(32'hbb55fcdf),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b3e41),
	.w1(32'hbc03c5f3),
	.w2(32'h3bec1653),
	.w3(32'hba596aa0),
	.w4(32'h3b0d2aea),
	.w5(32'h3b6d82aa),
	.w6(32'hbbcd185e),
	.w7(32'h3bcbf127),
	.w8(32'h3c5325e2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc096ddc),
	.w1(32'hbbee69a0),
	.w2(32'hba669e7f),
	.w3(32'hb7fa5f57),
	.w4(32'h39da13e7),
	.w5(32'hbbc12a1a),
	.w6(32'h3b13727f),
	.w7(32'hb8ae438b),
	.w8(32'hbc1fff06),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beea002),
	.w1(32'h3b9155e8),
	.w2(32'h3b6775ac),
	.w3(32'h39971212),
	.w4(32'hbb3a4d60),
	.w5(32'hbb9ff994),
	.w6(32'hbb6193cb),
	.w7(32'hbb0726e3),
	.w8(32'h3b4393a2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c0040c),
	.w1(32'h3bd23563),
	.w2(32'h3bb8e735),
	.w3(32'hbc112d07),
	.w4(32'hb9ba82cb),
	.w5(32'h3b21a460),
	.w6(32'hbc337639),
	.w7(32'h3a7dd4ed),
	.w8(32'h3b167181),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b837785),
	.w1(32'hbbb324b8),
	.w2(32'h3b43707f),
	.w3(32'h3ba3818b),
	.w4(32'h3b9c76d8),
	.w5(32'h3b164a47),
	.w6(32'h3c03c2ea),
	.w7(32'h3b689fd6),
	.w8(32'h3b30722b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba073b94),
	.w1(32'hbb6859ba),
	.w2(32'hbb48b939),
	.w3(32'h3b93f362),
	.w4(32'h3b520bf1),
	.w5(32'hbb55e63b),
	.w6(32'h3a4f41b1),
	.w7(32'h3b68c118),
	.w8(32'h3b1fb9ad),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae21eba),
	.w1(32'hbb240f25),
	.w2(32'h3b0b0cba),
	.w3(32'hba2e39d6),
	.w4(32'hb96926da),
	.w5(32'hba8599cf),
	.w6(32'h3ba2e0d5),
	.w7(32'h3c04e999),
	.w8(32'hbbb830a5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39819edc),
	.w1(32'h3b5528ed),
	.w2(32'hbbb4b1fc),
	.w3(32'hbbdfcde6),
	.w4(32'h3b50b943),
	.w5(32'hb992c4d3),
	.w6(32'h3bc5abf7),
	.w7(32'hbaba97ef),
	.w8(32'hbb091647),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51900e),
	.w1(32'h3b77922b),
	.w2(32'hbad6ee7d),
	.w3(32'hbb98b58e),
	.w4(32'hbaf3fba8),
	.w5(32'hbb262b11),
	.w6(32'h3b6c563c),
	.w7(32'hbb9a9986),
	.w8(32'hbb4bc921),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd73db),
	.w1(32'hb9ce3253),
	.w2(32'hbb41c835),
	.w3(32'hbba770ed),
	.w4(32'h3a93806e),
	.w5(32'hbb853f0e),
	.w6(32'h3acaaec8),
	.w7(32'hbb821e6b),
	.w8(32'hbbe51858),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bdab6),
	.w1(32'h3b531241),
	.w2(32'hbbdf506a),
	.w3(32'h3b75cd24),
	.w4(32'hbc1b5f67),
	.w5(32'hba71e216),
	.w6(32'h3bf1cd5a),
	.w7(32'hbc088967),
	.w8(32'hbb71936f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39698558),
	.w1(32'hbb294811),
	.w2(32'hbace332a),
	.w3(32'h3ab1b9d4),
	.w4(32'hbbbc642c),
	.w5(32'h3ac35e07),
	.w6(32'hbb00599d),
	.w7(32'hbb1fa4ba),
	.w8(32'h3b4ef6cf),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d1087),
	.w1(32'h3b8acbcd),
	.w2(32'hb9954726),
	.w3(32'hba95b860),
	.w4(32'h3b51e200),
	.w5(32'hbba1cccf),
	.w6(32'h3b5ac26e),
	.w7(32'h3a50b18a),
	.w8(32'hbba229b4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1077ab),
	.w1(32'hbb945a6c),
	.w2(32'hbb45e2d8),
	.w3(32'hbc2d468c),
	.w4(32'hbc00905e),
	.w5(32'hbb89c86d),
	.w6(32'hbb21061f),
	.w7(32'hbc0be60d),
	.w8(32'hba197dfe),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4757d),
	.w1(32'hb8ff49b9),
	.w2(32'h3a656ed0),
	.w3(32'hbc1b5912),
	.w4(32'h3b9ad468),
	.w5(32'hbb1c6dd9),
	.w6(32'h3c35fd8e),
	.w7(32'h3bb92be9),
	.w8(32'h3b789046),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b562382),
	.w1(32'hba7bfa33),
	.w2(32'hbbb284d1),
	.w3(32'hbb53ecf2),
	.w4(32'hbba9e87c),
	.w5(32'h3c1994e0),
	.w6(32'hbbc89c79),
	.w7(32'hbadce707),
	.w8(32'h3c728e99),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03e5e8),
	.w1(32'h3b390f4a),
	.w2(32'h3a85551f),
	.w3(32'h3bb6d5cb),
	.w4(32'h3b81a99f),
	.w5(32'hb96d212d),
	.w6(32'h3c8dc3fc),
	.w7(32'h3bf01d7b),
	.w8(32'h3bda8a1d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c127378),
	.w1(32'h3c243f4e),
	.w2(32'h3a3ac4aa),
	.w3(32'hba59c6be),
	.w4(32'hbb8b9141),
	.w5(32'h3b248229),
	.w6(32'h3c2e620a),
	.w7(32'hbb9ddda5),
	.w8(32'hbaf25407),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b214a96),
	.w1(32'h3bb7d159),
	.w2(32'hbb791aa9),
	.w3(32'h3a5e0fcc),
	.w4(32'hbb7768e9),
	.w5(32'hbb0faf58),
	.w6(32'h3b38e495),
	.w7(32'hbbd43461),
	.w8(32'h3ac4b2e6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba059e66),
	.w1(32'hbb1c4fb9),
	.w2(32'hbb4ee5cf),
	.w3(32'hb9824a5d),
	.w4(32'hba17e977),
	.w5(32'hb9c72d03),
	.w6(32'h3bb8c686),
	.w7(32'h3af92ae8),
	.w8(32'hbb78eef8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1eb104),
	.w1(32'h3b9da769),
	.w2(32'hbb91ba2e),
	.w3(32'hbab1dfd7),
	.w4(32'hbb68f045),
	.w5(32'hbbc6b5c2),
	.w6(32'hba609dea),
	.w7(32'hbb7d11c8),
	.w8(32'hbc29c419),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9384ad),
	.w1(32'hbb3d2553),
	.w2(32'h3bb35353),
	.w3(32'h3ab946fa),
	.w4(32'h3bc03f07),
	.w5(32'h3befea67),
	.w6(32'hbc1eaeb3),
	.w7(32'h3bc4cdae),
	.w8(32'h3a4fef91),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08c569),
	.w1(32'hbb86ab78),
	.w2(32'hbba73181),
	.w3(32'h3b68444e),
	.w4(32'h3c070ac7),
	.w5(32'hbae2f2b5),
	.w6(32'h396a26d5),
	.w7(32'h3a22928e),
	.w8(32'hbaff9024),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15ae2a),
	.w1(32'h3ac5959a),
	.w2(32'hbb0e06b9),
	.w3(32'hbb504cd6),
	.w4(32'hbb3de066),
	.w5(32'hbab90b33),
	.w6(32'h3b068f25),
	.w7(32'h3a8764a0),
	.w8(32'h386a9b49),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fc3b1),
	.w1(32'hb9fbccd9),
	.w2(32'h3b062485),
	.w3(32'h3b9e3622),
	.w4(32'h3b818e63),
	.w5(32'h3adf1032),
	.w6(32'hbad4f42e),
	.w7(32'h3b064010),
	.w8(32'h3b71c3b4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b877f3c),
	.w1(32'hbabf6c80),
	.w2(32'hb9f1c331),
	.w3(32'h3b9567e7),
	.w4(32'hbb1202e2),
	.w5(32'h3b14a53d),
	.w6(32'hb7e9941e),
	.w7(32'h3b8174ef),
	.w8(32'hbb0d8331),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba005dfb),
	.w1(32'hba48a864),
	.w2(32'hbb1b33f3),
	.w3(32'h3b6c732c),
	.w4(32'h3b38b7b4),
	.w5(32'hb9b08092),
	.w6(32'hbb6570f3),
	.w7(32'h3b5f088e),
	.w8(32'hbb1c6d0d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a450dd),
	.w1(32'hbb377717),
	.w2(32'hba2b0ffc),
	.w3(32'h3b772302),
	.w4(32'h39866ca8),
	.w5(32'hbb65a02e),
	.w6(32'hbab10eeb),
	.w7(32'h39dcb299),
	.w8(32'hbbbc166a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb824781d),
	.w1(32'hbaf0b0a4),
	.w2(32'hbb496372),
	.w3(32'hbb9f5dc2),
	.w4(32'h3a935f2d),
	.w5(32'hba8de20e),
	.w6(32'h3becc04a),
	.w7(32'hb9f752df),
	.w8(32'hbb8aa22a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba898306),
	.w1(32'h3a83458c),
	.w2(32'hbb86f28d),
	.w3(32'hbb6fb298),
	.w4(32'hbb8eb6d4),
	.w5(32'h3bba937b),
	.w6(32'hbb226b22),
	.w7(32'hbb6bcc3a),
	.w8(32'h3b8251bd),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cfc6e),
	.w1(32'h3be65ead),
	.w2(32'hbb94714b),
	.w3(32'hbba97c92),
	.w4(32'hbb9d3038),
	.w5(32'hbac15af9),
	.w6(32'h3aa50bcb),
	.w7(32'hbb83739e),
	.w8(32'hbb7171e4),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb126c1e),
	.w1(32'hba07547f),
	.w2(32'hbb15e7f6),
	.w3(32'hbb330d96),
	.w4(32'hba97b431),
	.w5(32'hbb8308c6),
	.w6(32'h3ac5cceb),
	.w7(32'hbb0cab81),
	.w8(32'h3a6a36dc),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12a249),
	.w1(32'h3ba1be90),
	.w2(32'hbb9e04cf),
	.w3(32'hbb8c0abb),
	.w4(32'hb98d73b1),
	.w5(32'hbb33d94a),
	.w6(32'h3b90a98a),
	.w7(32'h3a67a98c),
	.w8(32'h393a38fe),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81fc91),
	.w1(32'h3afd7fa9),
	.w2(32'h3a692eba),
	.w3(32'hbb490175),
	.w4(32'hba7c26fb),
	.w5(32'hbb4ab0bc),
	.w6(32'h396ae4a8),
	.w7(32'hbaa36c52),
	.w8(32'hbb95dc01),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb796488),
	.w1(32'hbb4364fb),
	.w2(32'hb6b5458b),
	.w3(32'h3b9a29b8),
	.w4(32'h3aa30d69),
	.w5(32'hba8b173d),
	.w6(32'hbabc94db),
	.w7(32'hbaf3c0e5),
	.w8(32'hbb18dc03),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912da6),
	.w1(32'hbbd5944e),
	.w2(32'hbb48ffe1),
	.w3(32'h3a6cba53),
	.w4(32'h3a4b7f91),
	.w5(32'hba8e8783),
	.w6(32'hbb474dcd),
	.w7(32'h3b9461f9),
	.w8(32'hba96a65f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafa146),
	.w1(32'h38d84ba8),
	.w2(32'hb9d34fca),
	.w3(32'hbaee5a12),
	.w4(32'hbbf983df),
	.w5(32'hbb07c190),
	.w6(32'h39416b2a),
	.w7(32'hb926aaca),
	.w8(32'hbb8c2134),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac53ae1),
	.w1(32'h3a6d662d),
	.w2(32'hbab712ae),
	.w3(32'h3a8da244),
	.w4(32'hbb2f4992),
	.w5(32'h3af27f76),
	.w6(32'h3bb2f848),
	.w7(32'hbb9c9c30),
	.w8(32'h3b81c0c1),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c59b0),
	.w1(32'h38bcf025),
	.w2(32'h3b72b457),
	.w3(32'h3b98de60),
	.w4(32'h3a44609a),
	.w5(32'h3a0467c6),
	.w6(32'h3c153bdb),
	.w7(32'h3ad5be15),
	.w8(32'hb9a5b136),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b81bac),
	.w1(32'hba7714fe),
	.w2(32'h3bf2fdd6),
	.w3(32'hba54dcd6),
	.w4(32'hbae72ef4),
	.w5(32'h3ac9585b),
	.w6(32'hbbd2c5c7),
	.w7(32'h3b8a59b6),
	.w8(32'h3ac1fc39),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39a94c),
	.w1(32'hba000308),
	.w2(32'h3aee6e47),
	.w3(32'hbb6be8ea),
	.w4(32'h3b58ce18),
	.w5(32'hbb64f43e),
	.w6(32'h3c1fc84f),
	.w7(32'h3b0620b3),
	.w8(32'hbb6de381),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd40c6),
	.w1(32'h3a0ac336),
	.w2(32'hb9aef063),
	.w3(32'hbb2ead51),
	.w4(32'h3aa2ab9b),
	.w5(32'h3b3d4399),
	.w6(32'h3ae5926f),
	.w7(32'hbaa96d7d),
	.w8(32'hbb7a052f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c3f55),
	.w1(32'h3ba1d835),
	.w2(32'h3a82f27b),
	.w3(32'hbaad97b8),
	.w4(32'h3a9e779a),
	.w5(32'hbb7dce9f),
	.w6(32'h3beb8823),
	.w7(32'h3b259700),
	.w8(32'hbb836591),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba977752),
	.w1(32'hbad13e11),
	.w2(32'hbb8c513e),
	.w3(32'hbbc1ca2a),
	.w4(32'hba9210d7),
	.w5(32'h3bc510d5),
	.w6(32'hbae5ddd7),
	.w7(32'hbab1c522),
	.w8(32'h3bfec1d6),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f43e7),
	.w1(32'hbbd51abe),
	.w2(32'h3a2bf579),
	.w3(32'h3c320e27),
	.w4(32'h3c17c28b),
	.w5(32'hbb4fd771),
	.w6(32'h3c7acc4a),
	.w7(32'h3bb9d465),
	.w8(32'hbaacc6f9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99e81a),
	.w1(32'h3b415a2d),
	.w2(32'hbb76f23c),
	.w3(32'hbb120456),
	.w4(32'hbb9c860f),
	.w5(32'hbb444dac),
	.w6(32'h3be53c3b),
	.w7(32'hbb4d19e2),
	.w8(32'h3a4b676f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0013e5),
	.w1(32'hbac9b228),
	.w2(32'h3b3d3d04),
	.w3(32'h3b99b4fa),
	.w4(32'hbadf054f),
	.w5(32'hbae09880),
	.w6(32'h3b2f6f64),
	.w7(32'h3a0eb9bf),
	.w8(32'hbb4954b7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b3408),
	.w1(32'hb9820fdd),
	.w2(32'hba30460c),
	.w3(32'hbb5b04af),
	.w4(32'hbb796969),
	.w5(32'h3b235ec5),
	.w6(32'h3a4857a7),
	.w7(32'hbb7da6a6),
	.w8(32'h3b0bdee1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a1324),
	.w1(32'hbb4fd7c9),
	.w2(32'hbb25c20a),
	.w3(32'hba06d0b7),
	.w4(32'hbbbebd7a),
	.w5(32'h3ba582c0),
	.w6(32'h3b652565),
	.w7(32'hba40b098),
	.w8(32'h3bb46380),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152eaf),
	.w1(32'h3c18de9b),
	.w2(32'h3b072886),
	.w3(32'h3bc9ed8f),
	.w4(32'hb858e33c),
	.w5(32'hb81bf111),
	.w6(32'h3c5f7f28),
	.w7(32'hbaba4f5e),
	.w8(32'hbb10c8ca),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96cca88),
	.w1(32'hbb0a7bba),
	.w2(32'hbafb5152),
	.w3(32'h3aef5a78),
	.w4(32'h3b13d216),
	.w5(32'hbba474fe),
	.w6(32'h3bd3f7ec),
	.w7(32'hb9d571f8),
	.w8(32'hbc014ad8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8b96c),
	.w1(32'hbbcf0a92),
	.w2(32'hbbaf0e88),
	.w3(32'hba2dffe9),
	.w4(32'hbbe666e8),
	.w5(32'hbba6136a),
	.w6(32'hbb0a17ec),
	.w7(32'hbb8cf577),
	.w8(32'h39fe0de6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994173),
	.w1(32'hbac3bf73),
	.w2(32'hbb76a9a4),
	.w3(32'hbbb32d27),
	.w4(32'hbbcf514f),
	.w5(32'hbaab7fa1),
	.w6(32'h3b43dba8),
	.w7(32'hba93f7f1),
	.w8(32'hba4a0fcd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e438ac),
	.w1(32'h3b337555),
	.w2(32'h3b5b772d),
	.w3(32'hbb3eb38a),
	.w4(32'hbaa457e1),
	.w5(32'h3b9d33f9),
	.w6(32'hbb48cecd),
	.w7(32'h394d30f0),
	.w8(32'h3b42fa3e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf26d65),
	.w1(32'h3c219465),
	.w2(32'h3c889fe1),
	.w3(32'h370611b6),
	.w4(32'h3b7892e3),
	.w5(32'hbb61f58d),
	.w6(32'h3c392665),
	.w7(32'h3b980777),
	.w8(32'h3a5617c1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb1b23),
	.w1(32'h3af7e656),
	.w2(32'h3bbc5810),
	.w3(32'hbb4822d6),
	.w4(32'hbb294f3f),
	.w5(32'h39994be1),
	.w6(32'hbb16dbe7),
	.w7(32'h3a714499),
	.w8(32'h3b1d1557),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b365fab),
	.w1(32'h3aba7486),
	.w2(32'h3bf7a461),
	.w3(32'hb921b1c0),
	.w4(32'h3b574b0d),
	.w5(32'hbb7b2ee9),
	.w6(32'h3be46be3),
	.w7(32'h3b8cf1b7),
	.w8(32'hbb8b272f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74f852),
	.w1(32'h3c3bf424),
	.w2(32'hbb5e68dd),
	.w3(32'hbbd9b4ae),
	.w4(32'hbb714674),
	.w5(32'h39fa3b84),
	.w6(32'h3b863c0a),
	.w7(32'hbbfb7548),
	.w8(32'hbb03f8fc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab85ddd),
	.w1(32'hbb775758),
	.w2(32'hb9ba8f49),
	.w3(32'h3a43a974),
	.w4(32'h3ad9d9d5),
	.w5(32'hba90bce6),
	.w6(32'hb9020104),
	.w7(32'hba458d55),
	.w8(32'hbb9d8afb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ca067),
	.w1(32'h3b50b682),
	.w2(32'hbb61b2fe),
	.w3(32'hb89bafc5),
	.w4(32'h3a989698),
	.w5(32'hbb66eba6),
	.w6(32'h3b4bd556),
	.w7(32'hbb2697ee),
	.w8(32'h3a348d9a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e71b46),
	.w1(32'hbb524853),
	.w2(32'h3b2b17e1),
	.w3(32'h3bf745ce),
	.w4(32'hba3adb08),
	.w5(32'h39c87243),
	.w6(32'hb8ac35d3),
	.w7(32'h3af02a53),
	.w8(32'h3ab9b153),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9a06b),
	.w1(32'hbbbd3580),
	.w2(32'hb9a5ae1f),
	.w3(32'h3b6b032f),
	.w4(32'hbaad3e54),
	.w5(32'hbb12eabe),
	.w6(32'h3acb4e10),
	.w7(32'h38a12213),
	.w8(32'h3c095970),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05554d),
	.w1(32'h3932b6f2),
	.w2(32'h3bbc8a2e),
	.w3(32'hbb897c44),
	.w4(32'h3c05b182),
	.w5(32'h3b4ae5ec),
	.w6(32'hbc02b338),
	.w7(32'h3c03efd8),
	.w8(32'h3b4d9081),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a6943),
	.w1(32'h3c404e25),
	.w2(32'h3ba8ca93),
	.w3(32'h3b7252e4),
	.w4(32'h3af6cd4f),
	.w5(32'hba87ba6a),
	.w6(32'hbc0756bc),
	.w7(32'h3b16323c),
	.w8(32'h3a02603d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb050084),
	.w1(32'hba9b56eb),
	.w2(32'hbb2080de),
	.w3(32'hb9f6e8be),
	.w4(32'h3b4ff628),
	.w5(32'h3ad4ccf7),
	.w6(32'h39e0a4d4),
	.w7(32'h3b1d93d6),
	.w8(32'h3b7de671),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a779798),
	.w1(32'h3b89a8f1),
	.w2(32'hba2eaa74),
	.w3(32'hbb4186b1),
	.w4(32'hbb408184),
	.w5(32'hbb358bd5),
	.w6(32'h39d9800e),
	.w7(32'hbab5e444),
	.w8(32'hbc398085),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba07028),
	.w1(32'h39135264),
	.w2(32'hbadb8177),
	.w3(32'hba923c75),
	.w4(32'hbba1172a),
	.w5(32'h3bb0a467),
	.w6(32'hbb4441d3),
	.w7(32'hbc1b3928),
	.w8(32'h3ba9a15c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78eb75),
	.w1(32'h3bacfba7),
	.w2(32'hbab632f3),
	.w3(32'h3c2c726c),
	.w4(32'h3a8602cc),
	.w5(32'h3a8753d0),
	.w6(32'h3c31d88d),
	.w7(32'hbb61550a),
	.w8(32'h3bfd9e17),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2b1ea),
	.w1(32'hbbad8cad),
	.w2(32'h3beefc0c),
	.w3(32'h3b88522a),
	.w4(32'hbaefe851),
	.w5(32'hb9ad482a),
	.w6(32'hbc029a32),
	.w7(32'h3b27d855),
	.w8(32'hbb67af09),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03f715),
	.w1(32'hba618962),
	.w2(32'h3b7a9667),
	.w3(32'hbb9d06a9),
	.w4(32'hbb183d3f),
	.w5(32'h3b9be016),
	.w6(32'hbb867780),
	.w7(32'h39c843e6),
	.w8(32'h3bc317d7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb586f),
	.w1(32'h3aacd54f),
	.w2(32'h3bf69836),
	.w3(32'hbbeb65a3),
	.w4(32'hbbf356bd),
	.w5(32'hbb92765b),
	.w6(32'hba4735a6),
	.w7(32'hbb442d5c),
	.w8(32'hbb092f37),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa19422),
	.w1(32'hbb9b1777),
	.w2(32'hbb70a042),
	.w3(32'h3903e6d3),
	.w4(32'hbbf1dbdb),
	.w5(32'h3b359c36),
	.w6(32'h3a8be7f4),
	.w7(32'hb8b8ddd3),
	.w8(32'hbc0ac8e6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25051b),
	.w1(32'hbc029d9b),
	.w2(32'hbb27aee3),
	.w3(32'h3c5bd116),
	.w4(32'hba239a5c),
	.w5(32'h3b8cae74),
	.w6(32'hbbfa02fd),
	.w7(32'hbb0fa67f),
	.w8(32'h3c1df812),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b476),
	.w1(32'hba6cb8ec),
	.w2(32'h3ad2522f),
	.w3(32'h3bb3ef21),
	.w4(32'h37e30ba1),
	.w5(32'h3bec78b1),
	.w6(32'hbb2c5d6e),
	.w7(32'hbb7af545),
	.w8(32'h3b49b17f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae560fa),
	.w1(32'h3b701dfd),
	.w2(32'h3bbd0b88),
	.w3(32'h3b94721c),
	.w4(32'h3abe182a),
	.w5(32'h3a26c6ed),
	.w6(32'hbb833b4d),
	.w7(32'h3afaa9d7),
	.w8(32'h3b171391),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6903d),
	.w1(32'h3a960e01),
	.w2(32'h3af9062b),
	.w3(32'h3bfae84e),
	.w4(32'h3b5d787b),
	.w5(32'h3acf8074),
	.w6(32'h3c4d091f),
	.w7(32'h3b54bf94),
	.w8(32'hbaff1e3c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb009129),
	.w1(32'hbb582ae7),
	.w2(32'hbb8df95e),
	.w3(32'h3a70b6b7),
	.w4(32'h3baa313d),
	.w5(32'h3c891429),
	.w6(32'hba8e36e9),
	.w7(32'hbb01c354),
	.w8(32'h3c31176d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e78c6),
	.w1(32'h3b583f80),
	.w2(32'hbb8337e3),
	.w3(32'h3c06f319),
	.w4(32'h3a82929f),
	.w5(32'hbb0fff61),
	.w6(32'hbc410f89),
	.w7(32'hbbcda454),
	.w8(32'hba955486),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6f0d6),
	.w1(32'h39f11698),
	.w2(32'hbac68638),
	.w3(32'hbb842dd0),
	.w4(32'hbac3935d),
	.w5(32'hbb4e8095),
	.w6(32'h3b9d7601),
	.w7(32'hbb212380),
	.w8(32'hbbcfe3e4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0163e1),
	.w1(32'h3ac34cfd),
	.w2(32'h3c0c1e6d),
	.w3(32'hbb4281f2),
	.w4(32'hb99b371a),
	.w5(32'hba7b456f),
	.w6(32'hbb5c9c42),
	.w7(32'h3afb4a65),
	.w8(32'hb906ee5e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba023955),
	.w1(32'h3a9f60e0),
	.w2(32'h3add726e),
	.w3(32'hb90585c8),
	.w4(32'h3a2a9972),
	.w5(32'h3b35db15),
	.w6(32'h3b5c7702),
	.w7(32'h3a083398),
	.w8(32'h3943938a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98ed93),
	.w1(32'h3b2281a7),
	.w2(32'h3abb1443),
	.w3(32'hbba031a5),
	.w4(32'hbb773bd6),
	.w5(32'hbb8ff2c2),
	.w6(32'h3b16965d),
	.w7(32'h3b3d1acb),
	.w8(32'hbad0a673),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20a78d),
	.w1(32'hbbb29059),
	.w2(32'hbc1c3f82),
	.w3(32'hbb9d8eb9),
	.w4(32'hbb99a1aa),
	.w5(32'hbbfb886e),
	.w6(32'hbbb601dc),
	.w7(32'hbbe8a439),
	.w8(32'hbbb9286c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90dcc0),
	.w1(32'h39ac1f12),
	.w2(32'hbb33fa42),
	.w3(32'hbb970f0f),
	.w4(32'hbb080eff),
	.w5(32'h3b0484e0),
	.w6(32'h3b1a5052),
	.w7(32'hbb014aff),
	.w8(32'h3b94d18b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe6caf),
	.w1(32'hbbf663c7),
	.w2(32'hbb3a8caa),
	.w3(32'h3bd50d9b),
	.w4(32'hba81aaaf),
	.w5(32'hbbe856ed),
	.w6(32'h3ba70ef2),
	.w7(32'h3b892cd4),
	.w8(32'h3c06e2d9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf16f6),
	.w1(32'h3b6d9c89),
	.w2(32'h3bc744c8),
	.w3(32'h3bb4a9fe),
	.w4(32'h3c0b8189),
	.w5(32'h3b7ce77a),
	.w6(32'h3bd49590),
	.w7(32'h3a1e3eb5),
	.w8(32'hba8150a6),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04ad71),
	.w1(32'hbbcd7f34),
	.w2(32'hbbfe1320),
	.w3(32'h3a933882),
	.w4(32'hbb8426c5),
	.w5(32'hbb03302c),
	.w6(32'hbbac6404),
	.w7(32'hbbf67189),
	.w8(32'hbb0fb5be),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4170f5),
	.w1(32'hbb8f7677),
	.w2(32'hbaaad245),
	.w3(32'hb9de168b),
	.w4(32'hbb1932b4),
	.w5(32'hbb863806),
	.w6(32'hbb012f50),
	.w7(32'hbacbaec5),
	.w8(32'hbc028552),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2acae6),
	.w1(32'hbb41e5de),
	.w2(32'h3ba83bf4),
	.w3(32'hb931c96c),
	.w4(32'hbb2b038a),
	.w5(32'h3b3292ba),
	.w6(32'hb992bcaa),
	.w7(32'hba922cba),
	.w8(32'h3a4b2082),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa71645),
	.w1(32'h3994cb8e),
	.w2(32'h3b5c50f3),
	.w3(32'hbb666a9c),
	.w4(32'hbb6ddef0),
	.w5(32'h3baed5ad),
	.w6(32'hb9b285f5),
	.w7(32'h3acca9ed),
	.w8(32'h3a3f73ad),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81237b),
	.w1(32'hbb9e511c),
	.w2(32'hbaa55184),
	.w3(32'hbbaab3a2),
	.w4(32'hbbe299a9),
	.w5(32'hbb773e26),
	.w6(32'hbc843065),
	.w7(32'hb9bdb7b0),
	.w8(32'h3b23bfea),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19b15e),
	.w1(32'hbbad7d36),
	.w2(32'hbbff2ab0),
	.w3(32'hb9fb1374),
	.w4(32'hbb37c1b0),
	.w5(32'hbb39864b),
	.w6(32'h3b620073),
	.w7(32'hbbaa93ac),
	.w8(32'hbbd2fb0c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4cc05),
	.w1(32'h3a1c8be5),
	.w2(32'h3b3dd480),
	.w3(32'hbb4549bb),
	.w4(32'hbacb9d20),
	.w5(32'hbb442c0c),
	.w6(32'h38a6cde6),
	.w7(32'h3ba9703f),
	.w8(32'hbb82344f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d8b2f),
	.w1(32'h3ab571f9),
	.w2(32'hbaadb545),
	.w3(32'h3b431b32),
	.w4(32'h3a98a36b),
	.w5(32'hbb0be881),
	.w6(32'hbba00f13),
	.w7(32'hbbb18c18),
	.w8(32'hba8454fd),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56fc0b),
	.w1(32'h3b023dc0),
	.w2(32'hba9a3c30),
	.w3(32'hb91bc4a8),
	.w4(32'h3996fbc4),
	.w5(32'hbaffeb03),
	.w6(32'h3aaecb5d),
	.w7(32'hbb80fc5e),
	.w8(32'hbbdbae7e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b527b),
	.w1(32'h3ba3fcc0),
	.w2(32'h3b1a320f),
	.w3(32'hbb3bd9db),
	.w4(32'hba333458),
	.w5(32'h3c61df2b),
	.w6(32'hbbca910d),
	.w7(32'hbb3c4c00),
	.w8(32'hbae78426),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc71180),
	.w1(32'hbbe0fe11),
	.w2(32'h3b7d3286),
	.w3(32'h3cb00c11),
	.w4(32'h3ba8e41a),
	.w5(32'hbb9229fe),
	.w6(32'h3c19a324),
	.w7(32'h3c96198d),
	.w8(32'hb8ca6155),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f8c80),
	.w1(32'h3a4427bc),
	.w2(32'hb9aef9e9),
	.w3(32'hba85c035),
	.w4(32'hba6b1bf5),
	.w5(32'hba1a32ef),
	.w6(32'h3baf1258),
	.w7(32'hbb88640d),
	.w8(32'hbb67950f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd4839),
	.w1(32'hbb8f7032),
	.w2(32'hbb2dcfd4),
	.w3(32'h3ad7be2b),
	.w4(32'hba1e4e98),
	.w5(32'hbad19c8b),
	.w6(32'hbb6ef909),
	.w7(32'h3b822fac),
	.w8(32'hba5984f9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule