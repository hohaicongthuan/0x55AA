module layer_10_featuremap_240(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fce2a2),
	.w1(32'h3838019b),
	.w2(32'h38a523d3),
	.w3(32'h390ad943),
	.w4(32'h381043a9),
	.w5(32'h38147602),
	.w6(32'h3911f442),
	.w7(32'h3802fd8c),
	.w8(32'h38a2b5f1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5f4f),
	.w1(32'hbab2f2c8),
	.w2(32'hbb4ba817),
	.w3(32'hbbc54399),
	.w4(32'h3aa8c15e),
	.w5(32'h39463308),
	.w6(32'hbbccc8cd),
	.w7(32'h39a7b00e),
	.w8(32'hbaf2cf78),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c25cfd),
	.w1(32'hb7af0cb5),
	.w2(32'h37ec7052),
	.w3(32'h37fc7034),
	.w4(32'h378b33d9),
	.w5(32'h380fcff7),
	.w6(32'h388e2790),
	.w7(32'h3823e001),
	.w8(32'h385ddb19),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f82e6),
	.w1(32'h3a075f22),
	.w2(32'h3a7beaf4),
	.w3(32'h398a9ce2),
	.w4(32'hb9e2ff14),
	.w5(32'h3910e548),
	.w6(32'h3a1f39f8),
	.w7(32'h39be0ad5),
	.w8(32'h39489a35),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78e86d2),
	.w1(32'hb9c35030),
	.w2(32'hba563437),
	.w3(32'h39a3acdc),
	.w4(32'hb88299e9),
	.w5(32'hb9e78b88),
	.w6(32'h39c1b35a),
	.w7(32'h39867059),
	.w8(32'h380ee3a4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c0a14),
	.w1(32'h3812508c),
	.w2(32'h3889c6bf),
	.w3(32'h390fa16e),
	.w4(32'h3815bd4e),
	.w5(32'h38a4689c),
	.w6(32'h391240ba),
	.w7(32'h37e0570e),
	.w8(32'h38da950b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b5329),
	.w1(32'hbb893c58),
	.w2(32'hbc0e540e),
	.w3(32'h3a8d4034),
	.w4(32'hbbb30b63),
	.w5(32'hbc26080c),
	.w6(32'h3b0c3f68),
	.w7(32'hbb6c5c62),
	.w8(32'hbc14ac54),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c537a),
	.w1(32'hbc0e30e0),
	.w2(32'hbc17ee16),
	.w3(32'hbc281107),
	.w4(32'hbc11a091),
	.w5(32'hbba80d4f),
	.w6(32'hbba03610),
	.w7(32'hbb885d9e),
	.w8(32'hbb4b1c38),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29f25b),
	.w1(32'h3a2e358d),
	.w2(32'hba381122),
	.w3(32'hb9af33ba),
	.w4(32'h3a2b151d),
	.w5(32'hba395e7f),
	.w6(32'hba8c4e9c),
	.w7(32'hb922d826),
	.w8(32'hba9a4d00),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51cbc0),
	.w1(32'hbaaa5689),
	.w2(32'hbc9e207d),
	.w3(32'hbbba27de),
	.w4(32'h3afd3a44),
	.w5(32'hbc57ab3b),
	.w6(32'hbc0e525a),
	.w7(32'h3b49a45d),
	.w8(32'hbc1e5f97),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf711ff),
	.w1(32'hbaa04288),
	.w2(32'hbb04c584),
	.w3(32'hbacc6be1),
	.w4(32'hba23d759),
	.w5(32'hba8cdb3d),
	.w6(32'hbad439b2),
	.w7(32'hbaa5bc64),
	.w8(32'hbad9b843),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafda52a),
	.w1(32'h3b739660),
	.w2(32'hbbd0f4f3),
	.w3(32'hbb0cfcab),
	.w4(32'h3b7a3569),
	.w5(32'hbbb25faf),
	.w6(32'hbb36c278),
	.w7(32'h3b69fde6),
	.w8(32'hbc50d3a8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b76d9),
	.w1(32'hbb2a50de),
	.w2(32'hbcab49d6),
	.w3(32'hb9907ae0),
	.w4(32'h3ab1c0e1),
	.w5(32'hbc77539b),
	.w6(32'h3a01aad7),
	.w7(32'h3b97e646),
	.w8(32'hbc1d83ff),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e5e26),
	.w1(32'hbbc1fa38),
	.w2(32'hbbb0bc3c),
	.w3(32'hbba164b9),
	.w4(32'hbb22c8ad),
	.w5(32'hbaeb9e2c),
	.w6(32'hbbb6fd9c),
	.w7(32'hbad9afa0),
	.w8(32'hbad14ca7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4901e6),
	.w1(32'h3b40e962),
	.w2(32'hbb858321),
	.w3(32'hba89d2cc),
	.w4(32'h3c050fe6),
	.w5(32'h3b1848dc),
	.w6(32'hbbd92646),
	.w7(32'h3b81b263),
	.w8(32'hbad7f4a6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ddfa8),
	.w1(32'hbb475f5a),
	.w2(32'hbc64242f),
	.w3(32'hbb720f3e),
	.w4(32'h3b48d24b),
	.w5(32'hbb984338),
	.w6(32'hbbcddc54),
	.w7(32'hba8b63f3),
	.w8(32'hbbbe18d3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d8ec1),
	.w1(32'h39d580d1),
	.w2(32'h3988d1ce),
	.w3(32'h3a1d2a2c),
	.w4(32'h3a3fcbe7),
	.w5(32'h39d0d56c),
	.w6(32'h3a159c01),
	.w7(32'h3a842f07),
	.w8(32'h3a1f3c3d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a76df),
	.w1(32'hbbac5108),
	.w2(32'hbc7d8bd1),
	.w3(32'hbbf91790),
	.w4(32'hbb8d43ff),
	.w5(32'hbc5f3ab9),
	.w6(32'hbbb29d9e),
	.w7(32'hbb76da98),
	.w8(32'hbc559efe),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba35356),
	.w1(32'hbb2c849c),
	.w2(32'hbc171939),
	.w3(32'hbab7653a),
	.w4(32'hbad4b0b2),
	.w5(32'hbbfe37fe),
	.w6(32'hbaad5bb7),
	.w7(32'hba726a0e),
	.w8(32'hbbdf01b3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f061cd),
	.w1(32'h393d8e43),
	.w2(32'h393a093d),
	.w3(32'h394a6b6b),
	.w4(32'h3984988e),
	.w5(32'h395df946),
	.w6(32'h396dc22b),
	.w7(32'h399f4d9b),
	.w8(32'h390af032),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7f1ad),
	.w1(32'h3925e590),
	.w2(32'h3981faf8),
	.w3(32'h399bf91b),
	.w4(32'h38add71d),
	.w5(32'h393608fb),
	.w6(32'h39e38898),
	.w7(32'h39527265),
	.w8(32'h39b51800),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14bee2),
	.w1(32'h3b7ab7e7),
	.w2(32'hbb217319),
	.w3(32'h3b5f7fe8),
	.w4(32'h3bc47414),
	.w5(32'hb9cdda64),
	.w6(32'h3a864d5a),
	.w7(32'h3b8aba7a),
	.w8(32'hba96fb52),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf5c510),
	.w1(32'hbc12a008),
	.w2(32'hbc9df6e3),
	.w3(32'hbccf251e),
	.w4(32'hbac04bbb),
	.w5(32'hbcaa5397),
	.w6(32'hbcec6eab),
	.w7(32'hbc2ded58),
	.w8(32'hbcf0e027),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc427714),
	.w1(32'h390cde2d),
	.w2(32'hbc8ea7c6),
	.w3(32'hbb2f6ae4),
	.w4(32'h3bf64688),
	.w5(32'hbc16e6b5),
	.w6(32'hbc0a7531),
	.w7(32'h3bc15d8d),
	.w8(32'hbc0e82a4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b3445),
	.w1(32'h3a95636e),
	.w2(32'hbc3bdb2e),
	.w3(32'hbc382fe9),
	.w4(32'h3c211366),
	.w5(32'hbb1ad465),
	.w6(32'hbc88a68e),
	.w7(32'h3be5e5af),
	.w8(32'hbba4a964),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941e73f),
	.w1(32'h3881089e),
	.w2(32'hb9ba1dc8),
	.w3(32'hb86988fa),
	.w4(32'hb8a60744),
	.w5(32'hba49aa4f),
	.w6(32'hb88e1611),
	.w7(32'h39b9c577),
	.w8(32'h39dff4e7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a188a01),
	.w1(32'h39865a31),
	.w2(32'h39ff8808),
	.w3(32'h39f2180a),
	.w4(32'h3903671e),
	.w5(32'h39cdc1d2),
	.w6(32'h3a189dec),
	.w7(32'h3993021f),
	.w8(32'h3a037dcd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba262fe),
	.w1(32'h3b70e31f),
	.w2(32'hba5c8aed),
	.w3(32'h3abd9ebc),
	.w4(32'h3bbbf232),
	.w5(32'h3be7ec8a),
	.w6(32'h3a372efc),
	.w7(32'h3b85aa7f),
	.w8(32'h3b9b4a74),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82dc71),
	.w1(32'hb99cf847),
	.w2(32'hbb8abf93),
	.w3(32'hbb16fa2f),
	.w4(32'h3ad94242),
	.w5(32'hbab69057),
	.w6(32'hbbadd88d),
	.w7(32'hb8bd97f7),
	.w8(32'hbb46ccf2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb878ebd),
	.w1(32'h3bc832e7),
	.w2(32'hbb8e138c),
	.w3(32'hbb03a4ec),
	.w4(32'h3be49a4f),
	.w5(32'hb841d15c),
	.w6(32'hbbb07e84),
	.w7(32'h3bee688d),
	.w8(32'h3aeef0f3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e2684),
	.w1(32'h392ae678),
	.w2(32'h392b00ab),
	.w3(32'h39523ed4),
	.w4(32'h3923643c),
	.w5(32'h38c128c6),
	.w6(32'h38dd6558),
	.w7(32'h38bbd616),
	.w8(32'h391dc2c9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e2c945),
	.w1(32'hb7426cc9),
	.w2(32'hb860b18f),
	.w3(32'h39295772),
	.w4(32'h3981f4a8),
	.w5(32'h393cfe06),
	.w6(32'h399845e9),
	.w7(32'h39af6d32),
	.w8(32'h393b72d6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb79d),
	.w1(32'hb80a66e1),
	.w2(32'hbc0a5bd2),
	.w3(32'h3abe83db),
	.w4(32'h3b75d7e6),
	.w5(32'hbb99dbc3),
	.w6(32'hbac313da),
	.w7(32'h3b2e8c69),
	.w8(32'hbb88b652),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8262b),
	.w1(32'h39aece14),
	.w2(32'hbb0e6437),
	.w3(32'hbb889804),
	.w4(32'h3afacf90),
	.w5(32'h3884c4c5),
	.w6(32'hbbaeda22),
	.w7(32'h39fd5975),
	.w8(32'hba9675e8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38db9ec3),
	.w1(32'h3999b052),
	.w2(32'hba1bb59a),
	.w3(32'h3a1fbde0),
	.w4(32'hb802949f),
	.w5(32'hb98c8e00),
	.w6(32'h395d5e3d),
	.w7(32'hb9bdbb3c),
	.w8(32'hbabf05bc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac412d8),
	.w1(32'hbb30b4cc),
	.w2(32'hbbaa4ba6),
	.w3(32'h3a8ca24e),
	.w4(32'hbabf5f86),
	.w5(32'hbb809a7f),
	.w6(32'h3aa1e78a),
	.w7(32'hba746b2b),
	.w8(32'hbb8b76d6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d6404),
	.w1(32'hbaf9b6f6),
	.w2(32'hbc75d35f),
	.w3(32'hbb88006b),
	.w4(32'h3b909ea2),
	.w5(32'hbbf2ee9d),
	.w6(32'h3abb1ac7),
	.w7(32'h3bfeec4f),
	.w8(32'hbc4adc5b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf319ae),
	.w1(32'h3b556490),
	.w2(32'h3a22a89b),
	.w3(32'hbca84e3a),
	.w4(32'h3c1c470b),
	.w5(32'h3c0034f6),
	.w6(32'hbd0fe9f2),
	.w7(32'hba418ba3),
	.w8(32'hbbdb5640),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc938ecf),
	.w1(32'h3bd85b98),
	.w2(32'hbb97e7f3),
	.w3(32'hbc8de8fa),
	.w4(32'h3c172277),
	.w5(32'hbad01ac3),
	.w6(32'hbcf1495e),
	.w7(32'hbb13c855),
	.w8(32'hbc68c9d0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba9778),
	.w1(32'h3a7f3828),
	.w2(32'h3b1b4c5b),
	.w3(32'hbb72409a),
	.w4(32'h3b24d905),
	.w5(32'h3b86462a),
	.w6(32'hbbb95557),
	.w7(32'h3a797dc4),
	.w8(32'h3a8b2dba),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b0d70),
	.w1(32'h37168a0c),
	.w2(32'h398f413f),
	.w3(32'h397af83b),
	.w4(32'hb8b5ed6a),
	.w5(32'h395bc9dc),
	.w6(32'h39f535d8),
	.w7(32'h3907b85c),
	.w8(32'h39cc5c29),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981eff6),
	.w1(32'hb7eaf848),
	.w2(32'h3a09acc7),
	.w3(32'h39ff844c),
	.w4(32'hb90a20b6),
	.w5(32'h39a4d1e7),
	.w6(32'h3a2179d1),
	.w7(32'h39389682),
	.w8(32'h39fb63f2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2618b0),
	.w1(32'hba014abf),
	.w2(32'hbb06418d),
	.w3(32'hbc100b27),
	.w4(32'h3a1f3ee6),
	.w5(32'hbb0f84c3),
	.w6(32'hbbf76560),
	.w7(32'hb986d4bc),
	.w8(32'hbb636af0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7725b9),
	.w1(32'hbb5f8654),
	.w2(32'hbc923877),
	.w3(32'hbc23fad6),
	.w4(32'hbb4393ab),
	.w5(32'hbc398a1f),
	.w6(32'hbc5fae89),
	.w7(32'hbbcf3a61),
	.w8(32'hbc578346),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc328602),
	.w1(32'h3afe41dd),
	.w2(32'hbc61115a),
	.w3(32'hbb23d511),
	.w4(32'h3c2c870f),
	.w5(32'hbb9aab17),
	.w6(32'hbc084ea9),
	.w7(32'h3c04b247),
	.w8(32'hbbab4db0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc706bbb),
	.w1(32'h3a36a5a4),
	.w2(32'hbc968d54),
	.w3(32'hbb81ce58),
	.w4(32'h3c141c81),
	.w5(32'hbc1aba06),
	.w6(32'hbc285a44),
	.w7(32'h3c106ee7),
	.w8(32'hbbec3773),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b426c),
	.w1(32'h3a9f1d7d),
	.w2(32'hbbd1b6b0),
	.w3(32'hbc21940e),
	.w4(32'h3b904b0a),
	.w5(32'hbb37c6f9),
	.w6(32'hbc471eff),
	.w7(32'h3aff03d6),
	.w8(32'hbbec6b68),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12487e),
	.w1(32'hbc142bfc),
	.w2(32'hbc80cf7e),
	.w3(32'hbbfe4abe),
	.w4(32'hbc351e9b),
	.w5(32'hbc878834),
	.w6(32'hbb25a827),
	.w7(32'hbb923f52),
	.w8(32'hbc4b66bb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919c841),
	.w1(32'h3896025b),
	.w2(32'h38a84ff0),
	.w3(32'hb94f03f9),
	.w4(32'hb98df0ba),
	.w5(32'h38185ba6),
	.w6(32'hb83d1dae),
	.w7(32'hb86ceca1),
	.w8(32'h396d3ecb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a5e6e1),
	.w1(32'h3a803de2),
	.w2(32'h3b109007),
	.w3(32'hb9cfc09c),
	.w4(32'hb9a9f3e4),
	.w5(32'h3a7fe2fd),
	.w6(32'hba8b3f0f),
	.w7(32'hba5b7c70),
	.w8(32'hb980cc20),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999589b),
	.w1(32'hb9be71c9),
	.w2(32'hb99ce987),
	.w3(32'hb689df1a),
	.w4(32'hb9b01b07),
	.w5(32'hb93a6f3b),
	.w6(32'h396d0d21),
	.w7(32'hb89e824a),
	.w8(32'hb982fa81),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaaf46),
	.w1(32'hba91c9da),
	.w2(32'hbc112fc2),
	.w3(32'hba252579),
	.w4(32'h3b958320),
	.w5(32'hbb7943bb),
	.w6(32'hba50596b),
	.w7(32'h3bb6f47b),
	.w8(32'hb98acd05),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2926aa),
	.w1(32'hba855079),
	.w2(32'hbb80f750),
	.w3(32'hbabb74f3),
	.w4(32'h377e1345),
	.w5(32'hbb4d5788),
	.w6(32'hbac2aaa5),
	.w7(32'h3994707e),
	.w8(32'hbb191e50),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23e791),
	.w1(32'hbb936518),
	.w2(32'hbc8d1616),
	.w3(32'hbb8e95ec),
	.w4(32'hbb2af87e),
	.w5(32'hbc524821),
	.w6(32'hbbac9061),
	.w7(32'h390d0f23),
	.w8(32'hbc1cf2cd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadafbfb),
	.w1(32'h39f8cd69),
	.w2(32'hba50b0cb),
	.w3(32'hbb05f3f5),
	.w4(32'hba2cd67a),
	.w5(32'hbacfea52),
	.w6(32'hbb353044),
	.w7(32'hba8b8293),
	.w8(32'hbb0a9bc5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d7fe3),
	.w1(32'hb930ac78),
	.w2(32'hb9bd0274),
	.w3(32'h3732dbcd),
	.w4(32'h38bc58b7),
	.w5(32'h38b4a614),
	.w6(32'h38ea6c4a),
	.w7(32'h39cc7621),
	.w8(32'h39b6bf1b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39029648),
	.w1(32'h38c32d7c),
	.w2(32'h3872a34e),
	.w3(32'h3917a890),
	.w4(32'h38b83892),
	.w5(32'h3893c3db),
	.w6(32'h391d6976),
	.w7(32'h38d5fe90),
	.w8(32'h38a1f7b5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39942f7e),
	.w1(32'h39c9b353),
	.w2(32'h39373e4f),
	.w3(32'h38994e55),
	.w4(32'h39aa8176),
	.w5(32'h39d8413b),
	.w6(32'hb86061ba),
	.w7(32'h396e8d7d),
	.w8(32'h3931d06a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2181ee),
	.w1(32'h3ade0ae5),
	.w2(32'hba1e5c81),
	.w3(32'h3988613d),
	.w4(32'h3b33a9b9),
	.w5(32'h3a1ca690),
	.w6(32'hbae8981b),
	.w7(32'h3a28cde3),
	.w8(32'hba82ee79),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8585e3),
	.w1(32'hb93ff7ff),
	.w2(32'hba49a94f),
	.w3(32'h38d1685e),
	.w4(32'h39873f17),
	.w5(32'hba30e500),
	.w6(32'hb9adf71c),
	.w7(32'hb99ffd37),
	.w8(32'hba8073a9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93815c),
	.w1(32'hba92f52e),
	.w2(32'hbbe45484),
	.w3(32'hbb16060c),
	.w4(32'hba1247cd),
	.w5(32'hbba3adfe),
	.w6(32'hba4695b9),
	.w7(32'h3a06298f),
	.w8(32'hbb9f9c53),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe29af3),
	.w1(32'hbb2cb9e4),
	.w2(32'hbb6f97b3),
	.w3(32'hbbacbe9d),
	.w4(32'hbb2d34f1),
	.w5(32'hbb935901),
	.w6(32'hbb879fec),
	.w7(32'hbb30ae6d),
	.w8(32'hbb9c8252),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395949a7),
	.w1(32'h37f75ec6),
	.w2(32'h391c6e45),
	.w3(32'h3928b0ba),
	.w4(32'hb6b71871),
	.w5(32'h38955c7a),
	.w6(32'h3937614b),
	.w7(32'h379edaa7),
	.w8(32'h3957d08e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a1f8c),
	.w1(32'h3859eb8b),
	.w2(32'h3925da18),
	.w3(32'h38f86fd9),
	.w4(32'hb7e2b2d4),
	.w5(32'h388622fe),
	.w6(32'h39528e64),
	.w7(32'h38895ce2),
	.w8(32'h392e56d7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3827191c),
	.w1(32'h388f1428),
	.w2(32'hb835c0c9),
	.w3(32'h392fba4a),
	.w4(32'h3946db5a),
	.w5(32'h392d0488),
	.w6(32'h3976a487),
	.w7(32'h398d7a5d),
	.w8(32'h3982be24),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0e263),
	.w1(32'h38c00740),
	.w2(32'h396d57fc),
	.w3(32'h39993d70),
	.w4(32'h387daa06),
	.w5(32'h3930a259),
	.w6(32'h39c55bc9),
	.w7(32'h3914db6b),
	.w8(32'h3988b250),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4ea76),
	.w1(32'hbb38b43e),
	.w2(32'hbbff1fab),
	.w3(32'hbbc713af),
	.w4(32'hbbc4d712),
	.w5(32'hbbab85ec),
	.w6(32'hbb7284fc),
	.w7(32'hbb9f35f8),
	.w8(32'hbbc6441c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55bcc6),
	.w1(32'hbadb9245),
	.w2(32'hbc96be33),
	.w3(32'hbb89d3a1),
	.w4(32'h3b6b29f1),
	.w5(32'hbc918ca1),
	.w6(32'hbc15103a),
	.w7(32'h3b5688fd),
	.w8(32'hbc814bd3),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc517675),
	.w1(32'hb8c643fa),
	.w2(32'hbc5623cb),
	.w3(32'hbbfb875f),
	.w4(32'h3ba16f84),
	.w5(32'hbc029b77),
	.w6(32'hbc7abfdb),
	.w7(32'hbb26df94),
	.w8(32'hbc59d5f0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc575d8f),
	.w1(32'h3c38869e),
	.w2(32'hbc908480),
	.w3(32'hbb00ee8f),
	.w4(32'h3cf3f14e),
	.w5(32'h3c01a7b9),
	.w6(32'hbc8785d7),
	.w7(32'h3ca8ad7d),
	.w8(32'hbbd718c3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1eb0d),
	.w1(32'h386da473),
	.w2(32'h3984754f),
	.w3(32'h39a55619),
	.w4(32'hb81fed8d),
	.w5(32'h390a5b05),
	.w6(32'h39e6f6f5),
	.w7(32'h38f21dd4),
	.w8(32'h399b12e2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e1702),
	.w1(32'h39341935),
	.w2(32'h3a074359),
	.w3(32'h39ea3301),
	.w4(32'h36a4eac1),
	.w5(32'h39ae88bb),
	.w6(32'h3a34265f),
	.w7(32'h398db64b),
	.w8(32'h3a1c1a36),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff3177),
	.w1(32'hb7db9565),
	.w2(32'h39a9760e),
	.w3(32'h39f3e3d2),
	.w4(32'hb90b23d7),
	.w5(32'h398951ca),
	.w6(32'h3a3513b9),
	.w7(32'h38f91d71),
	.w8(32'h39f0062f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e6665),
	.w1(32'h3aa7984d),
	.w2(32'hba6efbe7),
	.w3(32'hb99844c3),
	.w4(32'hb8a5dc8d),
	.w5(32'hbaf7a275),
	.w6(32'hb9a91691),
	.w7(32'hba2afb66),
	.w8(32'hbaec8300),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39909d2e),
	.w1(32'hb7859bd8),
	.w2(32'h39787b61),
	.w3(32'h39b1df8c),
	.w4(32'hb894525d),
	.w5(32'h391f240e),
	.w6(32'h3a01a494),
	.w7(32'h390d2dee),
	.w8(32'h39b6b635),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8936ba),
	.w1(32'hbac25943),
	.w2(32'hbb7bb44d),
	.w3(32'hbae4511b),
	.w4(32'hbb3bbc01),
	.w5(32'hbb5950b7),
	.w6(32'h3aabed27),
	.w7(32'h39ab3ade),
	.w8(32'hbac7d259),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d0eb1),
	.w1(32'hbb49e9c7),
	.w2(32'hbc261cb4),
	.w3(32'hbb932519),
	.w4(32'h3a716e6e),
	.w5(32'hba572531),
	.w6(32'hbba9e5e7),
	.w7(32'hba8717f9),
	.w8(32'hbc0379d2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23abb3),
	.w1(32'hbb2205a1),
	.w2(32'hbc27a656),
	.w3(32'hbb4c3825),
	.w4(32'h3bb9e8df),
	.w5(32'hbb06bd45),
	.w6(32'hbb57227b),
	.w7(32'h3bdf912a),
	.w8(32'hbae817c3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1de12),
	.w1(32'hbb2a2294),
	.w2(32'hbc208e64),
	.w3(32'hbb909f50),
	.w4(32'hb8cbf0d1),
	.w5(32'hbbceaa8a),
	.w6(32'hbbdab407),
	.w7(32'hbacc30dc),
	.w8(32'hbbe00541),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982ed57),
	.w1(32'h3a0f3c68),
	.w2(32'hbbbba950),
	.w3(32'hb965117d),
	.w4(32'h39f8cdd1),
	.w5(32'hbb54f442),
	.w6(32'h3a347a88),
	.w7(32'h3b746a2d),
	.w8(32'hbb290500),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb576ebb),
	.w1(32'h390fbdf3),
	.w2(32'hbbd3f24a),
	.w3(32'hbaa25f39),
	.w4(32'h3b0ab997),
	.w5(32'hbb43adae),
	.w6(32'hbb2aa831),
	.w7(32'h3af1ba25),
	.w8(32'hbae6e4f8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2b344),
	.w1(32'hbabd65a9),
	.w2(32'hbc145618),
	.w3(32'hba1ec28b),
	.w4(32'hbb298180),
	.w5(32'hbc20915a),
	.w6(32'hb989f2b4),
	.w7(32'h3938d255),
	.w8(32'hbbd4adfc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373b631f),
	.w1(32'h37c1ac3e),
	.w2(32'h388a374d),
	.w3(32'h380ff28d),
	.w4(32'h35b3f55b),
	.w5(32'h3835f0bf),
	.w6(32'h388b032e),
	.w7(32'h37c92da3),
	.w8(32'h38aeca13),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8308c),
	.w1(32'h38665038),
	.w2(32'h38c40e0d),
	.w3(32'h38b77286),
	.w4(32'h38481e8b),
	.w5(32'h38b5d7b7),
	.w6(32'h389e3ce4),
	.w7(32'h37b2db96),
	.w8(32'h38b54e4b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b04f5),
	.w1(32'h39025e1c),
	.w2(32'h3933d3fc),
	.w3(32'hb7961605),
	.w4(32'h3844c44d),
	.w5(32'h38d67dda),
	.w6(32'h3895d942),
	.w7(32'h390f31bb),
	.w8(32'h38ac2e34),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5b762),
	.w1(32'h3a53ce10),
	.w2(32'h3a49b72f),
	.w3(32'h39b8f258),
	.w4(32'h3a3f07de),
	.w5(32'h3a4e1695),
	.w6(32'h391bc4c9),
	.w7(32'h3a41cc0d),
	.w8(32'h3a340aa9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ce201),
	.w1(32'hba657f48),
	.w2(32'h39b26968),
	.w3(32'hbc4e7800),
	.w4(32'h3a99ca48),
	.w5(32'h3b941aee),
	.w6(32'hbc60d210),
	.w7(32'h3ad727b8),
	.w8(32'h3a68dacc),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a43d6),
	.w1(32'h3b03f4c4),
	.w2(32'hb95d07be),
	.w3(32'h3b056015),
	.w4(32'h3b6ee903),
	.w5(32'h3a31bef7),
	.w6(32'hb9bcfe5d),
	.w7(32'h3ade0f74),
	.w8(32'hba13bcd2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ffeff),
	.w1(32'hbb5efc38),
	.w2(32'hbc2a4901),
	.w3(32'hbb8ce1b7),
	.w4(32'h396b8040),
	.w5(32'hbbfd381c),
	.w6(32'hbbbb429b),
	.w7(32'h3a96b8ed),
	.w8(32'hbbc04609),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72fd93),
	.w1(32'hbbc0270f),
	.w2(32'hbc05cc47),
	.w3(32'hbca73d74),
	.w4(32'hbbdca7f1),
	.w5(32'hbc1ab6db),
	.w6(32'hbc99cef6),
	.w7(32'hbc145929),
	.w8(32'hbc2bcc69),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae493c),
	.w1(32'h3b36b93e),
	.w2(32'hbb1a8f65),
	.w3(32'hbba3eb93),
	.w4(32'h3b7c59d4),
	.w5(32'h3ae3653b),
	.w6(32'hbc233168),
	.w7(32'h3aadb3c9),
	.w8(32'hbb6fd46c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f386a),
	.w1(32'hbbcc2d71),
	.w2(32'hbc3c6461),
	.w3(32'hbbf90a0a),
	.w4(32'hbaabfe5b),
	.w5(32'hbbca7cb7),
	.w6(32'hbbd04286),
	.w7(32'hbb89caa6),
	.w8(32'hbc4ad77d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80cc3d),
	.w1(32'h3bcec438),
	.w2(32'hba9966e3),
	.w3(32'h3b02577c),
	.w4(32'h3c0a2a1f),
	.w5(32'h3abef05e),
	.w6(32'h39c56025),
	.w7(32'h3c1bacc7),
	.w8(32'h3b5887f2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc901dca),
	.w1(32'hbb46fb50),
	.w2(32'hbc059394),
	.w3(32'hbc6e3057),
	.w4(32'hbaab938a),
	.w5(32'hbb3a8276),
	.w6(32'hbc933461),
	.w7(32'hbb6558d2),
	.w8(32'hbbc92247),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21d20f),
	.w1(32'hbb14712f),
	.w2(32'hbb9ea460),
	.w3(32'hbbf288af),
	.w4(32'h3b1b2854),
	.w5(32'hb9c160aa),
	.w6(32'hbbdfdb0c),
	.w7(32'h3b280362),
	.w8(32'hbadf3885),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42a611),
	.w1(32'h3b55dbca),
	.w2(32'hba9f3830),
	.w3(32'hbbdc3e9b),
	.w4(32'h3beb9a8e),
	.w5(32'h3a9e1601),
	.w6(32'hbc311471),
	.w7(32'h3bc69adc),
	.w8(32'h3b2816e6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c712e8),
	.w1(32'hb93035a2),
	.w2(32'h39d3cc5f),
	.w3(32'hb680cd18),
	.w4(32'hb928555f),
	.w5(32'h39b3452f),
	.w6(32'h39e5cb10),
	.w7(32'h39a57535),
	.w8(32'h3a2f0f7d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc353f45),
	.w1(32'hbb092f12),
	.w2(32'hbc6c1177),
	.w3(32'hbbbc1345),
	.w4(32'h3b83d692),
	.w5(32'hbbea3454),
	.w6(32'hbc2dcbbd),
	.w7(32'hb986f500),
	.w8(32'hbc245e90),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e21d),
	.w1(32'hba98f5c3),
	.w2(32'hbbedd137),
	.w3(32'hbb9ecdc5),
	.w4(32'h3b486936),
	.w5(32'hba736b34),
	.w6(32'hbb86c685),
	.w7(32'hba207436),
	.w8(32'hbc191a53),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d35a0),
	.w1(32'hbb8b366a),
	.w2(32'hbc9d55ef),
	.w3(32'h389176ce),
	.w4(32'h3b612f4c),
	.w5(32'hbc23adfe),
	.w6(32'h3b4404c2),
	.w7(32'h3beaa786),
	.w8(32'hbc5e841a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd302946),
	.w1(32'hbb8971af),
	.w2(32'h3b9f3fc4),
	.w3(32'hbd08df77),
	.w4(32'h3ba1bbdd),
	.w5(32'h3b836997),
	.w6(32'hbd17cf18),
	.w7(32'hbbfbdd57),
	.w8(32'hbc4cbe8f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2293a8),
	.w1(32'h3ac3f287),
	.w2(32'hbc78e0fc),
	.w3(32'hbb3e08a3),
	.w4(32'h3be2a6a1),
	.w5(32'hbbfcee06),
	.w6(32'hbbe1af42),
	.w7(32'h3c0b6e3c),
	.w8(32'hbb75f2b8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc682028),
	.w1(32'hbba220f7),
	.w2(32'hbc1d2784),
	.w3(32'hbc0ace6d),
	.w4(32'hbb3ad29d),
	.w5(32'hbbf8abff),
	.w6(32'hbb0522b9),
	.w7(32'h3a809f19),
	.w8(32'hbc2f1ee6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2957e),
	.w1(32'h39b6ef34),
	.w2(32'h3a445f66),
	.w3(32'h3a5ea7ec),
	.w4(32'h3a409c9e),
	.w5(32'h3a00efb7),
	.w6(32'h3a827ab4),
	.w7(32'h3a9dc4e9),
	.w8(32'h3aa3db11),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc671942),
	.w1(32'hbc277923),
	.w2(32'hbc8e9a02),
	.w3(32'hbaec686b),
	.w4(32'hb99c23ed),
	.w5(32'hbc235602),
	.w6(32'h3a66b905),
	.w7(32'h3bc45827),
	.w8(32'hbbc2acf5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64f239),
	.w1(32'h3ae2e944),
	.w2(32'hbb780434),
	.w3(32'h3b63ffc0),
	.w4(32'h3b4f99a4),
	.w5(32'hbb4b7d2e),
	.w6(32'h3b2c22e6),
	.w7(32'h3bbce9ba),
	.w8(32'hbb63a4d1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc5a8d),
	.w1(32'h396598b3),
	.w2(32'hb980df71),
	.w3(32'h399c34e0),
	.w4(32'h3a4a5dab),
	.w5(32'hb956aac0),
	.w6(32'hb892bf04),
	.w7(32'h39eded75),
	.w8(32'hb85e2b08),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb291341),
	.w1(32'hbacaefa6),
	.w2(32'hbb16925b),
	.w3(32'hbac31f53),
	.w4(32'h390cb9fb),
	.w5(32'hba7082fc),
	.w6(32'hbb23989f),
	.w7(32'hba4df0ad),
	.w8(32'hbaadb92b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23ea96),
	.w1(32'hbb872ad6),
	.w2(32'hbc19f4f3),
	.w3(32'hbbb72b74),
	.w4(32'hbb471b32),
	.w5(32'hbbf5a59c),
	.w6(32'hbbe80469),
	.w7(32'hbb833b91),
	.w8(32'hbc061f7a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb865302),
	.w1(32'h3af50b6c),
	.w2(32'hbbd90e2e),
	.w3(32'h38cb2d5c),
	.w4(32'h3bd1940b),
	.w5(32'hba3eac95),
	.w6(32'hbb515d7c),
	.w7(32'h3bcdbc31),
	.w8(32'h3a617667),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc11b3),
	.w1(32'h3a126787),
	.w2(32'hb9a33220),
	.w3(32'hbbd3e670),
	.w4(32'h3b032f0f),
	.w5(32'h3a9bb674),
	.w6(32'hbc5137c0),
	.w7(32'hbb5e085d),
	.w8(32'hbb9206d8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf57208),
	.w1(32'hb9d61993),
	.w2(32'hbb8e89d8),
	.w3(32'hbba26235),
	.w4(32'h3b2b45d2),
	.w5(32'h3993b071),
	.w6(32'hbbbcfcdc),
	.w7(32'h39dd4270),
	.w8(32'hbaa4bb24),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb822934),
	.w1(32'h3b2dc05d),
	.w2(32'hbb285646),
	.w3(32'hbabb1655),
	.w4(32'h3b8f2c2f),
	.w5(32'hbaf3e88e),
	.w6(32'hbb92de9a),
	.w7(32'h3b32c557),
	.w8(32'hbb96f9d4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc1293),
	.w1(32'hba746264),
	.w2(32'hbbf431af),
	.w3(32'hbb96c865),
	.w4(32'h3adb1671),
	.w5(32'hbb58fdc2),
	.w6(32'hbb2b50c5),
	.w7(32'h3a0b2293),
	.w8(32'hbb6d5ec8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1f966),
	.w1(32'h3a3fc14a),
	.w2(32'hbb9fa534),
	.w3(32'hbb23e958),
	.w4(32'h3b247121),
	.w5(32'hbb373ef1),
	.w6(32'hbb96e651),
	.w7(32'h3b1978e0),
	.w8(32'hbb4bb779),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bb6591),
	.w1(32'hb880a641),
	.w2(32'hb83be5b9),
	.w3(32'hb8cb0687),
	.w4(32'h37de1125),
	.w5(32'h388bd823),
	.w6(32'hb87ef9bc),
	.w7(32'h3719bb3e),
	.w8(32'h3929c9a0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba323932),
	.w1(32'hb9786e6c),
	.w2(32'hb8fd90be),
	.w3(32'hb9b16643),
	.w4(32'h38b56b4b),
	.w5(32'h3960647d),
	.w6(32'hb9ff3738),
	.w7(32'h37eb1c07),
	.w8(32'hb753a25f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39403100),
	.w1(32'h397a9b4c),
	.w2(32'h397a20f2),
	.w3(32'hb8a45e82),
	.w4(32'h3855eb8b),
	.w5(32'h38ef0433),
	.w6(32'h3901cc20),
	.w7(32'h39066c17),
	.w8(32'h394521ac),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4b9d1),
	.w1(32'hb9846f7f),
	.w2(32'h38747a57),
	.w3(32'hb92eb711),
	.w4(32'h3a0951d2),
	.w5(32'h3a1b1c40),
	.w6(32'hb9ba067c),
	.w7(32'h39ba118a),
	.w8(32'h3a41af4f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92c094),
	.w1(32'h3b755923),
	.w2(32'hbbcce858),
	.w3(32'hb9800891),
	.w4(32'h3bd89577),
	.w5(32'hbb6b81f2),
	.w6(32'hbb517e45),
	.w7(32'h3be21dc5),
	.w8(32'hbab08d9f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10756d),
	.w1(32'hbace3309),
	.w2(32'hbb29bbe0),
	.w3(32'hbab0922b),
	.w4(32'hba08213d),
	.w5(32'hbabce57b),
	.w6(32'hbac06bad),
	.w7(32'hb9ea18ce),
	.w8(32'hba147d85),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6a69e),
	.w1(32'hbb236a65),
	.w2(32'hbb93934f),
	.w3(32'hbace3a64),
	.w4(32'hbacb5f5d),
	.w5(32'hbb4c3f36),
	.w6(32'h3a189431),
	.w7(32'hb98d4d5e),
	.w8(32'hbb3a13f5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b6715),
	.w1(32'hba8671eb),
	.w2(32'hb9b15230),
	.w3(32'hbc3188eb),
	.w4(32'h3ad837b7),
	.w5(32'h3adb8ed7),
	.w6(32'hbc5e69ac),
	.w7(32'h396aa827),
	.w8(32'hbadc741d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b025b),
	.w1(32'h394d7581),
	.w2(32'h396cfe13),
	.w3(32'h3a1ba080),
	.w4(32'h3a1e1711),
	.w5(32'h39c7aebb),
	.w6(32'h3a04feb5),
	.w7(32'h3a1c8bfb),
	.w8(32'h39a56c62),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38da7429),
	.w1(32'hb818cf02),
	.w2(32'hba5f6fc6),
	.w3(32'h3a1a5d1c),
	.w4(32'h3979e77f),
	.w5(32'hb94d9f19),
	.w6(32'h388d560f),
	.w7(32'hb911cf40),
	.w8(32'hba2d6645),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394629be),
	.w1(32'h39154ab0),
	.w2(32'h3929adac),
	.w3(32'h3992bb9c),
	.w4(32'h391146bb),
	.w5(32'h38cddf3b),
	.w6(32'h393e9a15),
	.w7(32'h38cdafe9),
	.w8(32'h38f420c1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749ddd),
	.w1(32'hbac10c09),
	.w2(32'hba2d9f65),
	.w3(32'hbb4477f7),
	.w4(32'hba249a79),
	.w5(32'h399290c8),
	.w6(32'hbb5b0332),
	.w7(32'hbb045862),
	.w8(32'hbaca2430),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5de7c8),
	.w1(32'hbb33d861),
	.w2(32'hbbe238e0),
	.w3(32'h3bb1465f),
	.w4(32'hbb290622),
	.w5(32'hbc496dbd),
	.w6(32'h3ad921b6),
	.w7(32'hbaa7c2e8),
	.w8(32'hbbf89da2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca8f5e),
	.w1(32'hba8ed342),
	.w2(32'hbc441702),
	.w3(32'hba1fbf33),
	.w4(32'h3aac6556),
	.w5(32'hbc18d625),
	.w6(32'hbb46121f),
	.w7(32'h3a0689dc),
	.w8(32'hbbec3746),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cecbf),
	.w1(32'hba17edb9),
	.w2(32'hb9ff02bb),
	.w3(32'hb9630428),
	.w4(32'hb9c2e97c),
	.w5(32'hb90ad2be),
	.w6(32'h39ea88de),
	.w7(32'hb8fe24c9),
	.w8(32'hba329f48),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c653d),
	.w1(32'hba87dc37),
	.w2(32'hbb853b65),
	.w3(32'hbb4706de),
	.w4(32'h39580887),
	.w5(32'hbafd16c4),
	.w6(32'hbb95efea),
	.w7(32'hbafea910),
	.w8(32'hbb7f5c27),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8464d6),
	.w1(32'h3a4361e7),
	.w2(32'hbb014853),
	.w3(32'hbb886629),
	.w4(32'h3a7aa4c8),
	.w5(32'hbab0ca44),
	.w6(32'hbb8e7587),
	.w7(32'h3b1b88f1),
	.w8(32'hba826e3e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e9776),
	.w1(32'hba0da60b),
	.w2(32'hbb98c7fa),
	.w3(32'hbad3df9f),
	.w4(32'h3ad32f0f),
	.w5(32'hbb0179d6),
	.w6(32'hbb864c27),
	.w7(32'h38c260ba),
	.w8(32'hbb2303fd),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc024fa),
	.w1(32'hbae4b830),
	.w2(32'hbbdeb837),
	.w3(32'hbb9dc58e),
	.w4(32'h3b40e43e),
	.w5(32'hbaf15353),
	.w6(32'hbb91b42a),
	.w7(32'h3b172d27),
	.w8(32'hbac2c20b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb823a03),
	.w1(32'hbb25ddc8),
	.w2(32'hbc4caed0),
	.w3(32'hbb615ff2),
	.w4(32'hbb20085c),
	.w5(32'hbc31d7de),
	.w6(32'hba4d83ba),
	.w7(32'hba5009d7),
	.w8(32'hbc3de808),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc240b6e),
	.w1(32'hba4de899),
	.w2(32'hbb375223),
	.w3(32'hbbc40698),
	.w4(32'h3b38a158),
	.w5(32'h3a112bdc),
	.w6(32'hbc0a6e77),
	.w7(32'h3ad14bff),
	.w8(32'hbb0f9772),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3856f0),
	.w1(32'hbb931d9c),
	.w2(32'hbbec1db9),
	.w3(32'hbb997ffe),
	.w4(32'h3a988a9a),
	.w5(32'hba9a550e),
	.w6(32'hbb90e40d),
	.w7(32'hbb1a8c7f),
	.w8(32'hbbb7fd5c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52d522),
	.w1(32'hbbe6b62d),
	.w2(32'hbc58faeb),
	.w3(32'hbc123940),
	.w4(32'hbb83c5b5),
	.w5(32'hbc541856),
	.w6(32'hbbf3382e),
	.w7(32'hbad88f91),
	.w8(32'hbc14ebd8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b9e0f),
	.w1(32'hbac621af),
	.w2(32'hbb06517c),
	.w3(32'hbbae82e1),
	.w4(32'h3af5ae22),
	.w5(32'h39807b98),
	.w6(32'hbbf97ffe),
	.w7(32'h3ae711f4),
	.w8(32'hbaa8d044),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3d03f),
	.w1(32'hb95df167),
	.w2(32'hbb9f6559),
	.w3(32'hbb7be3c2),
	.w4(32'h3a6b16d9),
	.w5(32'hbb3e4e7f),
	.w6(32'hbba53ae0),
	.w7(32'hba959e11),
	.w8(32'hbbc2f041),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7c4cc),
	.w1(32'h38332cfa),
	.w2(32'hbb41ebfb),
	.w3(32'h3949533b),
	.w4(32'h3aebdd9d),
	.w5(32'hba9aa13a),
	.w6(32'hba84fc0b),
	.w7(32'h3acdd12b),
	.w8(32'hba7a1e3c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dbea3),
	.w1(32'h3bdf2a33),
	.w2(32'h3ac75eb5),
	.w3(32'hbc2db407),
	.w4(32'h3bbe52f5),
	.w5(32'h3a83d45c),
	.w6(32'hbc5ffd2f),
	.w7(32'h3b89030c),
	.w8(32'hb9a5771e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc033051),
	.w1(32'hb9d58d99),
	.w2(32'h3afb4639),
	.w3(32'hbbe20418),
	.w4(32'h3993a138),
	.w5(32'h3b36598a),
	.w6(32'hbc15d073),
	.w7(32'hbad0d3c9),
	.w8(32'hb94553b9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8729328),
	.w1(32'h38fcf0df),
	.w2(32'h37e8c67f),
	.w3(32'h37cebda1),
	.w4(32'hb8f6ad34),
	.w5(32'hb8f2a766),
	.w6(32'h38c898a2),
	.w7(32'hb863001c),
	.w8(32'hb65f9a4f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e394a),
	.w1(32'h38c9827e),
	.w2(32'h3895af90),
	.w3(32'h3831567e),
	.w4(32'h381f6ff1),
	.w5(32'h381bff0c),
	.w6(32'h38e1a0d2),
	.w7(32'h38e749df),
	.w8(32'h39526827),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35306e),
	.w1(32'hba868ccb),
	.w2(32'hbb200da2),
	.w3(32'hbaf26ab1),
	.w4(32'h3a8b23b1),
	.w5(32'h3a6cdabc),
	.w6(32'hbab793ca),
	.w7(32'h3a021d77),
	.w8(32'hb9c4947f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48e36c),
	.w1(32'h3a49b8dc),
	.w2(32'h3aeafbdb),
	.w3(32'hbbc7f507),
	.w4(32'h3b881eb1),
	.w5(32'h3b895d5d),
	.w6(32'hbc1f585e),
	.w7(32'h3b3c6c4d),
	.w8(32'hb8d1580c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd8f8e),
	.w1(32'hbab64803),
	.w2(32'hbc58f1fa),
	.w3(32'hbaab3f89),
	.w4(32'h3b878598),
	.w5(32'hbc028b27),
	.w6(32'hbac5e005),
	.w7(32'h3b9e434b),
	.w8(32'hbbb77c55),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89465f8),
	.w1(32'h392873a3),
	.w2(32'h38e6b51f),
	.w3(32'h394f30df),
	.w4(32'h3830c0d5),
	.w5(32'h38d27fc2),
	.w6(32'h391d8716),
	.w7(32'h3711d3eb),
	.w8(32'h39069b2b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe736e7),
	.w1(32'hbac3a335),
	.w2(32'hbc4c65d7),
	.w3(32'hbb12e6f9),
	.w4(32'h3ac45f7b),
	.w5(32'hbc0e41ad),
	.w6(32'hbbaaea52),
	.w7(32'h3a37b033),
	.w8(32'hbbdaf5a9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8a66f),
	.w1(32'hb91f566c),
	.w2(32'hbbb73fcb),
	.w3(32'hbb3ed0d6),
	.w4(32'h3b2a45ad),
	.w5(32'hbb15b50a),
	.w6(32'hbb80f758),
	.w7(32'h3b0329ac),
	.w8(32'hbb306424),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb80108),
	.w1(32'hbb5e9556),
	.w2(32'hbc2401e2),
	.w3(32'hbb560e13),
	.w4(32'hbb25694a),
	.w5(32'hbc02cbd0),
	.w6(32'h3a633039),
	.w7(32'hb81c147b),
	.w8(32'hbc135fba),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baafe50),
	.w1(32'h3c25ffee),
	.w2(32'hbb8dda83),
	.w3(32'h3ba1ac37),
	.w4(32'h3c830c99),
	.w5(32'h3b980493),
	.w6(32'hb98de282),
	.w7(32'h3c7bfa41),
	.w8(32'h3b96466b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc287b6b),
	.w1(32'hbb15977d),
	.w2(32'hb9ca4aa5),
	.w3(32'hbc18b38a),
	.w4(32'hbb351000),
	.w5(32'hbac7981d),
	.w6(32'hbc23534c),
	.w7(32'hbb4b09b2),
	.w8(32'hbb8277a9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ca5d7),
	.w1(32'h3a5a2531),
	.w2(32'h3a814fcd),
	.w3(32'hb928586a),
	.w4(32'h39f2ba2b),
	.w5(32'h39644a67),
	.w6(32'h3983e915),
	.w7(32'h3a673cf2),
	.w8(32'h39d0ca43),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2e26d),
	.w1(32'h3b54fb19),
	.w2(32'h39b47d04),
	.w3(32'hbb3fe4aa),
	.w4(32'h3bb998da),
	.w5(32'h3b3af871),
	.w6(32'hbc092b85),
	.w7(32'h3b357b26),
	.w8(32'hb9a1b11e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e39af),
	.w1(32'hbac2b915),
	.w2(32'hba85bb2a),
	.w3(32'hbc64bc7d),
	.w4(32'hb96f1bdc),
	.w5(32'h38f47536),
	.w6(32'hbc8518d3),
	.w7(32'hbb1692c5),
	.w8(32'hbbb8b1c2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a15131),
	.w1(32'h3bb0bba1),
	.w2(32'hb993da59),
	.w3(32'hb90a2a8b),
	.w4(32'h3bdad3f2),
	.w5(32'h3aba791b),
	.w6(32'hbb5a86fc),
	.w7(32'h3b928565),
	.w8(32'hba50e53e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34a77a),
	.w1(32'hbaa55874),
	.w2(32'hbb072a69),
	.w3(32'hbab09017),
	.w4(32'hbb202825),
	.w5(32'hbb0d57f3),
	.w6(32'hb9e4c628),
	.w7(32'hba930545),
	.w8(32'hbb1f4a9a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97d42c),
	.w1(32'hba8ecd64),
	.w2(32'hba5ec850),
	.w3(32'hba7c7bc6),
	.w4(32'hba7dcddc),
	.w5(32'hba5a0985),
	.w6(32'hba8b9d29),
	.w7(32'hba974fb5),
	.w8(32'hba92cfe1),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2dd8d),
	.w1(32'hbb19b564),
	.w2(32'hbbd08ba4),
	.w3(32'hbb8952ae),
	.w4(32'hb9fb7cd1),
	.w5(32'hbbb57f81),
	.w6(32'hbbe2bab6),
	.w7(32'hbb105b7d),
	.w8(32'hbbd862d6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91e2bb),
	.w1(32'h39620590),
	.w2(32'hba1aaeb6),
	.w3(32'h3a70df0e),
	.w4(32'h38dba120),
	.w5(32'hb8df171c),
	.w6(32'h3a9aeda2),
	.w7(32'h3a22377d),
	.w8(32'hb49c34a0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ab0c6),
	.w1(32'h3afa149a),
	.w2(32'hbb23473a),
	.w3(32'h3947aa5c),
	.w4(32'h3b7c25f8),
	.w5(32'hba584e9a),
	.w6(32'hbb447da6),
	.w7(32'h3b7d57d8),
	.w8(32'h3a8595fb),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380dc83e),
	.w1(32'h38cfbbc4),
	.w2(32'hba4e43d2),
	.w3(32'h39e2ac72),
	.w4(32'h39582853),
	.w5(32'hba433925),
	.w6(32'h393cbc6d),
	.w7(32'h39a3ffbf),
	.w8(32'hb9df1813),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb00c38),
	.w1(32'h3b093aa8),
	.w2(32'hbc2057ab),
	.w3(32'h3b88d705),
	.w4(32'h3b61666a),
	.w5(32'hbbc0089d),
	.w6(32'h3a7ea601),
	.w7(32'h3b1e6376),
	.w8(32'hbbecbb57),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cafeee),
	.w1(32'hb8814b9c),
	.w2(32'h38914b3d),
	.w3(32'h36f55774),
	.w4(32'hb94d1755),
	.w5(32'hb92db9b3),
	.w6(32'h372e293d),
	.w7(32'hb94833e0),
	.w8(32'hb90dc633),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27adc8),
	.w1(32'hb9fb8b35),
	.w2(32'hba0fcdb5),
	.w3(32'hb9d7abca),
	.w4(32'hb999c4d5),
	.w5(32'hb9ed80f8),
	.w6(32'hba1f67e7),
	.w7(32'hba03cd53),
	.w8(32'hba042600),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36007d),
	.w1(32'h394bac68),
	.w2(32'hba21fca2),
	.w3(32'hbc0c41fd),
	.w4(32'h3a5fd345),
	.w5(32'h3a5054e1),
	.w6(32'hbc4ae188),
	.w7(32'hbb2b76a3),
	.w8(32'hbb2016fe),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc512ccb),
	.w1(32'h3a9739bd),
	.w2(32'hbc1e3c55),
	.w3(32'hbc0344c3),
	.w4(32'hbb19bd19),
	.w5(32'hbca28385),
	.w6(32'hbc238276),
	.w7(32'hb9af8876),
	.w8(32'hbc628d77),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d8a24),
	.w1(32'h3af6ce25),
	.w2(32'hbb1e191d),
	.w3(32'h38c8ca75),
	.w4(32'h3b5defdf),
	.w5(32'hbac0a063),
	.w6(32'hbb3e99ab),
	.w7(32'h3ae442c4),
	.w8(32'hbb36410a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bb6be),
	.w1(32'hbb20a5fa),
	.w2(32'hbc24d7be),
	.w3(32'hbbb7cd1e),
	.w4(32'h3a97a84f),
	.w5(32'hbbdd5d3e),
	.w6(32'hbbce532b),
	.w7(32'h3ac74384),
	.w8(32'hbbec5825),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94e925),
	.w1(32'hb9828bf4),
	.w2(32'hbac4f424),
	.w3(32'hbb12e503),
	.w4(32'h3927d582),
	.w5(32'hb8fdc9ee),
	.w6(32'hbae7b4e9),
	.w7(32'hb96da909),
	.w8(32'hba10ea3e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cbfaf),
	.w1(32'hbab99669),
	.w2(32'hbc9c8752),
	.w3(32'hbbc33f4e),
	.w4(32'h3bc9abbf),
	.w5(32'hbc0e9180),
	.w6(32'hbc116dad),
	.w7(32'hb92e7af5),
	.w8(32'hbc527ecd),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc252889),
	.w1(32'hbacbda85),
	.w2(32'hbc323f21),
	.w3(32'hbbd60cf7),
	.w4(32'h3b5247ef),
	.w5(32'hbb987895),
	.w6(32'hbc17237e),
	.w7(32'h3ac38137),
	.w8(32'hbbeb8193),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb673c3c),
	.w1(32'hb9e870c0),
	.w2(32'hbc5e1236),
	.w3(32'h3a1c8c2b),
	.w4(32'h3b019957),
	.w5(32'hbc339332),
	.w6(32'hba652fc8),
	.w7(32'h3b7b388a),
	.w8(32'hbbd42624),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984c290),
	.w1(32'h39890d66),
	.w2(32'hb8f22697),
	.w3(32'h3979f2c0),
	.w4(32'h3a1698e8),
	.w5(32'h39fb574b),
	.w6(32'h394e2d3c),
	.w7(32'h39f6e713),
	.w8(32'h39cd9a9f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3fc4d),
	.w1(32'hbabd9939),
	.w2(32'hbb90540f),
	.w3(32'hbb8cd56b),
	.w4(32'hba8e1480),
	.w5(32'hbb7d750e),
	.w6(32'hbb591fb2),
	.w7(32'h3a436f2a),
	.w8(32'hbae9afd7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398405d4),
	.w1(32'h38b65479),
	.w2(32'h3916fb9e),
	.w3(32'h397f71ce),
	.w4(32'h37937358),
	.w5(32'h38cff9a4),
	.w6(32'h39a9fb4d),
	.w7(32'h38f1df1b),
	.w8(32'h3938ba8d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b064497),
	.w1(32'h3a2b73bb),
	.w2(32'hbb9de208),
	.w3(32'h3b332eb9),
	.w4(32'h3b1f9108),
	.w5(32'hba269c06),
	.w6(32'h3ac3681f),
	.w7(32'h3a853c1f),
	.w8(32'hbb293c64),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dfe8f),
	.w1(32'h3ac20ecb),
	.w2(32'hb825d819),
	.w3(32'hbb049a1b),
	.w4(32'h3a5ee676),
	.w5(32'h393e2650),
	.w6(32'hbb124ffc),
	.w7(32'h3a31c06d),
	.w8(32'hb9a545a7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe67658),
	.w1(32'hba74303a),
	.w2(32'hbc0a8007),
	.w3(32'hbb8945ba),
	.w4(32'h3a97666f),
	.w5(32'hbb472b7d),
	.w6(32'hbba0902c),
	.w7(32'h3a2f5fb6),
	.w8(32'hbbb778aa),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39170239),
	.w1(32'hb90799c1),
	.w2(32'hb7067108),
	.w3(32'hb834d0a8),
	.w4(32'hb8c5f2eb),
	.w5(32'h3846c251),
	.w6(32'h38c8788a),
	.w7(32'h384b7da0),
	.w8(32'h39345eeb),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c3341e),
	.w1(32'h3848a151),
	.w2(32'hb845626d),
	.w3(32'hb6a4ec68),
	.w4(32'hb8f93433),
	.w5(32'h379067f6),
	.w6(32'h39592eba),
	.w7(32'h39326388),
	.w8(32'h390a448b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eff0c),
	.w1(32'h3a4b1259),
	.w2(32'hb9101804),
	.w3(32'hba7ac3ec),
	.w4(32'h3af85dc7),
	.w5(32'h3a572f2f),
	.w6(32'hbb069915),
	.w7(32'h3ace9421),
	.w8(32'h3a483c6c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc159daa),
	.w1(32'hbb3a1853),
	.w2(32'hbbd1b48f),
	.w3(32'hbbbb4462),
	.w4(32'hb90c863d),
	.w5(32'hbb175b12),
	.w6(32'hbbf36ebc),
	.w7(32'hbb108b5e),
	.w8(32'hbbcfd9c9),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84448c),
	.w1(32'h382454e5),
	.w2(32'hbab70546),
	.w3(32'hbb04aaf2),
	.w4(32'hba0ef262),
	.w5(32'hbaf0c25b),
	.w6(32'h3a7192d2),
	.w7(32'h3b3cd973),
	.w8(32'hbb462f8e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9828e),
	.w1(32'hba27a996),
	.w2(32'hbb0c26bc),
	.w3(32'hbaee907f),
	.w4(32'hba24dd5e),
	.w5(32'hbab753e4),
	.w6(32'hbaed2a0f),
	.w7(32'hb9be892d),
	.w8(32'hbb0c1d4b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20538f),
	.w1(32'hbb1de30a),
	.w2(32'hbcd65ddd),
	.w3(32'h3a8a7944),
	.w4(32'h3b080f8c),
	.w5(32'hbc8e3a4c),
	.w6(32'h3bcac192),
	.w7(32'h3b77dfb1),
	.w8(32'hbc660312),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3dfd1),
	.w1(32'hba968ac1),
	.w2(32'hbbc91f55),
	.w3(32'hbc915561),
	.w4(32'h3b8f0f4c),
	.w5(32'h3b8a46ef),
	.w6(32'hbc96c94a),
	.w7(32'h3b122faf),
	.w8(32'hbabe4aa6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ba044),
	.w1(32'hb9e4eebe),
	.w2(32'hba2db480),
	.w3(32'h3a9cdd9e),
	.w4(32'hba98d034),
	.w5(32'hba984506),
	.w6(32'h3aba119e),
	.w7(32'hb83a69a7),
	.w8(32'hbac2cafc),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a5cf6),
	.w1(32'h387bd2fb),
	.w2(32'h38983fc1),
	.w3(32'h37d253f4),
	.w4(32'hb90dcd38),
	.w5(32'hb87305cf),
	.w6(32'h38de3b22),
	.w7(32'hb7a80f60),
	.w8(32'h37693466),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378ed53b),
	.w1(32'h383160b3),
	.w2(32'hb88fb82b),
	.w3(32'hb7fecbad),
	.w4(32'hb896d94f),
	.w5(32'h38468b39),
	.w6(32'h3918d049),
	.w7(32'h38dbbe1c),
	.w8(32'h39610744),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967bdb5),
	.w1(32'h38913f51),
	.w2(32'h38fe5b5d),
	.w3(32'h39219e53),
	.w4(32'hb853795e),
	.w5(32'h389e0f01),
	.w6(32'h3994bdcd),
	.w7(32'h38253ad2),
	.w8(32'h394ab354),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf5c72),
	.w1(32'hbb062703),
	.w2(32'hbb2c1aa8),
	.w3(32'hb96f7fcd),
	.w4(32'hbb11183d),
	.w5(32'hbb2d9823),
	.w6(32'hba23d0f1),
	.w7(32'hbb301dbf),
	.w8(32'hbb8913ab),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc572b09),
	.w1(32'hbb7137a6),
	.w2(32'hbbd1775d),
	.w3(32'hbbd40f21),
	.w4(32'h3a25960b),
	.w5(32'hbb359650),
	.w6(32'hbc184fa6),
	.w7(32'hba513c4f),
	.w8(32'hbc06fbfc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cb628),
	.w1(32'hb9a4d372),
	.w2(32'hbc30f3ec),
	.w3(32'hbb52974d),
	.w4(32'h3bf5a1d7),
	.w5(32'hbadcd07a),
	.w6(32'hbbaae609),
	.w7(32'h3bf6c120),
	.w8(32'hba81a5e2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0932d8),
	.w1(32'h3b1e95d2),
	.w2(32'h38b2209e),
	.w3(32'hb99d0ce5),
	.w4(32'h3b15ae99),
	.w5(32'h3a2f2d34),
	.w6(32'hbb083de7),
	.w7(32'hb938fc76),
	.w8(32'hbb0084d2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e3567),
	.w1(32'hbbc636bb),
	.w2(32'hbc8457d5),
	.w3(32'hbb56d506),
	.w4(32'h3aded997),
	.w5(32'hbc164711),
	.w6(32'hbbbf02bb),
	.w7(32'h3a2be08e),
	.w8(32'hbc20091a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1966b),
	.w1(32'hbaa96959),
	.w2(32'hbb55fb96),
	.w3(32'h3a68d1ac),
	.w4(32'h373527b4),
	.w5(32'hbaffaf2e),
	.w6(32'h3a8f5095),
	.w7(32'h39a1ec50),
	.w8(32'hbb117116),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962a2eb),
	.w1(32'h39600638),
	.w2(32'h396d4b12),
	.w3(32'h39735ad9),
	.w4(32'h38a9abcc),
	.w5(32'h393cab8e),
	.w6(32'h39c37b0f),
	.w7(32'h390c345a),
	.w8(32'h395daa37),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d5e04),
	.w1(32'hbae38b07),
	.w2(32'hb807d885),
	.w3(32'hbac6ddca),
	.w4(32'hb9e91af3),
	.w5(32'h3a3e8207),
	.w6(32'h35bc6d34),
	.w7(32'h3889258a),
	.w8(32'h3a692cf6),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a373fe6),
	.w1(32'h3972a1c8),
	.w2(32'h3a2aa14b),
	.w3(32'h3a029082),
	.w4(32'h385185f4),
	.w5(32'h39c1db2c),
	.w6(32'h3a3f815e),
	.w7(32'h39a99eca),
	.w8(32'h3a26c4b4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd65d03),
	.w1(32'h3aac96d4),
	.w2(32'hba221552),
	.w3(32'hbb577f91),
	.w4(32'h3b8298da),
	.w5(32'h3b75e294),
	.w6(32'hbbb1c4b2),
	.w7(32'h3ac9da11),
	.w8(32'h3ade30dc),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc399171),
	.w1(32'h3b644190),
	.w2(32'hbb13e576),
	.w3(32'hbbfcab91),
	.w4(32'h3bc5d9b6),
	.w5(32'h3a0c6f52),
	.w6(32'hbc7b78cf),
	.w7(32'h3a99ad8c),
	.w8(32'hbbdbc8e4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ed4e7),
	.w1(32'hbad92e02),
	.w2(32'hbc0695e8),
	.w3(32'hbbdc686c),
	.w4(32'h3b564fbb),
	.w5(32'hbb4222f5),
	.w6(32'hbc2d2910),
	.w7(32'h38d54898),
	.w8(32'hbbe287ed),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fcd2d),
	.w1(32'hbad73ba9),
	.w2(32'hbac8bf42),
	.w3(32'hbb89f206),
	.w4(32'hbadab0c5),
	.w5(32'hbad925da),
	.w6(32'hbbb83834),
	.w7(32'hbb5fd625),
	.w8(32'hbb6a6196),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc666c37),
	.w1(32'hba6e71fd),
	.w2(32'hbbc799c3),
	.w3(32'hbc0b11ac),
	.w4(32'h3b989d83),
	.w5(32'h3a164f28),
	.w6(32'hbc5a93c6),
	.w7(32'hb86eee48),
	.w8(32'hbb9fe050),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81be9f),
	.w1(32'h3a1fdc99),
	.w2(32'hbbaa8312),
	.w3(32'hbb18daa9),
	.w4(32'h3a9143dc),
	.w5(32'hbb5a7203),
	.w6(32'hbb85f62a),
	.w7(32'h3979b5b0),
	.w8(32'hbb1aab32),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8021e),
	.w1(32'h3b22c076),
	.w2(32'hbc7f986a),
	.w3(32'h3a0fec5b),
	.w4(32'h3c0efecc),
	.w5(32'hbc0950c3),
	.w6(32'h3a2c5f5d),
	.w7(32'h3c14a85c),
	.w8(32'hbc1da21b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946be26),
	.w1(32'h380a3d4d),
	.w2(32'h37d0ddca),
	.w3(32'h390b435e),
	.w4(32'h36ea0c14),
	.w5(32'hb791d051),
	.w6(32'h392f1433),
	.w7(32'h38d0dd32),
	.w8(32'h383641b8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980aee6),
	.w1(32'h396f1a64),
	.w2(32'h3892a0b5),
	.w3(32'h3806b917),
	.w4(32'h3886b1ce),
	.w5(32'hb8666ad7),
	.w6(32'h388a02fd),
	.w7(32'h39572c37),
	.w8(32'h396715a8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a992e),
	.w1(32'h3a699fc1),
	.w2(32'hbc227ba0),
	.w3(32'hbb94ac51),
	.w4(32'h3b5b584b),
	.w5(32'hbc0a0eb2),
	.w6(32'hbc0797b2),
	.w7(32'h3a57e83c),
	.w8(32'hbc33695e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe117ad),
	.w1(32'h3b8637cf),
	.w2(32'hbc4e1160),
	.w3(32'hbb5a30cd),
	.w4(32'h3b87c6ae),
	.w5(32'hbc77e3cf),
	.w6(32'hbbd3c633),
	.w7(32'h3b8d79c2),
	.w8(32'hbc1a65b2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f9a02),
	.w1(32'hb9452288),
	.w2(32'hbc199e5d),
	.w3(32'hbb7862b1),
	.w4(32'h3bd07a7a),
	.w5(32'hbb6d1185),
	.w6(32'hbc0c295b),
	.w7(32'h3b9376d0),
	.w8(32'hbb7bc1b2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c7205),
	.w1(32'hba0c8af9),
	.w2(32'hb9c0f3b0),
	.w3(32'hbb67dbe8),
	.w4(32'hbb9ac8e1),
	.w5(32'hba154852),
	.w6(32'h3b7d674c),
	.w7(32'h39a12576),
	.w8(32'hbb72e754),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb800d87a),
	.w1(32'hb941cd54),
	.w2(32'h38a928bd),
	.w3(32'hb95cfbf6),
	.w4(32'hb974b739),
	.w5(32'h3908513d),
	.w6(32'hb80f4416),
	.w7(32'hb94abf28),
	.w8(32'h3925c838),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa7737),
	.w1(32'hba183730),
	.w2(32'h38ee6911),
	.w3(32'hba89c625),
	.w4(32'hba1d995d),
	.w5(32'hb8241dca),
	.w6(32'hba455212),
	.w7(32'hba297f5f),
	.w8(32'h386420fc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba12ffc),
	.w1(32'hb7954293),
	.w2(32'hbbb1a855),
	.w3(32'h3b951867),
	.w4(32'hbb6bfaee),
	.w5(32'hbc1de6f0),
	.w6(32'h3bafbcb7),
	.w7(32'h3a3c2ecb),
	.w8(32'hbc0b5412),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29bfd4),
	.w1(32'hbb92664c),
	.w2(32'hbc8419e9),
	.w3(32'hbb87f133),
	.w4(32'hba482dc9),
	.w5(32'hbc481dfb),
	.w6(32'hbb0d030f),
	.w7(32'h3976d69d),
	.w8(32'hbc4c45c1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b961f),
	.w1(32'hbb645a6f),
	.w2(32'hbb5bb6a0),
	.w3(32'hbb85e3d0),
	.w4(32'hbb9b20de),
	.w5(32'hbba25ccf),
	.w6(32'h3a2d5696),
	.w7(32'hbb0b1b4d),
	.w8(32'hbbd7d474),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8b80d),
	.w1(32'h3b7554b4),
	.w2(32'hb7a95ce1),
	.w3(32'hbbbb1a92),
	.w4(32'h3b9ba9e2),
	.w5(32'h3a9f688a),
	.w6(32'hbc1cc5e2),
	.w7(32'h3af0d0a5),
	.w8(32'hbacaad39),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc67704),
	.w1(32'h3a365ed0),
	.w2(32'hbbdcb6ed),
	.w3(32'hbbabaffa),
	.w4(32'h3bb0ccb1),
	.w5(32'hb9ebd206),
	.w6(32'hbc189f0b),
	.w7(32'h3b2aae0a),
	.w8(32'hbb2eaf23),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a30478),
	.w1(32'h37f09641),
	.w2(32'h38bf6089),
	.w3(32'h37b54431),
	.w4(32'hb6d2f880),
	.w5(32'h38963fab),
	.w6(32'h38327f38),
	.w7(32'h3755b8a6),
	.w8(32'h38048bda),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c8157),
	.w1(32'h38907ea9),
	.w2(32'h38b8fda5),
	.w3(32'h396deb42),
	.w4(32'h382ad2b9),
	.w5(32'h38c72f4e),
	.w6(32'h397d45d1),
	.w7(32'h38ac0edb),
	.w8(32'h38f2d998),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a764282),
	.w1(32'h3936e4ea),
	.w2(32'h39ea2707),
	.w3(32'h3aabc0de),
	.w4(32'hba10df20),
	.w5(32'hba58eda8),
	.w6(32'h397b2386),
	.w7(32'hba5363b4),
	.w8(32'hba0a18a6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dba2f7),
	.w1(32'hb884ac45),
	.w2(32'hb8097853),
	.w3(32'h3903d580),
	.w4(32'hb91247e0),
	.w5(32'hbb94e97d),
	.w6(32'h39596915),
	.w7(32'hb90a8310),
	.w8(32'hbb9722ff),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9414b3),
	.w1(32'hbc0b8076),
	.w2(32'hbbbe0eeb),
	.w3(32'hbbf30013),
	.w4(32'hb8283007),
	.w5(32'hbb1a4389),
	.w6(32'hbbd289fb),
	.w7(32'hbb0ce20e),
	.w8(32'h3a47f939),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03d33d),
	.w1(32'hbab19931),
	.w2(32'hbb808d5c),
	.w3(32'hba834df4),
	.w4(32'hbb1ea94b),
	.w5(32'hbb6fd908),
	.w6(32'h3aad5ef7),
	.w7(32'h39aef79d),
	.w8(32'hbc062588),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc7a42),
	.w1(32'hba0ad35b),
	.w2(32'hbbbb3d65),
	.w3(32'hbc1ee26b),
	.w4(32'h3a46275b),
	.w5(32'h3a12cba5),
	.w6(32'hbc6461f8),
	.w7(32'hbb179cde),
	.w8(32'h3b62a507),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf0d4d),
	.w1(32'hbbbd4a01),
	.w2(32'hbbb1eb2d),
	.w3(32'hba0bb19a),
	.w4(32'hbb8b8465),
	.w5(32'hbb6756d9),
	.w6(32'h3bb03f4a),
	.w7(32'hbc135362),
	.w8(32'h3a5e54f3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04f67c),
	.w1(32'h3c351149),
	.w2(32'hbc06b00f),
	.w3(32'h3c43feb6),
	.w4(32'h3c270233),
	.w5(32'hbc17cf55),
	.w6(32'h3c710711),
	.w7(32'h3be1ee4d),
	.w8(32'hbc336529),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b000b32),
	.w1(32'h3bbfcc82),
	.w2(32'hbbc661cd),
	.w3(32'h3ac24d94),
	.w4(32'hbbe8f9c2),
	.w5(32'hbb45e59e),
	.w6(32'h3bba5810),
	.w7(32'hbbc64a46),
	.w8(32'hbbc2c643),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa325ad),
	.w1(32'h3b852e9e),
	.w2(32'hbbadff83),
	.w3(32'hbb579a96),
	.w4(32'hba7dbf8f),
	.w5(32'hbb0faae8),
	.w6(32'hbaca557d),
	.w7(32'hb915babc),
	.w8(32'hba908e60),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d042d9),
	.w1(32'hba4e0f39),
	.w2(32'hbbd8eba4),
	.w3(32'h3b285e4e),
	.w4(32'hbb8c9605),
	.w5(32'hbbf8cf14),
	.w6(32'hbb1be4db),
	.w7(32'h3ade7dba),
	.w8(32'hbbff68b0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb466977),
	.w1(32'hba255bc1),
	.w2(32'h3b04d81a),
	.w3(32'h3b1bac4b),
	.w4(32'hbad2aab4),
	.w5(32'h3902c871),
	.w6(32'h3ba0700e),
	.w7(32'h3b75eaf3),
	.w8(32'hba949815),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d8945),
	.w1(32'hbb27cc6f),
	.w2(32'hb9cb121c),
	.w3(32'hbbd50b80),
	.w4(32'hbb3b6253),
	.w5(32'hbb4ef32a),
	.w6(32'hbbad8c40),
	.w7(32'hbb570639),
	.w8(32'hbc13692b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd106eb),
	.w1(32'hbb81cbc4),
	.w2(32'hbb61eef4),
	.w3(32'hbbfac84a),
	.w4(32'hb8970012),
	.w5(32'hba86263c),
	.w6(32'hbc0d7a2e),
	.w7(32'hbb80c35e),
	.w8(32'hbae70c88),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd2ddb),
	.w1(32'h39f54871),
	.w2(32'h3b048593),
	.w3(32'hbaf6e2a1),
	.w4(32'h3b26adb4),
	.w5(32'h3aa819c3),
	.w6(32'hb95539cc),
	.w7(32'h3a4bbfcf),
	.w8(32'hb994d6a2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a31d5),
	.w1(32'hba60817a),
	.w2(32'hbb209855),
	.w3(32'hbb83caf6),
	.w4(32'hbac4d057),
	.w5(32'hbb47aad7),
	.w6(32'hbbf664d1),
	.w7(32'hba82f883),
	.w8(32'hbc2406ac),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fc748),
	.w1(32'hbc4824b2),
	.w2(32'hbcf616d2),
	.w3(32'hbc2b3560),
	.w4(32'hbc381e77),
	.w5(32'hbc4a1153),
	.w6(32'hbbd01dd6),
	.w7(32'hbc31ee99),
	.w8(32'hbc167380),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc027f67),
	.w1(32'hba4b7cf7),
	.w2(32'hbc13c17e),
	.w3(32'h3b094441),
	.w4(32'h3b0abfac),
	.w5(32'hbc4faa6d),
	.w6(32'h3a34c60a),
	.w7(32'h3ae9c9ff),
	.w8(32'hbca29d39),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6ad22),
	.w1(32'hbc3e23f6),
	.w2(32'h3ac68f15),
	.w3(32'hbc213ee7),
	.w4(32'h3b164ed0),
	.w5(32'hbc3a7bd1),
	.w6(32'hbc008887),
	.w7(32'hbb6bf701),
	.w8(32'hbc43a0f9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4898a),
	.w1(32'hb9c7517e),
	.w2(32'hbb0652f8),
	.w3(32'hbb18ccfe),
	.w4(32'h3ba64cce),
	.w5(32'hbc5a0e7c),
	.w6(32'hbb624b55),
	.w7(32'hb8a12121),
	.w8(32'hbc315a7d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d6950),
	.w1(32'hbbd1a0fa),
	.w2(32'hbc9a436b),
	.w3(32'hbb7a588d),
	.w4(32'hbb175150),
	.w5(32'h3a87de31),
	.w6(32'hbbbc063a),
	.w7(32'hbbe60dd4),
	.w8(32'h3b8b6487),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73b6a9),
	.w1(32'hba5c031d),
	.w2(32'hbbb02e05),
	.w3(32'hbb25f7c4),
	.w4(32'hbba36720),
	.w5(32'hbaa50281),
	.w6(32'hb92e58db),
	.w7(32'hbba1785d),
	.w8(32'hb997e6fe),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af20cad),
	.w1(32'h3b8b35a9),
	.w2(32'hba90b9db),
	.w3(32'h3afae617),
	.w4(32'hba6ae2bf),
	.w5(32'hbaa105c8),
	.w6(32'h3af953dd),
	.w7(32'h3b06ccb7),
	.w8(32'hbb52f721),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fc35b),
	.w1(32'hbb85db7d),
	.w2(32'hbade99f1),
	.w3(32'hbb843290),
	.w4(32'h3c161cd4),
	.w5(32'hbc58e93e),
	.w6(32'hba5c52cf),
	.w7(32'h3b71d91f),
	.w8(32'hbc814ce6),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07d333),
	.w1(32'hbb9ffd48),
	.w2(32'hbb26f225),
	.w3(32'hbb9be989),
	.w4(32'h3aed7514),
	.w5(32'h3bd19fa0),
	.w6(32'hbb1879c2),
	.w7(32'hbb25a238),
	.w8(32'h3bdae90d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cea1f9a),
	.w1(32'h39b63392),
	.w2(32'h3c012654),
	.w3(32'hbc22f88e),
	.w4(32'h3ba50e20),
	.w5(32'hbb70a7cb),
	.w6(32'hbc936bed),
	.w7(32'h3c2dc30b),
	.w8(32'hbb9e9cb3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4da91),
	.w1(32'hbb241ec9),
	.w2(32'h3bb910b7),
	.w3(32'hbab57c92),
	.w4(32'h3b8fab67),
	.w5(32'hbb5b772e),
	.w6(32'h3aa4b201),
	.w7(32'h3b8d3da2),
	.w8(32'hbbc7d332),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e087d),
	.w1(32'hba65a06c),
	.w2(32'h3a5de8fa),
	.w3(32'hb7a62f5a),
	.w4(32'hbc469e79),
	.w5(32'h3b4db204),
	.w6(32'hbb4e0d06),
	.w7(32'hbbc5c9b8),
	.w8(32'h3b0d65c2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd989a6),
	.w1(32'h3a8b9a46),
	.w2(32'hbbc3a065),
	.w3(32'hbae79976),
	.w4(32'hbb861db5),
	.w5(32'hb9658caa),
	.w6(32'h3a0b00e4),
	.w7(32'hba5abeb1),
	.w8(32'hbb9fbc57),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29ab90),
	.w1(32'hba5e0225),
	.w2(32'h3a24734b),
	.w3(32'h3aaa11aa),
	.w4(32'hbb13dd6c),
	.w5(32'h3b9449b7),
	.w6(32'h3a89edbe),
	.w7(32'hbb6fafb1),
	.w8(32'hbc377ef3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f3c48),
	.w1(32'hbcbd4cae),
	.w2(32'hbc3fc116),
	.w3(32'hbc80ef77),
	.w4(32'hbc244a2e),
	.w5(32'hbc04f71f),
	.w6(32'hbc3877d1),
	.w7(32'hbca47eed),
	.w8(32'hbc57712d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2930b),
	.w1(32'hbbc6d448),
	.w2(32'hbb522937),
	.w3(32'hb9165b69),
	.w4(32'hbab13fb4),
	.w5(32'h3b8a70c8),
	.w6(32'hbb64bb08),
	.w7(32'hba269864),
	.w8(32'hbb3f7e60),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95b92),
	.w1(32'h3b67e3f0),
	.w2(32'h3b93c2e9),
	.w3(32'hbbad95a4),
	.w4(32'h3a524c5c),
	.w5(32'hb9765ef6),
	.w6(32'hbc0bcd00),
	.w7(32'hbba78a02),
	.w8(32'hbc2f3143),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule