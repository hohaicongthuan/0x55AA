module layer_10_featuremap_123(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c6be3),
	.w1(32'hbc96133a),
	.w2(32'h3d10954a),
	.w3(32'h3ba04847),
	.w4(32'hbc62b287),
	.w5(32'hbbecaf55),
	.w6(32'hbc113525),
	.w7(32'hbc34c085),
	.w8(32'hbc6b2a29),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80468e),
	.w1(32'hbc58068d),
	.w2(32'h3b9b92dd),
	.w3(32'hbc15d5ce),
	.w4(32'hbac4e49b),
	.w5(32'h3b669ce8),
	.w6(32'hbbe88df8),
	.w7(32'h3b225e22),
	.w8(32'hb980c4bb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf947e2),
	.w1(32'h39db1bab),
	.w2(32'h3a6fbcec),
	.w3(32'hbb813f5f),
	.w4(32'h3b09197a),
	.w5(32'h3b232e7d),
	.w6(32'h39d1142f),
	.w7(32'hba8efc5d),
	.w8(32'hbb3d93ac),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb302a23),
	.w1(32'hbcd19c6d),
	.w2(32'h3be523a9),
	.w3(32'hbadc3f51),
	.w4(32'hbaf9e35f),
	.w5(32'h398d1b3b),
	.w6(32'hbc131689),
	.w7(32'h3c3239ec),
	.w8(32'h3ca431e4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf28cf8),
	.w1(32'hbb959852),
	.w2(32'hbd1f7679),
	.w3(32'h3b171f18),
	.w4(32'hbc2171c4),
	.w5(32'hbc6e14eb),
	.w6(32'hbc2056bf),
	.w7(32'hbc04bc03),
	.w8(32'h3a2324a8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b347dd0),
	.w1(32'hbc7acf7a),
	.w2(32'hbbebd5d5),
	.w3(32'hbbce223b),
	.w4(32'hbc118f95),
	.w5(32'h3b1fef85),
	.w6(32'hbc156008),
	.w7(32'h3b738df6),
	.w8(32'h3c46462c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a82c6),
	.w1(32'hbc618aaa),
	.w2(32'hbc1034ce),
	.w3(32'h3c3eec1b),
	.w4(32'hbc0b15a0),
	.w5(32'hbb80fbeb),
	.w6(32'hbbd2df76),
	.w7(32'hba6ad092),
	.w8(32'hbb78af8a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9045a5),
	.w1(32'h3bca8d84),
	.w2(32'hbc428a5f),
	.w3(32'hbc1c89ef),
	.w4(32'hbb09e8ef),
	.w5(32'hbb80eec6),
	.w6(32'h3a8a521c),
	.w7(32'hbb853aed),
	.w8(32'hbb6905f4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e5b37),
	.w1(32'h3b7895b6),
	.w2(32'hb8f1e752),
	.w3(32'hbb2f990a),
	.w4(32'h3b9e4ebe),
	.w5(32'h38cb2792),
	.w6(32'h3bb2b9e2),
	.w7(32'hbadc08c6),
	.w8(32'h3a0aefb6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826417),
	.w1(32'hbc779a4c),
	.w2(32'h39339474),
	.w3(32'h3b3cc81c),
	.w4(32'h3aaa61a7),
	.w5(32'hb953b276),
	.w6(32'hbbf92eb4),
	.w7(32'h3a65f6ac),
	.w8(32'h39ff9b9d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c2d8f),
	.w1(32'h3b90bfc9),
	.w2(32'h3c1e2b37),
	.w3(32'hbab0fcd9),
	.w4(32'hbb71785f),
	.w5(32'h3b0e853f),
	.w6(32'h3b4f241b),
	.w7(32'h3bfdc6b6),
	.w8(32'hbab9a9b2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2da084),
	.w1(32'hbb05f0dc),
	.w2(32'hbbf44b18),
	.w3(32'h3a8286ee),
	.w4(32'hbb6e7b5f),
	.w5(32'hbc57b637),
	.w6(32'hbb88401d),
	.w7(32'hbb6b2166),
	.w8(32'hbc448e5f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc001731),
	.w1(32'h3bca44a4),
	.w2(32'hbc0939ca),
	.w3(32'hbc700160),
	.w4(32'h3a8a8749),
	.w5(32'hbbcfa5ec),
	.w6(32'h3bb23c53),
	.w7(32'hbb47982e),
	.w8(32'hbc16ccc4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42298d),
	.w1(32'h3d31d487),
	.w2(32'h3b490834),
	.w3(32'hbc2528dd),
	.w4(32'h3c39f8ea),
	.w5(32'hbbfd6fe8),
	.w6(32'h3cac22f2),
	.w7(32'hbbde25be),
	.w8(32'hbcb26091),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3ef956),
	.w1(32'h3b84616f),
	.w2(32'hbc15dbaf),
	.w3(32'hbccf6142),
	.w4(32'hba7bb748),
	.w5(32'hbbc6f879),
	.w6(32'hbc0584f0),
	.w7(32'h3bfcaaf4),
	.w8(32'h3b3a5de9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcba546),
	.w1(32'hbbb8d179),
	.w2(32'hbb66309d),
	.w3(32'hbca75f9e),
	.w4(32'hba813866),
	.w5(32'hba7fd2fa),
	.w6(32'hbb3a9626),
	.w7(32'hbb15777c),
	.w8(32'h399d001b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963f9c4),
	.w1(32'hbad83ec4),
	.w2(32'hba06e06b),
	.w3(32'h3b10dea3),
	.w4(32'hbb900d6a),
	.w5(32'h3a02ee5d),
	.w6(32'hbb191e17),
	.w7(32'h3ba78633),
	.w8(32'h3c048505),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaada9),
	.w1(32'hbc531b47),
	.w2(32'hbb1e456d),
	.w3(32'h3b1ce1d2),
	.w4(32'h3b1aec1f),
	.w5(32'hb7bfac40),
	.w6(32'hbb9e0ea2),
	.w7(32'h3b8be38b),
	.w8(32'hbb359857),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c363cac),
	.w1(32'hbb95bf00),
	.w2(32'hbafb5f87),
	.w3(32'hb9c97216),
	.w4(32'hb81d8a2a),
	.w5(32'hba23bfc2),
	.w6(32'hbb9103d8),
	.w7(32'h3ad394ca),
	.w8(32'hbb83ddf5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89050b),
	.w1(32'hbaa85ef2),
	.w2(32'hbb7e6402),
	.w3(32'hbb3dad80),
	.w4(32'hba8683b4),
	.w5(32'hbaac2b13),
	.w6(32'h388d5a6e),
	.w7(32'hbb38dda9),
	.w8(32'h3adf5649),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13127c),
	.w1(32'h3c0f2761),
	.w2(32'h3a33b9f2),
	.w3(32'h3ae4a318),
	.w4(32'h3b8799fe),
	.w5(32'h3a770d40),
	.w6(32'h3a904378),
	.w7(32'hbae5e906),
	.w8(32'hbb7f20d4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2d6b9),
	.w1(32'h3cda73fc),
	.w2(32'h39b414a2),
	.w3(32'hbb609739),
	.w4(32'h3bbeaa9d),
	.w5(32'h3b87b781),
	.w6(32'h3c5aae2d),
	.w7(32'hb956f924),
	.w8(32'hbc067075),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd048aa3),
	.w1(32'hbc956820),
	.w2(32'hbb8d987b),
	.w3(32'hbcb7ba1a),
	.w4(32'hbc1c91af),
	.w5(32'hbb1047ca),
	.w6(32'hbc546756),
	.w7(32'h3b784a68),
	.w8(32'hbbb1f131),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a333ffd),
	.w1(32'h3c39e0d6),
	.w2(32'hba883822),
	.w3(32'h3abca90d),
	.w4(32'h3af998b1),
	.w5(32'hbabd4e42),
	.w6(32'h3ba7de94),
	.w7(32'hbb2b626e),
	.w8(32'hbb6d3b8c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b376b),
	.w1(32'hbba5632a),
	.w2(32'h3b93ca4b),
	.w3(32'hbb378691),
	.w4(32'h3a795127),
	.w5(32'hbbe26910),
	.w6(32'hbbf3ddd5),
	.w7(32'hbba3b07b),
	.w8(32'hbad836da),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf996b),
	.w1(32'h3b350da1),
	.w2(32'h3bb1e56f),
	.w3(32'hbb890d30),
	.w4(32'h391bf0bc),
	.w5(32'h3bc02f1b),
	.w6(32'h3be46bfa),
	.w7(32'h3b16fc89),
	.w8(32'h3acaf234),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b754faa),
	.w1(32'hbaf06807),
	.w2(32'hbb46bedd),
	.w3(32'h3b5c2f30),
	.w4(32'hb8d37eb8),
	.w5(32'h39ab8265),
	.w6(32'h3992cb39),
	.w7(32'hba16f514),
	.w8(32'hba980c6b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19aac2),
	.w1(32'hbc1815cb),
	.w2(32'h3a287016),
	.w3(32'h3a37e8e1),
	.w4(32'hbc10aa56),
	.w5(32'hbc28c8f3),
	.w6(32'h3b734734),
	.w7(32'h3b2d0c46),
	.w8(32'h3bbd9e28),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4d966),
	.w1(32'hbb6085e2),
	.w2(32'hbbe2d218),
	.w3(32'hbadd5364),
	.w4(32'hba050e61),
	.w5(32'hbba038ef),
	.w6(32'hbb7a3b06),
	.w7(32'hbbbf2427),
	.w8(32'hba83c9ce),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42e3d2),
	.w1(32'h3b22bf53),
	.w2(32'hbb533837),
	.w3(32'h3b5e720d),
	.w4(32'h3a85a41f),
	.w5(32'hbb47c7a6),
	.w6(32'h3a3fcff1),
	.w7(32'hbc2ff63f),
	.w8(32'h3ae09a0c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb64b4a),
	.w1(32'h3b19b19f),
	.w2(32'hbade1965),
	.w3(32'h3b100197),
	.w4(32'hba375083),
	.w5(32'h395af13a),
	.w6(32'h3aa93056),
	.w7(32'hba5f1a5b),
	.w8(32'hbb0b9871),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ff5c7),
	.w1(32'hba7d68da),
	.w2(32'hbb8d1c1b),
	.w3(32'hbb1220af),
	.w4(32'hba73f214),
	.w5(32'hbb013b22),
	.w6(32'h3a6a121a),
	.w7(32'hbae1a643),
	.w8(32'hbb53c105),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc094cb1),
	.w1(32'hbc4346a9),
	.w2(32'hbc84633b),
	.w3(32'hbb135bf4),
	.w4(32'hbc0426b8),
	.w5(32'hbbfcf58a),
	.w6(32'hbb9dfd1a),
	.w7(32'hbc3046fb),
	.w8(32'hbb7b23d6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a718),
	.w1(32'hbcb19b3d),
	.w2(32'hbcf8c47e),
	.w3(32'hba57f0cc),
	.w4(32'hbc12df66),
	.w5(32'hbcb2a3ea),
	.w6(32'hbbf7385c),
	.w7(32'hbc8b2d63),
	.w8(32'hbbce2df1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba069372),
	.w1(32'hbcc0dd70),
	.w2(32'h3afd27fc),
	.w3(32'hbab05685),
	.w4(32'hbbd30b2a),
	.w5(32'hbba7ab21),
	.w6(32'hbc031098),
	.w7(32'hba7c828e),
	.w8(32'hb876ce4a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84407a),
	.w1(32'hbbcbd538),
	.w2(32'hbc1e4407),
	.w3(32'hbac50369),
	.w4(32'hbbb98281),
	.w5(32'hbbb63548),
	.w6(32'hbb727573),
	.w7(32'hbaa8d84d),
	.w8(32'hbb3ecb04),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23c917),
	.w1(32'hbcbc9df4),
	.w2(32'hba855400),
	.w3(32'hbad7bdd9),
	.w4(32'hbbc62a5c),
	.w5(32'h3b1d3145),
	.w6(32'hbc61caac),
	.w7(32'h3c075a61),
	.w8(32'hb9c2c74a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4decd),
	.w1(32'hbbea96db),
	.w2(32'h3b20a5f5),
	.w3(32'hba85bd4c),
	.w4(32'h3adb89de),
	.w5(32'h3bbf156f),
	.w6(32'hbbd3517a),
	.w7(32'hb8bfb239),
	.w8(32'hbb5d2c5d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb41f8e),
	.w1(32'h3b0b9d48),
	.w2(32'hba636cd2),
	.w3(32'hbb0e7ec8),
	.w4(32'hbb52abbe),
	.w5(32'hbb3b9156),
	.w6(32'h3b86570e),
	.w7(32'hbae7c4f9),
	.w8(32'h3a8becea),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e1212),
	.w1(32'hbbc87891),
	.w2(32'hba693ff8),
	.w3(32'h3ae7cda3),
	.w4(32'hbb1bbb58),
	.w5(32'h3a6f6aa6),
	.w6(32'hbbbb0ab6),
	.w7(32'h3ad98438),
	.w8(32'hb9909700),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf392c),
	.w1(32'h3baa8b32),
	.w2(32'hbb917358),
	.w3(32'hbb2308fc),
	.w4(32'h3b3f2598),
	.w5(32'hbb9f7e32),
	.w6(32'h38297236),
	.w7(32'hbbe21737),
	.w8(32'hbacd4798),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9717ff),
	.w1(32'hbbdaa8b5),
	.w2(32'hbbef43ce),
	.w3(32'hbbadf66f),
	.w4(32'hbb629a8a),
	.w5(32'hbc1cda8e),
	.w6(32'hbb1e87b4),
	.w7(32'h3aa0f2e4),
	.w8(32'hbbd498d0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaef732),
	.w1(32'h3a0fd1b1),
	.w2(32'hb8b586a8),
	.w3(32'hbc03195e),
	.w4(32'h39b017df),
	.w5(32'h3a169295),
	.w6(32'h3b060345),
	.w7(32'h3b3f823c),
	.w8(32'hbb56668b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d5a57),
	.w1(32'hbbe400f5),
	.w2(32'hbb7c6995),
	.w3(32'hbbc97c5f),
	.w4(32'h3b7df5e1),
	.w5(32'hbbadd977),
	.w6(32'hbb8b276e),
	.w7(32'hbb4d1bec),
	.w8(32'hbb6ce195),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c460365),
	.w1(32'h3c4626e8),
	.w2(32'h3bf03140),
	.w3(32'hba720322),
	.w4(32'h3b259d11),
	.w5(32'hbbe836bd),
	.w6(32'h3bbb91f1),
	.w7(32'hbc20fe9e),
	.w8(32'hbc53c474),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7ba9e),
	.w1(32'h3bdef1b9),
	.w2(32'hbc357d4f),
	.w3(32'hbbd13d10),
	.w4(32'h398f9cb2),
	.w5(32'hbb384445),
	.w6(32'hbb60b57d),
	.w7(32'hbb9c0dce),
	.w8(32'hbba8ed22),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36c511),
	.w1(32'hbc465859),
	.w2(32'hbc1ddfae),
	.w3(32'hbbc81611),
	.w4(32'h3b0d35af),
	.w5(32'hbba0bb96),
	.w6(32'hbbadb5d7),
	.w7(32'h3c247640),
	.w8(32'h3b08a97c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b420939),
	.w1(32'hbb32f33a),
	.w2(32'hbbf891c8),
	.w3(32'hbc4670e9),
	.w4(32'hba1143af),
	.w5(32'hbbe43523),
	.w6(32'hbbc3d300),
	.w7(32'hbae86583),
	.w8(32'hbc0657bd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d4182),
	.w1(32'hbbb6719b),
	.w2(32'hbb716b66),
	.w3(32'h3b698a2a),
	.w4(32'hbb290ca6),
	.w5(32'hba97614d),
	.w6(32'hbaa41d07),
	.w7(32'h3af14194),
	.w8(32'hb989dfbe),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1ba4d),
	.w1(32'h3cb79dcf),
	.w2(32'hb969312f),
	.w3(32'hbb37802a),
	.w4(32'h3ba57886),
	.w5(32'hbae01c91),
	.w6(32'h3c45c469),
	.w7(32'hba478846),
	.w8(32'hbbec7f0f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc952f67),
	.w1(32'h3cc16ff8),
	.w2(32'hbc287b98),
	.w3(32'hbc0a2400),
	.w4(32'h3c296136),
	.w5(32'hba88397c),
	.w6(32'h3bf20b0b),
	.w7(32'hbbb3eabd),
	.w8(32'hbc0aaa29),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93e37c),
	.w1(32'hbc8bf499),
	.w2(32'h3d5d9644),
	.w3(32'hbc172ce7),
	.w4(32'hbc7929c1),
	.w5(32'hbcc41270),
	.w6(32'hbc2fa356),
	.w7(32'hbc4bad4f),
	.w8(32'hbc441320),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29c357),
	.w1(32'hbc658ed0),
	.w2(32'h3c36a7eb),
	.w3(32'hbc8db549),
	.w4(32'hbaa4b148),
	.w5(32'h3b91dd76),
	.w6(32'hbc08edc7),
	.w7(32'h3b82099d),
	.w8(32'h3c069d10),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c154cdc),
	.w1(32'hbccff870),
	.w2(32'hbcb4e4fe),
	.w3(32'h3bbbe3e0),
	.w4(32'hbcbe5767),
	.w5(32'hbc3a9a51),
	.w6(32'hbcb879e5),
	.w7(32'hbc3d0878),
	.w8(32'hbc105f27),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c137254),
	.w1(32'hbc6a7d54),
	.w2(32'h3c1d368a),
	.w3(32'hbba50ba7),
	.w4(32'hba9e33ba),
	.w5(32'h3bf7598d),
	.w6(32'hbb91eb45),
	.w7(32'h3c01833d),
	.w8(32'h3b8430db),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8c663),
	.w1(32'hbb70f72a),
	.w2(32'hbb51b972),
	.w3(32'h3a86c7ff),
	.w4(32'hbb72da97),
	.w5(32'hba86ad3d),
	.w6(32'hbb1b8336),
	.w7(32'hbb9cca7e),
	.w8(32'hbc207cca),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d4e1e),
	.w1(32'h3c7594b0),
	.w2(32'h3ba397e9),
	.w3(32'hbc171dea),
	.w4(32'h3bcb5ada),
	.w5(32'h399f0d40),
	.w6(32'h3bc676db),
	.w7(32'h3aa28911),
	.w8(32'hbc23752a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85583f),
	.w1(32'hbc182230),
	.w2(32'hbcf8f872),
	.w3(32'hbc36ac0e),
	.w4(32'hbcc92383),
	.w5(32'hbc9e85d7),
	.w6(32'hbc89e946),
	.w7(32'hbc479791),
	.w8(32'hbcea7a9c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf8648a),
	.w1(32'hbc1bc390),
	.w2(32'h3b59eb40),
	.w3(32'hbcdb9375),
	.w4(32'hba9d1eff),
	.w5(32'hbae5baa3),
	.w6(32'hbbbf1df9),
	.w7(32'hbaed80ed),
	.w8(32'hbb6ee14a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39722802),
	.w1(32'h3ba1cf13),
	.w2(32'h3afdc526),
	.w3(32'hbb60a8d8),
	.w4(32'hbace99af),
	.w5(32'hbac7ba2e),
	.w6(32'h3b76a921),
	.w7(32'hba7184ab),
	.w8(32'hb863e348),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ae35c),
	.w1(32'hbba6fc54),
	.w2(32'h3a30159b),
	.w3(32'hba9fd8b2),
	.w4(32'h3ac609ef),
	.w5(32'h3a24a8e6),
	.w6(32'hbb1098e1),
	.w7(32'h3b807234),
	.w8(32'hbb0d6a76),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0797c6),
	.w1(32'h3c48be54),
	.w2(32'h3b011af6),
	.w3(32'hbba2b12a),
	.w4(32'h3a6fa761),
	.w5(32'hba4cfd49),
	.w6(32'h3c0830da),
	.w7(32'hb807c2c8),
	.w8(32'hbbe13eaa),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f57d2),
	.w1(32'hbc0362e0),
	.w2(32'hbcded9d6),
	.w3(32'hbb1c9509),
	.w4(32'hbaff9527),
	.w5(32'hbcbaad4a),
	.w6(32'hba99115e),
	.w7(32'hbcba52d5),
	.w8(32'hbb017e7a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82cf0a),
	.w1(32'hbc18d834),
	.w2(32'h3a5c9650),
	.w3(32'hbb433b1e),
	.w4(32'h39cc2b59),
	.w5(32'hbb240d95),
	.w6(32'hbb9dad26),
	.w7(32'hba860570),
	.w8(32'h3b06f381),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ca934),
	.w1(32'h3a2b9bee),
	.w2(32'h3b4a4e1f),
	.w3(32'h383c4bcf),
	.w4(32'h3c10a2e5),
	.w5(32'h3bf45d71),
	.w6(32'h3b9f3ae9),
	.w7(32'h3c088d37),
	.w8(32'h3af4f63d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a9e95),
	.w1(32'h3c19ebb8),
	.w2(32'hbcc4e6c7),
	.w3(32'h3ba6835e),
	.w4(32'hbbd91816),
	.w5(32'hbc20839e),
	.w6(32'hbbd97863),
	.w7(32'hbc30eb30),
	.w8(32'hbc5d485b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f987f),
	.w1(32'hbbd532a0),
	.w2(32'hbc213c8b),
	.w3(32'hbc89ae1f),
	.w4(32'hbb666850),
	.w5(32'hbb720d76),
	.w6(32'hbc0ae1d7),
	.w7(32'hbbdc2342),
	.w8(32'hbbcfe46d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e45d8),
	.w1(32'hbc0bb22b),
	.w2(32'h3aa7d7db),
	.w3(32'hbb54e4a3),
	.w4(32'hbb798f67),
	.w5(32'hba1c4df3),
	.w6(32'hbc3c3315),
	.w7(32'hbbb010dc),
	.w8(32'hbbfc5b1c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf55238),
	.w1(32'hbb1d17e4),
	.w2(32'h39610acf),
	.w3(32'hbbb64a84),
	.w4(32'h3aa46080),
	.w5(32'hbb85adb9),
	.w6(32'hbb0c89ba),
	.w7(32'h3a735323),
	.w8(32'hbb742a84),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a338379),
	.w1(32'h3d262854),
	.w2(32'hbcd770a1),
	.w3(32'h3b0466d9),
	.w4(32'h3c542de1),
	.w5(32'hbb787915),
	.w6(32'h3c2d8db3),
	.w7(32'hbbc7df6c),
	.w8(32'hbc9b4140),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcedadea),
	.w1(32'hbc36b70a),
	.w2(32'h3b59c370),
	.w3(32'hbc993f62),
	.w4(32'hb8d4d2a4),
	.w5(32'hbac88180),
	.w6(32'hbbc653cb),
	.w7(32'hbb1f9a22),
	.w8(32'hba4e4a93),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00c925),
	.w1(32'h3bb31dd5),
	.w2(32'hbbf3e68f),
	.w3(32'hbb2e53dc),
	.w4(32'h39bb9a42),
	.w5(32'hbb86ac72),
	.w6(32'h3b508ac2),
	.w7(32'hbaa064b7),
	.w8(32'hba46fde7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d6f39),
	.w1(32'h3b26dd74),
	.w2(32'h3b18dd1e),
	.w3(32'hba08661d),
	.w4(32'hbab70a4a),
	.w5(32'hb9ef3660),
	.w6(32'h3ae4f2c5),
	.w7(32'h3a5f4a75),
	.w8(32'h3b1f573a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb680b9c),
	.w1(32'hbafb2e3f),
	.w2(32'hbb6e19cf),
	.w3(32'h3ab0cacf),
	.w4(32'hbac1e25d),
	.w5(32'hbab17bb7),
	.w6(32'hba35277a),
	.w7(32'hb9ce842f),
	.w8(32'hbb36d752),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe30987),
	.w1(32'hbbf6bacb),
	.w2(32'h3c007a40),
	.w3(32'hbb1b6b3a),
	.w4(32'h3af4e41b),
	.w5(32'hbaf58094),
	.w6(32'hbae2710c),
	.w7(32'h3b3103c5),
	.w8(32'hbb6b6877),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388546e7),
	.w1(32'hbc1e4fa1),
	.w2(32'hbb6db424),
	.w3(32'hbbc773c9),
	.w4(32'hb9b363f3),
	.w5(32'hbc4f4e99),
	.w6(32'hbb443ad1),
	.w7(32'hbb3c4607),
	.w8(32'hbc53f90e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbea72e),
	.w1(32'h3c9f5323),
	.w2(32'hbc1f232d),
	.w3(32'hbcb84f87),
	.w4(32'h3b458fa9),
	.w5(32'hbb674ea5),
	.w6(32'h3c17a28d),
	.w7(32'hbb6560c9),
	.w8(32'hbbeb36e3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84e2b2),
	.w1(32'hbaaf0b8e),
	.w2(32'hbc6d9e64),
	.w3(32'hbb333e5b),
	.w4(32'h3b9a847f),
	.w5(32'hbc34b63e),
	.w6(32'h39adf738),
	.w7(32'hbc841b8d),
	.w8(32'hbc171014),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc087c53),
	.w1(32'hbc4e7cbd),
	.w2(32'h3c8ef34f),
	.w3(32'hbc068d9b),
	.w4(32'hba48e8ef),
	.w5(32'h3c9bb6f5),
	.w6(32'hbba710fe),
	.w7(32'h3c79d9f8),
	.w8(32'h3bf5ca23),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58e796),
	.w1(32'h3aebbf77),
	.w2(32'hbbb1fb7c),
	.w3(32'h3aeac265),
	.w4(32'hba0aa86c),
	.w5(32'h3a443380),
	.w6(32'hba6e5fd1),
	.w7(32'hbb0475f1),
	.w8(32'hbb40bb7c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdceeaf),
	.w1(32'hbba94cc7),
	.w2(32'h3acfdb9e),
	.w3(32'hbb6519b3),
	.w4(32'hbb5d959b),
	.w5(32'h39c9846d),
	.w6(32'hbc05a839),
	.w7(32'hbb09e0a3),
	.w8(32'hbb8a91c3),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82cef5),
	.w1(32'hbc0e6b10),
	.w2(32'hbb200b15),
	.w3(32'hbb96c7de),
	.w4(32'hbb13067a),
	.w5(32'hbb7c28ed),
	.w6(32'hbbb41159),
	.w7(32'hbaa665bb),
	.w8(32'hbbb40c7c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf1c7a),
	.w1(32'hbb193977),
	.w2(32'hbb797ef8),
	.w3(32'hbbca8a06),
	.w4(32'hbace858a),
	.w5(32'hbc3dae77),
	.w6(32'hbb5122ef),
	.w7(32'hbbaf106b),
	.w8(32'hbbd3af83),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd9562),
	.w1(32'hbbdf92dd),
	.w2(32'h3bbf3dc3),
	.w3(32'hbc03570c),
	.w4(32'h395030aa),
	.w5(32'h3b61a014),
	.w6(32'hbb374dbb),
	.w7(32'h3b1ab690),
	.w8(32'hbb6eaf50),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae68271),
	.w1(32'hbb3e859a),
	.w2(32'hbba8e10a),
	.w3(32'hba2ddff5),
	.w4(32'h3b0f8a5f),
	.w5(32'hb94554c0),
	.w6(32'hbb077952),
	.w7(32'h3a148887),
	.w8(32'h3b623c6b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5799ce),
	.w1(32'h3bb0041a),
	.w2(32'h3bb8ab2d),
	.w3(32'h3ba5f2ad),
	.w4(32'h3bdf7502),
	.w5(32'h3bc6dead),
	.w6(32'h3b847d16),
	.w7(32'h3b3c1e03),
	.w8(32'hbafc4470),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6e5b3),
	.w1(32'h3bf0f444),
	.w2(32'hbc10c4ca),
	.w3(32'hbaad2790),
	.w4(32'h3aaa5e63),
	.w5(32'hbc5ec573),
	.w6(32'hbb3fd76a),
	.w7(32'hbc8f70b4),
	.w8(32'hbca6f307),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae806e),
	.w1(32'h3b918e3f),
	.w2(32'h3a846bed),
	.w3(32'hbc79a49d),
	.w4(32'h3af1529c),
	.w5(32'h3add1b9c),
	.w6(32'h3b01b6d7),
	.w7(32'h398b0d08),
	.w8(32'hba9dd29d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae117f),
	.w1(32'hbc8c0f97),
	.w2(32'h3bd89ae5),
	.w3(32'hbb123451),
	.w4(32'hbb9905d2),
	.w5(32'h3b9ef504),
	.w6(32'hbc17e2e3),
	.w7(32'h3b248d06),
	.w8(32'h3ab65171),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b041a82),
	.w1(32'h3ae6233f),
	.w2(32'hbc0fe487),
	.w3(32'hbb95fb50),
	.w4(32'h3a2ec9c6),
	.w5(32'hbb4f419a),
	.w6(32'hba8d844b),
	.w7(32'hbb8adf6b),
	.w8(32'hbc241521),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed6b1),
	.w1(32'h3b8d072d),
	.w2(32'h3ac71dea),
	.w3(32'hbb8fa616),
	.w4(32'hb9d2cd9e),
	.w5(32'hb988e0aa),
	.w6(32'h3b590202),
	.w7(32'h399dee7f),
	.w8(32'hbb4221ae),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe78538),
	.w1(32'hbafd3df1),
	.w2(32'hbb53bb35),
	.w3(32'hbb13c17e),
	.w4(32'h3beabf65),
	.w5(32'h3acc7799),
	.w6(32'hbb132396),
	.w7(32'h3ac06efd),
	.w8(32'hbb8f94ab),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6436b9),
	.w1(32'hbc89ecdd),
	.w2(32'h3c380769),
	.w3(32'hbb866b2c),
	.w4(32'hbb53eed9),
	.w5(32'h3b9875a8),
	.w6(32'hbc295eab),
	.w7(32'h3b404a3b),
	.w8(32'h3b32a184),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1baedb),
	.w1(32'hbc32b59d),
	.w2(32'hbba14ff2),
	.w3(32'hbb78d033),
	.w4(32'hbbe66409),
	.w5(32'h3a82964b),
	.w6(32'hbc704bab),
	.w7(32'hbb7e94ba),
	.w8(32'hbb6bfe26),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd69ac),
	.w1(32'hbb211b53),
	.w2(32'h398b8209),
	.w3(32'hbb85491e),
	.w4(32'hbb306531),
	.w5(32'h3a4d4c30),
	.w6(32'hbb184c55),
	.w7(32'h37f1da16),
	.w8(32'h3a2f3eb2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1be2a1),
	.w1(32'hbca81ba9),
	.w2(32'hbc121f0c),
	.w3(32'h3aa75b55),
	.w4(32'hbc8289f4),
	.w5(32'hbaf58676),
	.w6(32'hbc27eb07),
	.w7(32'hbc0e4045),
	.w8(32'h39c3efa2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c621c4d),
	.w1(32'hbbbe7cf6),
	.w2(32'h3b7a5ab4),
	.w3(32'h3c46b1ac),
	.w4(32'hba8203cd),
	.w5(32'h3b18994a),
	.w6(32'hbb8b35f0),
	.w7(32'h3b53f267),
	.w8(32'h3bcc47d2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ef7c9),
	.w1(32'hbc15d891),
	.w2(32'hbc1b00fb),
	.w3(32'h3bcb852e),
	.w4(32'hbc0eee0b),
	.w5(32'hbcc00043),
	.w6(32'hbb28ad76),
	.w7(32'hbc7a1c1c),
	.w8(32'hbba72791),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3091b2),
	.w1(32'hbc14429a),
	.w2(32'h3a30d76d),
	.w3(32'h3ba83dd8),
	.w4(32'hbb5b3dc7),
	.w5(32'hbb3bdaaa),
	.w6(32'hbbaff79a),
	.w7(32'h3b01c66a),
	.w8(32'hbb8ac7fd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da47f2),
	.w1(32'hbccd6c3a),
	.w2(32'h3b550afe),
	.w3(32'hbbf64d41),
	.w4(32'hbb942e73),
	.w5(32'hbb13424b),
	.w6(32'hbc86a5ba),
	.w7(32'hb9195ecc),
	.w8(32'h3af2031b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57ccf6),
	.w1(32'h3c3c4a3d),
	.w2(32'hbc74e805),
	.w3(32'h3a52c5ca),
	.w4(32'hb80093fc),
	.w5(32'h3c3d8dcb),
	.w6(32'hbb605be7),
	.w7(32'h3b860ba0),
	.w8(32'hbc30c95b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc6b3f),
	.w1(32'h38dc4a59),
	.w2(32'hbced7fb9),
	.w3(32'hbbd90cbe),
	.w4(32'hbc297f30),
	.w5(32'hbb0667fd),
	.w6(32'hbae053d4),
	.w7(32'hbc510321),
	.w8(32'hbc458216),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d5757),
	.w1(32'h3d06317f),
	.w2(32'hbc44e3a8),
	.w3(32'hbb77be5f),
	.w4(32'h3c03aeb7),
	.w5(32'hbbb8c90d),
	.w6(32'h3ca27688),
	.w7(32'hbabee474),
	.w8(32'hbc2c48c3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccf2b29),
	.w1(32'h3b737530),
	.w2(32'hbc17c8a3),
	.w3(32'hbbd55d40),
	.w4(32'hba9e815d),
	.w5(32'hbb4802f8),
	.w6(32'h3b0bedd0),
	.w7(32'h3a66c3cd),
	.w8(32'hb9ec453d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50f5c5),
	.w1(32'h3bdc03a8),
	.w2(32'hbc1b57fd),
	.w3(32'hbbc1c76b),
	.w4(32'h3b9cadeb),
	.w5(32'hbb4a9945),
	.w6(32'h3b69f2ab),
	.w7(32'h3aac7651),
	.w8(32'hbba15f49),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012cb4),
	.w1(32'hbb106133),
	.w2(32'hbb8e0eb1),
	.w3(32'h39bd5a83),
	.w4(32'hbb51638d),
	.w5(32'hbb568871),
	.w6(32'hb9bf0cec),
	.w7(32'hbb1379d9),
	.w8(32'hbb784c35),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4488e6),
	.w1(32'hbadc8b03),
	.w2(32'h3b456cd9),
	.w3(32'hb874fdbd),
	.w4(32'h3b0bd8da),
	.w5(32'h3b2790c4),
	.w6(32'h3acffea3),
	.w7(32'h3abbdd7a),
	.w8(32'hb81abca6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385ec979),
	.w1(32'h3b184734),
	.w2(32'h3b7a1ac4),
	.w3(32'hbb315bfe),
	.w4(32'hbb11f3eb),
	.w5(32'h3af3292b),
	.w6(32'h3916f402),
	.w7(32'hba151b38),
	.w8(32'hbb434ba2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb422a17),
	.w1(32'h3cabed8c),
	.w2(32'hbbc12a7c),
	.w3(32'h39fd6854),
	.w4(32'h3be6e191),
	.w5(32'hba808279),
	.w6(32'h3c395080),
	.w7(32'hba164c2f),
	.w8(32'hbbbfca01),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b658a),
	.w1(32'h3bd56aa8),
	.w2(32'h3bfa3cd8),
	.w3(32'hbb314e0a),
	.w4(32'h3bcdfb2b),
	.w5(32'hbaf0e722),
	.w6(32'h3b569a33),
	.w7(32'hbc138d00),
	.w8(32'hbc205290),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5290e6),
	.w1(32'hbb813e74),
	.w2(32'h3c574581),
	.w3(32'hbb2e9ac0),
	.w4(32'hba9ff90d),
	.w5(32'h3b1a8254),
	.w6(32'hbad9ed12),
	.w7(32'h3b0a52a7),
	.w8(32'h3b8bdf3c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb913e5f5),
	.w1(32'hba1a764a),
	.w2(32'h3c9718a0),
	.w3(32'h3a38bf07),
	.w4(32'hbbd6dcbb),
	.w5(32'hbd01f834),
	.w6(32'hbba927f0),
	.w7(32'hbd1ccb87),
	.w8(32'hbcb74ff5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96057c),
	.w1(32'hbbb9a02f),
	.w2(32'h3bd9242e),
	.w3(32'hbc7e45b3),
	.w4(32'hbb4c04bf),
	.w5(32'h3add8d8a),
	.w6(32'hbb8790fe),
	.w7(32'h3b5a751b),
	.w8(32'h3bbd1660),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f6788),
	.w1(32'hbbb0f661),
	.w2(32'hbc3af699),
	.w3(32'hba92979a),
	.w4(32'hbb40b959),
	.w5(32'hbbe11a91),
	.w6(32'hbba957eb),
	.w7(32'hbbc56c10),
	.w8(32'hbb73f8b3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e7c95),
	.w1(32'h3c910d07),
	.w2(32'h3bea0113),
	.w3(32'hbbca248f),
	.w4(32'h3b040b5e),
	.w5(32'hbbb2a8c1),
	.w6(32'h3b2bcd10),
	.w7(32'hbad96718),
	.w8(32'hbc9c4efb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce3b819),
	.w1(32'h3cde3817),
	.w2(32'hbba51140),
	.w3(32'hbca5284f),
	.w4(32'h3bfe5243),
	.w5(32'hba032027),
	.w6(32'h3c8294e1),
	.w7(32'hb888ef34),
	.w8(32'hbb7d78f9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97c3f6),
	.w1(32'h3c0677da),
	.w2(32'hbb2ffc62),
	.w3(32'hbb9c35e4),
	.w4(32'h3ae71a25),
	.w5(32'h3a880d91),
	.w6(32'h3bb4dec3),
	.w7(32'h3a88e8bc),
	.w8(32'h3a9ae391),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50cd48),
	.w1(32'h3bca6ca7),
	.w2(32'hbb26e3f6),
	.w3(32'h3b0855db),
	.w4(32'h3a9e9358),
	.w5(32'h3aacb5f7),
	.w6(32'h3bb4eeab),
	.w7(32'h3b141065),
	.w8(32'h3b592f94),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39922ebc),
	.w1(32'h3bcf4392),
	.w2(32'h3ac25227),
	.w3(32'h3b8c51fd),
	.w4(32'hbc1b0cb4),
	.w5(32'hbba5c1f2),
	.w6(32'h3c03d5fa),
	.w7(32'hbb834391),
	.w8(32'hbc74ff68),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8eb646),
	.w1(32'h3a2bd105),
	.w2(32'hbb937c8c),
	.w3(32'hbbf20abb),
	.w4(32'h3a25ea27),
	.w5(32'h3b82809b),
	.w6(32'hbbe336a2),
	.w7(32'h3ab67589),
	.w8(32'hbb3940c5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc2388),
	.w1(32'hbc392983),
	.w2(32'hbbcc3bcd),
	.w3(32'hbb596ee3),
	.w4(32'hbc4df421),
	.w5(32'hbb936795),
	.w6(32'hbc0c1a6e),
	.w7(32'h3ad4f5e1),
	.w8(32'h3c13ae16),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b56fc),
	.w1(32'hbbe1df8f),
	.w2(32'hbb58c232),
	.w3(32'h3bae093f),
	.w4(32'hbba061c9),
	.w5(32'hbbb0de66),
	.w6(32'hbbe6be67),
	.w7(32'hbbd06e57),
	.w8(32'h3bb7f0cd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1457c),
	.w1(32'h3c178cef),
	.w2(32'h38e4ff20),
	.w3(32'h3bb7381a),
	.w4(32'h39c3c499),
	.w5(32'hb79526fa),
	.w6(32'h3b923876),
	.w7(32'hbb2ab8e5),
	.w8(32'hbb1d2ac4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25bc89),
	.w1(32'hbc41371b),
	.w2(32'hbc712f72),
	.w3(32'hba9f2508),
	.w4(32'hbbfd51a3),
	.w5(32'h3b1b34c9),
	.w6(32'hbb2c2250),
	.w7(32'hbbf9d767),
	.w8(32'hbc3b3023),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a71d9),
	.w1(32'hbca30e99),
	.w2(32'h3b6b4888),
	.w3(32'h3a85d46c),
	.w4(32'hbb5da85f),
	.w5(32'h3c1274dd),
	.w6(32'hbc297c80),
	.w7(32'h3ae8e9aa),
	.w8(32'h3c66d717),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce5198f),
	.w1(32'h3b16a524),
	.w2(32'hb91433d3),
	.w3(32'h3c78a100),
	.w4(32'h3b25f716),
	.w5(32'h3aac146f),
	.w6(32'h3a851e1f),
	.w7(32'h39b7b04c),
	.w8(32'h3b0d4303),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d2253),
	.w1(32'h398d44ea),
	.w2(32'hb774e683),
	.w3(32'h3aece317),
	.w4(32'h39026e73),
	.w5(32'hb93d1ad9),
	.w6(32'h39085fbe),
	.w7(32'h3844a56f),
	.w8(32'hb90ed944),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab88eb4),
	.w1(32'hbbb500ed),
	.w2(32'hbbbaa149),
	.w3(32'h39573484),
	.w4(32'hbba7762e),
	.w5(32'hbba89336),
	.w6(32'hbad4e1d3),
	.w7(32'hbb844942),
	.w8(32'hbb78bbb7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45f4f5),
	.w1(32'h382f6c0a),
	.w2(32'hbb3b5892),
	.w3(32'hb8b973a5),
	.w4(32'hba3b292d),
	.w5(32'hba9b8649),
	.w6(32'hb9bfbdb7),
	.w7(32'h39c1d26b),
	.w8(32'hbab03d74),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a456e9),
	.w1(32'hba3e8ab3),
	.w2(32'hba61165f),
	.w3(32'h38b7ea1b),
	.w4(32'hb94dde1a),
	.w5(32'hba023710),
	.w6(32'hba1d5129),
	.w7(32'hba0882bd),
	.w8(32'hba450ccd),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04f511),
	.w1(32'hbb0cd3f8),
	.w2(32'hbad3ff64),
	.w3(32'hba30bea2),
	.w4(32'hba014f42),
	.w5(32'hba1c2e35),
	.w6(32'hbae7480c),
	.w7(32'hbac98b93),
	.w8(32'hbaaf461b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f1ef06),
	.w1(32'h39a15649),
	.w2(32'h39ef74c3),
	.w3(32'h3a16b41c),
	.w4(32'h3a90785a),
	.w5(32'h3a814098),
	.w6(32'h388c9ed0),
	.w7(32'hb90f07ad),
	.w8(32'hb99e5884),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c7123),
	.w1(32'hb9ca4c79),
	.w2(32'hbae53690),
	.w3(32'hb9a54d64),
	.w4(32'h39a416dd),
	.w5(32'hb9321109),
	.w6(32'hbaaa6a2e),
	.w7(32'hb9a43288),
	.w8(32'hba0190b3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb299d7c),
	.w1(32'hbb0d9410),
	.w2(32'hbb19c905),
	.w3(32'hba62a04d),
	.w4(32'h3820ba8a),
	.w5(32'h3a1d2961),
	.w6(32'hb95c0cac),
	.w7(32'hb9a6f514),
	.w8(32'hb9ca8394),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb040828),
	.w1(32'hbb2aa73e),
	.w2(32'hbbaebebf),
	.w3(32'hba81f67e),
	.w4(32'hbb14ec04),
	.w5(32'hbb751e49),
	.w6(32'hbb18f88c),
	.w7(32'hbb00015d),
	.w8(32'hbb9d26a1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba408c21),
	.w1(32'h3a0c7f6a),
	.w2(32'h3a8edc27),
	.w3(32'h38f009c9),
	.w4(32'h3ad749ce),
	.w5(32'h3ad77b26),
	.w6(32'hb822625b),
	.w7(32'h39afb17a),
	.w8(32'h398c1c9f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba719f2a),
	.w1(32'hba7d198f),
	.w2(32'hbae3293f),
	.w3(32'hb9b85329),
	.w4(32'hb868fa4d),
	.w5(32'hb973287c),
	.w6(32'hbac42bb7),
	.w7(32'hb9042675),
	.w8(32'hbab2b870),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3fa2a),
	.w1(32'hbaf8a92c),
	.w2(32'hbb8f5634),
	.w3(32'h390cb52a),
	.w4(32'hba8cadb2),
	.w5(32'hbb3cb7fb),
	.w6(32'hba41ce24),
	.w7(32'hbac04f20),
	.w8(32'hbb6cd5e8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a433f),
	.w1(32'h398f3eba),
	.w2(32'h3ab46e35),
	.w3(32'hb9cdfc06),
	.w4(32'h3aa4314a),
	.w5(32'h3aea7883),
	.w6(32'hbae2a394),
	.w7(32'hb944c459),
	.w8(32'hb88bca54),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b50aa),
	.w1(32'hba5dbf25),
	.w2(32'hbab238bc),
	.w3(32'hb8de93de),
	.w4(32'hba81252b),
	.w5(32'hbac29188),
	.w6(32'hbad3f9c2),
	.w7(32'hbad67d1d),
	.w8(32'hbb017364),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387a3e06),
	.w1(32'h384115e6),
	.w2(32'hb906ff93),
	.w3(32'h38f04473),
	.w4(32'h394052dc),
	.w5(32'h385cff4d),
	.w6(32'hb98fb665),
	.w7(32'hb8e96014),
	.w8(32'hb9db9267),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af51c37),
	.w1(32'h3a63c211),
	.w2(32'h3b7e2873),
	.w3(32'h3b1a0442),
	.w4(32'hb941f6de),
	.w5(32'h3b21d1f1),
	.w6(32'h3a868ad9),
	.w7(32'hbb197364),
	.w8(32'h399cebb2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad42030),
	.w1(32'hbaadaeaa),
	.w2(32'hb9a0cd7a),
	.w3(32'hba5daa80),
	.w4(32'hb999c84f),
	.w5(32'hb87f55ac),
	.w6(32'hbaea1d3b),
	.w7(32'hba4794a7),
	.w8(32'hba0c7e18),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e882e),
	.w1(32'h37440eab),
	.w2(32'hb8fffac9),
	.w3(32'h38c8b0b5),
	.w4(32'h3913d45f),
	.w5(32'h37ca144b),
	.w6(32'h37ece30d),
	.w7(32'h38a4e269),
	.w8(32'h38f710b8),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38306668),
	.w1(32'h39a0688e),
	.w2(32'h38ccd365),
	.w3(32'h3815a171),
	.w4(32'h38a024be),
	.w5(32'h384d5d29),
	.w6(32'h3998d7a4),
	.w7(32'h396e48c4),
	.w8(32'h393d73e6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d97b20),
	.w1(32'h38e87b5a),
	.w2(32'hb91aaff3),
	.w3(32'h39858879),
	.w4(32'hb74748d4),
	.w5(32'hb957e2a6),
	.w6(32'hba03d59d),
	.w7(32'hb90ad751),
	.w8(32'hb9292fa8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fb1e6),
	.w1(32'hba341fb1),
	.w2(32'h3a273aa9),
	.w3(32'hba69fa0f),
	.w4(32'h3ab5572f),
	.w5(32'h3afbd766),
	.w6(32'hba6a4115),
	.w7(32'hb8ae014c),
	.w8(32'hb9b671c0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c7268),
	.w1(32'hb9c72f6a),
	.w2(32'hba199130),
	.w3(32'h3a37ea12),
	.w4(32'h3a262b55),
	.w5(32'h39863745),
	.w6(32'hbaa03405),
	.w7(32'hba80aef1),
	.w8(32'hbaedd209),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3847037e),
	.w1(32'hb90a9cb4),
	.w2(32'hb9ceb99e),
	.w3(32'hb6292059),
	.w4(32'hb82fb6a8),
	.w5(32'hb96ac4b6),
	.w6(32'hb8878e1a),
	.w7(32'hb966c320),
	.w8(32'hb98a0cc5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac10845),
	.w1(32'hb9af1633),
	.w2(32'hbac44a2c),
	.w3(32'hba2fd36f),
	.w4(32'hb7ca6f00),
	.w5(32'hb9e8c1f6),
	.w6(32'hb9f80786),
	.w7(32'hba0a9a9c),
	.w8(32'hbacf369c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00fc45),
	.w1(32'h3722ab89),
	.w2(32'hba128f74),
	.w3(32'h3acdf2c0),
	.w4(32'h3a36a0c9),
	.w5(32'h39b5eb0c),
	.w6(32'hb96bcab1),
	.w7(32'hb9dabcf8),
	.w8(32'hba912eac),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf39a04),
	.w1(32'hbb005f41),
	.w2(32'hbb65070b),
	.w3(32'hba806bb7),
	.w4(32'hbb09dc06),
	.w5(32'hbb4caed7),
	.w6(32'hba3f2219),
	.w7(32'hba231eec),
	.w8(32'hbb4d2e2a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a358e1a),
	.w1(32'hba54aee8),
	.w2(32'h38f7fb43),
	.w3(32'h3ac44d42),
	.w4(32'h39b5194a),
	.w5(32'h38cc9c6d),
	.w6(32'h3af7f599),
	.w7(32'hba82aebd),
	.w8(32'hbb08aa06),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba148435),
	.w1(32'hba75c106),
	.w2(32'hba8353b1),
	.w3(32'h32d42c00),
	.w4(32'hb97e16ad),
	.w5(32'hb9acf843),
	.w6(32'hb817389b),
	.w7(32'hb9ebc5ba),
	.w8(32'hba4cfb16),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9a680),
	.w1(32'h39ac0058),
	.w2(32'h39cf9bb8),
	.w3(32'h39c8a4ae),
	.w4(32'h397a20ce),
	.w5(32'h39a75e45),
	.w6(32'h3a05d8ef),
	.w7(32'h39efd1cc),
	.w8(32'h39e0cfa5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ade0c),
	.w1(32'h3a80fb07),
	.w2(32'h3a9a5106),
	.w3(32'h3a92295c),
	.w4(32'h3aa59772),
	.w5(32'h3ad16ee6),
	.w6(32'h396d688e),
	.w7(32'h3924a8c3),
	.w8(32'hb9f348b7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba350ceb),
	.w1(32'hb9f76870),
	.w2(32'hb9dd7297),
	.w3(32'h38cf569a),
	.w4(32'h3a822bfc),
	.w5(32'h3a39c7f4),
	.w6(32'hba21bfa4),
	.w7(32'hb9bf962b),
	.w8(32'hba8c6a52),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392332bd),
	.w1(32'h3a5f4aea),
	.w2(32'h3a466e69),
	.w3(32'h395b2cbb),
	.w4(32'h3a91ae6b),
	.w5(32'h3a7ce462),
	.w6(32'hb9b12981),
	.w7(32'h37ba3640),
	.w8(32'hb8f16746),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c87b0f),
	.w1(32'hba108ad0),
	.w2(32'hbaa132b5),
	.w3(32'hb9c6af3e),
	.w4(32'hba20f2d7),
	.w5(32'hbaa37889),
	.w6(32'hb9f74986),
	.w7(32'hba0e1986),
	.w8(32'hba9a2174),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91326a3),
	.w1(32'hb8937d70),
	.w2(32'hb993bf5f),
	.w3(32'hb981b198),
	.w4(32'hb8a8e3f4),
	.w5(32'hb9da3e60),
	.w6(32'hb7d53aab),
	.w7(32'hb8a4cf29),
	.w8(32'hb919b831),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5a642),
	.w1(32'hbafd2eb6),
	.w2(32'hbb111275),
	.w3(32'hb8aa31d6),
	.w4(32'hba1ea091),
	.w5(32'hba547ced),
	.w6(32'hbaa79f57),
	.w7(32'hba492212),
	.w8(32'hba9935f4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22de93),
	.w1(32'h38d0bc27),
	.w2(32'hba802072),
	.w3(32'h39c302af),
	.w4(32'hba071901),
	.w5(32'hbab20479),
	.w6(32'h3a56b35d),
	.w7(32'hb967f0de),
	.w8(32'hba88e39f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397377ed),
	.w1(32'hb875b3f8),
	.w2(32'h3a190015),
	.w3(32'hb93a6673),
	.w4(32'h38c1453c),
	.w5(32'h39a0cf49),
	.w6(32'hba329ee0),
	.w7(32'hba4c4981),
	.w8(32'hbaa1d9ac),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e5cbf4),
	.w1(32'h38fba14e),
	.w2(32'h3910de48),
	.w3(32'hb8244850),
	.w4(32'h394ee1b7),
	.w5(32'h38b5017d),
	.w6(32'h384d815b),
	.w7(32'h39070ebb),
	.w8(32'h3929a8db),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a263e60),
	.w1(32'hba154603),
	.w2(32'hb9d074db),
	.w3(32'h3a46ea9b),
	.w4(32'hba631c6c),
	.w5(32'hba101832),
	.w6(32'h388d677d),
	.w7(32'hba932c57),
	.w8(32'hba17dcc3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392385a4),
	.w1(32'hb9372c3a),
	.w2(32'hb94499c8),
	.w3(32'h39b052f8),
	.w4(32'h39099aa2),
	.w5(32'h3946cc9d),
	.w6(32'hb7730380),
	.w7(32'hb8b65af9),
	.w8(32'hb83aefff),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92556cb),
	.w1(32'h3942ae0e),
	.w2(32'h393bf3ba),
	.w3(32'hb8dcbe2f),
	.w4(32'h39358691),
	.w5(32'h3915cbc5),
	.w6(32'h393528a1),
	.w7(32'h398bfcb6),
	.w8(32'h397bdb7b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b3635),
	.w1(32'h38fa0b1b),
	.w2(32'h38dd1a96),
	.w3(32'h3a4b0a8d),
	.w4(32'h3abdf08f),
	.w5(32'h3a9e5d5c),
	.w6(32'h3a191ed4),
	.w7(32'h3a4602ff),
	.w8(32'hb8b085fb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb055ccf),
	.w1(32'hbaf9aecb),
	.w2(32'hbb70457b),
	.w3(32'hb9ec0f1e),
	.w4(32'hba2e6e04),
	.w5(32'hbb0afc32),
	.w6(32'hbb87cba9),
	.w7(32'hbb16db76),
	.w8(32'hbb7ad203),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed5922),
	.w1(32'h3949ac99),
	.w2(32'hb6ecdefe),
	.w3(32'h3994d5ed),
	.w4(32'h39e1f5b1),
	.w5(32'h38d98bdb),
	.w6(32'hb8c6eccb),
	.w7(32'hb90fefd4),
	.w8(32'hb94f4d61),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a8ef7),
	.w1(32'h38ca4aba),
	.w2(32'hb9cfe49d),
	.w3(32'h3a483bcc),
	.w4(32'h3a1e4987),
	.w5(32'h39b82b1a),
	.w6(32'h3a189a94),
	.w7(32'hb96b212a),
	.w8(32'hbae3e87b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919532d),
	.w1(32'hba49c4c7),
	.w2(32'hbadf49b7),
	.w3(32'hba13471c),
	.w4(32'hba119a48),
	.w5(32'hba81849a),
	.w6(32'h3a194ac8),
	.w7(32'hba0a18ba),
	.w8(32'hba0cfd0a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fc843),
	.w1(32'hba187272),
	.w2(32'hbb92c367),
	.w3(32'hbab40a84),
	.w4(32'h38e55df0),
	.w5(32'hbb28bf25),
	.w6(32'hbafbf8a9),
	.w7(32'hbaf835b7),
	.w8(32'hbb6f4f48),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35476b),
	.w1(32'hbb1cd50d),
	.w2(32'hbb6e9d13),
	.w3(32'hbaa19dfd),
	.w4(32'hb9bce9bc),
	.w5(32'hba06b575),
	.w6(32'hbad8e913),
	.w7(32'hba8935ed),
	.w8(32'hbadfe39a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2f9cf),
	.w1(32'hb8b72c40),
	.w2(32'hbb0339e1),
	.w3(32'hba16eeed),
	.w4(32'hb96ef59b),
	.w5(32'hbab1c540),
	.w6(32'hbacd84ac),
	.w7(32'hba82f252),
	.w8(32'hbb2ee898),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28d7e4),
	.w1(32'hb7e4c70b),
	.w2(32'hb801c76d),
	.w3(32'h3932e999),
	.w4(32'h3973022f),
	.w5(32'h38df6f4b),
	.w6(32'h3964fe4a),
	.w7(32'h393aa343),
	.w8(32'h39ad1f1f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa73485),
	.w1(32'hbaa94cf5),
	.w2(32'hbae6238e),
	.w3(32'hba0ddb4b),
	.w4(32'hba39d1dd),
	.w5(32'hb8d5efbe),
	.w6(32'hb9db2161),
	.w7(32'hb9281d94),
	.w8(32'hba304474),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86a00dc),
	.w1(32'h397fd8b6),
	.w2(32'h3904ae18),
	.w3(32'hb891393f),
	.w4(32'h3984c523),
	.w5(32'h393d4d28),
	.w6(32'h39659c5d),
	.w7(32'h3944bb3f),
	.w8(32'h39a3a597),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a65a73),
	.w1(32'h39a1d805),
	.w2(32'h38bfb5f7),
	.w3(32'h39c10b74),
	.w4(32'h39870d5c),
	.w5(32'h391accfd),
	.w6(32'hba09aaca),
	.w7(32'hb90f4725),
	.w8(32'h3898f264),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988ea0e),
	.w1(32'h39a59941),
	.w2(32'h39f9fe1a),
	.w3(32'hba270433),
	.w4(32'h39e66484),
	.w5(32'h3a1cd455),
	.w6(32'h3919ba9a),
	.w7(32'hb6f56dce),
	.w8(32'h394e48c8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bd4a9),
	.w1(32'hbaad7e64),
	.w2(32'hbb2ec71b),
	.w3(32'hbab0cf04),
	.w4(32'h39343125),
	.w5(32'h3a1a6f78),
	.w6(32'hbaeddcc7),
	.w7(32'hb9b27f98),
	.w8(32'hb9c1ae91),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8521f),
	.w1(32'h39adcb86),
	.w2(32'hb8f2a9dd),
	.w3(32'h39bfe011),
	.w4(32'h3989825b),
	.w5(32'h371fbf3a),
	.w6(32'h39a249fc),
	.w7(32'h39bbb800),
	.w8(32'h384f07e5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cba24d),
	.w1(32'h3882e999),
	.w2(32'hb9832c46),
	.w3(32'h37848c4b),
	.w4(32'h394e6919),
	.w5(32'hb7c58a23),
	.w6(32'h386a59ff),
	.w7(32'hb86a4132),
	.w8(32'h37a4f017),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f4807),
	.w1(32'hba2c206b),
	.w2(32'hb93df282),
	.w3(32'h3a1210c3),
	.w4(32'h3a109e45),
	.w5(32'h39f31d59),
	.w6(32'h3985756e),
	.w7(32'hb9af8e55),
	.w8(32'hb9cfd716),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e41a1),
	.w1(32'hbaed4c7f),
	.w2(32'hbb7154aa),
	.w3(32'hb9e9eddc),
	.w4(32'hba913860),
	.w5(32'hbb1fc5f1),
	.w6(32'hba8581c8),
	.w7(32'hbb0c8457),
	.w8(32'hbb80fdbc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c64dc),
	.w1(32'hbaef8a31),
	.w2(32'hbafd1187),
	.w3(32'hbae1fc28),
	.w4(32'hb872c7a6),
	.w5(32'hbadd5a22),
	.w6(32'hbac1e4e8),
	.w7(32'hba190d1c),
	.w8(32'hbaec2926),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a5738),
	.w1(32'hb9e847ff),
	.w2(32'hba5dbd8e),
	.w3(32'hb9d941b5),
	.w4(32'h391656df),
	.w5(32'hba0890df),
	.w6(32'hb90ba417),
	.w7(32'hba1d7ecb),
	.w8(32'hba63d1d5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1af5f3),
	.w1(32'hbb024940),
	.w2(32'hbb94ddc4),
	.w3(32'hba4dad7a),
	.w4(32'hba73a33e),
	.w5(32'hbb4cfaca),
	.w6(32'hbaf117ee),
	.w7(32'hba977bbc),
	.w8(32'hbb818e2e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2c900),
	.w1(32'hb99d7dc5),
	.w2(32'hbb24c451),
	.w3(32'h3ad84a9c),
	.w4(32'h3b0159b9),
	.w5(32'h3b077861),
	.w6(32'h3b21ae7c),
	.w7(32'h3a6546f3),
	.w8(32'hb9dcbedf),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fafe9a),
	.w1(32'hba34bb96),
	.w2(32'hbaf693ee),
	.w3(32'h3aa4f04e),
	.w4(32'hbaa384e9),
	.w5(32'hbb0cd0fd),
	.w6(32'h391d3af3),
	.w7(32'hba79e639),
	.w8(32'hbaa24f05),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fcbfd0),
	.w1(32'h3767aa88),
	.w2(32'hb9402bcf),
	.w3(32'h38cf5ac5),
	.w4(32'hb9a7dfbc),
	.w5(32'hb99df2b5),
	.w6(32'hb80c1b3a),
	.w7(32'hb9afa42f),
	.w8(32'hb8cd7a62),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9772e71),
	.w1(32'hb97ad08c),
	.w2(32'hb9aa3f40),
	.w3(32'hb776884b),
	.w4(32'h38161593),
	.w5(32'h386406e5),
	.w6(32'hb96297d3),
	.w7(32'hb9d66f9d),
	.w8(32'hb8c99d54),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b60546),
	.w1(32'hb9e0236d),
	.w2(32'hb9a1ed46),
	.w3(32'h39836a0f),
	.w4(32'hb91e3ec6),
	.w5(32'hb97351aa),
	.w6(32'hb96aa768),
	.w7(32'hb94c9abc),
	.w8(32'hb81a214d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7a36b),
	.w1(32'hba738a46),
	.w2(32'hbb11eeaa),
	.w3(32'h3a6f42fe),
	.w4(32'hbb0bc2a6),
	.w5(32'hbb4e83b6),
	.w6(32'h39c97bb2),
	.w7(32'hba4f3e57),
	.w8(32'hbacefc94),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9368ed),
	.w1(32'hba569325),
	.w2(32'hba76eeae),
	.w3(32'hb6a05f5d),
	.w4(32'h396382fb),
	.w5(32'hb8d73326),
	.w6(32'hba96fdb3),
	.w7(32'hba78c76f),
	.w8(32'hbb04aced),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6547e),
	.w1(32'hbabd0de4),
	.w2(32'h3a0522fb),
	.w3(32'hb9342922),
	.w4(32'h3ac21ee3),
	.w5(32'h3b1fb95d),
	.w6(32'hbab7067e),
	.w7(32'hba41455f),
	.w8(32'hba406e1e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3882836e),
	.w1(32'h3a0418c0),
	.w2(32'h39f7784c),
	.w3(32'h39bf88b1),
	.w4(32'h3a0d0262),
	.w5(32'h3a382a98),
	.w6(32'h399dcace),
	.w7(32'h396ef2f8),
	.w8(32'h38e5a1a5),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6404e9),
	.w1(32'hba6e529b),
	.w2(32'hbb3fb6c8),
	.w3(32'h3a9d5004),
	.w4(32'hb9969936),
	.w5(32'hbb229184),
	.w6(32'hbb0119f9),
	.w7(32'hbaf30cf8),
	.w8(32'hbb6f0ca0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e53992),
	.w1(32'hba8e45e9),
	.w2(32'hbad8a886),
	.w3(32'hba07a571),
	.w4(32'hba4f44e8),
	.w5(32'hbab0ec6f),
	.w6(32'hba1688e6),
	.w7(32'hb9ece420),
	.w8(32'hbadcb7a7),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a1c55),
	.w1(32'h39b88db7),
	.w2(32'h393ed403),
	.w3(32'h386264f9),
	.w4(32'h399d9fc9),
	.w5(32'h390900ed),
	.w6(32'h398bf21e),
	.w7(32'h397badf6),
	.w8(32'h396e2645),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a44fc),
	.w1(32'hbb4ea4ff),
	.w2(32'hbace01fe),
	.w3(32'hbb0ae07b),
	.w4(32'hba2e60de),
	.w5(32'hb90ff95f),
	.w6(32'hbaab9678),
	.w7(32'hb958fc86),
	.w8(32'h3a2f8798),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e27f0),
	.w1(32'h380d2c81),
	.w2(32'hb726f4f7),
	.w3(32'h395f8a8d),
	.w4(32'h3898bdb1),
	.w5(32'h38011aed),
	.w6(32'h39642c84),
	.w7(32'h392f7ad6),
	.w8(32'h38faadfb),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae86ec2),
	.w1(32'hba8c266c),
	.w2(32'hbaee6b62),
	.w3(32'hba3ae9e3),
	.w4(32'h39046bde),
	.w5(32'hba1da99c),
	.w6(32'hbad7b739),
	.w7(32'hba8cc0fd),
	.w8(32'hbafc064d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e7b6bd),
	.w1(32'h393fccc4),
	.w2(32'h3a9e36d7),
	.w3(32'h39d68846),
	.w4(32'h3a3a1eb5),
	.w5(32'h3a048faf),
	.w6(32'hba94f0d3),
	.w7(32'hba9d2cdf),
	.w8(32'hbb0221ad),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a195b74),
	.w1(32'h39acd8a5),
	.w2(32'hb9b8b2f3),
	.w3(32'h39ff7c07),
	.w4(32'h3a98a87c),
	.w5(32'h39b153bc),
	.w6(32'hba0aa525),
	.w7(32'hb9c93862),
	.w8(32'hbaaea335),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd679c),
	.w1(32'h3812a68e),
	.w2(32'hb901a7d8),
	.w3(32'h3992a01e),
	.w4(32'h3925aff6),
	.w5(32'h37f5c668),
	.w6(32'h3826062a),
	.w7(32'hb88ce845),
	.w8(32'hb8adb3ed),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d88fd),
	.w1(32'hba608398),
	.w2(32'hba9a9c85),
	.w3(32'h3a337ea4),
	.w4(32'h3abf8625),
	.w5(32'h3ab3f5cb),
	.w6(32'hb9a5a585),
	.w7(32'hba0d5f3e),
	.w8(32'hba9dd685),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba938296),
	.w1(32'hba42ecd2),
	.w2(32'hbac26890),
	.w3(32'hb9893937),
	.w4(32'hb96ebf71),
	.w5(32'hb9caa9d2),
	.w6(32'hbac0b14d),
	.w7(32'hba16b6cf),
	.w8(32'hba20b60e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba738268),
	.w1(32'hb99a0213),
	.w2(32'hba96893a),
	.w3(32'h3a2db29d),
	.w4(32'h39f46e47),
	.w5(32'hb9221ea7),
	.w6(32'hba8f164b),
	.w7(32'hbae5c851),
	.w8(32'hbb0cafc9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3809cfc8),
	.w1(32'hb83fd6ff),
	.w2(32'hb8f76e58),
	.w3(32'hb6e70259),
	.w4(32'h37fe843b),
	.w5(32'h397e381e),
	.w6(32'h38075b56),
	.w7(32'hb812f3c7),
	.w8(32'h376d4ff6),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b188b),
	.w1(32'h39345a7d),
	.w2(32'hb785da21),
	.w3(32'h39810b63),
	.w4(32'h38dd9bc9),
	.w5(32'hb8a61f50),
	.w6(32'h38d1254e),
	.w7(32'hb86a917a),
	.w8(32'hb7698ebd),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c35371),
	.w1(32'hbb27e113),
	.w2(32'hbb40a267),
	.w3(32'h3ae079fa),
	.w4(32'hb9ed6832),
	.w5(32'h3813ee45),
	.w6(32'hbb498b4a),
	.w7(32'hbb2b557a),
	.w8(32'hbb45b293),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb483c33),
	.w1(32'hbb6551b4),
	.w2(32'hbb9b30a5),
	.w3(32'hbaa120bb),
	.w4(32'hb8eebeac),
	.w5(32'hbad6f23e),
	.w6(32'hbb7017ff),
	.w7(32'hbb2ebaa4),
	.w8(32'hbb9b9253),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74f0e8),
	.w1(32'h3a11a2f8),
	.w2(32'h3a3d9e04),
	.w3(32'h3a9e9507),
	.w4(32'h3add90fe),
	.w5(32'h3b10c955),
	.w6(32'hba86705a),
	.w7(32'hb8e692ce),
	.w8(32'hba5ae253),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1c9ef),
	.w1(32'hbab61168),
	.w2(32'hba6e7c31),
	.w3(32'h3a9d5b34),
	.w4(32'hbb58f95f),
	.w5(32'hbb6a1b20),
	.w6(32'h3a012691),
	.w7(32'hbaac39a1),
	.w8(32'hbaff6a80),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59cb57),
	.w1(32'hba4a6aa5),
	.w2(32'hba431f1a),
	.w3(32'hba5a6317),
	.w4(32'hb9d2ef02),
	.w5(32'hb94c4177),
	.w6(32'hba121595),
	.w7(32'hb9caf9be),
	.w8(32'hb8951213),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaea66),
	.w1(32'hbab12675),
	.w2(32'hba970c18),
	.w3(32'hba2e9c00),
	.w4(32'hb97a60a2),
	.w5(32'h396e2bfc),
	.w6(32'hba294e61),
	.w7(32'hba14ac83),
	.w8(32'h37e06e36),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd6474),
	.w1(32'hbb0d890c),
	.w2(32'hbba036cc),
	.w3(32'h3aad90e6),
	.w4(32'hbb613d9b),
	.w5(32'hbbc30c12),
	.w6(32'hbb2000be),
	.w7(32'hbabbcaf6),
	.w8(32'hbb42b118),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13d7e3),
	.w1(32'hbb02feb1),
	.w2(32'hbb9938e5),
	.w3(32'hbaa151c2),
	.w4(32'hbad6710b),
	.w5(32'hbb33607f),
	.w6(32'hbad8ce7a),
	.w7(32'hba9348b2),
	.w8(32'hbb5b04b1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242f3f),
	.w1(32'hbb3b6ef4),
	.w2(32'hbb698b49),
	.w3(32'hba77f516),
	.w4(32'hbaa0dd01),
	.w5(32'hbb0fb5ec),
	.w6(32'hbb9d6759),
	.w7(32'hba3d6106),
	.w8(32'hbb6f9e19),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01cab4),
	.w1(32'h3a8e710a),
	.w2(32'h3ab5d4e8),
	.w3(32'h3998b7fd),
	.w4(32'h3a72e281),
	.w5(32'h3a803b95),
	.w6(32'hba1e2cc3),
	.w7(32'hba54517d),
	.w8(32'hba3b03ce),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4892b),
	.w1(32'hbaa703b6),
	.w2(32'hba96ab99),
	.w3(32'hb9553557),
	.w4(32'h3a4a32ec),
	.w5(32'h3a747a1f),
	.w6(32'hba5661d1),
	.w7(32'hba955217),
	.w8(32'hbae08155),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64daa15),
	.w1(32'hb81acc13),
	.w2(32'hb8e9c2fc),
	.w3(32'hb4edfe92),
	.w4(32'h394c51e6),
	.w5(32'h3971c658),
	.w6(32'h38f2d2be),
	.w7(32'hb819bbff),
	.w8(32'h38137dd4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3827cbc4),
	.w1(32'h3a7ee38c),
	.w2(32'h3a50b2e2),
	.w3(32'h3957ef24),
	.w4(32'h399f5db4),
	.w5(32'h389f50fc),
	.w6(32'h3a5b289d),
	.w7(32'h3a81f320),
	.w8(32'h3a3e3c5a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e057c),
	.w1(32'h3917335e),
	.w2(32'hb88d3e26),
	.w3(32'h3a54ae92),
	.w4(32'hb9a6cd25),
	.w5(32'hba2de615),
	.w6(32'hb89ea466),
	.w7(32'hb9c48f0b),
	.w8(32'hba089fe4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9847972),
	.w1(32'h37ece462),
	.w2(32'hb92de0b1),
	.w3(32'hb895950c),
	.w4(32'hb896124f),
	.w5(32'hb92b63ef),
	.w6(32'h39dde316),
	.w7(32'h3834a782),
	.w8(32'h3895b532),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83723d2),
	.w1(32'hbae7d66b),
	.w2(32'hbb3b7346),
	.w3(32'h39d6ad12),
	.w4(32'hbaf5ce56),
	.w5(32'hbb24cd7a),
	.w6(32'h39a2129b),
	.w7(32'hba9789fb),
	.w8(32'hbaaa502d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb405197),
	.w1(32'hbb4c0132),
	.w2(32'hbb5a5864),
	.w3(32'hb9b11533),
	.w4(32'hba4abde2),
	.w5(32'hbac0fee0),
	.w6(32'hbb0fbe11),
	.w7(32'hbaf1975c),
	.w8(32'hbb2fdec4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971d8a3),
	.w1(32'hba178011),
	.w2(32'hbacdb6c4),
	.w3(32'h3a82ca68),
	.w4(32'hb98f483d),
	.w5(32'hb92d84fe),
	.w6(32'hba823a6a),
	.w7(32'hba89df60),
	.w8(32'hba9755e6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7766e),
	.w1(32'h3a341f0a),
	.w2(32'h3a42d504),
	.w3(32'hb9596fb4),
	.w4(32'h38886274),
	.w5(32'h39b9acd3),
	.w6(32'h3a01c090),
	.w7(32'h3aad2ce8),
	.w8(32'h3a5d081c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c488),
	.w1(32'hbb823108),
	.w2(32'hbbcd0d19),
	.w3(32'hba6bde05),
	.w4(32'hbb04c986),
	.w5(32'hbb1542b7),
	.w6(32'hbb75fb6f),
	.w7(32'hbae56309),
	.w8(32'hbba17b6b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38034b33),
	.w1(32'hb7dc5846),
	.w2(32'hba87c5d8),
	.w3(32'h3a2070f6),
	.w4(32'h3958833a),
	.w5(32'hb9ee6ca2),
	.w6(32'hba25f44a),
	.w7(32'hba167376),
	.w8(32'hba98ef7c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c2150b),
	.w1(32'h3983dbec),
	.w2(32'h39518a82),
	.w3(32'h39163b35),
	.w4(32'h3952b652),
	.w5(32'h3853e279),
	.w6(32'h394b98fc),
	.w7(32'h394ea5c4),
	.w8(32'h398aa085),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9963c11),
	.w1(32'hba9f087e),
	.w2(32'hbb0866e5),
	.w3(32'h398094ad),
	.w4(32'hba4d15ad),
	.w5(32'hbabcb375),
	.w6(32'hba6bb806),
	.w7(32'hba4ae125),
	.w8(32'hbabf860d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e69893),
	.w1(32'hb93ea886),
	.w2(32'hb9020abd),
	.w3(32'hb7d9f3d7),
	.w4(32'h39148cbf),
	.w5(32'h3945182f),
	.w6(32'h38098f26),
	.w7(32'hb8bfee6b),
	.w8(32'hb8f5bc32),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920d4fe),
	.w1(32'hb7e4c866),
	.w2(32'hb9a2db72),
	.w3(32'h39a13f4e),
	.w4(32'h3714bf35),
	.w5(32'hb8dbedbb),
	.w6(32'hb956f170),
	.w7(32'hb99f4899),
	.w8(32'hb9bbf452),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9272382),
	.w1(32'h39913634),
	.w2(32'h39753ec9),
	.w3(32'hb90bc95c),
	.w4(32'h39625c05),
	.w5(32'h3908767a),
	.w6(32'h39610da5),
	.w7(32'h394e8265),
	.w8(32'h39aa1b93),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a889e4),
	.w1(32'hb9045b73),
	.w2(32'hb9929a8a),
	.w3(32'h397e6423),
	.w4(32'h3956346b),
	.w5(32'h389e67ff),
	.w6(32'hb99593be),
	.w7(32'hb9e3160a),
	.w8(32'hb92dd4e1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39942d93),
	.w1(32'h3aa63993),
	.w2(32'h39a7ec70),
	.w3(32'h399c0a3f),
	.w4(32'h3a90e697),
	.w5(32'h39afa454),
	.w6(32'hb9a89d96),
	.w7(32'h39b39837),
	.w8(32'hb86cc0a8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914b4b3),
	.w1(32'hba75a6c3),
	.w2(32'hbb7ed51b),
	.w3(32'hba83105d),
	.w4(32'hbb1b7521),
	.w5(32'hbb2c667f),
	.w6(32'hba7d6a48),
	.w7(32'hbaa4e035),
	.w8(32'hbb47a6c8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad39432),
	.w1(32'hba29f2af),
	.w2(32'hbb183904),
	.w3(32'hb9c52d9c),
	.w4(32'h39d0aa91),
	.w5(32'hb9aa0af0),
	.w6(32'hb9ee7177),
	.w7(32'h3927b34b),
	.w8(32'hba7623a8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1af59c),
	.w1(32'hb997bfe4),
	.w2(32'hbb0829de),
	.w3(32'h38de5e30),
	.w4(32'hba6a9aa0),
	.w5(32'hbafe328a),
	.w6(32'hba972b6a),
	.w7(32'hba857502),
	.w8(32'hbb1fd7b5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fdbf3d),
	.w1(32'h37d65a9b),
	.w2(32'hb8ad814d),
	.w3(32'h38e5eb9e),
	.w4(32'h393f9d74),
	.w5(32'h38b1344f),
	.w6(32'h37a48e06),
	.w7(32'hb77e2387),
	.w8(32'hb87c0c79),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22b6cc),
	.w1(32'hb98912b9),
	.w2(32'hb8679ed8),
	.w3(32'hb9a0e53e),
	.w4(32'h388ef1d0),
	.w5(32'h38e23fc2),
	.w6(32'h38bef602),
	.w7(32'h38a31fd4),
	.w8(32'h39d5dd00),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efa03a),
	.w1(32'h39a8e85b),
	.w2(32'h39b4787f),
	.w3(32'h39b4b8dc),
	.w4(32'h397a9f60),
	.w5(32'h394a88a6),
	.w6(32'h399d248c),
	.w7(32'h39bcf2a6),
	.w8(32'h39bb4219),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4f484),
	.w1(32'h39b73817),
	.w2(32'h39c322a9),
	.w3(32'h398d5639),
	.w4(32'h3994f77d),
	.w5(32'h39520713),
	.w6(32'h39baa4f6),
	.w7(32'h39dd6693),
	.w8(32'h39d8df56),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bfff4),
	.w1(32'hbb11443e),
	.w2(32'hbb86419b),
	.w3(32'hbafd4617),
	.w4(32'hba322d6b),
	.w5(32'hba9bd78a),
	.w6(32'hbb103391),
	.w7(32'hba24fddf),
	.w8(32'hbaf6d038),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81c1db4),
	.w1(32'hb962308f),
	.w2(32'hb88aa706),
	.w3(32'h398ced59),
	.w4(32'hb92bbd42),
	.w5(32'hb7f6f8d9),
	.w6(32'hb936e300),
	.w7(32'hb8cb988c),
	.w8(32'h39122859),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2edc2),
	.w1(32'h39be66ce),
	.w2(32'h39a3bdfd),
	.w3(32'h3881be85),
	.w4(32'h3a3f4bf6),
	.w5(32'h3a1db8f6),
	.w6(32'h398d9b26),
	.w7(32'h39aa91d5),
	.w8(32'h39e10c7b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad112c8),
	.w1(32'hbad9846d),
	.w2(32'hbac41730),
	.w3(32'hbad07c97),
	.w4(32'hba56f557),
	.w5(32'hb9ac29ec),
	.w6(32'hba232ef3),
	.w7(32'hb7be477a),
	.w8(32'hb9275ceb),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8501b3f),
	.w1(32'h39aff3a9),
	.w2(32'h398870bc),
	.w3(32'hb7928f95),
	.w4(32'h39a6dcf1),
	.w5(32'h3986d47f),
	.w6(32'h39a90a4c),
	.w7(32'h39ae7feb),
	.w8(32'h39a7620f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382595b3),
	.w1(32'hb96e5a36),
	.w2(32'hba775e1f),
	.w3(32'h39e48fd4),
	.w4(32'hb9026bb9),
	.w5(32'hb9ce1b8d),
	.w6(32'h39a1a7f2),
	.w7(32'h3a5826d3),
	.w8(32'hba0299fc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d31ba),
	.w1(32'h3908bc3f),
	.w2(32'hb932648a),
	.w3(32'hb6a0b613),
	.w4(32'h38b4d13e),
	.w5(32'h3734d76d),
	.w6(32'h390f8dd8),
	.w7(32'h391b2301),
	.w8(32'h38e4fae5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba297b7),
	.w1(32'hbb9f38ae),
	.w2(32'hbc01cd8e),
	.w3(32'hbb97ed26),
	.w4(32'hbb332e9f),
	.w5(32'hbb154bfa),
	.w6(32'hbaefcc45),
	.w7(32'h3901373c),
	.w8(32'hba1808d5),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967aaf0),
	.w1(32'h39d434bb),
	.w2(32'h3a4d8754),
	.w3(32'hb959e366),
	.w4(32'h3a82cb80),
	.w5(32'h389105fd),
	.w6(32'h3a8ec00e),
	.w7(32'h3a1b7c2c),
	.w8(32'hb8b736a5),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc2823),
	.w1(32'hba5d5788),
	.w2(32'hba4b70b5),
	.w3(32'hbaeb7e41),
	.w4(32'hba7e89e9),
	.w5(32'hbaa1be09),
	.w6(32'hbadc5ba0),
	.w7(32'hba84994d),
	.w8(32'hbb01d7ff),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule