module layer_10_featuremap_417(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75a49e),
	.w1(32'h3b1091a6),
	.w2(32'h3b1c8a6a),
	.w3(32'hbb0ddce2),
	.w4(32'hbb76d87c),
	.w5(32'h3a3dd7ef),
	.w6(32'h3a108403),
	.w7(32'hbbd093f2),
	.w8(32'hbabc572d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34fec7),
	.w1(32'h3b2f78bf),
	.w2(32'h3bf0e567),
	.w3(32'h3c0009c8),
	.w4(32'h39d40252),
	.w5(32'h3cc62daa),
	.w6(32'h3b40d500),
	.w7(32'hba1a971c),
	.w8(32'h3c8ed8e2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a00b8),
	.w1(32'h3b745b3a),
	.w2(32'h3af331a0),
	.w3(32'h3be90ea6),
	.w4(32'h3b49c120),
	.w5(32'h3b8e83ec),
	.w6(32'h3bd8c7b8),
	.w7(32'hbb22d4d3),
	.w8(32'h3b56f3e6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad91b9e),
	.w1(32'hbabf1b46),
	.w2(32'h3c1c523e),
	.w3(32'hbb90aaa7),
	.w4(32'hbb97b842),
	.w5(32'h3bbc3794),
	.w6(32'hbbb1a93d),
	.w7(32'hbb428215),
	.w8(32'h3b3473b2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac29247),
	.w1(32'hbadc154c),
	.w2(32'hbb84fbc7),
	.w3(32'h3995e125),
	.w4(32'h3b92491c),
	.w5(32'h3b152bd3),
	.w6(32'hbb40cec8),
	.w7(32'h3b4df8ab),
	.w8(32'h3bdaec6f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af29b20),
	.w1(32'h3b72e4d8),
	.w2(32'hba579598),
	.w3(32'h3a403196),
	.w4(32'h3b10e672),
	.w5(32'h3b664ef2),
	.w6(32'h3999d73c),
	.w7(32'h3b3247ac),
	.w8(32'h3b50484e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a76f),
	.w1(32'hbc06f4d0),
	.w2(32'hbb6a35e0),
	.w3(32'hbb32f706),
	.w4(32'hbc1f6b7f),
	.w5(32'hbc1a91d3),
	.w6(32'hbaca53e9),
	.w7(32'hbb9d115c),
	.w8(32'hbb65bff8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bbfb2),
	.w1(32'hbc1d82a1),
	.w2(32'hbc35707c),
	.w3(32'hbc1c1d4d),
	.w4(32'hbb72770a),
	.w5(32'hbac16ae5),
	.w6(32'hbc746ea8),
	.w7(32'h3bb6b092),
	.w8(32'h3ba823d4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7c0f3),
	.w1(32'h3b67e71a),
	.w2(32'h3b379297),
	.w3(32'h3a591f00),
	.w4(32'hba26374f),
	.w5(32'h3bf07918),
	.w6(32'h3b9337ae),
	.w7(32'h3b5bca39),
	.w8(32'h3b896d63),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26ee75),
	.w1(32'hbafed040),
	.w2(32'hbc16dfca),
	.w3(32'hbbeb271c),
	.w4(32'h3b4ea86c),
	.w5(32'hbbdcd3b2),
	.w6(32'hbad6c969),
	.w7(32'h3ba0dd6f),
	.w8(32'hba9bef30),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95f3f1),
	.w1(32'h3b01b21e),
	.w2(32'h3a460ab8),
	.w3(32'hbb68e434),
	.w4(32'h37c7c176),
	.w5(32'h3c0a5475),
	.w6(32'hba965a69),
	.w7(32'hbbfda439),
	.w8(32'hb9471fd1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35a8b6),
	.w1(32'h3a4ac748),
	.w2(32'h398c613f),
	.w3(32'hbb8ca429),
	.w4(32'h3bed0279),
	.w5(32'hbc059827),
	.w6(32'h3b909582),
	.w7(32'h3c2161c1),
	.w8(32'hba1ae0eb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a299e),
	.w1(32'hba677d45),
	.w2(32'h38f38d3e),
	.w3(32'hba6b5431),
	.w4(32'hbb5b6476),
	.w5(32'h3bcf533a),
	.w6(32'h3b3be295),
	.w7(32'h3c1934ca),
	.w8(32'h3c587f5a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb53026),
	.w1(32'hba27bfc8),
	.w2(32'hbc272f12),
	.w3(32'hbbfc815a),
	.w4(32'hbac6a81b),
	.w5(32'hbb93b70b),
	.w6(32'hbaf7b2e5),
	.w7(32'hbba03113),
	.w8(32'hb9ae4ce1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc051d7e),
	.w1(32'h3b48ecc6),
	.w2(32'h39a990ff),
	.w3(32'hbbcc7f75),
	.w4(32'h3b35e19c),
	.w5(32'h3c03a82f),
	.w6(32'hbb830631),
	.w7(32'h3be625f5),
	.w8(32'h3c09201f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb9c15),
	.w1(32'h396755e8),
	.w2(32'hbc0148fa),
	.w3(32'hbbd03e16),
	.w4(32'h3bb9eb72),
	.w5(32'hbb97078f),
	.w6(32'hbaf938fd),
	.w7(32'h3c40940b),
	.w8(32'h3b2433a9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b700455),
	.w1(32'hbb89b257),
	.w2(32'hbbbcfd91),
	.w3(32'hbb283389),
	.w4(32'hbad814b3),
	.w5(32'hbbb43074),
	.w6(32'hbb8e1d44),
	.w7(32'h3b4d9e67),
	.w8(32'hbaae300a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf780a8),
	.w1(32'h3b6baaa5),
	.w2(32'hbc18fbbb),
	.w3(32'hba9fb603),
	.w4(32'h3c35c29f),
	.w5(32'hbb552bec),
	.w6(32'hb9bfeac5),
	.w7(32'h3c669ddd),
	.w8(32'h3c083169),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8a709),
	.w1(32'h3b1bd28b),
	.w2(32'hbb48969f),
	.w3(32'h3a56bb90),
	.w4(32'h3b8dd6aa),
	.w5(32'h3b85067b),
	.w6(32'hba6a6fb2),
	.w7(32'h3bff39e4),
	.w8(32'h3ba346ca),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba524abf),
	.w1(32'hbbc230ba),
	.w2(32'h398989ef),
	.w3(32'hbb1dbb82),
	.w4(32'hbc07cdb1),
	.w5(32'h3bdc835d),
	.w6(32'h3a94de31),
	.w7(32'hbb16ad0f),
	.w8(32'h3a9fe6fe),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a50881),
	.w1(32'hbb56bedc),
	.w2(32'h3be30af8),
	.w3(32'h3aaae9ce),
	.w4(32'hbab2f3fa),
	.w5(32'h3ba4f492),
	.w6(32'h3b31556c),
	.w7(32'h3b005abd),
	.w8(32'h3b9ea657),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ea5bf),
	.w1(32'hbba1a683),
	.w2(32'h3c2f7ff1),
	.w3(32'hbb4c60cc),
	.w4(32'hbb8c8d62),
	.w5(32'h3c287a0d),
	.w6(32'hbb999f1e),
	.w7(32'h3843c027),
	.w8(32'h3c56f411),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd22089),
	.w1(32'hbbf46309),
	.w2(32'h398e2aca),
	.w3(32'hbcc6d638),
	.w4(32'hbba9ce50),
	.w5(32'hbb81c745),
	.w6(32'hbcd40449),
	.w7(32'hbc622732),
	.w8(32'hbbf88cf4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35cc45),
	.w1(32'hbbd6c712),
	.w2(32'hbb378c0d),
	.w3(32'h3b892489),
	.w4(32'hbb0e9163),
	.w5(32'h3ba268cd),
	.w6(32'h3be446e5),
	.w7(32'hbaa4467c),
	.w8(32'h3bd0b5d4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50ec32),
	.w1(32'hbb296192),
	.w2(32'hbc35a847),
	.w3(32'hbc4ca561),
	.w4(32'hbbda869c),
	.w5(32'hbb8fff55),
	.w6(32'hbca53ccc),
	.w7(32'hba1fb92e),
	.w8(32'hbb94ed10),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b9a9e),
	.w1(32'h3b8bfcb5),
	.w2(32'h3b973697),
	.w3(32'hbb98299e),
	.w4(32'h3bb3882c),
	.w5(32'hbbb73c9c),
	.w6(32'h3bd4ebc8),
	.w7(32'h3b567b31),
	.w8(32'hbb2e0817),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b891a05),
	.w1(32'hbbb6d045),
	.w2(32'h3c38e6a8),
	.w3(32'h3c40c111),
	.w4(32'hbbe8f916),
	.w5(32'h3c31436f),
	.w6(32'h3bcb6f77),
	.w7(32'h3a66db02),
	.w8(32'h3bb23172),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ca2cf),
	.w1(32'h3a41a3ae),
	.w2(32'h3b104bf8),
	.w3(32'hbaa65075),
	.w4(32'h3bb33534),
	.w5(32'h3be4ac4d),
	.w6(32'hbaed3e5e),
	.w7(32'h3c1775c9),
	.w8(32'h3c11b4ab),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d625b),
	.w1(32'hbb499b0f),
	.w2(32'h3b87dee3),
	.w3(32'hbc453a56),
	.w4(32'hbaab0cd8),
	.w5(32'hbab40198),
	.w6(32'hbc25fcb6),
	.w7(32'h3c0c00b8),
	.w8(32'hbc028923),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81ece0),
	.w1(32'hba9baa47),
	.w2(32'hbb598ae6),
	.w3(32'h398f7073),
	.w4(32'h3b8f2a1c),
	.w5(32'hbb3f4e86),
	.w6(32'hbbc240cf),
	.w7(32'h3b25c15c),
	.w8(32'hb9c353c1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397bdf60),
	.w1(32'hbb90395e),
	.w2(32'hbb0c5adf),
	.w3(32'hb8a80999),
	.w4(32'h3b4d1dee),
	.w5(32'hbbef35ba),
	.w6(32'hb9b435ac),
	.w7(32'hbaef6937),
	.w8(32'h3a5abd02),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ffa2),
	.w1(32'h3a8f3099),
	.w2(32'h39fc9846),
	.w3(32'h3bd99767),
	.w4(32'h3a3a13cb),
	.w5(32'h3bbd8e8b),
	.w6(32'h3b3503f1),
	.w7(32'h3ae07e55),
	.w8(32'h3b87ed6d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a3e42),
	.w1(32'h3bc703a0),
	.w2(32'hbb1d7552),
	.w3(32'h3a2bafb5),
	.w4(32'h3c583340),
	.w5(32'h3c5cfdd3),
	.w6(32'h3aadd2bc),
	.w7(32'h3a8e87fe),
	.w8(32'h3bc5ce7e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e48da),
	.w1(32'hba1a5ac6),
	.w2(32'hbb5c3479),
	.w3(32'hbb12efe6),
	.w4(32'h3baa1f10),
	.w5(32'hbb843fa3),
	.w6(32'hba4e8764),
	.w7(32'hbb2b9c17),
	.w8(32'hbbcd259e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85d08d),
	.w1(32'h393c8b69),
	.w2(32'hba50ac51),
	.w3(32'h3a839ee0),
	.w4(32'h3b3e7bdc),
	.w5(32'hbbc5a488),
	.w6(32'h3b7d22de),
	.w7(32'h3c22a42a),
	.w8(32'hbb1d547d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aafa3),
	.w1(32'hbb802ec5),
	.w2(32'hbc04c382),
	.w3(32'h3b835a55),
	.w4(32'hbb5ece18),
	.w5(32'hbb9e4028),
	.w6(32'h3b36a373),
	.w7(32'h3bcf1f8d),
	.w8(32'h3b07e887),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8965ca),
	.w1(32'hbba7a362),
	.w2(32'h3b77df7e),
	.w3(32'hbc89718a),
	.w4(32'hbb3956ac),
	.w5(32'h3c92fbbd),
	.w6(32'hbb19f502),
	.w7(32'hbb7f02fb),
	.w8(32'hbbb1e845),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f1645),
	.w1(32'hbb11a9b6),
	.w2(32'h3a51b832),
	.w3(32'hbc94740c),
	.w4(32'hbbe71a11),
	.w5(32'h3c1a4bbc),
	.w6(32'hbc8796c0),
	.w7(32'hbc7e63f1),
	.w8(32'h3b9285dc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e68a3),
	.w1(32'hba41c754),
	.w2(32'h3b97332c),
	.w3(32'hbc9699fe),
	.w4(32'hbc3cba3e),
	.w5(32'h3b6658db),
	.w6(32'hbcd5a775),
	.w7(32'hbc880acb),
	.w8(32'hbbce7f1c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9d750),
	.w1(32'hbbcc6769),
	.w2(32'hbb5581c4),
	.w3(32'h3b8706e1),
	.w4(32'hbbeb1a40),
	.w5(32'hbaaafe91),
	.w6(32'h3a94174b),
	.w7(32'hbbc9e0ee),
	.w8(32'hbb924ef7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba3756),
	.w1(32'hbbc1400c),
	.w2(32'h3b075ac2),
	.w3(32'hbbcdad27),
	.w4(32'hbad2a162),
	.w5(32'hbc0be764),
	.w6(32'hbb12c54d),
	.w7(32'hbb60a8cd),
	.w8(32'hbb37bed4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b820136),
	.w1(32'hbb0fe786),
	.w2(32'hb9ed4be9),
	.w3(32'h3a96d64f),
	.w4(32'hbba0d899),
	.w5(32'h3c1222ee),
	.w6(32'hbba3fe9b),
	.w7(32'hbaef5f92),
	.w8(32'h3b9ec137),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc481dc),
	.w1(32'hbb432b10),
	.w2(32'h3aae508a),
	.w3(32'hbc04c34a),
	.w4(32'hbc0cfab7),
	.w5(32'h3b302487),
	.w6(32'hbc28273e),
	.w7(32'hbb4c1313),
	.w8(32'hbabb6aac),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f44af),
	.w1(32'hbba7bd7b),
	.w2(32'hb99f8dfc),
	.w3(32'hbc410311),
	.w4(32'hbbe746ae),
	.w5(32'h3c031635),
	.w6(32'hbb80268c),
	.w7(32'hbbf56d6d),
	.w8(32'h3c8d328b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ad17a),
	.w1(32'h3c1391fc),
	.w2(32'hbb8a58f3),
	.w3(32'hb990d4d7),
	.w4(32'h3c3030b1),
	.w5(32'h39bd093f),
	.w6(32'hbb79a699),
	.w7(32'h3c73f659),
	.w8(32'hbb462e96),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3e54a),
	.w1(32'h3bafef2c),
	.w2(32'hba9f7afc),
	.w3(32'h3ae2f533),
	.w4(32'h3c02cdee),
	.w5(32'h3ab52756),
	.w6(32'h3be96e35),
	.w7(32'h3c97e18b),
	.w8(32'h3b911195),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ef45e),
	.w1(32'hbb51f0f6),
	.w2(32'h3b0dfd88),
	.w3(32'hbb75a620),
	.w4(32'hbb99c6e2),
	.w5(32'h3940fc76),
	.w6(32'hbc12e6d5),
	.w7(32'hbb08cab2),
	.w8(32'h3b565def),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e4d74),
	.w1(32'hbb467375),
	.w2(32'hbaff6153),
	.w3(32'hbc497402),
	.w4(32'hbb36e300),
	.w5(32'h3bcd5399),
	.w6(32'hbba310a4),
	.w7(32'h3a744911),
	.w8(32'h3bb67705),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa5f79),
	.w1(32'hbbb69261),
	.w2(32'hbb03a185),
	.w3(32'hbb25eed4),
	.w4(32'hba2bf854),
	.w5(32'hbc54e2df),
	.w6(32'hbba9b9e4),
	.w7(32'hbb4b346b),
	.w8(32'hbbe96b7a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387bde4f),
	.w1(32'hbbe5b7ee),
	.w2(32'hbc1d9df5),
	.w3(32'hbbd4c07a),
	.w4(32'hb9db1fea),
	.w5(32'hbcbc979d),
	.w6(32'hbc022f6b),
	.w7(32'h3ac56ca3),
	.w8(32'hbc4f3347),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07ff2d),
	.w1(32'hbbb9e5c0),
	.w2(32'hbb69e5ce),
	.w3(32'hbc1408fe),
	.w4(32'hbb6c2c08),
	.w5(32'hbbdcb7d7),
	.w6(32'hbc19aa3b),
	.w7(32'hbb8d055d),
	.w8(32'hbbc7b157),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d11f1),
	.w1(32'h3bd05610),
	.w2(32'h3cb55cb3),
	.w3(32'hbc392867),
	.w4(32'h3b4a25ea),
	.w5(32'h3d3cf472),
	.w6(32'hbc1e00a5),
	.w7(32'h3b49643e),
	.w8(32'h3d2c19be),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c371e21),
	.w1(32'hbb015b13),
	.w2(32'hbbb2d6ed),
	.w3(32'h3c84c70b),
	.w4(32'h3adefe71),
	.w5(32'hbc1cf9df),
	.w6(32'h3c1c2739),
	.w7(32'h3b04fe09),
	.w8(32'hbbeb7353),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb999c18),
	.w1(32'h39328546),
	.w2(32'hbc14b965),
	.w3(32'hbb9e5234),
	.w4(32'h3bf8568d),
	.w5(32'h3bc8d2d7),
	.w6(32'h39d16368),
	.w7(32'h3c12e526),
	.w8(32'h3b99914e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b911796),
	.w1(32'h39bf5d7e),
	.w2(32'hbc622cbc),
	.w3(32'h3b815c74),
	.w4(32'h3b80f7b9),
	.w5(32'hbbbf0f9c),
	.w6(32'h3b2d3ef9),
	.w7(32'h3c348d91),
	.w8(32'hbb864e37),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb8d1d),
	.w1(32'h3bc56394),
	.w2(32'h3a7cc2c1),
	.w3(32'hbc07ca5b),
	.w4(32'h39e9eee7),
	.w5(32'h3c86d7fb),
	.w6(32'hbb99a6f2),
	.w7(32'h3b1e7ce4),
	.w8(32'h3b83ec62),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d3c5b),
	.w1(32'hbbee7395),
	.w2(32'hb926ee3e),
	.w3(32'h3a289924),
	.w4(32'hbbdef836),
	.w5(32'hbb0aae10),
	.w6(32'hbabb456c),
	.w7(32'hbb8b6a26),
	.w8(32'hbaa55413),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64de44),
	.w1(32'hbbd6306d),
	.w2(32'hbad6c9a4),
	.w3(32'h3b92b032),
	.w4(32'hbb42e29b),
	.w5(32'h3b376e65),
	.w6(32'h3b92b11a),
	.w7(32'hbb90dc3a),
	.w8(32'h3c2292d6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1905c6),
	.w1(32'hb9d29c17),
	.w2(32'hbb05e1fa),
	.w3(32'h3a56e5ae),
	.w4(32'hbbf8660b),
	.w5(32'h3a9baea8),
	.w6(32'hbb470c0c),
	.w7(32'hbacbae12),
	.w8(32'hbb363710),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb1ad8),
	.w1(32'hbb895e66),
	.w2(32'hbc1c2af5),
	.w3(32'hbbc0d437),
	.w4(32'hbbc523f4),
	.w5(32'hbab42f88),
	.w6(32'hbb1a3174),
	.w7(32'hba0d53e6),
	.w8(32'h3a583c26),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b474998),
	.w1(32'hbb824f82),
	.w2(32'h3a262d55),
	.w3(32'hbb82f008),
	.w4(32'h3bc0ff53),
	.w5(32'hba62ac82),
	.w6(32'hbb8d90ea),
	.w7(32'h3bcf3f85),
	.w8(32'h3c09b20b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb7a8f),
	.w1(32'hba143d05),
	.w2(32'hbbbc07a1),
	.w3(32'hbc0b7532),
	.w4(32'hb89fd0c0),
	.w5(32'h3a75fc60),
	.w6(32'hbbd64770),
	.w7(32'h3b86e820),
	.w8(32'h3b410dff),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb05d14),
	.w1(32'hbbc04fa9),
	.w2(32'h3be4d4da),
	.w3(32'hbbf460a1),
	.w4(32'hbc3570d9),
	.w5(32'h3c6e8381),
	.w6(32'hbb652ac7),
	.w7(32'hbbf2c9cc),
	.w8(32'h3b931834),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11d830),
	.w1(32'h3ae1c24b),
	.w2(32'hbbaae63b),
	.w3(32'hbbd428fa),
	.w4(32'h3b57e05b),
	.w5(32'hbc26bda2),
	.w6(32'hbc0b5ba4),
	.w7(32'h3b13214b),
	.w8(32'hbb23bef4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf89a7),
	.w1(32'hbbd4c5ca),
	.w2(32'h39a22a1b),
	.w3(32'h3b430ce9),
	.w4(32'hbbbfa68a),
	.w5(32'hbb2121b3),
	.w6(32'h3b459b38),
	.w7(32'hbbc4ec66),
	.w8(32'hbaae4cdf),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cc115),
	.w1(32'h3bf5ddb4),
	.w2(32'h3a8a0b7f),
	.w3(32'h39fe495f),
	.w4(32'h3b09c5fc),
	.w5(32'h3b49e3f9),
	.w6(32'h3b0d14f2),
	.w7(32'h3b89dab7),
	.w8(32'h3b29d123),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e604a),
	.w1(32'hbb5ef498),
	.w2(32'hbc5339f2),
	.w3(32'hb9a5e89b),
	.w4(32'h3b2151fa),
	.w5(32'h3a53de2e),
	.w6(32'h3be26dc7),
	.w7(32'hba88b1a3),
	.w8(32'h3ba81200),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27b3c7),
	.w1(32'hbb863506),
	.w2(32'hbbf719c0),
	.w3(32'h3b55b590),
	.w4(32'h3c73cbcc),
	.w5(32'h3b65b7a0),
	.w6(32'hbac1ae0c),
	.w7(32'h3bc05ff3),
	.w8(32'h3c4c6607),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbeed28),
	.w1(32'h3a0a226e),
	.w2(32'h3bdde4fa),
	.w3(32'hbc7c04b4),
	.w4(32'h3b47d45d),
	.w5(32'h3c8c2b53),
	.w6(32'hbc822980),
	.w7(32'h3b1b22df),
	.w8(32'h3c07dd6e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9eebf),
	.w1(32'h3c0cf4fe),
	.w2(32'h3c24a168),
	.w3(32'h3c2d492e),
	.w4(32'h3c00d8dd),
	.w5(32'h3ba6c75c),
	.w6(32'hba3048d4),
	.w7(32'h3c05b977),
	.w8(32'h3bad510b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b0a1f),
	.w1(32'hba61990f),
	.w2(32'h39ef28ff),
	.w3(32'h3b9e4113),
	.w4(32'h3aade81d),
	.w5(32'hb82f5448),
	.w6(32'h3b8dfc69),
	.w7(32'h3b50c609),
	.w8(32'h3ab2f7a4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914d635),
	.w1(32'hbbd42f85),
	.w2(32'hbb02ffa2),
	.w3(32'h3a903271),
	.w4(32'hb8b469e6),
	.w5(32'h3b99b185),
	.w6(32'h3bcf00de),
	.w7(32'hb96987c2),
	.w8(32'hbb560b08),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a784101),
	.w1(32'h3b8a9234),
	.w2(32'h3a96a14b),
	.w3(32'h3b32893b),
	.w4(32'h3b49741b),
	.w5(32'hb8f7fd44),
	.w6(32'hbb7ecd17),
	.w7(32'hb9e0df5e),
	.w8(32'hb7fd60e1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9a8a6),
	.w1(32'h3bb28358),
	.w2(32'h3b1c476f),
	.w3(32'hbbfabfd0),
	.w4(32'h3b4b8bbc),
	.w5(32'h3ab4e7ec),
	.w6(32'hbb98ee33),
	.w7(32'h39ad2335),
	.w8(32'hbb40e92a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae32cd7),
	.w1(32'hbadb2c84),
	.w2(32'h3b215211),
	.w3(32'h3ad1bb36),
	.w4(32'h3a482644),
	.w5(32'h3b6e6eb0),
	.w6(32'hbb6b84ba),
	.w7(32'hbb0ef5de),
	.w8(32'h3ba72bdb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a9e24),
	.w1(32'hbc5094eb),
	.w2(32'hbc413347),
	.w3(32'hbae8d583),
	.w4(32'hbb9c129c),
	.w5(32'hbb15b81b),
	.w6(32'h3c0b472e),
	.w7(32'h3b42f5e3),
	.w8(32'h3c112157),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8f75c),
	.w1(32'hbb0d3546),
	.w2(32'hbb67a3aa),
	.w3(32'hbc237673),
	.w4(32'hba4baa50),
	.w5(32'h3b7832a5),
	.w6(32'hbbe542db),
	.w7(32'h3a9c2f85),
	.w8(32'h3bd3c648),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf11757),
	.w1(32'hb989ba1c),
	.w2(32'hbbf26af6),
	.w3(32'h3b0d8095),
	.w4(32'h3b51fc6e),
	.w5(32'h3b264667),
	.w6(32'hba354750),
	.w7(32'hba2a5496),
	.w8(32'hbb723557),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a5b8d),
	.w1(32'h3a3be9a9),
	.w2(32'h39d43d2c),
	.w3(32'h3c0166e4),
	.w4(32'h3a9b4df4),
	.w5(32'h3ab75be9),
	.w6(32'hbb6a2fb4),
	.w7(32'hb9277a1b),
	.w8(32'hbb7e75e0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04f886),
	.w1(32'hbb7e4e8f),
	.w2(32'hbbcf3ac6),
	.w3(32'h3b879838),
	.w4(32'hbb2a7146),
	.w5(32'h3a4f1722),
	.w6(32'h39e093be),
	.w7(32'h3ad74357),
	.w8(32'h3b24a3f3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d9e2),
	.w1(32'h3ba7465b),
	.w2(32'h3b3d1b54),
	.w3(32'hbabf9b63),
	.w4(32'h3b87b151),
	.w5(32'h3ad0564b),
	.w6(32'hb8350058),
	.w7(32'h3b6c24c6),
	.w8(32'h3a35da74),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42cd6b),
	.w1(32'hb9eeddc8),
	.w2(32'hbbf8740c),
	.w3(32'hbbe57797),
	.w4(32'h3aa0bb75),
	.w5(32'hbb5079c5),
	.w6(32'hbc1de731),
	.w7(32'h3b2a09d0),
	.w8(32'h3b83ffd7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0c798),
	.w1(32'hb9005c41),
	.w2(32'hbac7bbbe),
	.w3(32'hba749d4e),
	.w4(32'hba3ca100),
	.w5(32'h39e1c162),
	.w6(32'h39fd93ab),
	.w7(32'hbafc4b6d),
	.w8(32'hbc00108f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2a760),
	.w1(32'hbb59678e),
	.w2(32'hbb95d599),
	.w3(32'hbb8e9238),
	.w4(32'h3b420dcc),
	.w5(32'hbaf46489),
	.w6(32'hbbe545a8),
	.w7(32'h3b8e709c),
	.w8(32'h3ab930b3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cf339),
	.w1(32'h3ac660be),
	.w2(32'hbaadfd09),
	.w3(32'h3b3ba1cc),
	.w4(32'hbaf43b8f),
	.w5(32'h3a7d49ec),
	.w6(32'h3b02494e),
	.w7(32'hbba9afcf),
	.w8(32'hbb4bbbb1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f5e3),
	.w1(32'hbbb3e4fa),
	.w2(32'h38e4c2bf),
	.w3(32'h3bd03e28),
	.w4(32'hbb24d563),
	.w5(32'hbb9af07f),
	.w6(32'h3b65e47a),
	.w7(32'h3ace6247),
	.w8(32'hbb194b6e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd0bab),
	.w1(32'hbb738903),
	.w2(32'h399f2dc3),
	.w3(32'hbc4c2294),
	.w4(32'hbba3ac8a),
	.w5(32'h3bb8f324),
	.w6(32'hbc000806),
	.w7(32'h3ab4459a),
	.w8(32'hba5307bb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af22f79),
	.w1(32'h3c15cf8a),
	.w2(32'hbb819244),
	.w3(32'h3c16d3d9),
	.w4(32'h3c7432ca),
	.w5(32'h3c8fb85d),
	.w6(32'h3c01d169),
	.w7(32'h3c1bae57),
	.w8(32'h3b9c2e5c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a3344),
	.w1(32'hbb43754d),
	.w2(32'hbc2b2d7f),
	.w3(32'h3c95aff9),
	.w4(32'hb9f7160c),
	.w5(32'hbb304a6f),
	.w6(32'h3c7b993a),
	.w7(32'h3bca3993),
	.w8(32'hb9bb47f3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc199ba9),
	.w1(32'hbc1df6e8),
	.w2(32'hbc3a68bb),
	.w3(32'hbb21cb55),
	.w4(32'hbc2c6e04),
	.w5(32'hbbcf9a89),
	.w6(32'hbb855b94),
	.w7(32'hbbf61813),
	.w8(32'hbadc36e0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7be1ec),
	.w1(32'hbbb585ae),
	.w2(32'h3962a99d),
	.w3(32'h3b4da543),
	.w4(32'hbb963133),
	.w5(32'hb9d3c414),
	.w6(32'hbb5b1bef),
	.w7(32'hbbce9a2c),
	.w8(32'hbab717b6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a7286),
	.w1(32'h3a44d089),
	.w2(32'h3b1564ee),
	.w3(32'hbb82fe73),
	.w4(32'h3c11055d),
	.w5(32'h3b1a1ad7),
	.w6(32'h3c130109),
	.w7(32'h3b831547),
	.w8(32'hb9b7dda2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3159f),
	.w1(32'h3b9154b2),
	.w2(32'h3b79fc8e),
	.w3(32'h3b98a1a9),
	.w4(32'h3b204bd7),
	.w5(32'h3c025dc5),
	.w6(32'hbb8b7e0f),
	.w7(32'h3bc01bc2),
	.w8(32'h3c6ef6ab),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bbe05),
	.w1(32'hbb2b3896),
	.w2(32'hbbbf8cd2),
	.w3(32'hbadfb493),
	.w4(32'hba569b9c),
	.w5(32'hbb0b1541),
	.w6(32'h3c0324dd),
	.w7(32'h3ab2149e),
	.w8(32'h3bf5ca3b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffb06e),
	.w1(32'hba504f89),
	.w2(32'hbb9d761e),
	.w3(32'hbbadfff1),
	.w4(32'hb9fb2444),
	.w5(32'hbb99d088),
	.w6(32'hba2f8b29),
	.w7(32'h3a670520),
	.w8(32'hbb1b1505),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2f1d5),
	.w1(32'h3b882d44),
	.w2(32'h3b9b7bce),
	.w3(32'hbc0da5de),
	.w4(32'h3b914229),
	.w5(32'h3c1ea642),
	.w6(32'hbbd4e284),
	.w7(32'hb95c37b4),
	.w8(32'h3ba1bafb),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5f6ba),
	.w1(32'h3ac4b93d),
	.w2(32'h3b96389d),
	.w3(32'hbb6aff80),
	.w4(32'h3bbd7e4a),
	.w5(32'h3c5e054a),
	.w6(32'hbaec1f4e),
	.w7(32'h3b4db8f5),
	.w8(32'h3c132317),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a735643),
	.w1(32'h39b180dd),
	.w2(32'hbaa6129b),
	.w3(32'h3b8201d3),
	.w4(32'h3b40a0c6),
	.w5(32'hbade41f9),
	.w6(32'h3babdf1c),
	.w7(32'h3b77c926),
	.w8(32'hbb4e34d1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb428e93),
	.w1(32'h3c0208eb),
	.w2(32'h3b6defd4),
	.w3(32'hbc37d03d),
	.w4(32'h3bbf7538),
	.w5(32'hbaf7af12),
	.w6(32'hbc16ada6),
	.w7(32'hb92acc40),
	.w8(32'h3a2641d6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91a699),
	.w1(32'hbc497038),
	.w2(32'hb8786c28),
	.w3(32'hbc2f7ff7),
	.w4(32'hb9705212),
	.w5(32'hbb90f8b2),
	.w6(32'h3b2cdf70),
	.w7(32'hbb863cbc),
	.w8(32'hb96f7dde),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca06f26),
	.w1(32'hbc476185),
	.w2(32'h3be2bee6),
	.w3(32'hbce20fc0),
	.w4(32'hbc3fd73b),
	.w5(32'h3baf6867),
	.w6(32'hbd058b10),
	.w7(32'hbc26cbe3),
	.w8(32'h3a8809b0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b456e20),
	.w1(32'h3c0ad6e3),
	.w2(32'h3b0e4ef4),
	.w3(32'h3bed9197),
	.w4(32'h3b35ab17),
	.w5(32'h3c6b881d),
	.w6(32'h3c2ea0cb),
	.w7(32'h3c2c2e05),
	.w8(32'h3c84c5fa),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc359b15),
	.w1(32'hbc6342f4),
	.w2(32'hbc40374b),
	.w3(32'hbc1ef02e),
	.w4(32'hbc2a6d31),
	.w5(32'h3c3ab9fe),
	.w6(32'h3b313da2),
	.w7(32'hb8e2ef36),
	.w8(32'h3b0fba57),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38daa9),
	.w1(32'hbc62db5d),
	.w2(32'hbc2f72da),
	.w3(32'hbae52c19),
	.w4(32'hbb6c609c),
	.w5(32'hbba219c4),
	.w6(32'h3b5cd211),
	.w7(32'h3b716657),
	.w8(32'hbadae135),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd6ed52),
	.w1(32'hbbe74928),
	.w2(32'h390f4b32),
	.w3(32'hbc019b29),
	.w4(32'hba838129),
	.w5(32'h38ba0cdb),
	.w6(32'hbbe42a08),
	.w7(32'hbb5dfeb9),
	.w8(32'hbbb3250b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddf70f),
	.w1(32'hbabcc140),
	.w2(32'h3c0e3a83),
	.w3(32'hbc18cdd1),
	.w4(32'hbab57e67),
	.w5(32'h3ac6a6fd),
	.w6(32'hbbc916c5),
	.w7(32'h3b04cc5b),
	.w8(32'h3beae21a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff69f9),
	.w1(32'h3bf92fbc),
	.w2(32'h3af01b15),
	.w3(32'hbb851e6e),
	.w4(32'h3b9d2b09),
	.w5(32'hbb3e76aa),
	.w6(32'hb935517c),
	.w7(32'h3aeece1b),
	.w8(32'hbbf10f1b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6afe7d),
	.w1(32'h3a85120c),
	.w2(32'h3aed1043),
	.w3(32'hbbdc3302),
	.w4(32'hbb786ccd),
	.w5(32'hbafad6a1),
	.w6(32'hbc182db7),
	.w7(32'hbbd69766),
	.w8(32'hba562479),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb1f46),
	.w1(32'hbad77b88),
	.w2(32'h3ba2690d),
	.w3(32'hbc14ec0b),
	.w4(32'hbafd4b1b),
	.w5(32'h3b8d57df),
	.w6(32'hbb979f6f),
	.w7(32'h3b4b712f),
	.w8(32'h3c573c1b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84a194),
	.w1(32'h393232b3),
	.w2(32'hbb26369c),
	.w3(32'h3adbc5f4),
	.w4(32'hbc0cedb0),
	.w5(32'hb953a437),
	.w6(32'h3bf80cfa),
	.w7(32'hbbbaa4ed),
	.w8(32'h3c29d138),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08514f),
	.w1(32'hbbd1c089),
	.w2(32'hbb8b9487),
	.w3(32'hbbd4fac1),
	.w4(32'hbb56e9d9),
	.w5(32'hbc4769c5),
	.w6(32'hbadca209),
	.w7(32'hbbb46e6a),
	.w8(32'hbb8dc323),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c8d6d),
	.w1(32'h3a8df2c1),
	.w2(32'hba672038),
	.w3(32'hbc2122eb),
	.w4(32'hbb9dc064),
	.w5(32'hbb14a5e2),
	.w6(32'hbb7b9133),
	.w7(32'hbb6174a4),
	.w8(32'hbb19d8a9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fa3da),
	.w1(32'h3b610b91),
	.w2(32'h3bcf8f55),
	.w3(32'h3aa20e3e),
	.w4(32'h3b562b72),
	.w5(32'h3c6a42e3),
	.w6(32'hbb040dbf),
	.w7(32'h3b2c2fa1),
	.w8(32'h3c86913d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4b7e3),
	.w1(32'hbc4d5d0c),
	.w2(32'hbaff5226),
	.w3(32'hb9b4a799),
	.w4(32'hba833a9a),
	.w5(32'h3c62200f),
	.w6(32'h3b9ba168),
	.w7(32'h3c79d872),
	.w8(32'h3cac67b4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87b992),
	.w1(32'hbb8f1a7f),
	.w2(32'hbb4a60a5),
	.w3(32'h3c5bc418),
	.w4(32'hbb1250da),
	.w5(32'hba4e1a83),
	.w6(32'h3c52e4ce),
	.w7(32'hba92ea31),
	.w8(32'h3bb5b875),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac736e),
	.w1(32'h3b0d3a87),
	.w2(32'h3a811854),
	.w3(32'h3bd46722),
	.w4(32'h39d28b7f),
	.w5(32'h3ace0989),
	.w6(32'h3c10458c),
	.w7(32'h3ae2326e),
	.w8(32'h3b065576),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab02b2e),
	.w1(32'hbb0e54c8),
	.w2(32'h3aace7f0),
	.w3(32'h38e44e4e),
	.w4(32'hba8b6d9a),
	.w5(32'h3bce14c7),
	.w6(32'h3b73b2b9),
	.w7(32'hbb1bb769),
	.w8(32'h3ba3c339),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0386a8),
	.w1(32'h3b71106d),
	.w2(32'hbbaa5be1),
	.w3(32'h3ab5be05),
	.w4(32'h3b8e8c55),
	.w5(32'hbb0c9b13),
	.w6(32'h3b4bbc19),
	.w7(32'h3c35288e),
	.w8(32'h3c2e428a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d46b2),
	.w1(32'h3b9b4bb4),
	.w2(32'h3b41f3b8),
	.w3(32'hb969fb01),
	.w4(32'h3bf24902),
	.w5(32'h3c834ec9),
	.w6(32'h3b60b021),
	.w7(32'hba21f03c),
	.w8(32'h3b66f272),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31a1e3),
	.w1(32'hbc019e45),
	.w2(32'hbc180575),
	.w3(32'h3c7a0ab4),
	.w4(32'h394e5a8b),
	.w5(32'h3c3ac0b3),
	.w6(32'h3bfb0b10),
	.w7(32'h38da3919),
	.w8(32'h3c1b54e5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc024f93),
	.w1(32'hba24af61),
	.w2(32'hbb98cadd),
	.w3(32'hbc4ed393),
	.w4(32'hbb074274),
	.w5(32'hbb7b8002),
	.w6(32'hbc3f1db5),
	.w7(32'hbb2d2942),
	.w8(32'hbb762a7e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97fc52),
	.w1(32'hbc1daa59),
	.w2(32'hbb3e9557),
	.w3(32'hbb33fd82),
	.w4(32'hbb8fec05),
	.w5(32'h3b6aea63),
	.w6(32'hb9ae8921),
	.w7(32'h3b4f509b),
	.w8(32'h3b99c187),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd31160),
	.w1(32'h3ad41c44),
	.w2(32'hbb3223a5),
	.w3(32'hbb65d5ce),
	.w4(32'h3aa84748),
	.w5(32'h3ba2f0d4),
	.w6(32'hbc0c40eb),
	.w7(32'hbb813e1a),
	.w8(32'hba02f8a9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e38d6),
	.w1(32'h3bc01648),
	.w2(32'h3b6b82ac),
	.w3(32'h3ad4728a),
	.w4(32'hb912e902),
	.w5(32'h3b591403),
	.w6(32'h3bd685e6),
	.w7(32'hba438cc1),
	.w8(32'h3ba7e6b8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe590e),
	.w1(32'h3ba2469e),
	.w2(32'h3b628b4e),
	.w3(32'hbb0e8679),
	.w4(32'hba0adc1e),
	.w5(32'h3bd12b4d),
	.w6(32'h3b48a820),
	.w7(32'h3b3551d1),
	.w8(32'h3c0be971),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be85b18),
	.w1(32'hbb93c26a),
	.w2(32'hbbef8970),
	.w3(32'h3bee862f),
	.w4(32'hbb8825bf),
	.w5(32'hbba71952),
	.w6(32'h3c1a8207),
	.w7(32'h3a6bb6f8),
	.w8(32'h3be11335),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8fc02),
	.w1(32'hb8634e99),
	.w2(32'hbb2a659a),
	.w3(32'h3a231c8e),
	.w4(32'h3a7fc90d),
	.w5(32'hb9f3ce85),
	.w6(32'h3c9b153b),
	.w7(32'h3b91c58f),
	.w8(32'h3b24cc20),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a3ced),
	.w1(32'hbbe0338c),
	.w2(32'hbc0950e5),
	.w3(32'h3add1bfb),
	.w4(32'h3baf4fc4),
	.w5(32'h3b7f459e),
	.w6(32'h3bf87c31),
	.w7(32'h3c1c4f4c),
	.w8(32'h3c1a4bf2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4c04f),
	.w1(32'hbb72a18d),
	.w2(32'hbbd62cba),
	.w3(32'hbac6a586),
	.w4(32'h3ab8f06e),
	.w5(32'h3b2aa9bc),
	.w6(32'h39b41d64),
	.w7(32'h3bce42e9),
	.w8(32'h3c1dbcee),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a422f5e),
	.w1(32'hbc399078),
	.w2(32'hbbe3d1c8),
	.w3(32'hbade6d5f),
	.w4(32'hbc033ae4),
	.w5(32'hba0575af),
	.w6(32'h3b10c5bf),
	.w7(32'hbb10c8dd),
	.w8(32'h39d0a765),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17ab5f),
	.w1(32'hbc196b7a),
	.w2(32'hbabd7775),
	.w3(32'h3ad5b46a),
	.w4(32'hbbd0a0d9),
	.w5(32'h3bc2ae83),
	.w6(32'h3bc0f327),
	.w7(32'hbb18c5c2),
	.w8(32'h3c14ae3f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0d177),
	.w1(32'hbadb7782),
	.w2(32'h3b3b1642),
	.w3(32'h3bb52880),
	.w4(32'h3a924351),
	.w5(32'h3b88d4a9),
	.w6(32'hbaa9c2b5),
	.w7(32'h3b29290f),
	.w8(32'h3b58cb4c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc23ba),
	.w1(32'h3be99bf8),
	.w2(32'h3bb39f82),
	.w3(32'h3c16d8a3),
	.w4(32'h3c08f9b2),
	.w5(32'h3c0463ca),
	.w6(32'h3bc31cfe),
	.w7(32'h3c0c5bcf),
	.w8(32'h3c09835c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c1c05),
	.w1(32'hbb76514c),
	.w2(32'hbc3594ef),
	.w3(32'hbaae60d7),
	.w4(32'hbb8e822c),
	.w5(32'hbbafc042),
	.w6(32'hba83ce83),
	.w7(32'hba1f7402),
	.w8(32'h3a563d39),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc623b2a),
	.w1(32'hbb557aff),
	.w2(32'hbc1bc46c),
	.w3(32'hbc001e09),
	.w4(32'h3b91deb8),
	.w5(32'h3b09155e),
	.w6(32'h3a99c4bf),
	.w7(32'h3aa24542),
	.w8(32'hb9a0e1a9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3a6b0),
	.w1(32'h3c27c9a2),
	.w2(32'h3b9cc961),
	.w3(32'hbbab7319),
	.w4(32'h3ba12aaf),
	.w5(32'h3b477be9),
	.w6(32'hbc5c147a),
	.w7(32'h3b8b2df2),
	.w8(32'h3b35ec5a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f4887),
	.w1(32'hbaf18566),
	.w2(32'hbbbd72e2),
	.w3(32'h3b89959d),
	.w4(32'h3a761d4a),
	.w5(32'hbc5cd81c),
	.w6(32'h3ae79664),
	.w7(32'h3b6874c7),
	.w8(32'hbc2aba99),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80b5f5),
	.w1(32'hba0f9705),
	.w2(32'hbbf3f51b),
	.w3(32'hbc580532),
	.w4(32'h3b548c94),
	.w5(32'hbbb07000),
	.w6(32'hbc394721),
	.w7(32'h3b4254d4),
	.w8(32'hbb3e19a1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d75d9b),
	.w1(32'h3bb82c68),
	.w2(32'h3c4c103e),
	.w3(32'h3b47bdd8),
	.w4(32'h384748f4),
	.w5(32'h3bab3204),
	.w6(32'h3b62c688),
	.w7(32'hbbf66c5b),
	.w8(32'hbc2a9e81),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b025242),
	.w1(32'h3a8a7aa7),
	.w2(32'hba4c6871),
	.w3(32'hbac843f3),
	.w4(32'hba56c053),
	.w5(32'hba1d2a62),
	.w6(32'hbbe52aa3),
	.w7(32'h3b9faef6),
	.w8(32'h3b6e4d0a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a921c03),
	.w1(32'hbad78d37),
	.w2(32'hbb82bb19),
	.w3(32'h3ac045bf),
	.w4(32'hbaa96cba),
	.w5(32'hbb81df78),
	.w6(32'h3b8746d3),
	.w7(32'h3b830b9d),
	.w8(32'hbb60c9d7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24bc00),
	.w1(32'hbbcf55b4),
	.w2(32'hba100639),
	.w3(32'hbbe2f669),
	.w4(32'hbb8ca174),
	.w5(32'hbb442ce3),
	.w6(32'hbb2c0223),
	.w7(32'hbb074db6),
	.w8(32'hbc13a0be),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39742e),
	.w1(32'h3b6e1109),
	.w2(32'hb984bffc),
	.w3(32'h3a848829),
	.w4(32'hba979fba),
	.w5(32'h3b977c1d),
	.w6(32'hbc17d68d),
	.w7(32'hbaaafb3a),
	.w8(32'h3bc656bb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e5faa),
	.w1(32'hba7c45d2),
	.w2(32'hbb4d6cdd),
	.w3(32'hbb2271ee),
	.w4(32'hba1237fa),
	.w5(32'hbbb41e9c),
	.w6(32'h3a062932),
	.w7(32'hb9d364ec),
	.w8(32'hbb2f721a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab03e13),
	.w1(32'hbafd41fc),
	.w2(32'hbb202948),
	.w3(32'hbb8d7f34),
	.w4(32'hbb3947c3),
	.w5(32'hbb6f1030),
	.w6(32'h39b9d447),
	.w7(32'hbbaa1072),
	.w8(32'hbbb6076d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee6d7),
	.w1(32'h3a12eaed),
	.w2(32'h3b81500d),
	.w3(32'hbb8526bd),
	.w4(32'h39966cd2),
	.w5(32'h3b5885e3),
	.w6(32'hbbf5131f),
	.w7(32'h3a2e0abc),
	.w8(32'h3b81b70e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b2326),
	.w1(32'h3899cc15),
	.w2(32'h3b296d3d),
	.w3(32'hbbaf6997),
	.w4(32'h3ade9b8b),
	.w5(32'h3bcf7be4),
	.w6(32'hbbd34eaa),
	.w7(32'h3b760928),
	.w8(32'h3a531200),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4401ed),
	.w1(32'h3b7ad4ad),
	.w2(32'hbba27b8a),
	.w3(32'h3bc0391e),
	.w4(32'h3b8001b6),
	.w5(32'hbb653e47),
	.w6(32'h3c1c458c),
	.w7(32'h3c13237a),
	.w8(32'h3b0a1a86),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd0792),
	.w1(32'hbb00cd94),
	.w2(32'hbb8a4e80),
	.w3(32'hbb071a2e),
	.w4(32'hba9b289d),
	.w5(32'h3a5bd2aa),
	.w6(32'h3b40fbdd),
	.w7(32'h3b579cb2),
	.w8(32'h3ba962ff),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab83855),
	.w1(32'hbb3dca5f),
	.w2(32'hb905faef),
	.w3(32'h3aeee53b),
	.w4(32'hb843dc66),
	.w5(32'h3b141467),
	.w6(32'h3be0f815),
	.w7(32'h3ba8ad02),
	.w8(32'h3bdecd79),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6da697),
	.w1(32'hbb04aa8b),
	.w2(32'h3b1ae04c),
	.w3(32'h3aa42c67),
	.w4(32'h3a985db5),
	.w5(32'hbb243163),
	.w6(32'h3c0e3d58),
	.w7(32'h3b0cc46b),
	.w8(32'h3bb7826a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfb44f),
	.w1(32'h3ad6271b),
	.w2(32'hba39dd98),
	.w3(32'hbb434b9f),
	.w4(32'h3b407925),
	.w5(32'h3a8ee0c8),
	.w6(32'h3b581f54),
	.w7(32'hb9cec75e),
	.w8(32'h3b66b86b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04bcdc),
	.w1(32'h3bfdb1f1),
	.w2(32'h3c015665),
	.w3(32'h3b19494d),
	.w4(32'h3c3258fc),
	.w5(32'h3b99ddb5),
	.w6(32'hb9081261),
	.w7(32'h3c12ce33),
	.w8(32'h3bfce477),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9475b4),
	.w1(32'hbc640f28),
	.w2(32'hbbd5e4d3),
	.w3(32'hbb8a4fea),
	.w4(32'hbc086f39),
	.w5(32'hbbcd7e28),
	.w6(32'hbb8ad97b),
	.w7(32'hbbbfb031),
	.w8(32'hbb9e7847),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7ed84),
	.w1(32'hbb319461),
	.w2(32'h3bcda9e4),
	.w3(32'h3b196585),
	.w4(32'h3bc98342),
	.w5(32'h3b485dbc),
	.w6(32'h3a28e1e6),
	.w7(32'h3bb17476),
	.w8(32'hbaa0b6e6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15b1df),
	.w1(32'hbbd57e40),
	.w2(32'h3a655628),
	.w3(32'hbb20fd42),
	.w4(32'hbaf79306),
	.w5(32'h3c03ae2c),
	.w6(32'hbbf74497),
	.w7(32'hbaadc0de),
	.w8(32'h3b82a8ed),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c58c4),
	.w1(32'hbbe60f41),
	.w2(32'hba937e9b),
	.w3(32'hbc09ac70),
	.w4(32'hbb53429c),
	.w5(32'h38de2ec2),
	.w6(32'hbc03aede),
	.w7(32'hbbca42c7),
	.w8(32'hbbb13cec),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba064ca0),
	.w1(32'h3b777097),
	.w2(32'h3b670318),
	.w3(32'hba0ba87c),
	.w4(32'h3a458a11),
	.w5(32'hb8662d70),
	.w6(32'hba39c541),
	.w7(32'h3a7bacdc),
	.w8(32'h3a91dea7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b652a59),
	.w1(32'hbb633d33),
	.w2(32'hbb80e3a5),
	.w3(32'h3b76e061),
	.w4(32'hbbc23fce),
	.w5(32'hbb759084),
	.w6(32'h3b5033a7),
	.w7(32'hbb63be9e),
	.w8(32'hbb783fd5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42263f),
	.w1(32'h3a047f56),
	.w2(32'hbb19be0d),
	.w3(32'hbb876878),
	.w4(32'h389b9097),
	.w5(32'h3807d7e1),
	.w6(32'hbbc26352),
	.w7(32'hbb9dd7f8),
	.w8(32'hba48bd5f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf34f48),
	.w1(32'hbb9218d7),
	.w2(32'hbbb26ad7),
	.w3(32'hbc06e7ec),
	.w4(32'h3b12492e),
	.w5(32'h39bab2d9),
	.w6(32'hbc0dfb59),
	.w7(32'h3acbb908),
	.w8(32'hbb97bb3b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab60285),
	.w1(32'h3a628c46),
	.w2(32'h3b6c3320),
	.w3(32'hba89c9f3),
	.w4(32'h3aa9d044),
	.w5(32'h3b87b2d4),
	.w6(32'hbb3d5c29),
	.w7(32'hb869efb4),
	.w8(32'hb98a9963),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa8344),
	.w1(32'h3916c30b),
	.w2(32'hbacd21cb),
	.w3(32'h3b15c1db),
	.w4(32'hb986bfcf),
	.w5(32'h3b989f1f),
	.w6(32'hb9ab3b0e),
	.w7(32'h3bf00f53),
	.w8(32'hbac4693c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b250cc8),
	.w1(32'hbb933987),
	.w2(32'h3ade5b65),
	.w3(32'h3b9f8311),
	.w4(32'hbb7cac21),
	.w5(32'hbb0811ee),
	.w6(32'hbb9a30da),
	.w7(32'hbb4a4bc8),
	.w8(32'hbb3daeb4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62be4e4),
	.w1(32'hbc59fa21),
	.w2(32'hbc03407f),
	.w3(32'h3bd5d1fa),
	.w4(32'hbbf77191),
	.w5(32'h3b3fa7ba),
	.w6(32'h3b3cf5c4),
	.w7(32'hbb9290c5),
	.w8(32'hba969f8e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0173ab),
	.w1(32'h3b30c6c0),
	.w2(32'hbae7cb9d),
	.w3(32'h3abc5506),
	.w4(32'h39a787dd),
	.w5(32'h3ac7c074),
	.w6(32'hba09cacc),
	.w7(32'h3b29e6a7),
	.w8(32'hbbd9ca96),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd474dc),
	.w1(32'h3b87f9e6),
	.w2(32'h3ba9c0ad),
	.w3(32'hbbb2a23f),
	.w4(32'h39c908c2),
	.w5(32'h3ae02694),
	.w6(32'hbc3476d7),
	.w7(32'hb89f01d2),
	.w8(32'h3ba49931),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c014d),
	.w1(32'hbb629059),
	.w2(32'h3abd2899),
	.w3(32'hbc27b687),
	.w4(32'hbb45f6dd),
	.w5(32'h3b11462c),
	.w6(32'hbc10ca29),
	.w7(32'hbb5908e6),
	.w8(32'hbb6ff8d3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b3477),
	.w1(32'hbba60f2a),
	.w2(32'hbbdd46a6),
	.w3(32'hbb5d758a),
	.w4(32'h38e37db4),
	.w5(32'h3c49726d),
	.w6(32'hbb936352),
	.w7(32'h3b8fc564),
	.w8(32'h3c31264d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f8a4b8),
	.w1(32'h3bd05cce),
	.w2(32'h3c15ba16),
	.w3(32'h3b9ea088),
	.w4(32'h3c03e919),
	.w5(32'h3cab0f03),
	.w6(32'h39dde774),
	.w7(32'h3c111e9a),
	.w8(32'h3c833130),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3bcd9),
	.w1(32'hbad4af49),
	.w2(32'hbab09a6f),
	.w3(32'h3a1f3c43),
	.w4(32'hbafa28f6),
	.w5(32'h3b01841f),
	.w6(32'hb98c78b3),
	.w7(32'h3a4ea315),
	.w8(32'h3b545034),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59767b),
	.w1(32'hbb0e7cf0),
	.w2(32'h3b856343),
	.w3(32'h3c0f4d37),
	.w4(32'h3a9ce1ca),
	.w5(32'h3bbfba5d),
	.w6(32'h3c575705),
	.w7(32'h3b34cfc3),
	.w8(32'h3bb25098),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb67a4d),
	.w1(32'h3bc4dc3f),
	.w2(32'h3a77011b),
	.w3(32'hbbb788b1),
	.w4(32'h3c0d7c88),
	.w5(32'h3be22c61),
	.w6(32'hbc1ad7b7),
	.w7(32'h3bfab5f3),
	.w8(32'h3c6d29ff),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908eaf1),
	.w1(32'hb9b7a9b7),
	.w2(32'hbb99f8c1),
	.w3(32'hba647ad7),
	.w4(32'h3a15297c),
	.w5(32'hbb98c3cb),
	.w6(32'h3b6208e4),
	.w7(32'h3af6d0f0),
	.w8(32'hb9f2a8f9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1bd0a),
	.w1(32'h3b5e5b27),
	.w2(32'hbc198282),
	.w3(32'hbb4f0f7d),
	.w4(32'h3a36cc6a),
	.w5(32'hbbfe00f9),
	.w6(32'h3a9a6577),
	.w7(32'h3b697ee5),
	.w8(32'hbae6f655),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f5184),
	.w1(32'h3a9c87b0),
	.w2(32'h3b376b9b),
	.w3(32'hbbe726df),
	.w4(32'h3c0993f1),
	.w5(32'h3bbf4d0e),
	.w6(32'hb80f73bb),
	.w7(32'h3bb2a154),
	.w8(32'h3a0aca71),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e7119),
	.w1(32'h3b796de1),
	.w2(32'hbba4acee),
	.w3(32'hbc3a4f01),
	.w4(32'h3b8557cd),
	.w5(32'hbb1af825),
	.w6(32'hbc779377),
	.w7(32'h3b468831),
	.w8(32'hbaa62a9c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb94401),
	.w1(32'hba6bb75d),
	.w2(32'hbba7a863),
	.w3(32'h3bcd1598),
	.w4(32'hbb662917),
	.w5(32'h3ab08a86),
	.w6(32'h3ba433f9),
	.w7(32'hbbdd68f7),
	.w8(32'h3b75c9fa),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac25b88),
	.w1(32'h3be08033),
	.w2(32'h39c9144e),
	.w3(32'hbb30cb9c),
	.w4(32'h3b9271c5),
	.w5(32'h3c057c70),
	.w6(32'h3a4f2b22),
	.w7(32'h3b77dc28),
	.w8(32'h3b96d668),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeabc00),
	.w1(32'h3ba73f05),
	.w2(32'h3bbcc25c),
	.w3(32'h3b223a73),
	.w4(32'hba09f7ae),
	.w5(32'hba90f038),
	.w6(32'hbafb3451),
	.w7(32'h3b6cb1a9),
	.w8(32'hba609d88),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe58d47),
	.w1(32'h3c1d8c18),
	.w2(32'h3b0c1cf5),
	.w3(32'hbc467cb1),
	.w4(32'h3bbc8de6),
	.w5(32'h3bb9d7c9),
	.w6(32'hbbef75f8),
	.w7(32'hbac7c7d7),
	.w8(32'hba34ad61),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5ee79),
	.w1(32'h3bfc8ea3),
	.w2(32'h37ee84f2),
	.w3(32'h3c074045),
	.w4(32'h3bfd79bf),
	.w5(32'h3acf26d7),
	.w6(32'h3ad09602),
	.w7(32'h3c605bec),
	.w8(32'hbaf48306),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83d735),
	.w1(32'h3c07c850),
	.w2(32'h3b0001da),
	.w3(32'h3bfc34e0),
	.w4(32'h3b8a1d7b),
	.w5(32'h3b9a0e0f),
	.w6(32'h3b5ddbbb),
	.w7(32'h3b212a0c),
	.w8(32'hbb0de750),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae22313),
	.w1(32'hbb8ad720),
	.w2(32'hbb2cb16f),
	.w3(32'h3bb44867),
	.w4(32'h3a45c90d),
	.w5(32'h3b48a1f7),
	.w6(32'h3b8f553e),
	.w7(32'h3c0fc87f),
	.w8(32'h3ba7f529),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a5182),
	.w1(32'hbaf558d4),
	.w2(32'h3b8dbe24),
	.w3(32'h3bc5d13a),
	.w4(32'h3a3e9430),
	.w5(32'h3bba29f4),
	.w6(32'h3b9c3533),
	.w7(32'hbb82f794),
	.w8(32'h3ad13f8e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a4732),
	.w1(32'hbba7927a),
	.w2(32'h3a3f4a5e),
	.w3(32'hbbca6012),
	.w4(32'hbbaddb2d),
	.w5(32'hbb2b0d66),
	.w6(32'hbb034d6c),
	.w7(32'hbbd06d60),
	.w8(32'hbb89ff36),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb595884),
	.w1(32'h3aa24f06),
	.w2(32'hbc05e7bb),
	.w3(32'hbb385f42),
	.w4(32'h3bf205d3),
	.w5(32'h387c17d2),
	.w6(32'hbb979997),
	.w7(32'h3c29fe6c),
	.w8(32'h3b7b4884),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca38481),
	.w1(32'h3b8eed4f),
	.w2(32'hbc29a5fe),
	.w3(32'hb8b9d060),
	.w4(32'h3bfb555d),
	.w5(32'hba08c03e),
	.w6(32'h3c5f7184),
	.w7(32'h3c6b4f89),
	.w8(32'h3c7f5ec3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc092080),
	.w1(32'h3bb61367),
	.w2(32'h3aaf497d),
	.w3(32'hbc0fa719),
	.w4(32'h3c27f6c5),
	.w5(32'h3b6f5d31),
	.w6(32'hbc87084d),
	.w7(32'h39fd25c5),
	.w8(32'hba68288b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03c5a0),
	.w1(32'hbb277dcd),
	.w2(32'h3b3f0328),
	.w3(32'hbb52c26b),
	.w4(32'hb9f56641),
	.w5(32'h3c2e3ad4),
	.w6(32'hbbff3ae7),
	.w7(32'h3a93be59),
	.w8(32'h3c9a1733),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3291ab),
	.w1(32'hbb8c89d9),
	.w2(32'hbb90730a),
	.w3(32'h3a2c2751),
	.w4(32'hbb9dac60),
	.w5(32'hba54d0dd),
	.w6(32'h3bfee79e),
	.w7(32'hbc058a21),
	.w8(32'hba89511f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b366845),
	.w1(32'h3b23f19a),
	.w2(32'h3b3baf5e),
	.w3(32'h3be7b1f7),
	.w4(32'h3b24f24e),
	.w5(32'h3b7252a6),
	.w6(32'h3bfc1d95),
	.w7(32'h3b1e2f7b),
	.w8(32'h3b24719f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b641054),
	.w1(32'h3c142249),
	.w2(32'h3bc3f045),
	.w3(32'h3adc061b),
	.w4(32'h3bcc2dbb),
	.w5(32'hbb0890e5),
	.w6(32'h3b5b8f48),
	.w7(32'h3b78275e),
	.w8(32'hbbb98f05),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3b60b),
	.w1(32'h3b479ee4),
	.w2(32'h3b0eaa90),
	.w3(32'hbbf80ae4),
	.w4(32'hb7cdc127),
	.w5(32'h3b9a9449),
	.w6(32'hbc29a95b),
	.w7(32'hbb141d2b),
	.w8(32'h3bc1bde2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab577b2),
	.w1(32'hbc62cbb4),
	.w2(32'hbc857279),
	.w3(32'hbb435740),
	.w4(32'hbc2414e9),
	.w5(32'hbc2949b4),
	.w6(32'hbbb20e88),
	.w7(32'hbb133e4d),
	.w8(32'h3a9a7997),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e8311),
	.w1(32'hbb9665d5),
	.w2(32'hbb1c4674),
	.w3(32'hbb858384),
	.w4(32'h39430bfa),
	.w5(32'h3b09043b),
	.w6(32'hbb126855),
	.w7(32'hba90ba48),
	.w8(32'h3c0a661f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffff5d),
	.w1(32'hbb9c300b),
	.w2(32'hbb268fa4),
	.w3(32'h3b504de1),
	.w4(32'h3af5b5e1),
	.w5(32'h3b5e1bc0),
	.w6(32'h3bea3790),
	.w7(32'h3aa38d49),
	.w8(32'h3b54add2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41b630),
	.w1(32'h3ba8ad4d),
	.w2(32'hba9c6c49),
	.w3(32'hb9f85095),
	.w4(32'hb93af080),
	.w5(32'h3a831908),
	.w6(32'h3acf0219),
	.w7(32'h3b5f5d64),
	.w8(32'h3bad2a14),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984ce9a),
	.w1(32'hbc17df1f),
	.w2(32'hbb7ca652),
	.w3(32'hb95b0037),
	.w4(32'hbb9a1095),
	.w5(32'hba9042b9),
	.w6(32'h3ba2f95d),
	.w7(32'h3aa1e76a),
	.w8(32'h3a7a3db2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9afa56),
	.w1(32'h3b09fefa),
	.w2(32'h3c3fcd6b),
	.w3(32'hbb904ff9),
	.w4(32'h3ad6c82b),
	.w5(32'h3c71005b),
	.w6(32'hba9867a7),
	.w7(32'hbbc3b415),
	.w8(32'h3ba315cc),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4fe82),
	.w1(32'hbbee0408),
	.w2(32'hbb130290),
	.w3(32'h3b1d1ae5),
	.w4(32'hbc294936),
	.w5(32'hbb92939f),
	.w6(32'hbbb457da),
	.w7(32'hbc3fef0a),
	.w8(32'hbb667047),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40f308),
	.w1(32'h3aa8f4c6),
	.w2(32'h3a8f1de4),
	.w3(32'hbc03aa20),
	.w4(32'hba575c39),
	.w5(32'h3b139f8f),
	.w6(32'hbb1b87b1),
	.w7(32'h3af0e50c),
	.w8(32'h3b76830d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306e02),
	.w1(32'hbbd77519),
	.w2(32'h3c2677b4),
	.w3(32'hba295d78),
	.w4(32'hbb724525),
	.w5(32'h3c9ce208),
	.w6(32'h3accc937),
	.w7(32'hbbeb6e15),
	.w8(32'h3cafa8b1),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cc7b1),
	.w1(32'h3a25d221),
	.w2(32'hbacd922f),
	.w3(32'hbbd2fd94),
	.w4(32'h3a57f824),
	.w5(32'hbb6d7bc4),
	.w6(32'hbb0ef64e),
	.w7(32'hbb1f981a),
	.w8(32'hbb7833d7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9c857),
	.w1(32'hbb612f7a),
	.w2(32'hbafbb031),
	.w3(32'hbb66b631),
	.w4(32'hbac3dcda),
	.w5(32'h3b2170e9),
	.w6(32'hbbe70e60),
	.w7(32'hbb43d5e4),
	.w8(32'hb87a42bb),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9330a7),
	.w1(32'hbc4aacec),
	.w2(32'h3b8d5469),
	.w3(32'h3a08c010),
	.w4(32'hbc6a1121),
	.w5(32'h3bd6d9e4),
	.w6(32'hbb3ccb4c),
	.w7(32'hbbb264b7),
	.w8(32'h3c4c6023),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19a9a8),
	.w1(32'hbbae920d),
	.w2(32'hba76236b),
	.w3(32'hbbfbc2a2),
	.w4(32'hbc1189bd),
	.w5(32'hbb5fd414),
	.w6(32'hbc0ecc54),
	.w7(32'hbb5f732d),
	.w8(32'hb97b43f5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6fc66),
	.w1(32'h3a809e41),
	.w2(32'hbaf4a839),
	.w3(32'hbb04aaf1),
	.w4(32'h3bef2ecc),
	.w5(32'h3bd359cf),
	.w6(32'hba0992ca),
	.w7(32'h3c0daf9c),
	.w8(32'h3c3fbc60),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb169e2),
	.w1(32'h3c331942),
	.w2(32'h3bd04be0),
	.w3(32'hbb7099fb),
	.w4(32'h3c14d62a),
	.w5(32'h3ae397e2),
	.w6(32'hb97cc839),
	.w7(32'h3c2902b6),
	.w8(32'h3b4690d3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b958fc1),
	.w1(32'hba0a4e57),
	.w2(32'h3a05dce3),
	.w3(32'hbb83d44b),
	.w4(32'hbb34869b),
	.w5(32'hb94337c2),
	.w6(32'hbc01c7f2),
	.w7(32'hbb38fe76),
	.w8(32'hbab5d486),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003657),
	.w1(32'h3a803f2e),
	.w2(32'h3bb84cfc),
	.w3(32'hbb1a8bfe),
	.w4(32'hba7c90c6),
	.w5(32'h388a5be5),
	.w6(32'hbb173d31),
	.w7(32'hbb5d95be),
	.w8(32'hbb433f8a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d6e63),
	.w1(32'hbb06df97),
	.w2(32'hba47195b),
	.w3(32'hba69c8b4),
	.w4(32'h3b7887cc),
	.w5(32'h3c2e29f8),
	.w6(32'hbbee7ec7),
	.w7(32'h3c24c3aa),
	.w8(32'h3be4c3be),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3951b2),
	.w1(32'h3a610061),
	.w2(32'hbb3894dc),
	.w3(32'hbb310e3c),
	.w4(32'h3b4fd9e8),
	.w5(32'h3c1f4e1c),
	.w6(32'hbac61021),
	.w7(32'h3bde5760),
	.w8(32'h3c1b1fca),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe59e7b),
	.w1(32'hbb380270),
	.w2(32'hbb9be969),
	.w3(32'h3abcdf79),
	.w4(32'h3bc07fb5),
	.w5(32'hbba04093),
	.w6(32'hbb06737e),
	.w7(32'h3b3924b8),
	.w8(32'hbaa8dc75),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb473a29),
	.w1(32'hbbe61ae2),
	.w2(32'hbb98a06c),
	.w3(32'hbb814e3b),
	.w4(32'hbb122805),
	.w5(32'h3b1be40e),
	.w6(32'hbab97f53),
	.w7(32'h3bd608b5),
	.w8(32'h3c1d26c0),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1f127),
	.w1(32'hbc3b3c6b),
	.w2(32'h3a85639c),
	.w3(32'hbbdd4e62),
	.w4(32'hbbdea9e7),
	.w5(32'h3c15c1e6),
	.w6(32'hb9a67b6b),
	.w7(32'hbb58b625),
	.w8(32'h3c5f09c9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc357b7f),
	.w1(32'hbb8039e3),
	.w2(32'hbb75eb11),
	.w3(32'hbb65f0fa),
	.w4(32'hbbe17f56),
	.w5(32'h3b5f4593),
	.w6(32'h3b83ee90),
	.w7(32'hb9f74673),
	.w8(32'h3b327b65),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc364136),
	.w1(32'hbc840a2a),
	.w2(32'hbb6fb57f),
	.w3(32'hbbb505ef),
	.w4(32'hbb8153a5),
	.w5(32'h3bbf5866),
	.w6(32'hbacbe1ef),
	.w7(32'hbb34a5bc),
	.w8(32'h3b04680a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b9df5),
	.w1(32'hbbd1a3fc),
	.w2(32'hbc624691),
	.w3(32'h3b2fd8ba),
	.w4(32'hba09730f),
	.w5(32'hbb2560b7),
	.w6(32'hbb9063b8),
	.w7(32'h3bfb414c),
	.w8(32'h3b90d5c7),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9387cc),
	.w1(32'hbbf2707b),
	.w2(32'hbb46c51b),
	.w3(32'hbc00b2e6),
	.w4(32'h3b357ba0),
	.w5(32'h3baa7222),
	.w6(32'hbbf3ae1f),
	.w7(32'hbb53761a),
	.w8(32'hbb972cdc),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03f9f8),
	.w1(32'hbb8142ec),
	.w2(32'h3b67c87f),
	.w3(32'h3b8be5bc),
	.w4(32'h3a275426),
	.w5(32'h3b9cdb71),
	.w6(32'hbb8fdd0c),
	.w7(32'hbb783aad),
	.w8(32'h3b6c9458),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba138539),
	.w1(32'h3a837142),
	.w2(32'hbb2e450b),
	.w3(32'hba24ab7d),
	.w4(32'hbabdfde7),
	.w5(32'hbbc06ee3),
	.w6(32'hbc26f9d3),
	.w7(32'hbb24293d),
	.w8(32'hbbef5cc8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4638c5),
	.w1(32'hb9ff983c),
	.w2(32'h3b0efb03),
	.w3(32'hbbc2831b),
	.w4(32'h3af1c6de),
	.w5(32'h3aef9c48),
	.w6(32'hbbdc110b),
	.w7(32'h3b72a978),
	.w8(32'h3be5a08f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5fca4),
	.w1(32'hbb631623),
	.w2(32'hbbd0aeb3),
	.w3(32'h3b2089c8),
	.w4(32'hbb9f1b2f),
	.w5(32'h3b1650a4),
	.w6(32'h3bb8d757),
	.w7(32'hbc29b23e),
	.w8(32'hba4284ff),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3614ac),
	.w1(32'h399db6d9),
	.w2(32'hba5c2c28),
	.w3(32'h3c9ae921),
	.w4(32'h3b06c838),
	.w5(32'h3b0b82ba),
	.w6(32'h3c83e898),
	.w7(32'hbae57ba6),
	.w8(32'h3bb3cb36),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb606589),
	.w1(32'h3b13ab8c),
	.w2(32'h3b83c731),
	.w3(32'h3b1e2340),
	.w4(32'h3b88d01d),
	.w5(32'h3ab9f1bd),
	.w6(32'h3b1ba333),
	.w7(32'h3b996856),
	.w8(32'h3b6e3997),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e34a4),
	.w1(32'hbc0f3d89),
	.w2(32'hbc0fe3b2),
	.w3(32'hbb0513b1),
	.w4(32'hbc312b27),
	.w5(32'hbc43b489),
	.w6(32'hbad62438),
	.w7(32'hbbc832a6),
	.w8(32'hbb4e641b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8964ad),
	.w1(32'hbb8a84ce),
	.w2(32'hbbe6b25c),
	.w3(32'hbbdfce8a),
	.w4(32'h3b7cadab),
	.w5(32'hbb05878c),
	.w6(32'hbbafa9eb),
	.w7(32'h3b1a73f0),
	.w8(32'h3b0f248f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36b2a8),
	.w1(32'h3a22e146),
	.w2(32'h3b61d4eb),
	.w3(32'hbb929f87),
	.w4(32'hbb3c9702),
	.w5(32'h3b3d54c5),
	.w6(32'hbbb0b4a3),
	.w7(32'h3a305755),
	.w8(32'h3b87b433),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8380a0),
	.w1(32'hbc4cf360),
	.w2(32'hba94d57b),
	.w3(32'h3b4f4cb0),
	.w4(32'hba48389f),
	.w5(32'h3c82527d),
	.w6(32'h3badb6dc),
	.w7(32'hbbc7d663),
	.w8(32'h3bc437d7),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60c8f5),
	.w1(32'hbc80702a),
	.w2(32'hba80effe),
	.w3(32'h3c73f842),
	.w4(32'hbb8a1655),
	.w5(32'h3bc82f2d),
	.w6(32'h3b94fc30),
	.w7(32'hbbf44062),
	.w8(32'h3bc9d701),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36648e),
	.w1(32'h3b2c13a3),
	.w2(32'h3b2d9adc),
	.w3(32'h3b83a648),
	.w4(32'h3b894ed9),
	.w5(32'h3c60c097),
	.w6(32'h3be4be20),
	.w7(32'h3aba084f),
	.w8(32'h3bccb7dc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e74ec),
	.w1(32'h39999a6a),
	.w2(32'h3c129556),
	.w3(32'h3c20fc91),
	.w4(32'h3a895ed3),
	.w5(32'h3c05fd04),
	.w6(32'hbb07c325),
	.w7(32'hbb47df65),
	.w8(32'hb98bcb16),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3d475),
	.w1(32'hbba1aed3),
	.w2(32'hbbdbee45),
	.w3(32'h3b058510),
	.w4(32'hbb9359cc),
	.w5(32'hbb627994),
	.w6(32'hbbd0c517),
	.w7(32'hbb35c601),
	.w8(32'hba9fa243),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacefa1d),
	.w1(32'h3abfa237),
	.w2(32'hbab83f01),
	.w3(32'hb849792e),
	.w4(32'hbac7da79),
	.w5(32'hbc3ad2e8),
	.w6(32'hbb7c2dd8),
	.w7(32'h3a1ed6cd),
	.w8(32'hbbcc0135),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43639f),
	.w1(32'h3b8bb1f9),
	.w2(32'h3bc62866),
	.w3(32'hbc05bc44),
	.w4(32'hba9244ed),
	.w5(32'h3c1f19f8),
	.w6(32'hbb433c29),
	.w7(32'hbb409f99),
	.w8(32'h3ace710f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d7221),
	.w1(32'hbaa043b6),
	.w2(32'h3ba94baf),
	.w3(32'h3c049ae5),
	.w4(32'hbb10d954),
	.w5(32'h3b927dda),
	.w6(32'h3b451941),
	.w7(32'hb868c5f2),
	.w8(32'h3aeaf067),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfd425),
	.w1(32'hbc52b2ba),
	.w2(32'h3b11e393),
	.w3(32'h3c21e312),
	.w4(32'h3b7d189f),
	.w5(32'h3cafa762),
	.w6(32'h3b1b5e8d),
	.w7(32'hbbdbf0f4),
	.w8(32'h3b3e729e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fdccb),
	.w1(32'hbaea5d65),
	.w2(32'h3bb7827a),
	.w3(32'h3cc015b2),
	.w4(32'hb75bffd4),
	.w5(32'hbbba80b8),
	.w6(32'hbbf463ad),
	.w7(32'hbbf218a1),
	.w8(32'hbbab5de7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd31a7),
	.w1(32'hbb9a098a),
	.w2(32'hbc27f715),
	.w3(32'hbbc91341),
	.w4(32'hbb7f82ce),
	.w5(32'hbc4c722b),
	.w6(32'hba56b211),
	.w7(32'hbb643cac),
	.w8(32'hbba3c7bc),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21958f),
	.w1(32'hbaf55f71),
	.w2(32'hba52be70),
	.w3(32'hbb035534),
	.w4(32'h3b39a5e1),
	.w5(32'h3ae57713),
	.w6(32'hbb420e40),
	.w7(32'h3b4fb107),
	.w8(32'h3b829c1a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc071f67),
	.w1(32'hbc08252e),
	.w2(32'hbc23b24d),
	.w3(32'h3b98ef0b),
	.w4(32'h3ab33fb8),
	.w5(32'h3b68a21e),
	.w6(32'h3a9a4bef),
	.w7(32'hba9fe9f9),
	.w8(32'h3c2339f4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7c609),
	.w1(32'hbb248b37),
	.w2(32'hba1afe60),
	.w3(32'h3a979e7f),
	.w4(32'h3b49c980),
	.w5(32'hba13799a),
	.w6(32'h3ba1dcd0),
	.w7(32'hbb7add43),
	.w8(32'hbb347a29),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46e1dd),
	.w1(32'hba97e9ab),
	.w2(32'hb8c3e0c8),
	.w3(32'hb8a84242),
	.w4(32'hbb4099bf),
	.w5(32'h3c15ffc6),
	.w6(32'hbb3f4dee),
	.w7(32'hbaeb4bc7),
	.w8(32'h3bd25c27),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58b2a7),
	.w1(32'hbb4afafa),
	.w2(32'hbbe40e04),
	.w3(32'h3bfb746d),
	.w4(32'h39ffe685),
	.w5(32'hbbb83555),
	.w6(32'h3bbe8100),
	.w7(32'hb930b46d),
	.w8(32'hbb502e88),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0b8b9),
	.w1(32'h3ba8b1b9),
	.w2(32'hb8d1cfa0),
	.w3(32'h3b1b881a),
	.w4(32'hbad067fa),
	.w5(32'hbc6c24f3),
	.w6(32'hbbcdf71c),
	.w7(32'h3a0d511e),
	.w8(32'hbc07e0fa),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5ef7e),
	.w1(32'hbc24fff0),
	.w2(32'hbbf2b8a5),
	.w3(32'hbc8c2661),
	.w4(32'hbc355eac),
	.w5(32'hba7d9cc3),
	.w6(32'hbc7307cc),
	.w7(32'hbb9b4fff),
	.w8(32'h3c317f22),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b6bfd),
	.w1(32'h39e744c8),
	.w2(32'h3b82046e),
	.w3(32'hba58eaf7),
	.w4(32'h3c0a6990),
	.w5(32'h3b863d35),
	.w6(32'h3bb42467),
	.w7(32'hbac52e54),
	.w8(32'hba807a96),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7795e5),
	.w1(32'hbafa5498),
	.w2(32'hbad4210b),
	.w3(32'hbaeb2cf0),
	.w4(32'hba66f5d4),
	.w5(32'h3b3db924),
	.w6(32'hbbdba98c),
	.w7(32'hbb5f1fce),
	.w8(32'hba853418),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803c30),
	.w1(32'hbb97f648),
	.w2(32'hbb93f2d6),
	.w3(32'hb841d6b6),
	.w4(32'hbb9d86ea),
	.w5(32'h3b0807cd),
	.w6(32'hbb548195),
	.w7(32'hbaf01af9),
	.w8(32'h3a9ed1e3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b988bc5),
	.w1(32'hbbbf883c),
	.w2(32'hbc03a536),
	.w3(32'h3b7c8749),
	.w4(32'hbbc32786),
	.w5(32'hbc6259fe),
	.w6(32'h3b29e640),
	.w7(32'hbbbbb955),
	.w8(32'hbbaf3adf),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ce6cb),
	.w1(32'hbbfce259),
	.w2(32'h3a82c964),
	.w3(32'hbba45e03),
	.w4(32'hbb479379),
	.w5(32'h3b718638),
	.w6(32'hb8963d2f),
	.w7(32'hbba8286e),
	.w8(32'h3b09cff5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44efa1),
	.w1(32'hbb8208f7),
	.w2(32'h3b7d6911),
	.w3(32'h3bbbd896),
	.w4(32'hba61c4f2),
	.w5(32'h3be82b1b),
	.w6(32'hbb86bc5e),
	.w7(32'hbb89270e),
	.w8(32'hb9db3391),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91dd46b),
	.w1(32'hbc329042),
	.w2(32'hbc4c955b),
	.w3(32'h3b1b7161),
	.w4(32'h3b36303b),
	.w5(32'h3c6fb4c0),
	.w6(32'hbc1b09af),
	.w7(32'hbb3ee6ae),
	.w8(32'h3c4f4a31),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1642ba),
	.w1(32'hbb9a0eea),
	.w2(32'hbb745e99),
	.w3(32'h3bd0e0f5),
	.w4(32'h3b1be608),
	.w5(32'h3b4e475e),
	.w6(32'h3b079dc1),
	.w7(32'hbb3abf5c),
	.w8(32'h38c8e78e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a34c8),
	.w1(32'h39de9f0f),
	.w2(32'h3ba7785c),
	.w3(32'hbb4ef1ec),
	.w4(32'hbb87540a),
	.w5(32'h3b30fa64),
	.w6(32'hbb9d6971),
	.w7(32'hbbcd6541),
	.w8(32'hbb3e489a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule