module layer_8_featuremap_216(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85f45f),
	.w1(32'hbbca4d1a),
	.w2(32'hbc61d931),
	.w3(32'h3a2f22a8),
	.w4(32'h3cf6ab99),
	.w5(32'h3c9ecf1f),
	.w6(32'h3c9ab122),
	.w7(32'h3ccf4b93),
	.w8(32'h3c30901d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1d4bc),
	.w1(32'h380dbec6),
	.w2(32'h3b5621fa),
	.w3(32'hbaf1d0fe),
	.w4(32'hba1ec75c),
	.w5(32'hb9b36686),
	.w6(32'hba932e01),
	.w7(32'h39c0101a),
	.w8(32'h3818f2f8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b278208),
	.w1(32'hbaa48af2),
	.w2(32'h3b183c4c),
	.w3(32'hba8d0b6e),
	.w4(32'h3cb429f6),
	.w5(32'h3cc84e3b),
	.w6(32'h3b5f4e81),
	.w7(32'h3c3f4050),
	.w8(32'h3c15317e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2822d),
	.w1(32'h3b1a302a),
	.w2(32'h39b0a9d2),
	.w3(32'h3c1a7d8d),
	.w4(32'h3cd6e5ea),
	.w5(32'h3cc7d023),
	.w6(32'h3bb78185),
	.w7(32'h3c67355f),
	.w8(32'h3c94787b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58c0e0),
	.w1(32'hb9ddc06f),
	.w2(32'hbb88d903),
	.w3(32'h3ca0c5e7),
	.w4(32'h3a96b72d),
	.w5(32'h3a974797),
	.w6(32'hba4362d0),
	.w7(32'hb916d7b5),
	.w8(32'hb9cc33be),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab1ee2),
	.w1(32'hbb77ea5b),
	.w2(32'hbb00ee3a),
	.w3(32'hba39579b),
	.w4(32'hbc14f42d),
	.w5(32'hbc8a7d39),
	.w6(32'hbb215502),
	.w7(32'hbc3750a9),
	.w8(32'hbc93d7cc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aaa92),
	.w1(32'hbadd8ce3),
	.w2(32'hbbb00f7a),
	.w3(32'hb9a0c3da),
	.w4(32'hbb83a8f3),
	.w5(32'hbb9efbac),
	.w6(32'h394b9868),
	.w7(32'hba9d60fb),
	.w8(32'hbb7406d6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb880eb0),
	.w1(32'hbc960808),
	.w2(32'hbcf7fd51),
	.w3(32'hbb8d678e),
	.w4(32'h3d2af228),
	.w5(32'h3d1f9141),
	.w6(32'h3c0816e6),
	.w7(32'h3cab6c93),
	.w8(32'h3ca7066a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb355ee),
	.w1(32'h3ba2dfab),
	.w2(32'hbb102d1e),
	.w3(32'h3ccd4821),
	.w4(32'h3bcbffe0),
	.w5(32'h3b63af55),
	.w6(32'h3a8572d8),
	.w7(32'hb9aaf3af),
	.w8(32'hba6e3433),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52fc02),
	.w1(32'h3aa456e2),
	.w2(32'hbb939464),
	.w3(32'hb904703e),
	.w4(32'hbc487f4b),
	.w5(32'hbc8412c4),
	.w6(32'hbcb26028),
	.w7(32'hbcd64892),
	.w8(32'hbca883d1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe46329),
	.w1(32'hbc05b6cb),
	.w2(32'h39a68a03),
	.w3(32'hb979322a),
	.w4(32'h3a1b4a0e),
	.w5(32'hbc38bec0),
	.w6(32'hbbcaf6b7),
	.w7(32'hbb386ebf),
	.w8(32'hbbe7ec50),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2247b),
	.w1(32'h3a1f2b3f),
	.w2(32'hbab0314e),
	.w3(32'hbbf2e08f),
	.w4(32'h3a8d775b),
	.w5(32'hbbaa5a67),
	.w6(32'h3a989093),
	.w7(32'hbb52507d),
	.w8(32'hb9fcd80f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb846153),
	.w1(32'hbbdff092),
	.w2(32'hb9b938e4),
	.w3(32'hbc193bd5),
	.w4(32'hbb83089a),
	.w5(32'hbc95c95c),
	.w6(32'h3b383698),
	.w7(32'h3a2476cc),
	.w8(32'h3bc59fd2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b139d83),
	.w1(32'h3b9d7875),
	.w2(32'hba8c4f65),
	.w3(32'hbb348afa),
	.w4(32'h3c845c9a),
	.w5(32'h3cbce281),
	.w6(32'h391e2d06),
	.w7(32'h3c15ca7a),
	.w8(32'h39fc4be0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee2a8e),
	.w1(32'hb88fd497),
	.w2(32'hbb14d20b),
	.w3(32'h3cb3c714),
	.w4(32'h3a534904),
	.w5(32'h3afceacd),
	.w6(32'hba24131a),
	.w7(32'h39f26bab),
	.w8(32'h3b1a6478),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ab927),
	.w1(32'h3b45e304),
	.w2(32'h3c1b0333),
	.w3(32'h3b3a6619),
	.w4(32'hbbdab78a),
	.w5(32'hbcc41ebc),
	.w6(32'h3bced04b),
	.w7(32'h3bf98e39),
	.w8(32'hbbe7d586),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d793e),
	.w1(32'h3c868b0b),
	.w2(32'h3cae436a),
	.w3(32'hbc9e72b1),
	.w4(32'hbc466702),
	.w5(32'hbb65265b),
	.w6(32'h3c917563),
	.w7(32'h3c11a661),
	.w8(32'h3b64f1a1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48ebf2),
	.w1(32'h3bd4e3d3),
	.w2(32'h3bc58e14),
	.w3(32'hbb2f34f0),
	.w4(32'h3bda2790),
	.w5(32'h3b3ea2b0),
	.w6(32'h3c9faf5b),
	.w7(32'h3cac3635),
	.w8(32'h3c23f283),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd48f07),
	.w1(32'hbc8b2476),
	.w2(32'hba4abad9),
	.w3(32'hbbd3daf7),
	.w4(32'h3b1c5e70),
	.w5(32'hbad680f5),
	.w6(32'hba8165a5),
	.w7(32'hbb2ad9a7),
	.w8(32'h3aea36db),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb467e44),
	.w1(32'h3b9273bb),
	.w2(32'hb9dc058b),
	.w3(32'hbaa659d7),
	.w4(32'h3a516b14),
	.w5(32'hbb6255b0),
	.w6(32'h3b904ee0),
	.w7(32'h3a19e99c),
	.w8(32'hb98ccd70),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f9581),
	.w1(32'h3b428368),
	.w2(32'hb8d67565),
	.w3(32'hbb8aef54),
	.w4(32'hbc9fd27c),
	.w5(32'hbc583a7e),
	.w6(32'hba131a56),
	.w7(32'hbc756a2c),
	.w8(32'hbc314734),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c3404),
	.w1(32'hbbb38c89),
	.w2(32'h3bb29268),
	.w3(32'hbb95dc7c),
	.w4(32'hbc457749),
	.w5(32'hbc812504),
	.w6(32'hb79cfe4b),
	.w7(32'hbc4b1a64),
	.w8(32'hbc82c28d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74043c),
	.w1(32'h3b4ef6f0),
	.w2(32'h3b94c0d1),
	.w3(32'hbbd34935),
	.w4(32'hbc972156),
	.w5(32'hbc4367b5),
	.w6(32'hbc4096b5),
	.w7(32'hbbba9c18),
	.w8(32'hbaedae8b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ec5f6),
	.w1(32'h3c521d82),
	.w2(32'h3cdeb32f),
	.w3(32'hbc15664b),
	.w4(32'hbb5daa7c),
	.w5(32'hba6f7c11),
	.w6(32'h3bd1f7ca),
	.w7(32'hbbd39fdc),
	.w8(32'h3a864a3e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf90d8),
	.w1(32'h3c2a68ea),
	.w2(32'h3b897566),
	.w3(32'h3c26a53b),
	.w4(32'hbc54c8bc),
	.w5(32'hbc25e061),
	.w6(32'hbbefc4cd),
	.w7(32'hbbc42b3a),
	.w8(32'hba24782b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19b616),
	.w1(32'h3bf058bc),
	.w2(32'hbc17ba26),
	.w3(32'hbaa595ef),
	.w4(32'h3b8b6a60),
	.w5(32'h3b46dac9),
	.w6(32'h3b06753b),
	.w7(32'hbba80083),
	.w8(32'h3c2cdebe),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca5ac5),
	.w1(32'hbc4a295f),
	.w2(32'hbc84b3be),
	.w3(32'hbab3c871),
	.w4(32'h3c90cc69),
	.w5(32'h3c6d66b4),
	.w6(32'h3c205925),
	.w7(32'h3c3d49f7),
	.w8(32'h3b946664),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cafc4),
	.w1(32'hbb396e48),
	.w2(32'hbc7bac61),
	.w3(32'hbc46c779),
	.w4(32'h3abe4ea1),
	.w5(32'hbb65d248),
	.w6(32'hba26cb8a),
	.w7(32'hbbd9f1c5),
	.w8(32'hba609a78),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d241c),
	.w1(32'h3bb9dbe9),
	.w2(32'h3a600cd0),
	.w3(32'h3c15ed76),
	.w4(32'h3be26386),
	.w5(32'hba882833),
	.w6(32'h3a229b1f),
	.w7(32'h3983c3c2),
	.w8(32'hbb6ed7e1),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26c34d),
	.w1(32'hbaa1813f),
	.w2(32'hbbbc16cb),
	.w3(32'hbc0e3ea0),
	.w4(32'h3b79f680),
	.w5(32'h3b4007d1),
	.w6(32'h3ab605b3),
	.w7(32'h3a07a549),
	.w8(32'hbacc1ffc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb27a97),
	.w1(32'hba9e1159),
	.w2(32'hbb84b0f9),
	.w3(32'h39ae8239),
	.w4(32'hbaa7b33e),
	.w5(32'h3a0d42a2),
	.w6(32'h3b089cbe),
	.w7(32'h3b8f76e8),
	.w8(32'h3ba26bde),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb806de2),
	.w1(32'h3bc16579),
	.w2(32'h3c4dd4f3),
	.w3(32'hba894f3a),
	.w4(32'hbc377862),
	.w5(32'hbc57a3ff),
	.w6(32'hbb7aeaba),
	.w7(32'hbc1adb05),
	.w8(32'hbc014ac9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c031ac6),
	.w1(32'hbc8f9447),
	.w2(32'hbcdfaf01),
	.w3(32'hbc7da1e0),
	.w4(32'hbbc81326),
	.w5(32'hbbec6519),
	.w6(32'hbbb1beed),
	.w7(32'h3a426cce),
	.w8(32'hba91a620),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb294dd),
	.w1(32'h3b110847),
	.w2(32'hbb8b87f3),
	.w3(32'hbc020e3f),
	.w4(32'hbb327bdb),
	.w5(32'hbb8efe83),
	.w6(32'h3b155963),
	.w7(32'h3c546589),
	.w8(32'h3c7755a5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5e029),
	.w1(32'hbb9c6f0c),
	.w2(32'hbc187cf7),
	.w3(32'h3b85d4c9),
	.w4(32'hbb79f929),
	.w5(32'hbb2613bd),
	.w6(32'hba2d9c58),
	.w7(32'hbb25f1fc),
	.w8(32'hbabc1cdf),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01c77a),
	.w1(32'hbbcc54c6),
	.w2(32'hbcaf5f6e),
	.w3(32'hbbc24351),
	.w4(32'h3bccef19),
	.w5(32'h3b76e9a4),
	.w6(32'h3b9cc087),
	.w7(32'h3b166eab),
	.w8(32'h3be824d0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e689f),
	.w1(32'h3b6de3fc),
	.w2(32'h3a692eff),
	.w3(32'hbbd876ab),
	.w4(32'hbab8dc3a),
	.w5(32'hbb4ecaec),
	.w6(32'h3a771c5f),
	.w7(32'hbae923b6),
	.w8(32'h39742bd3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f93854),
	.w1(32'hbb47ebe9),
	.w2(32'hbb349f16),
	.w3(32'hbb0663a7),
	.w4(32'h3b84d5dc),
	.w5(32'h3c0c11f4),
	.w6(32'hbb639138),
	.w7(32'hba8113c4),
	.w8(32'h3bd721dd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e2df),
	.w1(32'hbbada76e),
	.w2(32'h3bff0d03),
	.w3(32'h3c3a537e),
	.w4(32'hbc0f07db),
	.w5(32'hbc814f99),
	.w6(32'hbbee5ff5),
	.w7(32'hbbdc15ce),
	.w8(32'hbbc0c7ab),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00234c),
	.w1(32'h3bcb389f),
	.w2(32'h3c7f6fc9),
	.w3(32'hbc1d45f0),
	.w4(32'hbbb1f908),
	.w5(32'hbb79bd51),
	.w6(32'h3c36bcfd),
	.w7(32'hba9f17fa),
	.w8(32'hbb312776),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2a385),
	.w1(32'h3b6aa078),
	.w2(32'hbb332cd0),
	.w3(32'h3be536e9),
	.w4(32'h3ba55cf3),
	.w5(32'h3a77a1ba),
	.w6(32'hb8d0067e),
	.w7(32'hbaa6e818),
	.w8(32'h3a591992),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb74b3f),
	.w1(32'hbbce1dfc),
	.w2(32'h3b1dd352),
	.w3(32'hbba6cce5),
	.w4(32'h3b199b22),
	.w5(32'hbbbe6bde),
	.w6(32'h385dc5a3),
	.w7(32'h3b520803),
	.w8(32'h3a84c085),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76a407),
	.w1(32'h39a5e725),
	.w2(32'h3c04f30c),
	.w3(32'h3b383523),
	.w4(32'h3a65070e),
	.w5(32'hb98fa629),
	.w6(32'h3b42a0cf),
	.w7(32'h3a9d2675),
	.w8(32'hbbfc1ddb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9950b),
	.w1(32'hbb34aca2),
	.w2(32'hbb27a28c),
	.w3(32'hba99ae84),
	.w4(32'hbb834a7a),
	.w5(32'hba59c5ec),
	.w6(32'h3c05073b),
	.w7(32'h3c7e349c),
	.w8(32'h3b0fa14e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddb289),
	.w1(32'h39510dc1),
	.w2(32'hbb461a96),
	.w3(32'hbbc4ba4a),
	.w4(32'h3bcb9d02),
	.w5(32'h3ce5ad89),
	.w6(32'hbc698c84),
	.w7(32'hbc788c27),
	.w8(32'hbc322c5f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc925ab5),
	.w1(32'h3baf604a),
	.w2(32'h3b27fcf9),
	.w3(32'h3c868b77),
	.w4(32'hbad9278c),
	.w5(32'hbb9d8f8e),
	.w6(32'h3b6d1846),
	.w7(32'h3b5212cc),
	.w8(32'h3aaf8340),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb334b54),
	.w1(32'h3b4dc8fe),
	.w2(32'h3b25d09e),
	.w3(32'hbbd963b7),
	.w4(32'hbba09819),
	.w5(32'hbb9bdc10),
	.w6(32'h3b1c94ed),
	.w7(32'hb9188fa4),
	.w8(32'hbae48da6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a586),
	.w1(32'h3b70daf1),
	.w2(32'h3c3650c8),
	.w3(32'hbbbd566b),
	.w4(32'hbc00af78),
	.w5(32'h3c06288e),
	.w6(32'h3a55cf43),
	.w7(32'hbb3bc203),
	.w8(32'hba8aa6e2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97e771),
	.w1(32'hba8b0aa2),
	.w2(32'hbc41b210),
	.w3(32'hba7929a0),
	.w4(32'hbc02439b),
	.w5(32'hbb58b6fd),
	.w6(32'hbb996408),
	.w7(32'hbcc6cf52),
	.w8(32'hbc44c569),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6258da),
	.w1(32'hbb29a458),
	.w2(32'hbbfc27cd),
	.w3(32'hbbcab650),
	.w4(32'h3bf15085),
	.w5(32'hb776e49a),
	.w6(32'h3bcbde2d),
	.w7(32'h3c4de542),
	.w8(32'h3c5e635b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2519c7),
	.w1(32'h3bc2c487),
	.w2(32'h3bdc351e),
	.w3(32'h3a16d1b2),
	.w4(32'h3b842384),
	.w5(32'h3b62bf99),
	.w6(32'h3aa73ba0),
	.w7(32'h3b47c1a8),
	.w8(32'h3b97cb11),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99dae6),
	.w1(32'hbb65d0f8),
	.w2(32'h3b78d3ae),
	.w3(32'h3a9306fa),
	.w4(32'hb99940b9),
	.w5(32'hb8f6656a),
	.w6(32'hb9abb50b),
	.w7(32'h3b15621e),
	.w8(32'h3a27e37b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5accb0),
	.w1(32'hbb3aeefc),
	.w2(32'h388ffce9),
	.w3(32'hbb4d0dc0),
	.w4(32'hbb793131),
	.w5(32'hba7c2f8b),
	.w6(32'hbb713b00),
	.w7(32'hbb035a64),
	.w8(32'hbab0cf64),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba469a5),
	.w1(32'h3c322125),
	.w2(32'h3c05003f),
	.w3(32'h3b6bde5e),
	.w4(32'h3c4bba46),
	.w5(32'h3ba0e7e1),
	.w6(32'h3bfd9b14),
	.w7(32'h3c2fffa7),
	.w8(32'h3c16cdf2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8e12a),
	.w1(32'hbbb2567a),
	.w2(32'hbc82a43b),
	.w3(32'h3a72bcee),
	.w4(32'h3bb7da4a),
	.w5(32'hba2d755b),
	.w6(32'h3bfd1cb0),
	.w7(32'h3b5f1349),
	.w8(32'h3c19d9c4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1cf73),
	.w1(32'h3bee7a49),
	.w2(32'h3b26685b),
	.w3(32'hba6e673b),
	.w4(32'h3c4aac78),
	.w5(32'hbb566b18),
	.w6(32'h3bfe6e4d),
	.w7(32'h3c8111a5),
	.w8(32'h3c07a367),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00f58a),
	.w1(32'hbc3e4ac9),
	.w2(32'hbc024159),
	.w3(32'hbc0fa1a8),
	.w4(32'hbbe4a13a),
	.w5(32'hbc3c4d7c),
	.w6(32'hbb3d812a),
	.w7(32'hbbc76e72),
	.w8(32'h3b098be2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee63f2),
	.w1(32'h3b1b7c84),
	.w2(32'hbb2f599f),
	.w3(32'hbc05a3bb),
	.w4(32'h3a5caf5c),
	.w5(32'hbb9214f8),
	.w6(32'h3aec0c42),
	.w7(32'hba835785),
	.w8(32'h39ad956d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64ac5c),
	.w1(32'hb9cfa93f),
	.w2(32'h3ad45a1a),
	.w3(32'hbb46d13e),
	.w4(32'h39252385),
	.w5(32'h3a0430d0),
	.w6(32'hbb954737),
	.w7(32'hbb10f69d),
	.w8(32'hbabb1f74),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b963040),
	.w1(32'h3ca87487),
	.w2(32'h3d1f7228),
	.w3(32'h3aff1f6d),
	.w4(32'h3b4c8154),
	.w5(32'hbb6bdb96),
	.w6(32'h3c0d5bcb),
	.w7(32'h3b7d77fc),
	.w8(32'hbb492724),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8c347),
	.w1(32'h3b82a18f),
	.w2(32'hbbeec42d),
	.w3(32'h3b677a05),
	.w4(32'hbc12b93b),
	.w5(32'hbc1369a4),
	.w6(32'hbb70d77b),
	.w7(32'hbc7e20bf),
	.w8(32'hbc079bba),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4730c1),
	.w1(32'h3b83f9c3),
	.w2(32'h3b867008),
	.w3(32'h3b85a090),
	.w4(32'hbc25ba9f),
	.w5(32'hbc0e2e7e),
	.w6(32'hba96da52),
	.w7(32'hbb71ab87),
	.w8(32'hba2c63c7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d61c1),
	.w1(32'h3c364c59),
	.w2(32'h3c2bf631),
	.w3(32'h3a98dbb4),
	.w4(32'h3b6128d3),
	.w5(32'h3a3cfe2a),
	.w6(32'hba7bc876),
	.w7(32'hbb592f35),
	.w8(32'hbad8209f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9729d),
	.w1(32'hba824e67),
	.w2(32'hbb4db8b2),
	.w3(32'h3a634eaa),
	.w4(32'h39627deb),
	.w5(32'hb9fbdca4),
	.w6(32'h3a1fb576),
	.w7(32'hba94ceb5),
	.w8(32'hba626a20),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb880753),
	.w1(32'h3af3e88f),
	.w2(32'h3bc5ada0),
	.w3(32'hbb01ea51),
	.w4(32'hbb22455b),
	.w5(32'hba661d18),
	.w6(32'hbad44dd1),
	.w7(32'h3afaa265),
	.w8(32'h3b294c21),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c217f12),
	.w1(32'h3bec2941),
	.w2(32'h3c82d589),
	.w3(32'h3a0acc14),
	.w4(32'hba760b25),
	.w5(32'h3ba286e6),
	.w6(32'h3b48e76e),
	.w7(32'hbbc6a277),
	.w8(32'h3aeb0802),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c725b64),
	.w1(32'h3ce62180),
	.w2(32'h3cc26aad),
	.w3(32'h3c27712c),
	.w4(32'hbc9961be),
	.w5(32'hbc0856ac),
	.w6(32'h3bd8e29f),
	.w7(32'hbc7906fb),
	.w8(32'hbca658bd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5e42c),
	.w1(32'h3b3528ff),
	.w2(32'hba666ff3),
	.w3(32'h3bcf1296),
	.w4(32'h3c789a3f),
	.w5(32'h3ba552e4),
	.w6(32'h3b9f9a08),
	.w7(32'hb9e6ca70),
	.w8(32'hbb389de0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec3fe4),
	.w1(32'hba3ec60b),
	.w2(32'hbc672c01),
	.w3(32'hbbbf87a8),
	.w4(32'hbb91a99c),
	.w5(32'h3c05d03b),
	.w6(32'h3b1036c0),
	.w7(32'h3cb418d2),
	.w8(32'h3bede867),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d0c12),
	.w1(32'h3b338190),
	.w2(32'hbbcc422a),
	.w3(32'h3baa8498),
	.w4(32'hbc617d3c),
	.w5(32'hbc0956d0),
	.w6(32'hbc51ca3d),
	.w7(32'hbc1b7ac2),
	.w8(32'hbc27a342),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc032f0a),
	.w1(32'hbbd038c2),
	.w2(32'h3b2682a0),
	.w3(32'h3b4f1f0f),
	.w4(32'hbb04a14f),
	.w5(32'h3bdba92f),
	.w6(32'h391b4f5b),
	.w7(32'h3b00c3c9),
	.w8(32'hba08615b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96857b),
	.w1(32'h3bcc4dfd),
	.w2(32'hbb43bd22),
	.w3(32'h3bbbe853),
	.w4(32'h3c61e493),
	.w5(32'h3c86fe7f),
	.w6(32'hbba0c74a),
	.w7(32'h3b19da62),
	.w8(32'h3a8a3aff),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a25ba),
	.w1(32'hbc5cebdc),
	.w2(32'hbc633e54),
	.w3(32'h3a16c671),
	.w4(32'hbb753cb2),
	.w5(32'h3b8847f6),
	.w6(32'hba8a61fe),
	.w7(32'h3ab060e7),
	.w8(32'h3ae15180),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b0b52),
	.w1(32'hba9fe131),
	.w2(32'h3b03faf5),
	.w3(32'h3c0a951f),
	.w4(32'hbb8a2898),
	.w5(32'h3bb6f946),
	.w6(32'h3b30f1c0),
	.w7(32'h3b823b2f),
	.w8(32'h3ad4dd08),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade9b1a),
	.w1(32'h3b9c6818),
	.w2(32'h3b1c711c),
	.w3(32'hbb6d2e1a),
	.w4(32'hbc28c758),
	.w5(32'hbc13c9f6),
	.w6(32'hbac3dcb0),
	.w7(32'hba31847a),
	.w8(32'hbb50c677),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df13de),
	.w1(32'hb9c79c93),
	.w2(32'h3bce3612),
	.w3(32'hbb94819e),
	.w4(32'hbb9ffef3),
	.w5(32'hbc4f538c),
	.w6(32'hbb91d85c),
	.w7(32'h3bd48732),
	.w8(32'h3aca677b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa6a5b),
	.w1(32'h3b7db317),
	.w2(32'h3b5b2921),
	.w3(32'hbb87c9ef),
	.w4(32'hbb081602),
	.w5(32'hbaedad14),
	.w6(32'hb9c15bcf),
	.w7(32'h3982a7b8),
	.w8(32'hbbfc3b5b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b601ce1),
	.w1(32'h3bda0a59),
	.w2(32'h3ba6cd77),
	.w3(32'hbbbf92bb),
	.w4(32'h3bea09af),
	.w5(32'h3b6af9bf),
	.w6(32'h3ae026a3),
	.w7(32'h3b6f9014),
	.w8(32'hba9356f1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07d874),
	.w1(32'hbac17a07),
	.w2(32'hbb1af2c0),
	.w3(32'h3b6bff95),
	.w4(32'h3c1fd4df),
	.w5(32'h3b13adc1),
	.w6(32'h3b0a0708),
	.w7(32'h3c08bec6),
	.w8(32'h3bffa472),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7a58c),
	.w1(32'hbbc9e6df),
	.w2(32'hbc35bb40),
	.w3(32'h3a8266e2),
	.w4(32'hbabeaf5c),
	.w5(32'hbb909d5b),
	.w6(32'hbb192562),
	.w7(32'h3c43f874),
	.w8(32'h3af1fa03),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ce1c9),
	.w1(32'hbc17abfb),
	.w2(32'hbc6f7605),
	.w3(32'hbb553f9c),
	.w4(32'h3bb9e21a),
	.w5(32'h3c4e1f0a),
	.w6(32'h3a3a320d),
	.w7(32'h3afcf9db),
	.w8(32'h3b75b2d4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55c355),
	.w1(32'hbb0c3aca),
	.w2(32'hbc490514),
	.w3(32'h3c15b7cd),
	.w4(32'hba65892f),
	.w5(32'hbac1405c),
	.w6(32'hbc0d2d83),
	.w7(32'h3af07aaf),
	.w8(32'hbb3cd93d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b34f4),
	.w1(32'hb973ddc4),
	.w2(32'h3bcd23b3),
	.w3(32'h3b85fa25),
	.w4(32'hbabf0043),
	.w5(32'hbc1a7ccb),
	.w6(32'h3b061bc4),
	.w7(32'hbb29796f),
	.w8(32'hbc049150),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb9e951),
	.w1(32'h3c4cdcf8),
	.w2(32'h3c946fe2),
	.w3(32'hbb1fead3),
	.w4(32'h3cad909f),
	.w5(32'h3c4209e0),
	.w6(32'h3c450c16),
	.w7(32'hbb79a0b9),
	.w8(32'h3c18bb8b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c953db6),
	.w1(32'hbab176d2),
	.w2(32'hbc2fd6a2),
	.w3(32'h3b08bd42),
	.w4(32'h3c0587e0),
	.w5(32'h3c09125c),
	.w6(32'hbb5973c8),
	.w7(32'h3bc67d25),
	.w8(32'h3b09b9a0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb865b7d),
	.w1(32'hb9f5b3a0),
	.w2(32'hbc8a3290),
	.w3(32'h3bf91127),
	.w4(32'h3c085dab),
	.w5(32'h3c80b117),
	.w6(32'h3c0d0062),
	.w7(32'h3ca83659),
	.w8(32'h3c40ff21),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e4d24),
	.w1(32'hba883f69),
	.w2(32'hbb1167e7),
	.w3(32'h3c539499),
	.w4(32'h3bd0d94a),
	.w5(32'h3b746782),
	.w6(32'hbb0dfc34),
	.w7(32'hbaea63e8),
	.w8(32'hbac77c23),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc812b2),
	.w1(32'h3c22dc35),
	.w2(32'h3be55088),
	.w3(32'h3b690b65),
	.w4(32'hbbfa175f),
	.w5(32'hbc136da2),
	.w6(32'hbbee7870),
	.w7(32'hbc156be7),
	.w8(32'hbba92859),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60397a),
	.w1(32'hbb8cf13c),
	.w2(32'hbc1255a1),
	.w3(32'hbbe1cc83),
	.w4(32'h3be3f177),
	.w5(32'h3b98b132),
	.w6(32'h3b7d6344),
	.w7(32'h3b639268),
	.w8(32'h39eb2465),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc440cac),
	.w1(32'h39b33b2e),
	.w2(32'h39b6fcd8),
	.w3(32'hbb017b40),
	.w4(32'hbbd6c2f1),
	.w5(32'h3beb79ca),
	.w6(32'hbb885563),
	.w7(32'hbb91ef4c),
	.w8(32'h3c2254ed),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c6bab),
	.w1(32'hbc7112bd),
	.w2(32'hbc820ea9),
	.w3(32'hba50d5f6),
	.w4(32'h3c449432),
	.w5(32'h3c7bcb41),
	.w6(32'hba9e008c),
	.w7(32'h3b1d56aa),
	.w8(32'h3bd14c63),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb175a7),
	.w1(32'h3b427359),
	.w2(32'h3b3ff90e),
	.w3(32'h3bb64bb4),
	.w4(32'hbb37b355),
	.w5(32'hbb22346f),
	.w6(32'h3becb1cc),
	.w7(32'h3c03a416),
	.w8(32'h3bc8bfa7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98e434),
	.w1(32'h39a1df9c),
	.w2(32'hbad07676),
	.w3(32'hbbee38db),
	.w4(32'hbb576c02),
	.w5(32'hbb91bbb1),
	.w6(32'h38fe0069),
	.w7(32'hbb4a8c1c),
	.w8(32'hbb68ca12),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf731c0),
	.w1(32'h3aa3e8da),
	.w2(32'h3aad10b4),
	.w3(32'hbb05ef71),
	.w4(32'hbaeb811a),
	.w5(32'hbb5c4d0d),
	.w6(32'h39983a23),
	.w7(32'hbad628b1),
	.w8(32'hbad336f2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b328e07),
	.w1(32'h3ac1041f),
	.w2(32'hbb34e181),
	.w3(32'hb9322e64),
	.w4(32'h3cb56ecd),
	.w5(32'h3c40139b),
	.w6(32'h3b58a825),
	.w7(32'h3b6ee3cb),
	.w8(32'h3c024f70),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a843f23),
	.w1(32'hbb10e19b),
	.w2(32'hbbd3838a),
	.w3(32'hbbd7b475),
	.w4(32'h3b97a92e),
	.w5(32'hbab62b35),
	.w6(32'hba5ab6a3),
	.w7(32'hbaa61453),
	.w8(32'hba6b8262),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb123c85),
	.w1(32'h3bc25748),
	.w2(32'h3c5442dc),
	.w3(32'hbb7b75f0),
	.w4(32'hbbc26367),
	.w5(32'hbc96a6cd),
	.w6(32'hbb2d721e),
	.w7(32'hbaac287d),
	.w8(32'hbbc8695f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6044fd),
	.w1(32'hbc0e08bc),
	.w2(32'h3b8eb877),
	.w3(32'hbcb0030e),
	.w4(32'hba880038),
	.w5(32'hbc7411f0),
	.w6(32'h3b389a66),
	.w7(32'h3b4862f6),
	.w8(32'hbc826902),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc80e8),
	.w1(32'hbbb73ded),
	.w2(32'h3c0a8fa2),
	.w3(32'hbcab0251),
	.w4(32'hbba5e6e7),
	.w5(32'hbc1f05f6),
	.w6(32'h3bdd5713),
	.w7(32'h3afef2ba),
	.w8(32'hbb6150f6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbffaae),
	.w1(32'hbc3ba162),
	.w2(32'hbb2e7648),
	.w3(32'hbc489c21),
	.w4(32'hbc5539f9),
	.w5(32'hbc4fd273),
	.w6(32'hb8ab126e),
	.w7(32'hbc0b0ec0),
	.w8(32'hbc1b0e8d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b046c77),
	.w1(32'h3b482eb2),
	.w2(32'hbbccf821),
	.w3(32'h3ba69a89),
	.w4(32'hbc0fc58e),
	.w5(32'hb910b231),
	.w6(32'hbb110a41),
	.w7(32'h3b6efffe),
	.w8(32'hbbbfb4e2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf96409),
	.w1(32'hbc1bd1df),
	.w2(32'hbc486eb5),
	.w3(32'h3b8e0c70),
	.w4(32'hbb433a60),
	.w5(32'h3b222f11),
	.w6(32'hbc60a64b),
	.w7(32'hbc5d864c),
	.w8(32'hbb0f3446),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5381e8),
	.w1(32'hba2241a9),
	.w2(32'h3b4da345),
	.w3(32'h3c3423b6),
	.w4(32'h3ba4c9a3),
	.w5(32'h3c653381),
	.w6(32'h3bdaa9c0),
	.w7(32'h3c37b964),
	.w8(32'h3b92c9ec),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc278692),
	.w1(32'h3c59cac8),
	.w2(32'h3c83417c),
	.w3(32'h3c390032),
	.w4(32'h3bd6e1b2),
	.w5(32'h3c12bdc2),
	.w6(32'h3b970a52),
	.w7(32'hba840c84),
	.w8(32'h3b4d5eda),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be63d43),
	.w1(32'h3d12f6d6),
	.w2(32'h3d37c60f),
	.w3(32'hbb2023c1),
	.w4(32'h3b0b58db),
	.w5(32'hbb97321f),
	.w6(32'h3c52d2e2),
	.w7(32'h3c558924),
	.w8(32'h3be7799d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb0f68),
	.w1(32'hbb0a10a6),
	.w2(32'hbb6ad161),
	.w3(32'h3924134c),
	.w4(32'hbc21f219),
	.w5(32'hbc36efed),
	.w6(32'hbbadde4f),
	.w7(32'hbb5536e0),
	.w8(32'hbbba409b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f20aa),
	.w1(32'h3be471cc),
	.w2(32'hbb7db7c6),
	.w3(32'hbb8af500),
	.w4(32'h3b92301b),
	.w5(32'h3b21de7d),
	.w6(32'h3b751e12),
	.w7(32'h3b49fc3c),
	.w8(32'h3b84e346),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd889f1),
	.w1(32'h3b29bf64),
	.w2(32'h3a3a9f47),
	.w3(32'hba8da971),
	.w4(32'hbb0663da),
	.w5(32'hbb1bd168),
	.w6(32'hba63ebdb),
	.w7(32'hbb52cb39),
	.w8(32'hbba937b8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe00401),
	.w1(32'hbb91848e),
	.w2(32'hbbd9a907),
	.w3(32'h3a21a3d6),
	.w4(32'h3b97c902),
	.w5(32'h392e23b6),
	.w6(32'hba922dac),
	.w7(32'h3acaa5e4),
	.w8(32'h3b8c5fe6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0b4fb),
	.w1(32'hbb810238),
	.w2(32'h37e4938d),
	.w3(32'hba981e20),
	.w4(32'hbb73b907),
	.w5(32'hbb58eb0f),
	.w6(32'hbb50d357),
	.w7(32'hbb0ffcf9),
	.w8(32'hbb1bc500),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54c5f1),
	.w1(32'h3b5faaab),
	.w2(32'h39b2be9d),
	.w3(32'hba056bd9),
	.w4(32'h3ce43e1d),
	.w5(32'h3d0674fb),
	.w6(32'h3c191f9c),
	.w7(32'h3c8b3b83),
	.w8(32'h3c05ba28),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0095f6),
	.w1(32'h3b23ab12),
	.w2(32'h3aa4ea21),
	.w3(32'h3c03987e),
	.w4(32'h3af1c0be),
	.w5(32'h3a43c4b2),
	.w6(32'h3b189429),
	.w7(32'h39f7caa8),
	.w8(32'h3a5b7e88),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedbe65),
	.w1(32'h3b86e3e8),
	.w2(32'h3b4859b8),
	.w3(32'hbab69160),
	.w4(32'hbb11fb06),
	.w5(32'h3ac1761b),
	.w6(32'h3b86fb72),
	.w7(32'h39223f94),
	.w8(32'h3a9c17a2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb294a44),
	.w1(32'h3c8b7bfc),
	.w2(32'h3cd9326c),
	.w3(32'h3c1d3136),
	.w4(32'hbcbb3e09),
	.w5(32'hbcaaae41),
	.w6(32'h3c0c5550),
	.w7(32'h3bab70b0),
	.w8(32'hba8355cb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ede19),
	.w1(32'hbb584169),
	.w2(32'hbbd322ef),
	.w3(32'hbc5a3c32),
	.w4(32'h3b9df993),
	.w5(32'h398acfec),
	.w6(32'hb6523ea8),
	.w7(32'h3b1196ec),
	.w8(32'hb99fcf6d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebf5c1),
	.w1(32'hbb32fcc3),
	.w2(32'h3a0e3509),
	.w3(32'hbb20f083),
	.w4(32'hbba5da0b),
	.w5(32'hbb82a80a),
	.w6(32'hbba2e630),
	.w7(32'hbb619540),
	.w8(32'hbb5bb80c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b232dfd),
	.w1(32'h3b7117d7),
	.w2(32'h3b810e39),
	.w3(32'hb9e98064),
	.w4(32'hbb885826),
	.w5(32'hbb9475d9),
	.w6(32'hbb449806),
	.w7(32'hbb339d3a),
	.w8(32'hb9daead1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fd08e),
	.w1(32'h3b251b63),
	.w2(32'hba8bed09),
	.w3(32'h3c015a84),
	.w4(32'h3b60b2d7),
	.w5(32'h3a2a8ed9),
	.w6(32'h3b11648c),
	.w7(32'h3be5a4ae),
	.w8(32'h3b5c5634),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05c92f),
	.w1(32'hbc69cdc5),
	.w2(32'hbccea094),
	.w3(32'h3b957464),
	.w4(32'hbc83213c),
	.w5(32'hbc34dcc3),
	.w6(32'hbcc94378),
	.w7(32'hbc38f9c3),
	.w8(32'hbbd450d8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1bb3e),
	.w1(32'h3b6c8ec5),
	.w2(32'h3ba98b44),
	.w3(32'hbbcf0295),
	.w4(32'h3a23828e),
	.w5(32'hb95c6eac),
	.w6(32'h3b6d0dd0),
	.w7(32'h3b1759a2),
	.w8(32'h3a22f0e4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b858d8e),
	.w1(32'hbb4c85a8),
	.w2(32'hbc45bc8f),
	.w3(32'h3b1d9ac2),
	.w4(32'hb9b7d108),
	.w5(32'hbbdb41c1),
	.w6(32'h3ba2762d),
	.w7(32'h3c85e69c),
	.w8(32'h3c08b893),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6cbd1),
	.w1(32'hbc3b46ea),
	.w2(32'hbc4d31fb),
	.w3(32'hbbeef26b),
	.w4(32'hba79e17a),
	.w5(32'hbb814228),
	.w6(32'hbbbfc050),
	.w7(32'hbb919b5d),
	.w8(32'hbb7d6926),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba748530),
	.w1(32'h3b80fac7),
	.w2(32'h3b630fda),
	.w3(32'hbbf4e6fe),
	.w4(32'h3aadc51e),
	.w5(32'h39a7cedf),
	.w6(32'h3b3b917b),
	.w7(32'h3afb8145),
	.w8(32'h3a0245b3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac792fb),
	.w1(32'hbabf6ef3),
	.w2(32'h3babe8f7),
	.w3(32'hbb664e56),
	.w4(32'hba5fbd92),
	.w5(32'hbb1dc1ee),
	.w6(32'hbba403df),
	.w7(32'h3b8c1291),
	.w8(32'hbab9c2b9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0278d),
	.w1(32'h3d4b0f75),
	.w2(32'h3d469460),
	.w3(32'h3b15c1ce),
	.w4(32'h3a10fa3b),
	.w5(32'h3ca061db),
	.w6(32'hbb896291),
	.w7(32'h3970669e),
	.w8(32'h3a028eb1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca616f1),
	.w1(32'h3c167612),
	.w2(32'h3beca117),
	.w3(32'h3cf221d9),
	.w4(32'hbb861fb5),
	.w5(32'hbaf93809),
	.w6(32'h3b8c4552),
	.w7(32'hbb9dfc59),
	.w8(32'hbbdb4d9f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcefd77),
	.w1(32'h3a2a9c2f),
	.w2(32'hb943be2d),
	.w3(32'h39daf91f),
	.w4(32'h3a1cefec),
	.w5(32'h39312847),
	.w6(32'hba5c0ff4),
	.w7(32'hb9cc9b9e),
	.w8(32'h3a53cc71),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52d489),
	.w1(32'h3b90877b),
	.w2(32'h3b9ab27e),
	.w3(32'hbaa1c0db),
	.w4(32'h3b4fd6c7),
	.w5(32'h3b9a0441),
	.w6(32'h3b24e5b4),
	.w7(32'h3b3c003f),
	.w8(32'h3b8c8c10),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule