module layer_10_featuremap_352(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e3f38),
	.w1(32'h3b616245),
	.w2(32'h3999a7cf),
	.w3(32'h3a9af828),
	.w4(32'h3b4cb643),
	.w5(32'hbc00d04c),
	.w6(32'h3bc5d9f4),
	.w7(32'h3b982fe6),
	.w8(32'hbbc08d9c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70e949),
	.w1(32'hbc15e2d0),
	.w2(32'hbc229d12),
	.w3(32'hbc03bda3),
	.w4(32'hbc038e87),
	.w5(32'hbb0fee48),
	.w6(32'hbb5eb20c),
	.w7(32'hbbfa0d4c),
	.w8(32'h39b554e4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c89fd),
	.w1(32'hb981eab2),
	.w2(32'hbbcce690),
	.w3(32'h3b0bac06),
	.w4(32'h39ba67f4),
	.w5(32'hbc0c2ea7),
	.w6(32'h3ac3bc5b),
	.w7(32'hbba735f8),
	.w8(32'hbc04af53),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc180c32),
	.w1(32'hbc1dffe2),
	.w2(32'hbc1df4a1),
	.w3(32'hbc498f0e),
	.w4(32'hbc2ebacd),
	.w5(32'h3bab284c),
	.w6(32'hbc174688),
	.w7(32'hbc1bce98),
	.w8(32'h3be16733),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bae1d),
	.w1(32'hbbbea9c6),
	.w2(32'hbb051465),
	.w3(32'hbb8c715d),
	.w4(32'hba3d92a0),
	.w5(32'h3a4be1da),
	.w6(32'hbb8583f5),
	.w7(32'hbb62c4ca),
	.w8(32'h3abb68b3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c3ba7),
	.w1(32'h3ba56317),
	.w2(32'h3b418a45),
	.w3(32'h3ba2a595),
	.w4(32'h3b99dd24),
	.w5(32'hbbef2d14),
	.w6(32'h3bd7978c),
	.w7(32'h3aca7709),
	.w8(32'hbb1cfeba),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3b623),
	.w1(32'hba870ec1),
	.w2(32'hbbf90800),
	.w3(32'hbbacde28),
	.w4(32'hbb0f0dfc),
	.w5(32'hbbbdacda),
	.w6(32'h3b815e48),
	.w7(32'hbbbd6636),
	.w8(32'h3b91a8e5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9859d3),
	.w1(32'h3c1785ab),
	.w2(32'h3c273499),
	.w3(32'h3bcfc22b),
	.w4(32'hb815706e),
	.w5(32'hbb65116f),
	.w6(32'h3bdad54d),
	.w7(32'h3c0279e2),
	.w8(32'hbb42fddb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04b44d),
	.w1(32'h3b215673),
	.w2(32'hba7e7dd2),
	.w3(32'h3a755288),
	.w4(32'hba4eeb77),
	.w5(32'h3a86e97d),
	.w6(32'h3b19b843),
	.w7(32'h39fa2370),
	.w8(32'hba8ce5f2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0553f6),
	.w1(32'h3b52594c),
	.w2(32'h3af620df),
	.w3(32'h3bd41209),
	.w4(32'h3bb67c2e),
	.w5(32'hbb053367),
	.w6(32'h3c0cb199),
	.w7(32'h3b170733),
	.w8(32'hbb3e53ea),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e83cf),
	.w1(32'hba444eaa),
	.w2(32'hbb9c0671),
	.w3(32'hbac2b58e),
	.w4(32'hbb86be72),
	.w5(32'hbaeecb7a),
	.w6(32'hb70bd61d),
	.w7(32'hbc24b10a),
	.w8(32'h38fd63ea),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cbd14),
	.w1(32'h3a6e0377),
	.w2(32'hbb45a907),
	.w3(32'h3ba30222),
	.w4(32'h3b35ea9f),
	.w5(32'h3b508925),
	.w6(32'h3b33066c),
	.w7(32'hbac5eb91),
	.w8(32'hba063c10),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baba0f9),
	.w1(32'hb8e3c7d2),
	.w2(32'h3af31256),
	.w3(32'h3c33eedc),
	.w4(32'h3bea957f),
	.w5(32'h3b6b5480),
	.w6(32'h3b26fd34),
	.w7(32'h3b545bc5),
	.w8(32'hb9954bf6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa40104),
	.w1(32'h3b6855c4),
	.w2(32'hba997721),
	.w3(32'h3a4cff46),
	.w4(32'hbb85a6b2),
	.w5(32'hbc25db16),
	.w6(32'h3c117a18),
	.w7(32'hba88c597),
	.w8(32'hbbf9ec9b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42aa15),
	.w1(32'hbc1feb3c),
	.w2(32'hbc13cd4f),
	.w3(32'hbbfd19d0),
	.w4(32'hbc33e47d),
	.w5(32'hbb7a62a8),
	.w6(32'hbb2df59d),
	.w7(32'hbc0e8500),
	.w8(32'hbb8408d2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18d729),
	.w1(32'hbb332736),
	.w2(32'hba2b496a),
	.w3(32'hbb65a42b),
	.w4(32'hbabe0588),
	.w5(32'h38ec0ac7),
	.w6(32'h3bf1cdc8),
	.w7(32'h3b5b8b7f),
	.w8(32'h3b4c1ceb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fadad),
	.w1(32'hbacdf768),
	.w2(32'h39b8c976),
	.w3(32'h39cd8757),
	.w4(32'h3aa3498c),
	.w5(32'h3aaf7a92),
	.w6(32'h3a918214),
	.w7(32'h3b340124),
	.w8(32'h3a8ccd96),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad19767),
	.w1(32'hbb8deadd),
	.w2(32'hbbc30fd2),
	.w3(32'hb9ef08f4),
	.w4(32'hbbc708e3),
	.w5(32'hbb26bb6d),
	.w6(32'hbb2d1a46),
	.w7(32'hbbef1c80),
	.w8(32'h3ad8bf62),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae20c17),
	.w1(32'hbb1f44d9),
	.w2(32'hbb8eb63b),
	.w3(32'hbaaafd92),
	.w4(32'hbbc39e21),
	.w5(32'hba74d5b4),
	.w6(32'hba8b817e),
	.w7(32'hbb626109),
	.w8(32'hbaa40650),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d8ff0),
	.w1(32'hb8761049),
	.w2(32'hba926d97),
	.w3(32'hbb289212),
	.w4(32'hbabfa5a5),
	.w5(32'hbbeca72b),
	.w6(32'h3aea0dfc),
	.w7(32'hbb396feb),
	.w8(32'hbc2f62b2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d8653),
	.w1(32'hbb9bf23e),
	.w2(32'hb9b11bb3),
	.w3(32'hbb527b39),
	.w4(32'hbb6b44dd),
	.w5(32'hba91dda7),
	.w6(32'h3bafdfa7),
	.w7(32'h3b888f31),
	.w8(32'h3ac14b80),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c82364),
	.w1(32'h3bb2b409),
	.w2(32'h3c0c4dfe),
	.w3(32'hba647e1f),
	.w4(32'h3b6c6ef4),
	.w5(32'hbb884be3),
	.w6(32'h3ace5dfb),
	.w7(32'h3c0b6fca),
	.w8(32'hbb86191c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48db5f),
	.w1(32'hbb1b8937),
	.w2(32'hbbd56029),
	.w3(32'hbb04b294),
	.w4(32'hbb334766),
	.w5(32'hbc110378),
	.w6(32'hbbf239ca),
	.w7(32'hbc3126f7),
	.w8(32'hbc5138c3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc495e16),
	.w1(32'hbbc12f46),
	.w2(32'hbb3f29e1),
	.w3(32'hbb90726c),
	.w4(32'hbb611c27),
	.w5(32'h3b140660),
	.w6(32'h3c6ddcf4),
	.w7(32'hbb3e3c9d),
	.w8(32'h399f3d9a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13d6f9),
	.w1(32'h3a8458c7),
	.w2(32'hb9ed1ac9),
	.w3(32'h39c9e096),
	.w4(32'h3ae20686),
	.w5(32'hbb175c75),
	.w6(32'hba431dbf),
	.w7(32'hbb0a0a4d),
	.w8(32'hba039f4a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3305ec),
	.w1(32'h3ae254b9),
	.w2(32'h3a0fe35d),
	.w3(32'h3b72b2d1),
	.w4(32'hbba5df89),
	.w5(32'hbbfdbe3d),
	.w6(32'h3c1cd690),
	.w7(32'h3a0a6988),
	.w8(32'hbbed2d17),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5f26a),
	.w1(32'hbb33d83a),
	.w2(32'hbaed0b1a),
	.w3(32'hbb7b02d6),
	.w4(32'hbbac0388),
	.w5(32'h3b52f5d0),
	.w6(32'hbab257d4),
	.w7(32'hbacbf362),
	.w8(32'h3b57b487),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa8df1),
	.w1(32'h3c592171),
	.w2(32'h3c1adc4c),
	.w3(32'h3c7be7a1),
	.w4(32'h3c400e5a),
	.w5(32'hb9c3cfba),
	.w6(32'h3cb02c1a),
	.w7(32'h3c6adcf7),
	.w8(32'hbb0abe77),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0bc58),
	.w1(32'hba3ce3ea),
	.w2(32'h3b730fad),
	.w3(32'hbb9c1f3f),
	.w4(32'hbb94c19e),
	.w5(32'hba475202),
	.w6(32'h3ac663ff),
	.w7(32'hb7214d5a),
	.w8(32'hbb461249),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad718c8),
	.w1(32'hbaf7c996),
	.w2(32'hba5819a4),
	.w3(32'hbae11c1f),
	.w4(32'h3b758969),
	.w5(32'h3afded32),
	.w6(32'h3aa75591),
	.w7(32'h3bb6780d),
	.w8(32'hb8319b7f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b996a03),
	.w1(32'h3c34207e),
	.w2(32'h3b2bbcb0),
	.w3(32'h3bb164bb),
	.w4(32'hb8c8dc25),
	.w5(32'h3b0bbd13),
	.w6(32'h3b9c60a3),
	.w7(32'hbaabd7a2),
	.w8(32'h3b2eb29b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b00ba),
	.w1(32'hbb238ca4),
	.w2(32'h3b8e4c26),
	.w3(32'h3b8d4534),
	.w4(32'h3c454d37),
	.w5(32'h3b83b6d6),
	.w6(32'h38272a72),
	.w7(32'h3b9e73b0),
	.w8(32'h3c0f2e46),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba4a7d),
	.w1(32'hbbe39355),
	.w2(32'hbb8c3f81),
	.w3(32'h38899cd7),
	.w4(32'hbba7cae5),
	.w5(32'h3b270edd),
	.w6(32'hbba5b45b),
	.w7(32'hbb87aed1),
	.w8(32'h3b392d03),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ac42c),
	.w1(32'hbade639e),
	.w2(32'hbbc73e27),
	.w3(32'hbb02be2a),
	.w4(32'hbbb90e92),
	.w5(32'hba50003f),
	.w6(32'hbb0fdf2d),
	.w7(32'hbc0ad692),
	.w8(32'hbb29361e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a3b20),
	.w1(32'h3a5edd34),
	.w2(32'h3993dd8b),
	.w3(32'hbaeb227c),
	.w4(32'h3a36ec24),
	.w5(32'hbb45b137),
	.w6(32'hba93d935),
	.w7(32'hbae453ca),
	.w8(32'hbbdc6d25),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb806e2f2),
	.w1(32'h38bc039e),
	.w2(32'hbb87bff4),
	.w3(32'hbb718f75),
	.w4(32'hbb0b260d),
	.w5(32'hba07ef80),
	.w6(32'hba37fd24),
	.w7(32'hba405af4),
	.w8(32'h3b45af0b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb24822),
	.w1(32'h3b49946f),
	.w2(32'hbbbae34f),
	.w3(32'hba86575d),
	.w4(32'hbaa35c9a),
	.w5(32'hbc1b2afb),
	.w6(32'h3a2974a5),
	.w7(32'hbb67bc2d),
	.w8(32'hbc5a0ce6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac669e),
	.w1(32'h3c12ea7f),
	.w2(32'hbb77a8f6),
	.w3(32'h3ac274ac),
	.w4(32'hbb60fb1e),
	.w5(32'h3a1841fa),
	.w6(32'h3bcf3e25),
	.w7(32'hbb8376d6),
	.w8(32'hba8610fc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ea881),
	.w1(32'hbb0df3b9),
	.w2(32'hbbcade84),
	.w3(32'hba9a1dbd),
	.w4(32'hbaa16c8b),
	.w5(32'hbc0b6219),
	.w6(32'hbbab9d81),
	.w7(32'hbc134994),
	.w8(32'hbbf5de11),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2cb69),
	.w1(32'h39f74ff3),
	.w2(32'h3b03f1f6),
	.w3(32'hba738ef8),
	.w4(32'h3ac11d3d),
	.w5(32'h3b86eb83),
	.w6(32'h3acbea1c),
	.w7(32'h3b7572e8),
	.w8(32'h3b4e01a5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f9039),
	.w1(32'hba1c0a15),
	.w2(32'h3ad68430),
	.w3(32'hbb8f967a),
	.w4(32'hb98a97c9),
	.w5(32'hbb6f1401),
	.w6(32'hba1a4c7d),
	.w7(32'h3ab93a69),
	.w8(32'h3a82fa47),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d8758),
	.w1(32'h3b4dfd1a),
	.w2(32'hba803ed2),
	.w3(32'h3a6a6a11),
	.w4(32'hbaf0d144),
	.w5(32'h3c103692),
	.w6(32'h3c0955ba),
	.w7(32'h3af6946b),
	.w8(32'h3bb39a0e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c478fa9),
	.w1(32'h3bafe3f2),
	.w2(32'h3b16c4f0),
	.w3(32'h3b978a2d),
	.w4(32'h3afbe1b9),
	.w5(32'hbb8ec0ba),
	.w6(32'h3b419ee1),
	.w7(32'h3b4c768f),
	.w8(32'hbb8c70cf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf176cf),
	.w1(32'hbbde29b3),
	.w2(32'hbc0adb0f),
	.w3(32'hbb535779),
	.w4(32'hbb332c90),
	.w5(32'hbb43a228),
	.w6(32'hba758934),
	.w7(32'hbb9340fc),
	.w8(32'hbb08d520),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97434d),
	.w1(32'hbbcaacc7),
	.w2(32'hbaec3390),
	.w3(32'hbc02853c),
	.w4(32'hbb817f9c),
	.w5(32'h3c099cbf),
	.w6(32'hbbad08a7),
	.w7(32'hbaab719a),
	.w8(32'h3c84f2e6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46165a),
	.w1(32'h3c704e6e),
	.w2(32'h3c2e0d45),
	.w3(32'h3c5ca2c8),
	.w4(32'h3c20b8c2),
	.w5(32'hbbc1ba39),
	.w6(32'h3c81f73f),
	.w7(32'h3c21635b),
	.w8(32'hbb1a303c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40ca6c),
	.w1(32'hb9f56055),
	.w2(32'h3a6c2c56),
	.w3(32'hbae74a70),
	.w4(32'hba41bc06),
	.w5(32'hba9325f7),
	.w6(32'hba16900c),
	.w7(32'hba716cd0),
	.w8(32'hbb3a33db),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0127ba),
	.w1(32'hbad2a108),
	.w2(32'h3a04cff6),
	.w3(32'h3b1f5017),
	.w4(32'h3a4186c1),
	.w5(32'hb9147db8),
	.w6(32'hbac2c53c),
	.w7(32'h3b157bd3),
	.w8(32'hbad2b0ba),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a274772),
	.w1(32'hbbb4f288),
	.w2(32'hbbdc15bf),
	.w3(32'hbb6371bf),
	.w4(32'hbb1446f6),
	.w5(32'hbba24a98),
	.w6(32'hbb14fc89),
	.w7(32'hbbb73f6d),
	.w8(32'h3b39c8d5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb649a17),
	.w1(32'h3badf880),
	.w2(32'h3bd42336),
	.w3(32'hb92c01f1),
	.w4(32'h3ae3619f),
	.w5(32'h3c128cad),
	.w6(32'h3c093bf4),
	.w7(32'h3c080104),
	.w8(32'h3bb6506a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5ece0),
	.w1(32'h39f0b39d),
	.w2(32'hb8b801c4),
	.w3(32'h3b30ca55),
	.w4(32'h3bc3492d),
	.w5(32'hba6bc3dd),
	.w6(32'h3ac80c84),
	.w7(32'h3b13c06e),
	.w8(32'h3a3dafbd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4eb34c),
	.w1(32'hba41fb67),
	.w2(32'hbb6e29ea),
	.w3(32'hb9caf428),
	.w4(32'hbb35ee81),
	.w5(32'h3b696e84),
	.w6(32'h387c7fb0),
	.w7(32'hbb16071d),
	.w8(32'h3ab2a02d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48f794),
	.w1(32'h39f6a75b),
	.w2(32'hbab31d5b),
	.w3(32'hbb08c100),
	.w4(32'h3ad94eac),
	.w5(32'hbb0cacdf),
	.w6(32'hba61ccab),
	.w7(32'hbab60ef1),
	.w8(32'h3b5abcd4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adeec21),
	.w1(32'h3bae5e75),
	.w2(32'hbb13af09),
	.w3(32'h3b610382),
	.w4(32'hbb35c7fa),
	.w5(32'hbb7f684d),
	.w6(32'h3c0ce780),
	.w7(32'hb9eaf633),
	.w8(32'hbaf16bce),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0874d6),
	.w1(32'hba9ef748),
	.w2(32'hbb0bdf0e),
	.w3(32'hbb1b5fcd),
	.w4(32'hbab16d0a),
	.w5(32'hba6ebb05),
	.w6(32'hb9f5249e),
	.w7(32'hbb5e2737),
	.w8(32'hba4a229a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90a632),
	.w1(32'hb9f4ddfc),
	.w2(32'hbb402955),
	.w3(32'hbb317763),
	.w4(32'h37ad0486),
	.w5(32'h3b08e772),
	.w6(32'h3af79523),
	.w7(32'hbb068940),
	.w8(32'h3ab84aa5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb7362),
	.w1(32'h3a86a0b9),
	.w2(32'h3a8d6234),
	.w3(32'hbb471854),
	.w4(32'h3b38c950),
	.w5(32'h3926f8b1),
	.w6(32'hba950006),
	.w7(32'h3b470ac4),
	.w8(32'h39c4a8d4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb504fee6),
	.w1(32'h3a50130e),
	.w2(32'hb7bd8937),
	.w3(32'hbb1d0c6d),
	.w4(32'h3abe9e60),
	.w5(32'hbc0934dc),
	.w6(32'hbb26b0aa),
	.w7(32'h3b60caf5),
	.w8(32'hbb89fe23),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd33fa),
	.w1(32'h3b766c7d),
	.w2(32'h3b807810),
	.w3(32'h38d5c40a),
	.w4(32'h3a96ca2e),
	.w5(32'h3c0e8c8c),
	.w6(32'h3c276ce2),
	.w7(32'h3bd223df),
	.w8(32'h3cac84b6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ac9f0),
	.w1(32'hbbc8d4e9),
	.w2(32'hbc44e07b),
	.w3(32'hbbd5003b),
	.w4(32'hbc5d67fd),
	.w5(32'hbb064171),
	.w6(32'hbc14e644),
	.w7(32'hbc68f9b1),
	.w8(32'h3afe6b6e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fe32d),
	.w1(32'hba792b00),
	.w2(32'hbb969500),
	.w3(32'h3aa4d331),
	.w4(32'hb99ec56e),
	.w5(32'hba356a39),
	.w6(32'h3b100c6b),
	.w7(32'hbb4a6b84),
	.w8(32'h3bcfa682),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82985a),
	.w1(32'hb97a325d),
	.w2(32'hba52ea92),
	.w3(32'hb97efdf5),
	.w4(32'hbb820801),
	.w5(32'h3a7a3c1b),
	.w6(32'h3c0c8924),
	.w7(32'hbac24465),
	.w8(32'h3b8648a3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54d02f),
	.w1(32'hbb7fbee2),
	.w2(32'hbb2f2ba2),
	.w3(32'hbad3cb02),
	.w4(32'h3ada5089),
	.w5(32'hb9f053f6),
	.w6(32'hbad38e39),
	.w7(32'hbb44cf31),
	.w8(32'hbb05d398),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fa8ea),
	.w1(32'h3b3a9ed9),
	.w2(32'hb9471dbb),
	.w3(32'h3a24e381),
	.w4(32'hb95cb8ee),
	.w5(32'hba50e2a5),
	.w6(32'h3ba07c1b),
	.w7(32'h3a7777e6),
	.w8(32'hb97898bc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bacdcc),
	.w1(32'h3b1468b1),
	.w2(32'hba822b18),
	.w3(32'hbb216926),
	.w4(32'hbb95dd54),
	.w5(32'hbb837852),
	.w6(32'h3a2fe3f0),
	.w7(32'hbb904905),
	.w8(32'hb903013b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cd120),
	.w1(32'hbbcd8367),
	.w2(32'hbbe6f94d),
	.w3(32'hbbe1c633),
	.w4(32'hbb4c7c67),
	.w5(32'hbb5a69d6),
	.w6(32'hbb9a74b1),
	.w7(32'hbbfdc1fb),
	.w8(32'h3bdfc207),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39261546),
	.w1(32'h3c0c8315),
	.w2(32'h3a9a97f7),
	.w3(32'h3b33fa2c),
	.w4(32'hbb3dc080),
	.w5(32'h3c0f5227),
	.w6(32'h3c082cd8),
	.w7(32'hbaf35668),
	.w8(32'h3b8373f1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae06f7a),
	.w1(32'hbbe40079),
	.w2(32'hbc01a0f1),
	.w3(32'h39b54852),
	.w4(32'hbbfa5b88),
	.w5(32'h3be04af1),
	.w6(32'hbb906a2b),
	.w7(32'hbbbee88a),
	.w8(32'h3c469cd4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdcbe6),
	.w1(32'hbb00793d),
	.w2(32'hbbc87964),
	.w3(32'hb90482f6),
	.w4(32'hbbb5ba24),
	.w5(32'hbbbc9b5b),
	.w6(32'hbb0c9102),
	.w7(32'hbbffafb0),
	.w8(32'hbb9efd12),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c0bb1),
	.w1(32'hba33e429),
	.w2(32'hbb0e8276),
	.w3(32'hbafc28fd),
	.w4(32'hbb28cf3d),
	.w5(32'hba482b9d),
	.w6(32'hbbf1a7af),
	.w7(32'hbb821fd1),
	.w8(32'hbb9d7f7c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b3016),
	.w1(32'hbaa717d5),
	.w2(32'hbb562de2),
	.w3(32'hba504c24),
	.w4(32'hbb42cc1b),
	.w5(32'hbbae429c),
	.w6(32'h3a6a4c86),
	.w7(32'hba8f1303),
	.w8(32'hbbd39684),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21183d),
	.w1(32'h3b029516),
	.w2(32'hbae759a8),
	.w3(32'hbb39954a),
	.w4(32'hba69c415),
	.w5(32'h3becfd08),
	.w6(32'h3b34bc05),
	.w7(32'h3a8a9e6c),
	.w8(32'hb96dd5f0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8fd5a),
	.w1(32'hbb9daeeb),
	.w2(32'hbc14e8bf),
	.w3(32'hba98420d),
	.w4(32'hbaf779af),
	.w5(32'h3b49c863),
	.w6(32'hb790e5c0),
	.w7(32'hbbbb8065),
	.w8(32'h3b47cd4a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2d5b),
	.w1(32'hbb526e04),
	.w2(32'hba75dd7d),
	.w3(32'h3b71586f),
	.w4(32'hba616225),
	.w5(32'hba879ac6),
	.w6(32'hba7e86c2),
	.w7(32'hba9906c1),
	.w8(32'h3ac3674e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cf7d9),
	.w1(32'h3bdcf97a),
	.w2(32'hbaae7ddd),
	.w3(32'h3bf6d6a2),
	.w4(32'hb9ed61da),
	.w5(32'h3b5f3d26),
	.w6(32'h3bfd003f),
	.w7(32'hbb81f831),
	.w8(32'hb8b66a0f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bbd1e),
	.w1(32'hbbd1c265),
	.w2(32'hbb994c58),
	.w3(32'h3a2d7976),
	.w4(32'hbaa953e9),
	.w5(32'hba5c838f),
	.w6(32'hbb92c12f),
	.w7(32'hbba0f311),
	.w8(32'h3a27fe4d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af65b32),
	.w1(32'hba4d33d2),
	.w2(32'hbbbc21fb),
	.w3(32'h3afe2289),
	.w4(32'hba11c1f7),
	.w5(32'hbb7efcd8),
	.w6(32'h3aa84270),
	.w7(32'hbba731d5),
	.w8(32'hbbe54e9b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb670915),
	.w1(32'hbb733491),
	.w2(32'hbb386d37),
	.w3(32'hbb872c09),
	.w4(32'hbb0df5a3),
	.w5(32'h3b044c63),
	.w6(32'hbb846f43),
	.w7(32'hba939fe2),
	.w8(32'h3b8de4b9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae66197),
	.w1(32'h3a04a173),
	.w2(32'hbbaf2957),
	.w3(32'hbb0eefc8),
	.w4(32'hbb9d2d88),
	.w5(32'hba2eb9c6),
	.w6(32'h39861337),
	.w7(32'hbb99ff54),
	.w8(32'h3bca9f1f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1603ce),
	.w1(32'h396aeb2d),
	.w2(32'hbb9ca5df),
	.w3(32'h3b17fd8a),
	.w4(32'hba1aa93e),
	.w5(32'hbbde005f),
	.w6(32'h3b847da7),
	.w7(32'hbb755936),
	.w8(32'hbc588e84),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc017541),
	.w1(32'hbb4f9fda),
	.w2(32'hbae9929e),
	.w3(32'hbb84a216),
	.w4(32'hba90dd3b),
	.w5(32'h3b458db8),
	.w6(32'hba9a5004),
	.w7(32'hb88e7531),
	.w8(32'h3b2dffc7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf1c79),
	.w1(32'hb9fe3750),
	.w2(32'hbb697c2b),
	.w3(32'h3b126624),
	.w4(32'hbb11d46c),
	.w5(32'h3b28a1cd),
	.w6(32'h3a12d987),
	.w7(32'hbb14a62d),
	.w8(32'h3ace10f1),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b005755),
	.w1(32'h3a21ad43),
	.w2(32'hbb5920ba),
	.w3(32'h3ab028b1),
	.w4(32'h3b1e659c),
	.w5(32'hbba9f97e),
	.w6(32'h3b1ae523),
	.w7(32'hba7df894),
	.w8(32'hbb8b4e16),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e2ecf),
	.w1(32'hbc370994),
	.w2(32'hbc54a4c9),
	.w3(32'hbbc1a239),
	.w4(32'hbc541412),
	.w5(32'hbafbd5df),
	.w6(32'hbb95237b),
	.w7(32'hbc43f732),
	.w8(32'hbacbbf85),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96da98),
	.w1(32'hb98028a0),
	.w2(32'h39939216),
	.w3(32'hb9330709),
	.w4(32'h3a818062),
	.w5(32'h3b10139e),
	.w6(32'h3986bbc2),
	.w7(32'h39347645),
	.w8(32'h3be8ff42),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25905c),
	.w1(32'h3b92ecfd),
	.w2(32'h3b81622a),
	.w3(32'h3bd3610a),
	.w4(32'h3b7e6b62),
	.w5(32'hbb748713),
	.w6(32'h3c302540),
	.w7(32'hbafe7981),
	.w8(32'hbb298663),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40ee01),
	.w1(32'h3bd74206),
	.w2(32'h3b223baa),
	.w3(32'h3b3f8499),
	.w4(32'h3bb23c8e),
	.w5(32'hbace5c0f),
	.w6(32'h3bd77343),
	.w7(32'h3b99d28c),
	.w8(32'h3a60e82a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ba0fb),
	.w1(32'hbb6f4dba),
	.w2(32'hbb0b44c0),
	.w3(32'hba36e5c5),
	.w4(32'hbb34159e),
	.w5(32'hbb9887a1),
	.w6(32'h399d46a4),
	.w7(32'hbb2c1670),
	.w8(32'h3b2cd2ae),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb341398),
	.w1(32'h3b1a1157),
	.w2(32'h3aa652bc),
	.w3(32'hb93bc4ba),
	.w4(32'hba4e0364),
	.w5(32'h3b2025c9),
	.w6(32'h3b5c6ba0),
	.w7(32'h3ad9adcb),
	.w8(32'hbc11f8fd),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13916a),
	.w1(32'hbb88425e),
	.w2(32'h3a6ed508),
	.w3(32'h3af8f38e),
	.w4(32'h3b9c615c),
	.w5(32'hbc3e52b0),
	.w6(32'h3a9a825d),
	.w7(32'h3b8b45e2),
	.w8(32'hbbfdfd2b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36d466),
	.w1(32'hba83f8de),
	.w2(32'h3a44ade7),
	.w3(32'h3aa198c6),
	.w4(32'h3b8d4e91),
	.w5(32'h3a804ce4),
	.w6(32'h3c0cb988),
	.w7(32'hbaa46e5d),
	.w8(32'h3a8486e8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ef32a),
	.w1(32'hbb825ea2),
	.w2(32'hbc1a94fd),
	.w3(32'hba192ef2),
	.w4(32'hbbc2347a),
	.w5(32'h3b3c75d7),
	.w6(32'hbb3941bb),
	.w7(32'hbc3efcc4),
	.w8(32'h3bac6bd0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e4973),
	.w1(32'hbb228c42),
	.w2(32'hbbb1d891),
	.w3(32'hbb742fc0),
	.w4(32'hbae4e2e5),
	.w5(32'hbaf03a39),
	.w6(32'hba193448),
	.w7(32'hbb7bfc04),
	.w8(32'h3ad3974a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c72e6),
	.w1(32'h3b1c79da),
	.w2(32'hb9d8cfcf),
	.w3(32'h3a981026),
	.w4(32'hba12a1dc),
	.w5(32'hbb238fdb),
	.w6(32'h3b86210f),
	.w7(32'h3a9596bd),
	.w8(32'hbc03f217),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6efe28),
	.w1(32'h3be00750),
	.w2(32'h38bdd10f),
	.w3(32'h3bb57bfd),
	.w4(32'h3a85fad5),
	.w5(32'h3b07aa13),
	.w6(32'h3c34d004),
	.w7(32'h3b8d8679),
	.w8(32'h3a2f55c7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88231b),
	.w1(32'h3b9ad9b8),
	.w2(32'hbadab048),
	.w3(32'h3ae0381f),
	.w4(32'hbbd0378f),
	.w5(32'h3a7054dc),
	.w6(32'h3b63b8f0),
	.w7(32'hbbeac65d),
	.w8(32'hba00e89a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558077),
	.w1(32'hbbfc4322),
	.w2(32'hbc0329d6),
	.w3(32'hbba275ac),
	.w4(32'hbbaa9989),
	.w5(32'h3c50371e),
	.w6(32'hbbbe7736),
	.w7(32'hbbd37363),
	.w8(32'h3c594d86),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2948cd),
	.w1(32'hbaebc604),
	.w2(32'hbb3a9c8f),
	.w3(32'h3b36f019),
	.w4(32'hbae83975),
	.w5(32'h3a860da8),
	.w6(32'h3b073784),
	.w7(32'hba7f0a49),
	.w8(32'hba4d9a70),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d72d3),
	.w1(32'hb972e15d),
	.w2(32'hba06576c),
	.w3(32'h3b8043d4),
	.w4(32'h3a355640),
	.w5(32'h3a7589a9),
	.w6(32'h3b142e11),
	.w7(32'hbba723d9),
	.w8(32'h3b57dee6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b030b),
	.w1(32'hbc079f89),
	.w2(32'hbb07513a),
	.w3(32'hbbcec1c9),
	.w4(32'hbbab5400),
	.w5(32'h3ac720de),
	.w6(32'hbb647910),
	.w7(32'hbadd42da),
	.w8(32'hb949e31e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd034),
	.w1(32'h3aca7770),
	.w2(32'h3a4876a7),
	.w3(32'h3991bdac),
	.w4(32'h3b2738b0),
	.w5(32'hbb8f7761),
	.w6(32'hbb1b1cd7),
	.w7(32'hbba8e353),
	.w8(32'hbc213ce3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7b761),
	.w1(32'hbb6d3629),
	.w2(32'h39431395),
	.w3(32'hbadda370),
	.w4(32'h3b717d79),
	.w5(32'h3b50b3d0),
	.w6(32'hbbac5ad3),
	.w7(32'h3a814f0a),
	.w8(32'h3ba10d2b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bb403),
	.w1(32'hbb2e2276),
	.w2(32'hbb54820c),
	.w3(32'hbab52729),
	.w4(32'hbb805fd8),
	.w5(32'hbbd8c023),
	.w6(32'hbb476a88),
	.w7(32'hbbff313f),
	.w8(32'hbc81f219),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41e43b),
	.w1(32'hbb3b51de),
	.w2(32'hb8f0d3b3),
	.w3(32'h3ba667cf),
	.w4(32'h3b8b13a0),
	.w5(32'hbaff976e),
	.w6(32'h3aebfb2e),
	.w7(32'h3a8aef2b),
	.w8(32'h3bb3e050),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82cd85),
	.w1(32'hbb3461d7),
	.w2(32'hbc0317da),
	.w3(32'hba991197),
	.w4(32'hbbd0f04e),
	.w5(32'hbb66c614),
	.w6(32'hbb0980f4),
	.w7(32'hbbee7bfa),
	.w8(32'hbb4688dc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba674ce),
	.w1(32'h3b9ada66),
	.w2(32'h3bf99aec),
	.w3(32'h3bd61b92),
	.w4(32'h3c141462),
	.w5(32'h3ba4c28d),
	.w6(32'h3ba761eb),
	.w7(32'h3c4f49fd),
	.w8(32'h3c30e8c8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b717c55),
	.w1(32'hbbe066ab),
	.w2(32'hbbea7722),
	.w3(32'hbbc80c2e),
	.w4(32'hbc44481f),
	.w5(32'h3a9376c4),
	.w6(32'hbc1c4053),
	.w7(32'hbc0f948f),
	.w8(32'h3b447a40),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba9a3e),
	.w1(32'hba7773cd),
	.w2(32'h3a5faf10),
	.w3(32'hbb30332e),
	.w4(32'hba9340d2),
	.w5(32'h3a4fe48d),
	.w6(32'hb9f9e5ad),
	.w7(32'hba993827),
	.w8(32'h3aaa926d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9157a),
	.w1(32'h3b252020),
	.w2(32'h3b98c204),
	.w3(32'h3be39ef4),
	.w4(32'h3b94ad9a),
	.w5(32'hba486ab8),
	.w6(32'h3bacd98f),
	.w7(32'hbb48588c),
	.w8(32'hbb279200),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6dcf0),
	.w1(32'hba80a2e1),
	.w2(32'h393d5037),
	.w3(32'hba4f6652),
	.w4(32'hb91de42a),
	.w5(32'hbae3918c),
	.w6(32'hbab6522e),
	.w7(32'hbab05443),
	.w8(32'hbab681be),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba813810),
	.w1(32'hbb9b97ba),
	.w2(32'hbaf9d03e),
	.w3(32'hbbda3e32),
	.w4(32'hbba7288c),
	.w5(32'h3b2ca9b8),
	.w6(32'hbbcf7c0a),
	.w7(32'hbba20882),
	.w8(32'h3ac1c9e3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7754f7),
	.w1(32'hba9891a4),
	.w2(32'h3a76c2a0),
	.w3(32'hbade594e),
	.w4(32'hba9d6668),
	.w5(32'hbbae5f40),
	.w6(32'hbb156d2c),
	.w7(32'hbac6f97a),
	.w8(32'hbbd2dea1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4226b2),
	.w1(32'hb95ce49a),
	.w2(32'hba97a71f),
	.w3(32'hbb016f93),
	.w4(32'hbad332cf),
	.w5(32'h3a7fb191),
	.w6(32'hbbc199db),
	.w7(32'hbb74e5ce),
	.w8(32'hbbaa1a70),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88191e),
	.w1(32'hba06d1dd),
	.w2(32'hb8ff5b16),
	.w3(32'h3bbcc835),
	.w4(32'h35db7d60),
	.w5(32'h3a127fc6),
	.w6(32'hbaea6053),
	.w7(32'h3ad9398b),
	.w8(32'h3b678107),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d6bad),
	.w1(32'h3ab8aae6),
	.w2(32'hbb46338f),
	.w3(32'hbb845f24),
	.w4(32'h391ad818),
	.w5(32'hbb2fe066),
	.w6(32'h3bdacfc5),
	.w7(32'h39fdf39f),
	.w8(32'hbb323816),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72897f),
	.w1(32'hbae79c47),
	.w2(32'hbaadab73),
	.w3(32'hbb14cc63),
	.w4(32'hbada61ba),
	.w5(32'hbb0f71eb),
	.w6(32'hbad16770),
	.w7(32'h39d02bd2),
	.w8(32'hbaa48fa1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e3f3a),
	.w1(32'hbab12621),
	.w2(32'hbb0c1ada),
	.w3(32'hbac3bb76),
	.w4(32'hb9b9e8fb),
	.w5(32'hb9b97a51),
	.w6(32'hbaa4dec5),
	.w7(32'hbb6e9119),
	.w8(32'h3b0ab540),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393300b4),
	.w1(32'hbb88d654),
	.w2(32'hbbc24b55),
	.w3(32'hbbd009ca),
	.w4(32'hbbe3a39b),
	.w5(32'hbbae86a0),
	.w6(32'hbbb24ec1),
	.w7(32'hbb174025),
	.w8(32'hbb477481),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf81056),
	.w1(32'hbba07401),
	.w2(32'hba77cfac),
	.w3(32'hbb049ffd),
	.w4(32'hb8960531),
	.w5(32'hbb9dbaf7),
	.w6(32'hbbb14cc0),
	.w7(32'hbad8a531),
	.w8(32'hbc248fa7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc035520),
	.w1(32'h3b6abd4c),
	.w2(32'h3a8e5f8b),
	.w3(32'h3bf7cf2c),
	.w4(32'hb956fda1),
	.w5(32'h3b31926b),
	.w6(32'h3b44cd79),
	.w7(32'hbb437987),
	.w8(32'h3afb79ff),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a84a4),
	.w1(32'hba10eafb),
	.w2(32'hb9ae4317),
	.w3(32'h3b447022),
	.w4(32'h3b00fe38),
	.w5(32'h3aae91d3),
	.w6(32'h3b242285),
	.w7(32'hb9b4658c),
	.w8(32'h3b134dcc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7de454),
	.w1(32'h3b90056c),
	.w2(32'hbb9ffffc),
	.w3(32'h3b9b4c7c),
	.w4(32'hbb046946),
	.w5(32'hbaf54923),
	.w6(32'h3ba2a38b),
	.w7(32'hbb675855),
	.w8(32'hbb873286),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92b61b),
	.w1(32'h3a60ea84),
	.w2(32'hb9f6caac),
	.w3(32'hbb1d558d),
	.w4(32'h39b7bdc5),
	.w5(32'h3b43aea2),
	.w6(32'hb8e98af8),
	.w7(32'h3b09502a),
	.w8(32'h3b0709a9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6b5f3),
	.w1(32'hbb32b3b4),
	.w2(32'hbab4329f),
	.w3(32'hba91bbc6),
	.w4(32'hba744ae1),
	.w5(32'hb9c2a321),
	.w6(32'hbb145c4a),
	.w7(32'hbaff709f),
	.w8(32'hbb7c7212),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55913e),
	.w1(32'h393a62ca),
	.w2(32'hbb115a81),
	.w3(32'hbac3a7cf),
	.w4(32'h39d484b5),
	.w5(32'hb9fde9ce),
	.w6(32'hbae7d941),
	.w7(32'hbab5417b),
	.w8(32'hbc03d42c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f9f3a),
	.w1(32'hbb3f164d),
	.w2(32'h38d1cfb3),
	.w3(32'h3b47d267),
	.w4(32'h3b2dadf4),
	.w5(32'h3b0c0336),
	.w6(32'hbb9c2b60),
	.w7(32'h38fd13df),
	.w8(32'h3b7d2360),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7060ac),
	.w1(32'h3a8aa311),
	.w2(32'hbb0135d6),
	.w3(32'hbb158f76),
	.w4(32'hbb558373),
	.w5(32'h3b649878),
	.w6(32'hba2dc7c7),
	.w7(32'hbb708cce),
	.w8(32'h3af5f534),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e0cdc),
	.w1(32'h3ac3ace0),
	.w2(32'hb9451d7e),
	.w3(32'h3b6b87e8),
	.w4(32'h3bf54cc1),
	.w5(32'hbaf61c20),
	.w6(32'h3ad6f30f),
	.w7(32'h3abb5684),
	.w8(32'hba88422b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3813cf83),
	.w1(32'h39ae23a5),
	.w2(32'h3b05183f),
	.w3(32'h3a58fbc6),
	.w4(32'h3b4d74d5),
	.w5(32'h3a9f5496),
	.w6(32'h3b005e6e),
	.w7(32'h3aa08fa7),
	.w8(32'h3b355579),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92d3ff),
	.w1(32'h3afb0980),
	.w2(32'hbaed0fbf),
	.w3(32'hbacb5997),
	.w4(32'h3a64a8d9),
	.w5(32'h3bb8beb4),
	.w6(32'h3a2e4f6c),
	.w7(32'hba25e8d4),
	.w8(32'h3b3d6324),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94b6d4),
	.w1(32'hbb4673d9),
	.w2(32'hba817797),
	.w3(32'h3b97ae87),
	.w4(32'h3a6edd34),
	.w5(32'hbb375e16),
	.w6(32'hbb85c57d),
	.w7(32'hb9878ff0),
	.w8(32'hbb0197bb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef89a2),
	.w1(32'h3b27d840),
	.w2(32'h3a833365),
	.w3(32'h3a628cc4),
	.w4(32'h3ae67b76),
	.w5(32'hbbb20927),
	.w6(32'h3b85d92d),
	.w7(32'hb9faabeb),
	.w8(32'hba8870b7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86da0e),
	.w1(32'hbbe95636),
	.w2(32'hbb59c519),
	.w3(32'hbb8ca5c4),
	.w4(32'h394b2512),
	.w5(32'hbb1a160e),
	.w6(32'hbb90ee5f),
	.w7(32'h3abd7bce),
	.w8(32'hbb545165),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5c2b3),
	.w1(32'hbb5e018c),
	.w2(32'hba6382ae),
	.w3(32'hbb78f17d),
	.w4(32'hbb1b2bf2),
	.w5(32'hba86ff62),
	.w6(32'hbb6a91d5),
	.w7(32'hbaebae5b),
	.w8(32'h39b17b4e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ce0f9),
	.w1(32'hbb414e58),
	.w2(32'hbb149dd8),
	.w3(32'hba466020),
	.w4(32'hbafec626),
	.w5(32'hbaae920e),
	.w6(32'hbafe8a6b),
	.w7(32'hbb395094),
	.w8(32'hb985b57b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e5ae6),
	.w1(32'h3a713e43),
	.w2(32'hb9ea6866),
	.w3(32'h3ac8ec59),
	.w4(32'h3a4d8120),
	.w5(32'hbb8123c0),
	.w6(32'h3a980951),
	.w7(32'hbae3d4ad),
	.w8(32'hbbb33658),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb782ec1),
	.w1(32'hbb36b5dd),
	.w2(32'hbad24e1e),
	.w3(32'hbb1d2b48),
	.w4(32'hba3c4efd),
	.w5(32'hbad5521a),
	.w6(32'hbb953c0a),
	.w7(32'hbb76b5fa),
	.w8(32'hbb0007d0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac32f6a),
	.w1(32'hbb80dbe3),
	.w2(32'hbb54f83b),
	.w3(32'hba90d528),
	.w4(32'hbb1972e8),
	.w5(32'hbb0d1eb7),
	.w6(32'hbad76776),
	.w7(32'hbb7e3c0b),
	.w8(32'hbb40505f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba441ccf),
	.w1(32'h3a0b6018),
	.w2(32'h3aa64d3b),
	.w3(32'hb9988fc5),
	.w4(32'h3a9a54fc),
	.w5(32'h3b67a555),
	.w6(32'hbaeb6d83),
	.w7(32'hba927547),
	.w8(32'h3ba752ba),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba16967),
	.w1(32'hbb00ffd8),
	.w2(32'hbb77ec52),
	.w3(32'h3bbd7e01),
	.w4(32'hbb3e64e4),
	.w5(32'h3babba17),
	.w6(32'hbbbf5a2d),
	.w7(32'hbad66239),
	.w8(32'h3b8667a5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cf99a),
	.w1(32'h3a0c522d),
	.w2(32'hb917cb39),
	.w3(32'h3a406cb2),
	.w4(32'hbabc138b),
	.w5(32'h3ad0350c),
	.w6(32'h3b2affc9),
	.w7(32'h3b1cff05),
	.w8(32'h3bb32ad2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dafe9),
	.w1(32'hbb63ef47),
	.w2(32'h3ab02596),
	.w3(32'hbbac0654),
	.w4(32'h3a988b17),
	.w5(32'h3999e15a),
	.w6(32'hbafaf4e8),
	.w7(32'h3b3e685e),
	.w8(32'h3a368d54),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a90c7),
	.w1(32'hba924084),
	.w2(32'hba908bc7),
	.w3(32'hbb63b642),
	.w4(32'hbb014d89),
	.w5(32'hbb4b6b02),
	.w6(32'hbaf0354b),
	.w7(32'hbb019b5b),
	.w8(32'hbac2fc1d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e8fad),
	.w1(32'hbae0cb19),
	.w2(32'h38a7cf25),
	.w3(32'hbb5d23b4),
	.w4(32'hbb20aad8),
	.w5(32'hbad8e7bb),
	.w6(32'hbb1c0c3c),
	.w7(32'hbaba0f9c),
	.w8(32'hb998c551),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb041cf5),
	.w1(32'hbb20318c),
	.w2(32'hbaf23c9c),
	.w3(32'hbb861a28),
	.w4(32'hbbb466c9),
	.w5(32'hbbd97f0e),
	.w6(32'hbb68d44c),
	.w7(32'hbb1fa48c),
	.w8(32'hbc388d7d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce7a7e),
	.w1(32'hbb0e9961),
	.w2(32'hbaf739a1),
	.w3(32'hbb0c9d11),
	.w4(32'h39de31cc),
	.w5(32'hbc250ee5),
	.w6(32'hbb809535),
	.w7(32'h39ead400),
	.w8(32'hbc78e990),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5046c),
	.w1(32'hbb7aef28),
	.w2(32'h3a3e13a3),
	.w3(32'hbb36ca83),
	.w4(32'h3adb8270),
	.w5(32'hbb33071d),
	.w6(32'hbbb7207a),
	.w7(32'hbb713244),
	.w8(32'hbb329615),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4059ab),
	.w1(32'hb9d93525),
	.w2(32'hbaa619fb),
	.w3(32'h3ae90cca),
	.w4(32'hb9e8b514),
	.w5(32'h3a75815f),
	.w6(32'hbacf14c4),
	.w7(32'h3a44efd9),
	.w8(32'h3ade422e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3085a),
	.w1(32'hba49488e),
	.w2(32'h3a8b2b97),
	.w3(32'h3a904813),
	.w4(32'h397ccce8),
	.w5(32'hbb1fefbd),
	.w6(32'h3b86993e),
	.w7(32'h3ac137f1),
	.w8(32'hba548a18),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba998651),
	.w1(32'hbb87811d),
	.w2(32'hbba3fe66),
	.w3(32'hbaace55b),
	.w4(32'hbb410057),
	.w5(32'h3b229380),
	.w6(32'h39819b9e),
	.w7(32'hbb92bacc),
	.w8(32'h3b2a1497),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7308fb),
	.w1(32'h3b701eaf),
	.w2(32'h3a252dbc),
	.w3(32'h3be74297),
	.w4(32'hbb18aa83),
	.w5(32'hb98e912c),
	.w6(32'h3af62886),
	.w7(32'hbb376319),
	.w8(32'h3b84ba87),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d3c8),
	.w1(32'hba89f6ca),
	.w2(32'hb9461a85),
	.w3(32'hbb3ca2af),
	.w4(32'h3aa7ffae),
	.w5(32'h3a392df3),
	.w6(32'hb99029ea),
	.w7(32'h3a86c9eb),
	.w8(32'hbbc490a8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb7272),
	.w1(32'h3a6e6407),
	.w2(32'h3b5181b9),
	.w3(32'hbaff7371),
	.w4(32'h3b48e7b3),
	.w5(32'h3a4c8496),
	.w6(32'hbb4911c5),
	.w7(32'h3b528f57),
	.w8(32'h3aab90c2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4cddab),
	.w1(32'hbb171736),
	.w2(32'hb89846f4),
	.w3(32'hbbad80c2),
	.w4(32'hbaddfef9),
	.w5(32'h38a98842),
	.w6(32'hbb3565ce),
	.w7(32'hb9d2ca5f),
	.w8(32'h3b1d1703),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba059dc9),
	.w1(32'hbb3b838e),
	.w2(32'hbb4db98e),
	.w3(32'hbb67f0a8),
	.w4(32'hbb402115),
	.w5(32'hbaf01add),
	.w6(32'hbaf5ecbd),
	.w7(32'hba944688),
	.w8(32'hbb550ce5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c44ec),
	.w1(32'hb9e2188a),
	.w2(32'h3aac8f67),
	.w3(32'hba913f8e),
	.w4(32'h3a383f60),
	.w5(32'h3b9e3daf),
	.w6(32'hbb9677df),
	.w7(32'hbb4a8f16),
	.w8(32'h3b88c904),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b971242),
	.w1(32'hba7f7c3f),
	.w2(32'hbb19e4b4),
	.w3(32'hbb25a1c1),
	.w4(32'hb8af58d0),
	.w5(32'h374e1167),
	.w6(32'hbb83ab8a),
	.w7(32'hbb032e24),
	.w8(32'h3b1326d2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa97865),
	.w1(32'hbb08c683),
	.w2(32'hbb2089f1),
	.w3(32'hb82e05b8),
	.w4(32'hbab7676c),
	.w5(32'hbbb51304),
	.w6(32'h3a65cc24),
	.w7(32'h3a3122bf),
	.w8(32'hbbdfc9ce),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac0007),
	.w1(32'hbbf5741a),
	.w2(32'hba10727a),
	.w3(32'hbba77ee1),
	.w4(32'h3b039d8f),
	.w5(32'h3ab7b1e8),
	.w6(32'hbbb59fcf),
	.w7(32'hbb1fa2e4),
	.w8(32'hbba34e04),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87ae8db),
	.w1(32'h3aac0708),
	.w2(32'hbb30db4b),
	.w3(32'h3a1a6116),
	.w4(32'h3a90ad49),
	.w5(32'hbbbfee37),
	.w6(32'hbb972f31),
	.w7(32'hbb0849f7),
	.w8(32'hbb9be3c6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babf6e8),
	.w1(32'h3af7b64c),
	.w2(32'h3b80f0f0),
	.w3(32'hbb43b4f3),
	.w4(32'h3bbbfe43),
	.w5(32'hbaa64282),
	.w6(32'hbad40d6a),
	.w7(32'hb9997088),
	.w8(32'hba2acf91),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93cd4a),
	.w1(32'h3a8d4ceb),
	.w2(32'hbb658be7),
	.w3(32'hbb95ccfa),
	.w4(32'hbb81fe50),
	.w5(32'hba07438b),
	.w6(32'hbb656fde),
	.w7(32'hbb57af37),
	.w8(32'hbb8c5fa4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb8434),
	.w1(32'h3a187518),
	.w2(32'hbacd2ad8),
	.w3(32'hbb476193),
	.w4(32'hbb6e509e),
	.w5(32'h3ad3a3e7),
	.w6(32'hbba507db),
	.w7(32'hbb8f4787),
	.w8(32'h3b28505c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d2a7b),
	.w1(32'hbb7ecc3f),
	.w2(32'h3b20bc9c),
	.w3(32'hbaf91d34),
	.w4(32'h39f4e913),
	.w5(32'hbbfae0b1),
	.w6(32'hb8b52c42),
	.w7(32'h3ba6b224),
	.w8(32'hbbbc9a27),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ab0c6),
	.w1(32'hbb67ce79),
	.w2(32'hba40e098),
	.w3(32'hbb88da9f),
	.w4(32'hbb7e3947),
	.w5(32'h3a5c1fbc),
	.w6(32'hbbf4be03),
	.w7(32'hbb21ad5f),
	.w8(32'h3a10cf0d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9835997),
	.w1(32'h3b2aa484),
	.w2(32'h3ad74f50),
	.w3(32'h3b2e6397),
	.w4(32'h3b538667),
	.w5(32'hbb5a5f76),
	.w6(32'h3b58b587),
	.w7(32'h3b41de06),
	.w8(32'hbaaebfde),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992b0aa),
	.w1(32'hb8f41b02),
	.w2(32'h3aa0f8ee),
	.w3(32'hbb3f149a),
	.w4(32'hba76b312),
	.w5(32'hbbd72d33),
	.w6(32'hbbbd4063),
	.w7(32'hbb16dd42),
	.w8(32'hbb0904df),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd28756),
	.w1(32'h3b8464cc),
	.w2(32'h3bb344e0),
	.w3(32'h3b86b5ce),
	.w4(32'h3bbf4c45),
	.w5(32'hba9733b7),
	.w6(32'h3c018573),
	.w7(32'h3afa17c2),
	.w8(32'h3b5e9b49),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc2fee),
	.w1(32'hb8ff8e2c),
	.w2(32'hbb406ccb),
	.w3(32'h3a446dd6),
	.w4(32'hbb40b848),
	.w5(32'h3af0a887),
	.w6(32'hb930cbf3),
	.w7(32'hbba906a7),
	.w8(32'h3b83759b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b91a9),
	.w1(32'hb8e5046d),
	.w2(32'hbafc6f1c),
	.w3(32'hbb08d586),
	.w4(32'hbb2cc3c7),
	.w5(32'hbc4dfca8),
	.w6(32'hba5cb0a5),
	.w7(32'hbaf20817),
	.w8(32'hbcb057a4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6518cb),
	.w1(32'hba0e1ac6),
	.w2(32'h3b11205f),
	.w3(32'h3a038f72),
	.w4(32'h3c1aee34),
	.w5(32'hbba010d3),
	.w6(32'h3a6fcd1c),
	.w7(32'h3bfbb9f2),
	.w8(32'hbb1a81cb),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96feed),
	.w1(32'hbbb8fafe),
	.w2(32'hbbac9993),
	.w3(32'hbc1d513a),
	.w4(32'hbc17a80e),
	.w5(32'hbb302e8b),
	.w6(32'hbbf433a1),
	.w7(32'hbb9537a3),
	.w8(32'hbb50a9e6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba67873),
	.w1(32'hbae7e009),
	.w2(32'hbb12953a),
	.w3(32'h3bab2016),
	.w4(32'h3b83c99a),
	.w5(32'h3b5c0b91),
	.w6(32'h3b9e7ff0),
	.w7(32'hba9e2224),
	.w8(32'h3be03a9b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59c5d),
	.w1(32'hbb36fd51),
	.w2(32'hbbebd29f),
	.w3(32'hbb858eb1),
	.w4(32'hbc348c4c),
	.w5(32'h3c00b230),
	.w6(32'hbc0e9fa3),
	.w7(32'hbc31297c),
	.w8(32'h3c74b039),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb6d80),
	.w1(32'hbb8859cb),
	.w2(32'hbb9b66ba),
	.w3(32'hbb0fcf5b),
	.w4(32'hbc0baf30),
	.w5(32'hbb6fa230),
	.w6(32'hbb5712d4),
	.w7(32'hbbb0a1ba),
	.w8(32'hbb8cd330),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb053604),
	.w1(32'hbbad68ba),
	.w2(32'hbb6e4776),
	.w3(32'hbbbd27ee),
	.w4(32'hbb6e8cae),
	.w5(32'h3b5bf3ce),
	.w6(32'hbbadaae8),
	.w7(32'hbbb664fc),
	.w8(32'h39c11bb9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac01fd5),
	.w1(32'h3a936336),
	.w2(32'h3bbafa7e),
	.w3(32'h3b40aa11),
	.w4(32'h3c028370),
	.w5(32'hbaf28a59),
	.w6(32'h3b31d63a),
	.w7(32'h3bccadb1),
	.w8(32'h39b506fd),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7c2a5),
	.w1(32'hbb22b528),
	.w2(32'hbb64f599),
	.w3(32'hbb443e16),
	.w4(32'hbb52caf7),
	.w5(32'hbbc28a41),
	.w6(32'hbb4cafad),
	.w7(32'hbb7b5204),
	.w8(32'hbaf0a38c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f71ea),
	.w1(32'hbc18df75),
	.w2(32'h3a4cf502),
	.w3(32'hbc1b8510),
	.w4(32'hbb4eacf8),
	.w5(32'h3a3446d5),
	.w6(32'hbbda71a2),
	.w7(32'hba17063b),
	.w8(32'h39c2a467),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9685e0),
	.w1(32'h3ad4aa19),
	.w2(32'hb9e00dd4),
	.w3(32'hbb4a5ede),
	.w4(32'hbb8e577b),
	.w5(32'h3ad9f6de),
	.w6(32'hbb8a2636),
	.w7(32'hb8ba6d35),
	.w8(32'h3bd2ab64),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a8d4f),
	.w1(32'hbb4c3e43),
	.w2(32'hba2f96fd),
	.w3(32'h3b085e03),
	.w4(32'h3a5aae23),
	.w5(32'hba3b3e29),
	.w6(32'hbb5059be),
	.w7(32'hbb0e7984),
	.w8(32'h3c22d056),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5ded),
	.w1(32'hbba395c1),
	.w2(32'hbb842faf),
	.w3(32'hbbc4073f),
	.w4(32'hbbb59b16),
	.w5(32'hbaed27ee),
	.w6(32'hbbeb0399),
	.w7(32'hbb2282f5),
	.w8(32'hba19ce5f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f0e5f),
	.w1(32'hbb35b8dc),
	.w2(32'h3a83d0a4),
	.w3(32'hba99c9cc),
	.w4(32'h38a01610),
	.w5(32'h3b094a4d),
	.w6(32'hbbeec46c),
	.w7(32'h3b2010b5),
	.w8(32'h3b2031a1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b760a3e),
	.w1(32'hbb04de34),
	.w2(32'hbb1221d2),
	.w3(32'hbbbbb928),
	.w4(32'hbb6c40e9),
	.w5(32'h3aa638af),
	.w6(32'hbbbe4f81),
	.w7(32'hbbb34c97),
	.w8(32'h3b160d43),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32c7ce),
	.w1(32'hbae4fdb2),
	.w2(32'hba3cc12b),
	.w3(32'hba93f952),
	.w4(32'hbab3e4b4),
	.w5(32'h38a960c4),
	.w6(32'hbacbd536),
	.w7(32'hbb982469),
	.w8(32'h3b8e263f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ff0f7),
	.w1(32'hbb0c09cc),
	.w2(32'h3a42ca8b),
	.w3(32'hbaed4032),
	.w4(32'hbaa75586),
	.w5(32'hbac0268b),
	.w6(32'hbb6b6e23),
	.w7(32'hba413ba0),
	.w8(32'h3a8de0a7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af95047),
	.w1(32'hba050979),
	.w2(32'hba56ee40),
	.w3(32'hba865c6a),
	.w4(32'hba091463),
	.w5(32'h3bbad706),
	.w6(32'hbb0d9c40),
	.w7(32'hbb1f494b),
	.w8(32'hbb9104da),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81c826),
	.w1(32'hba253119),
	.w2(32'h3b19006e),
	.w3(32'h3c309f4b),
	.w4(32'h3c43b3e0),
	.w5(32'h3a92334e),
	.w6(32'hbb19adfd),
	.w7(32'h3b744e8d),
	.w8(32'hb90c7da7),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fe66e),
	.w1(32'h3ad54f94),
	.w2(32'h3b3427e8),
	.w3(32'hba866398),
	.w4(32'hbadc56c0),
	.w5(32'h3b867c1a),
	.w6(32'hbb5411c1),
	.w7(32'hbb1782c3),
	.w8(32'h3b92830a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf136c),
	.w1(32'h3a1dedfc),
	.w2(32'hbaf15362),
	.w3(32'hbb54672d),
	.w4(32'hbb9f4ede),
	.w5(32'hba82558e),
	.w6(32'hba04ffed),
	.w7(32'hbb3e40a7),
	.w8(32'hbbdb1dd7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9687dd),
	.w1(32'hbb01f7ab),
	.w2(32'hb97dea1f),
	.w3(32'hbb19d9b6),
	.w4(32'h3a0ef084),
	.w5(32'h3b5bc2d6),
	.w6(32'hbb8aac9e),
	.w7(32'h3ac58362),
	.w8(32'h3bdf576e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13fc2c),
	.w1(32'hba8dbeb1),
	.w2(32'hbb6eabe5),
	.w3(32'hbb6fb26b),
	.w4(32'hbbe5d311),
	.w5(32'h3b32cb9a),
	.w6(32'hba0cf45f),
	.w7(32'hbbadedcf),
	.w8(32'h3b64603b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3713db),
	.w1(32'hbba1ab61),
	.w2(32'hbab57f16),
	.w3(32'hbb239ccc),
	.w4(32'hbbbf55e1),
	.w5(32'hbbc299fb),
	.w6(32'hbb8eba1e),
	.w7(32'hbb681ac1),
	.w8(32'hbb90b120),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73a6c2),
	.w1(32'hb9e7dfc9),
	.w2(32'h3ac6943e),
	.w3(32'h3b1b741c),
	.w4(32'h3af3614a),
	.w5(32'h3a533bbd),
	.w6(32'hbba2c0d6),
	.w7(32'h3aaa7f46),
	.w8(32'h3aa52fa9),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a889c),
	.w1(32'h3aa9b3e8),
	.w2(32'h398bbae0),
	.w3(32'h3ae73e16),
	.w4(32'hb99e4dd8),
	.w5(32'hbba8c7b0),
	.w6(32'hb9a027c9),
	.w7(32'h3aee5c16),
	.w8(32'hbbcf1212),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e7657),
	.w1(32'h3b354a51),
	.w2(32'hb9d29811),
	.w3(32'hba899aac),
	.w4(32'hba9b1057),
	.w5(32'hb96b6e59),
	.w6(32'h3b639399),
	.w7(32'hba33d172),
	.w8(32'h3b18cc88),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a115e35),
	.w1(32'hbbfa9623),
	.w2(32'h3a454bf5),
	.w3(32'hbbce5663),
	.w4(32'hba040fbc),
	.w5(32'hb9e10887),
	.w6(32'hbbabd2ce),
	.w7(32'h3b0e5aba),
	.w8(32'h3b5c82b4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b486535),
	.w1(32'h3a77cb06),
	.w2(32'h3ac8c438),
	.w3(32'hba07818f),
	.w4(32'h3967d4f4),
	.w5(32'hbb88ad13),
	.w6(32'h3b968cf6),
	.w7(32'h3b5b5794),
	.w8(32'hbb817beb),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ca23b),
	.w1(32'h3b6e1b00),
	.w2(32'hbad2298b),
	.w3(32'h3bbe840c),
	.w4(32'h3b142d52),
	.w5(32'h38852af0),
	.w6(32'h3be87d6f),
	.w7(32'hb9163889),
	.w8(32'h3b57c681),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00ee68),
	.w1(32'hbb8036c7),
	.w2(32'hba92c2ec),
	.w3(32'hbb829bab),
	.w4(32'hbba48eea),
	.w5(32'hbb0354db),
	.w6(32'hbbb9d7a5),
	.w7(32'h3976c266),
	.w8(32'hbb180629),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e5d2),
	.w1(32'hbb6e9a63),
	.w2(32'h3a7ffe77),
	.w3(32'hbb66d1b6),
	.w4(32'hb9c2769c),
	.w5(32'h3b8d607a),
	.w6(32'hba83bc6e),
	.w7(32'h3b0d20b4),
	.w8(32'h3b40b941),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22aa1f),
	.w1(32'h3ba62b3d),
	.w2(32'h3b3277c3),
	.w3(32'h3add73ff),
	.w4(32'h3b5ee851),
	.w5(32'hb8894f9e),
	.w6(32'h3b8c5588),
	.w7(32'h3be401ca),
	.w8(32'hbaa6f4ed),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f3a1a),
	.w1(32'h3b2bd4de),
	.w2(32'h3b41f21c),
	.w3(32'h3b12e62d),
	.w4(32'h3ae6fb1b),
	.w5(32'h3ba46296),
	.w6(32'h387b47b4),
	.w7(32'h3af0537c),
	.w8(32'hbb62562e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886f18),
	.w1(32'h3aa9d6d2),
	.w2(32'h3b8c5f35),
	.w3(32'h3b72c65b),
	.w4(32'h3bd1653c),
	.w5(32'hbb90d89f),
	.w6(32'h3b174820),
	.w7(32'h3bcfca4b),
	.w8(32'hbb3749ce),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f205d),
	.w1(32'hbac6fe44),
	.w2(32'h3a6819e4),
	.w3(32'h3a131023),
	.w4(32'hbb596e6f),
	.w5(32'hbae10176),
	.w6(32'hbb4bbb66),
	.w7(32'hbb906606),
	.w8(32'hb9ffee50),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb02730),
	.w1(32'hbb8c81ba),
	.w2(32'hbb7ff37c),
	.w3(32'hbb7d912e),
	.w4(32'hbbd40281),
	.w5(32'hbb3c93cd),
	.w6(32'hbb8e1729),
	.w7(32'hbbcec938),
	.w8(32'hbb55f2f5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4297f7),
	.w1(32'h3bb08d38),
	.w2(32'h3ba04f0c),
	.w3(32'h3c261d1a),
	.w4(32'h3b48cd82),
	.w5(32'hbb3a2b3f),
	.w6(32'h3c1ddf1b),
	.w7(32'h3bb5cdca),
	.w8(32'hbb6317a2),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93f6ce),
	.w1(32'hba22b8af),
	.w2(32'hba091fca),
	.w3(32'hbb5024e7),
	.w4(32'hbb862465),
	.w5(32'hbb8280e3),
	.w6(32'hbb86694f),
	.w7(32'hbb12cf96),
	.w8(32'hbab3a333),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd560eb),
	.w1(32'h3c1aeb80),
	.w2(32'h3c0150fa),
	.w3(32'h3c8fb418),
	.w4(32'h3c9769a4),
	.w5(32'hbb994d6e),
	.w6(32'h3cd06158),
	.w7(32'h3c8abd26),
	.w8(32'hbc8623c9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bca08),
	.w1(32'hbbb75257),
	.w2(32'h3b9735da),
	.w3(32'h3a9e03f3),
	.w4(32'h3c1e3153),
	.w5(32'h3b07862b),
	.w6(32'hbba8bae9),
	.w7(32'h3bf4aaef),
	.w8(32'h3a957946),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacdfc3),
	.w1(32'hbac067e6),
	.w2(32'h39f33a56),
	.w3(32'hba591449),
	.w4(32'hbb046d4a),
	.w5(32'hbb2be3ea),
	.w6(32'hba21ad1b),
	.w7(32'hba9272a3),
	.w8(32'hb9f7f912),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa3ab3),
	.w1(32'hbba899f4),
	.w2(32'hbb8b4017),
	.w3(32'hbac0edc1),
	.w4(32'hbbc2c63e),
	.w5(32'h3ae002e8),
	.w6(32'hbb81971e),
	.w7(32'hbc03c635),
	.w8(32'hbb457745),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb500d77),
	.w1(32'h3a5a901b),
	.w2(32'hbb32b71c),
	.w3(32'h3b0de653),
	.w4(32'hba4c86b1),
	.w5(32'h3ab5e26b),
	.w6(32'hbb102131),
	.w7(32'hbb6fb662),
	.w8(32'h3aa9558b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5126bf),
	.w1(32'h3a5f1cf5),
	.w2(32'h3a93b8ac),
	.w3(32'h383191e3),
	.w4(32'hbad942f9),
	.w5(32'hbaedaaa9),
	.w6(32'hbb623b8e),
	.w7(32'hbae1524f),
	.w8(32'h3b69f6ef),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac68490),
	.w1(32'hbbf26e6b),
	.w2(32'hbb399497),
	.w3(32'hbafa8a0d),
	.w4(32'hbba8e4a1),
	.w5(32'hbb67bac6),
	.w6(32'hbba70975),
	.w7(32'hbb326ba0),
	.w8(32'hbbe34e53),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18ca5f),
	.w1(32'h3b1eeb09),
	.w2(32'h3acf8c83),
	.w3(32'h3ac0b77f),
	.w4(32'h3a711f88),
	.w5(32'hbb2704de),
	.w6(32'hbb7c7364),
	.w7(32'h3a578347),
	.w8(32'hbb0a005c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa41f81),
	.w1(32'hba54aa6d),
	.w2(32'hba557b8d),
	.w3(32'hbb4a1273),
	.w4(32'hbb4a91b7),
	.w5(32'hbad5e59f),
	.w6(32'hbb85cd19),
	.w7(32'hbb0b85b2),
	.w8(32'h3a35e9cc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87583c),
	.w1(32'hbb48a7a7),
	.w2(32'hba1989a0),
	.w3(32'h3b8e23ff),
	.w4(32'h3bc424db),
	.w5(32'hbb1f8109),
	.w6(32'h3b00e0d8),
	.w7(32'hb94afbdd),
	.w8(32'h3aa2667a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a240f82),
	.w1(32'h3bad6356),
	.w2(32'hbaab4693),
	.w3(32'h3b4b2768),
	.w4(32'h3b95c99c),
	.w5(32'hbab8d1b8),
	.w6(32'h3b9ab792),
	.w7(32'h3ba9fbc6),
	.w8(32'h3aa8a1cc),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2af34c),
	.w1(32'hbb42df6b),
	.w2(32'hba5d7e6b),
	.w3(32'hba60ac49),
	.w4(32'hba970440),
	.w5(32'h39906658),
	.w6(32'hbb437bac),
	.w7(32'h39dd2e42),
	.w8(32'h39bdf526),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1382e),
	.w1(32'hbc1a1b01),
	.w2(32'hbc03e9c7),
	.w3(32'hbc063a2c),
	.w4(32'hbb2c3b6d),
	.w5(32'h3b08d8fe),
	.w6(32'hbbf17bb3),
	.w7(32'hbbce2709),
	.w8(32'h3ac40622),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22974e),
	.w1(32'h3b2465be),
	.w2(32'h3bc292a3),
	.w3(32'h3895067e),
	.w4(32'h3b391abc),
	.w5(32'h3a1fa92f),
	.w6(32'h39835447),
	.w7(32'h3b77ab89),
	.w8(32'h3b0205f7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8e26),
	.w1(32'h3a2ac9b0),
	.w2(32'h3b40ecef),
	.w3(32'h3abff945),
	.w4(32'h3b89c9b3),
	.w5(32'hbc01bf57),
	.w6(32'h3b616b72),
	.w7(32'h3b92bab3),
	.w8(32'hbc206aee),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44bbb),
	.w1(32'h3b8f274c),
	.w2(32'h3baf04ac),
	.w3(32'h3af96930),
	.w4(32'h3b7c0e95),
	.w5(32'hbb0d9da7),
	.w6(32'hbb405640),
	.w7(32'h3b0e8429),
	.w8(32'hbbd84b33),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fac06),
	.w1(32'h3c36ff3f),
	.w2(32'h3bbb5f1f),
	.w3(32'h3c2ca1eb),
	.w4(32'h3bb4c9e0),
	.w5(32'hbbddc038),
	.w6(32'h3c2ee03c),
	.w7(32'h3ba68119),
	.w8(32'hbac58b89),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba337bcc),
	.w1(32'hbb7040b7),
	.w2(32'hb8b1089d),
	.w3(32'hbbbd260b),
	.w4(32'h3a2b9ef0),
	.w5(32'hb9ef4d29),
	.w6(32'hb951ec28),
	.w7(32'hbb8fde22),
	.w8(32'hba386a44),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce46ed),
	.w1(32'hba60b4cc),
	.w2(32'hba8ad753),
	.w3(32'hb9102326),
	.w4(32'hb9507cbf),
	.w5(32'h3b263c11),
	.w6(32'hba869bd8),
	.w7(32'hba58a9ca),
	.w8(32'h3b4765c2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa77726),
	.w1(32'h3a637bd0),
	.w2(32'h3ade4f66),
	.w3(32'h3b14ab8a),
	.w4(32'h3a32d91c),
	.w5(32'hba00d090),
	.w6(32'h39ab7c95),
	.w7(32'h3ac1daa6),
	.w8(32'hb9c3fe50),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39806f95),
	.w1(32'h3a6108f0),
	.w2(32'h3a0a470d),
	.w3(32'h37ee5149),
	.w4(32'h39eb098c),
	.w5(32'hba3b6fa1),
	.w6(32'hbb0eaa3a),
	.w7(32'hba98c861),
	.w8(32'hbb191f16),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48eba3),
	.w1(32'hba941898),
	.w2(32'hba24dfc8),
	.w3(32'hbac50c05),
	.w4(32'hbab854a0),
	.w5(32'h37853a43),
	.w6(32'hba8c72e6),
	.w7(32'hba96b409),
	.w8(32'hb9362546),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac663a2),
	.w1(32'hba433214),
	.w2(32'hbb50a78d),
	.w3(32'h3acff048),
	.w4(32'h39de6927),
	.w5(32'h3a48f8ce),
	.w6(32'hba164378),
	.w7(32'hbac10c8f),
	.w8(32'h3a018e41),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c35bb),
	.w1(32'hb899aca5),
	.w2(32'h3a094afe),
	.w3(32'h3aafa404),
	.w4(32'h3ab367e2),
	.w5(32'h3a9b5354),
	.w6(32'h39f1dbc8),
	.w7(32'h3a62dc2d),
	.w8(32'hba4cd869),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a348b49),
	.w1(32'hb7e2ba88),
	.w2(32'hb89b25c3),
	.w3(32'h38aa3ce9),
	.w4(32'hba4a8dcc),
	.w5(32'h38cec4a1),
	.w6(32'hba85eabf),
	.w7(32'hb9b58e68),
	.w8(32'hb91d1fa7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c283da),
	.w1(32'hbaee12b4),
	.w2(32'hbb1ae8ba),
	.w3(32'h3a1861b6),
	.w4(32'hba8fc0ff),
	.w5(32'h3adc5819),
	.w6(32'hb9add3cc),
	.w7(32'hbb126b0a),
	.w8(32'h398e5fdc),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bd1a2),
	.w1(32'h3adb8fa7),
	.w2(32'h3b0b4ef5),
	.w3(32'h3a6b7199),
	.w4(32'h3a91ed7c),
	.w5(32'h39ff35cb),
	.w6(32'h3b20b21e),
	.w7(32'h3ad54293),
	.w8(32'h3a273aaf),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c92a5),
	.w1(32'hba24915c),
	.w2(32'hb7a3ee99),
	.w3(32'hb9adfe0e),
	.w4(32'h389623ca),
	.w5(32'hba0d8745),
	.w6(32'hb9d9a542),
	.w7(32'h38f08a55),
	.w8(32'hba8d4f6c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba089c8f),
	.w1(32'hba15b4ae),
	.w2(32'h3a4e486c),
	.w3(32'hba8e9c3c),
	.w4(32'h39f45d34),
	.w5(32'hba95c4e1),
	.w6(32'hbb03240f),
	.w7(32'hb83ada65),
	.w8(32'hba84fdf2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba777e53),
	.w1(32'hbac4a4ce),
	.w2(32'hba845969),
	.w3(32'hbaac35c8),
	.w4(32'hba25611b),
	.w5(32'h3868d416),
	.w6(32'hbb009a46),
	.w7(32'hba98bcc0),
	.w8(32'h3a36e3fa),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72e6aa),
	.w1(32'h3a412b34),
	.w2(32'hb9239c25),
	.w3(32'h3a40fe52),
	.w4(32'hb82e6c1f),
	.w5(32'hb704d7c0),
	.w6(32'h3a24b873),
	.w7(32'h395f407d),
	.w8(32'hba9c6e95),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb302e51),
	.w1(32'hbb4edc7c),
	.w2(32'hbac2e4a8),
	.w3(32'hbaad67ef),
	.w4(32'hbabfa1c9),
	.w5(32'hba5355b2),
	.w6(32'hba516b11),
	.w7(32'hbae32adf),
	.w8(32'hbb191a8f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfe134),
	.w1(32'hbb468bdc),
	.w2(32'hbb55ca72),
	.w3(32'hba9e8939),
	.w4(32'hbb075251),
	.w5(32'hb9ad9bcd),
	.w6(32'hbb036311),
	.w7(32'hbb3a67ec),
	.w8(32'hba4d947e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b59619),
	.w1(32'hba9e78b7),
	.w2(32'hbac11f46),
	.w3(32'h3a65b0e1),
	.w4(32'h39e7f80d),
	.w5(32'h3a0fe4e7),
	.w6(32'h3a0f617d),
	.w7(32'hb745c3e5),
	.w8(32'h3aadfedb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b39a),
	.w1(32'hb91fedda),
	.w2(32'hba30a275),
	.w3(32'hba742aa5),
	.w4(32'hba48ab72),
	.w5(32'hb9b65072),
	.w6(32'hba5c8133),
	.w7(32'hbad14c2c),
	.w8(32'hba79e3b5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b535b),
	.w1(32'hbab00b08),
	.w2(32'hb90c018c),
	.w3(32'hba695466),
	.w4(32'hba7c9910),
	.w5(32'hb9cad3c5),
	.w6(32'hb98a5e6f),
	.w7(32'hba49940a),
	.w8(32'hb9a04d0d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944af1e),
	.w1(32'hb98340f0),
	.w2(32'hba085f64),
	.w3(32'hb8c2cb5d),
	.w4(32'h397c8928),
	.w5(32'hba1ff6db),
	.w6(32'hb976fdf3),
	.w7(32'h3817fbb4),
	.w8(32'hbaaee1b6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba827e6e),
	.w1(32'hbab942bc),
	.w2(32'h37a444ef),
	.w3(32'hba5aab26),
	.w4(32'h3a807e45),
	.w5(32'hb97e7a57),
	.w6(32'hbad388c3),
	.w7(32'h3749e375),
	.w8(32'hb999e82f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf28c4c),
	.w1(32'hbb11d372),
	.w2(32'hbaa9f663),
	.w3(32'hbb01d55b),
	.w4(32'hba04a20b),
	.w5(32'hba5dc30b),
	.w6(32'hbb214dff),
	.w7(32'hbab32dd4),
	.w8(32'hbae70542),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6802e7),
	.w1(32'hbb040c22),
	.w2(32'hbb01a28e),
	.w3(32'hbab67e3c),
	.w4(32'hba80d793),
	.w5(32'hbab2b1fb),
	.w6(32'hbb1727ff),
	.w7(32'hbae6755d),
	.w8(32'hba8eb990),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed5128),
	.w1(32'h38b9f661),
	.w2(32'hba0ee318),
	.w3(32'hbac92217),
	.w4(32'hba6bef18),
	.w5(32'h38c6594c),
	.w6(32'hb8ac08b0),
	.w7(32'hb9a14530),
	.w8(32'h385b9b63),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b2bad),
	.w1(32'hba89cfb7),
	.w2(32'hba11786b),
	.w3(32'hba3dab8a),
	.w4(32'hba8d86f9),
	.w5(32'hba15cf54),
	.w6(32'hb67b77ac),
	.w7(32'hbab04181),
	.w8(32'hba7c984e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98cb67),
	.w1(32'hba561008),
	.w2(32'hb8ed7a9b),
	.w3(32'h3987117d),
	.w4(32'h38520607),
	.w5(32'hba880b42),
	.w6(32'h3822ab5a),
	.w7(32'hba9083a6),
	.w8(32'hba617679),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c9a4c),
	.w1(32'hba85aa6b),
	.w2(32'hbaa77f52),
	.w3(32'hba948c71),
	.w4(32'hba1a9178),
	.w5(32'h39c84827),
	.w6(32'hba662deb),
	.w7(32'hba667559),
	.w8(32'hba106f6e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d9fc5),
	.w1(32'hbaa875f6),
	.w2(32'hb9d0b81f),
	.w3(32'h3a073523),
	.w4(32'h3a107e1a),
	.w5(32'hbab48aca),
	.w6(32'h3a972e4e),
	.w7(32'hb9b34fdd),
	.w8(32'hbac51344),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77b814),
	.w1(32'hbb8459e2),
	.w2(32'hbae68129),
	.w3(32'hbb79591f),
	.w4(32'hbb1bdeb7),
	.w5(32'h3a8d568d),
	.w6(32'hbb70065c),
	.w7(32'hbb10161e),
	.w8(32'h39d621dd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d55a0c),
	.w1(32'hba7291c1),
	.w2(32'hb9d7e5fe),
	.w3(32'h3916d8c2),
	.w4(32'h39f2ca52),
	.w5(32'hb892883d),
	.w6(32'hba78c08d),
	.w7(32'h37e62ea8),
	.w8(32'h3a264d08),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a876ef6),
	.w1(32'h3af94f98),
	.w2(32'h39597b8a),
	.w3(32'h39859bc2),
	.w4(32'hbaa0d97e),
	.w5(32'hbad2c21f),
	.w6(32'hbb2d2e6c),
	.w7(32'hbb6997e7),
	.w8(32'hbb6730a4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule