module layer_10_featuremap_431(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9b1e),
	.w1(32'hbb8d32a5),
	.w2(32'hbae3263d),
	.w3(32'hbb7300f3),
	.w4(32'h3bac4167),
	.w5(32'h3c24568b),
	.w6(32'hbb8ce6ff),
	.w7(32'hba0b487c),
	.w8(32'h3aca5b78),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7a9cc),
	.w1(32'h3ac1e55d),
	.w2(32'hbb0fdf78),
	.w3(32'h3c20fa6e),
	.w4(32'hbbd1c3bd),
	.w5(32'hbb8bc6b3),
	.w6(32'h3a89f38b),
	.w7(32'hbb23b211),
	.w8(32'hbb83ed5c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1051c6),
	.w1(32'hbb66d1ae),
	.w2(32'hbb380228),
	.w3(32'h3b236ca5),
	.w4(32'hba9322e6),
	.w5(32'h3b22d72f),
	.w6(32'hb8bc35b4),
	.w7(32'h3a4ad2e8),
	.w8(32'h3a0d22fb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2266a),
	.w1(32'h3c09586a),
	.w2(32'h3b813e93),
	.w3(32'hbb32e511),
	.w4(32'hbb439b3e),
	.w5(32'hbac3243f),
	.w6(32'hbbd15931),
	.w7(32'h3b0f81f5),
	.w8(32'h3bbbe2f9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba896022),
	.w1(32'h3968e98c),
	.w2(32'h3b106c17),
	.w3(32'h3b927ffe),
	.w4(32'h3ada969f),
	.w5(32'h3aedb657),
	.w6(32'h3b84e88f),
	.w7(32'hbaaa2ca0),
	.w8(32'h3a0bca01),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa46888),
	.w1(32'hbb06a2bc),
	.w2(32'hbb8cde26),
	.w3(32'hb9d861e6),
	.w4(32'hb926ad89),
	.w5(32'hbbc35202),
	.w6(32'h3b4dff90),
	.w7(32'h3ba33cc4),
	.w8(32'h3b83f94b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdedb4d),
	.w1(32'h3bcfff23),
	.w2(32'h3c096a17),
	.w3(32'h3a8473a7),
	.w4(32'h3c2421cb),
	.w5(32'h3c7bc4ba),
	.w6(32'h3bca82e0),
	.w7(32'h3bc3ac47),
	.w8(32'h3ad6a8f6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f0232),
	.w1(32'hbc0a4cbd),
	.w2(32'hbc242a96),
	.w3(32'hbc16f6ca),
	.w4(32'hbbf5696e),
	.w5(32'hbc8cd06d),
	.w6(32'hbb0334c8),
	.w7(32'h3c1cef8d),
	.w8(32'h3c021fd9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05f748),
	.w1(32'hbb024374),
	.w2(32'h3a95bfd8),
	.w3(32'hbb78a1d9),
	.w4(32'hbb72bea8),
	.w5(32'hbb60e01e),
	.w6(32'h3ac8afbf),
	.w7(32'hbc16ce88),
	.w8(32'h393fc4cf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a36bc),
	.w1(32'hbba74246),
	.w2(32'hbb9d2c84),
	.w3(32'hbb0fea82),
	.w4(32'hba893090),
	.w5(32'h3ba2406f),
	.w6(32'hb78b89db),
	.w7(32'h3c31b964),
	.w8(32'h3ac34d9d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76e34b),
	.w1(32'h3b5f9af5),
	.w2(32'h3c27a47b),
	.w3(32'h3b0aecc1),
	.w4(32'h3b53e870),
	.w5(32'h3bee1c05),
	.w6(32'h3ac0fd8f),
	.w7(32'hbb3aaaa1),
	.w8(32'hbb1d5c09),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8d8c0),
	.w1(32'h3bc371c9),
	.w2(32'hbaa986e4),
	.w3(32'h3b476917),
	.w4(32'h3bcaae0d),
	.w5(32'h3c0e6bdb),
	.w6(32'h3b583b1e),
	.w7(32'h3bf942e2),
	.w8(32'h3c21dd55),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d8afc),
	.w1(32'h3b8ab592),
	.w2(32'hbc12911d),
	.w3(32'hba82d6b0),
	.w4(32'hbb3476c2),
	.w5(32'h3bd7d0f3),
	.w6(32'h3aca2a7b),
	.w7(32'h3b9b2188),
	.w8(32'h3c0608ac),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13ec8b),
	.w1(32'hba447ce9),
	.w2(32'hbb4f121f),
	.w3(32'h3c1b7114),
	.w4(32'hb7e8a4a0),
	.w5(32'h3b82dc08),
	.w6(32'h3b97c8d7),
	.w7(32'h3b5680ca),
	.w8(32'hba5bc024),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05ac8f),
	.w1(32'hbbae0ea6),
	.w2(32'hbb52927c),
	.w3(32'h38f11d37),
	.w4(32'hbb998f3c),
	.w5(32'hbb2b68bf),
	.w6(32'h3b5881b2),
	.w7(32'h3b2777b4),
	.w8(32'h3b07c15b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51a0f1),
	.w1(32'hbc26803d),
	.w2(32'hbbca3f91),
	.w3(32'hbaff9d3d),
	.w4(32'hbc8abf54),
	.w5(32'hbc382ea5),
	.w6(32'h3bdf3b3f),
	.w7(32'hbb4e314b),
	.w8(32'hbbd68b55),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb628167),
	.w1(32'h3a241245),
	.w2(32'h3abb293c),
	.w3(32'hbba2975f),
	.w4(32'hbb144c5f),
	.w5(32'hba3a2f4f),
	.w6(32'hba236f82),
	.w7(32'hbbbdf2e0),
	.w8(32'hbb2300a4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fcf11),
	.w1(32'hbc233e55),
	.w2(32'h39e6eae7),
	.w3(32'hbb20f488),
	.w4(32'hbb2f00b7),
	.w5(32'hbbb93297),
	.w6(32'hb8a88043),
	.w7(32'h3bad23a6),
	.w8(32'h3bcfbd03),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4fdce),
	.w1(32'hbbb4a258),
	.w2(32'hb955f63e),
	.w3(32'hbbd0c0d4),
	.w4(32'h3a937584),
	.w5(32'h3b54d3ec),
	.w6(32'hb96d42f3),
	.w7(32'h3bada391),
	.w8(32'h3b3c3943),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ba658),
	.w1(32'h3b63ee1f),
	.w2(32'h390fba83),
	.w3(32'h3b31107d),
	.w4(32'hbbaf9e3b),
	.w5(32'hba4d1b11),
	.w6(32'hbaed8229),
	.w7(32'h3a4a352e),
	.w8(32'hbb57e519),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90a338),
	.w1(32'hba1c3735),
	.w2(32'hbb102ecd),
	.w3(32'hbb8e2d9c),
	.w4(32'h3b541696),
	.w5(32'h3a4bb466),
	.w6(32'h3aacd46e),
	.w7(32'h3b383fc9),
	.w8(32'h3aa75cb9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2d9c3),
	.w1(32'h3ba9e967),
	.w2(32'h3b2bb5ef),
	.w3(32'h3bbc8b53),
	.w4(32'h3b54e489),
	.w5(32'h3b1bf532),
	.w6(32'h3abbd3d6),
	.w7(32'h3b2a180e),
	.w8(32'hbb3477de),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28d265),
	.w1(32'hbc3ded05),
	.w2(32'hbc7fdd4c),
	.w3(32'hb9802e5a),
	.w4(32'hbb0f2377),
	.w5(32'hbb42407e),
	.w6(32'h3b1dec3e),
	.w7(32'h3c241f7e),
	.w8(32'h3c5503f8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987b1e),
	.w1(32'h3b5b94aa),
	.w2(32'hb89c141b),
	.w3(32'h3ac52b54),
	.w4(32'hbb1cde36),
	.w5(32'hbbb94f4c),
	.w6(32'h3a797041),
	.w7(32'h3bbdb585),
	.w8(32'hba86bf42),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c681b),
	.w1(32'h3c6d5bd2),
	.w2(32'h3c063743),
	.w3(32'h3bc68ff8),
	.w4(32'h3c0ae047),
	.w5(32'hba07366f),
	.w6(32'h3b8bb287),
	.w7(32'h3a91f0c1),
	.w8(32'hbb7cf861),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc7c09),
	.w1(32'h3aeca844),
	.w2(32'hbbaa237e),
	.w3(32'h3bb1a41d),
	.w4(32'h3a88c94a),
	.w5(32'hbb168c79),
	.w6(32'h3aa2e2ec),
	.w7(32'h3bd0c874),
	.w8(32'h3a8ac8e4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb384623),
	.w1(32'h3bd19b42),
	.w2(32'h3b801373),
	.w3(32'h3b42f065),
	.w4(32'h3ba95e6f),
	.w5(32'h3b8c96c0),
	.w6(32'h3b9377e2),
	.w7(32'hbb98e0dd),
	.w8(32'hb9b34438),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90094df),
	.w1(32'h3a9d5fb6),
	.w2(32'h3c4fe36f),
	.w3(32'h3b07396d),
	.w4(32'hbbbeb0b5),
	.w5(32'hba77afa8),
	.w6(32'h3b1416ea),
	.w7(32'hbb551213),
	.w8(32'hbc1282aa),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12839a),
	.w1(32'hbb4d184b),
	.w2(32'hb9d032e1),
	.w3(32'h3b519aa8),
	.w4(32'hbaba4dc7),
	.w5(32'h3b494e4d),
	.w6(32'h3b110dbe),
	.w7(32'h3b51e052),
	.w8(32'h39f6fb57),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c722eef),
	.w1(32'h3c6d0bef),
	.w2(32'h3c56a968),
	.w3(32'h3be74022),
	.w4(32'hbabf7165),
	.w5(32'h3b178c24),
	.w6(32'h3b91735c),
	.w7(32'hbac36588),
	.w8(32'hbb416826),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3edee),
	.w1(32'hbb593a96),
	.w2(32'hbb6d6e39),
	.w3(32'h3b300ccf),
	.w4(32'hbaa5f1f8),
	.w5(32'h3b1cf055),
	.w6(32'h39af4474),
	.w7(32'hb97aec29),
	.w8(32'h3b0e0d91),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd504b5),
	.w1(32'hbb78b7d5),
	.w2(32'hbbb53c26),
	.w3(32'h3bc227c1),
	.w4(32'hbb3d6c2f),
	.w5(32'hbbcee0f3),
	.w6(32'h3979b069),
	.w7(32'h3b08f39e),
	.w8(32'hbb4cb6a2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab8bae),
	.w1(32'h3a6ad9b9),
	.w2(32'h3b5fda75),
	.w3(32'hbb3fa7d2),
	.w4(32'h3bffdc4a),
	.w5(32'h3c971396),
	.w6(32'hb9aa00ba),
	.w7(32'h388e7d0f),
	.w8(32'hbbc0634a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26a989),
	.w1(32'h3a85b42a),
	.w2(32'hb936f819),
	.w3(32'h3bacabfc),
	.w4(32'h3afa80d1),
	.w5(32'h3be2e697),
	.w6(32'hbb732e49),
	.w7(32'h3a90ddba),
	.w8(32'hbb5b95e5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02d35f),
	.w1(32'hbace1652),
	.w2(32'hbbc30cf3),
	.w3(32'hbbb69d21),
	.w4(32'hbb579d05),
	.w5(32'hbc0330d8),
	.w6(32'hb7caa670),
	.w7(32'hba8dc89c),
	.w8(32'h3ada5beb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cf82c),
	.w1(32'h3b6bb9ac),
	.w2(32'hbb1bc50b),
	.w3(32'hbc405531),
	.w4(32'hbad91395),
	.w5(32'hbbbe8a18),
	.w6(32'h3b6d1fe2),
	.w7(32'h3b01f663),
	.w8(32'h3b9604a0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6169c1),
	.w1(32'hbc425a34),
	.w2(32'hbc16c9d6),
	.w3(32'hbbc37ceb),
	.w4(32'h3c311ea8),
	.w5(32'h3ca2cade),
	.w6(32'h3a677a1f),
	.w7(32'h3c0f972a),
	.w8(32'h3c92fcdb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3572e3),
	.w1(32'h3c6fa189),
	.w2(32'hba227054),
	.w3(32'h3c390f15),
	.w4(32'hbb22ed38),
	.w5(32'hbb5b669e),
	.w6(32'h3c5e07b8),
	.w7(32'h3b76a606),
	.w8(32'hbb90b2f7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6ddf6),
	.w1(32'h3c5e399c),
	.w2(32'h3c33a214),
	.w3(32'h3c6f4d75),
	.w4(32'h3b929ca4),
	.w5(32'h3b9b3a81),
	.w6(32'h3c10db96),
	.w7(32'hbb49de12),
	.w8(32'hbba02eb1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dc7ba),
	.w1(32'h3b5b72eb),
	.w2(32'hba2295d6),
	.w3(32'h3b31b590),
	.w4(32'hbad72e83),
	.w5(32'hbb804393),
	.w6(32'hb9e640b0),
	.w7(32'h3b0079f8),
	.w8(32'hbac2731b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1858bf),
	.w1(32'hbbc5090b),
	.w2(32'hbbea6998),
	.w3(32'h3a3f7a96),
	.w4(32'h3b5c4d9b),
	.w5(32'h3c31a0a6),
	.w6(32'hbb085103),
	.w7(32'h3a453416),
	.w8(32'hbb8e3c73),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ca2329),
	.w1(32'h3b8712a3),
	.w2(32'h3b223107),
	.w3(32'h3ab8d812),
	.w4(32'h3b98b77f),
	.w5(32'h3bd14545),
	.w6(32'h3b622c78),
	.w7(32'hbb152044),
	.w8(32'hbb1ba58d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fcf8a),
	.w1(32'h3aeef6d7),
	.w2(32'h3ae093fc),
	.w3(32'hba0c2534),
	.w4(32'hbaa9730c),
	.w5(32'hb926ea6f),
	.w6(32'h397429ab),
	.w7(32'h3b53f49a),
	.w8(32'hb9801703),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61d6cd),
	.w1(32'hbb72ebf4),
	.w2(32'h3b09e412),
	.w3(32'hbb860122),
	.w4(32'hba99a111),
	.w5(32'hbbb6dc20),
	.w6(32'h3a7e5212),
	.w7(32'h3c06a9c6),
	.w8(32'h3af81610),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f7eba),
	.w1(32'hbbb6b748),
	.w2(32'h3aeefc20),
	.w3(32'hbad2941d),
	.w4(32'h3b74b5ec),
	.w5(32'h3b858b76),
	.w6(32'h3b040c65),
	.w7(32'h3abdf09a),
	.w8(32'hbb2d2686),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace5999),
	.w1(32'hbbe068c3),
	.w2(32'hbafd9e50),
	.w3(32'hbb218fce),
	.w4(32'hbbc12cce),
	.w5(32'hbbcf689f),
	.w6(32'hb9b18b3f),
	.w7(32'h3a95c26a),
	.w8(32'h3bae3fb4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf7229),
	.w1(32'hbb2b3e17),
	.w2(32'hbb9c4738),
	.w3(32'hbbd660b6),
	.w4(32'hbba8814e),
	.w5(32'h3bd37b69),
	.w6(32'h3ba6d166),
	.w7(32'h3a3a5a14),
	.w8(32'h3b631ae0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0984fa),
	.w1(32'hbbf6ed31),
	.w2(32'h3a8e21bf),
	.w3(32'hbba76f95),
	.w4(32'h3af857f9),
	.w5(32'h3bb50347),
	.w6(32'h3bc6832e),
	.w7(32'h3c5a4254),
	.w8(32'h3c1b22b9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64e5b1),
	.w1(32'h3b637a9f),
	.w2(32'h3b18052c),
	.w3(32'hbab3c34f),
	.w4(32'hba375a48),
	.w5(32'hbb466b3f),
	.w6(32'hbadc3c9b),
	.w7(32'h39a44cae),
	.w8(32'hba652c1c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03f49e),
	.w1(32'h3b47e787),
	.w2(32'hbaa1ab19),
	.w3(32'hbabbeeb8),
	.w4(32'hba13d5c9),
	.w5(32'hbbd3a73c),
	.w6(32'hbad225f6),
	.w7(32'hbb3a3ab1),
	.w8(32'hbbb1006a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58c300),
	.w1(32'hb420fb28),
	.w2(32'hbb91e9a4),
	.w3(32'h3b0d105b),
	.w4(32'hb95f0095),
	.w5(32'hbb5f939c),
	.w6(32'h3b1ceb3e),
	.w7(32'hba01f4f8),
	.w8(32'h3ae4cda9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb541be3),
	.w1(32'hbc039f08),
	.w2(32'hbb5c7ef0),
	.w3(32'h3b82314e),
	.w4(32'hbbb96d08),
	.w5(32'hba014db1),
	.w6(32'h3b42f3dc),
	.w7(32'hbbb5ee0e),
	.w8(32'hbae5938e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb1dcd),
	.w1(32'hbad4369a),
	.w2(32'hbb440e86),
	.w3(32'hbb7c0343),
	.w4(32'hb95c3d2e),
	.w5(32'hba707e58),
	.w6(32'hbb4b9bd9),
	.w7(32'h3b2b8d5b),
	.w8(32'hbafb903d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f3aed),
	.w1(32'hbc0d7c01),
	.w2(32'hbb506ba3),
	.w3(32'hbbcfe496),
	.w4(32'h3a858977),
	.w5(32'hb91b0948),
	.w6(32'hb8293a27),
	.w7(32'h3c8655c7),
	.w8(32'h3c1f0285),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad41bfc),
	.w1(32'h3b857fd9),
	.w2(32'hbb0a31ea),
	.w3(32'hbb7b7fb7),
	.w4(32'h39d1bfe7),
	.w5(32'hbae4a75e),
	.w6(32'hbb1b75e1),
	.w7(32'h3b6d9fbc),
	.w8(32'hbb2c5cee),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bf971),
	.w1(32'h3bc71244),
	.w2(32'hbae5d55f),
	.w3(32'h3bcf237d),
	.w4(32'hbb35d42e),
	.w5(32'hbb2e7e5d),
	.w6(32'hbadfb90f),
	.w7(32'hbb8b45e7),
	.w8(32'hbb9d6dc3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5254e),
	.w1(32'hba77c67c),
	.w2(32'h3a2ab1b2),
	.w3(32'h3b300673),
	.w4(32'h3b7096ae),
	.w5(32'h3c0a1f03),
	.w6(32'hbba67840),
	.w7(32'hba49a6a1),
	.w8(32'h3b564339),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e754f),
	.w1(32'h3b06e947),
	.w2(32'h3a960741),
	.w3(32'h3bea44f9),
	.w4(32'hbaa27180),
	.w5(32'hba156e06),
	.w6(32'h3b699dc6),
	.w7(32'hbb8cf76b),
	.w8(32'h3b427223),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77b5fe),
	.w1(32'hbb228440),
	.w2(32'h3ab940d6),
	.w3(32'h3b5c5219),
	.w4(32'h3a1d28e1),
	.w5(32'h3af61f48),
	.w6(32'h3a864b5b),
	.w7(32'h39dcc73c),
	.w8(32'hba34e3d1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb617769),
	.w1(32'h3bed7da2),
	.w2(32'hbafb5191),
	.w3(32'hbb1a9570),
	.w4(32'h3b3097ce),
	.w5(32'h396c0f5e),
	.w6(32'hbb8b5f5f),
	.w7(32'h3c213865),
	.w8(32'h3bc0526a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb439557),
	.w1(32'h3b64c712),
	.w2(32'h3baf1764),
	.w3(32'h3c13c513),
	.w4(32'hbb3c93c3),
	.w5(32'hbbd4e93f),
	.w6(32'h3bf77b6a),
	.w7(32'h3b803107),
	.w8(32'h3b3df8f4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc98c14),
	.w1(32'hbc4f5af8),
	.w2(32'hbad9ca7d),
	.w3(32'hbb322659),
	.w4(32'hbc16f89e),
	.w5(32'hbbc81e54),
	.w6(32'h3a8dda33),
	.w7(32'hbba21167),
	.w8(32'hbb99a826),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf991bd),
	.w1(32'h3c01e1ef),
	.w2(32'hbaac8bc3),
	.w3(32'hbad49e8e),
	.w4(32'h3b4ab392),
	.w5(32'hbbea1506),
	.w6(32'h3a42ef4d),
	.w7(32'hba9b6025),
	.w8(32'hbc1a709d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cbb94),
	.w1(32'hba8a73bf),
	.w2(32'hbb9ef3a0),
	.w3(32'hbb9d318b),
	.w4(32'h3b04f3bb),
	.w5(32'h3c4a82b5),
	.w6(32'hbbc872f9),
	.w7(32'hbb671698),
	.w8(32'hb9b44745),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74d6a4),
	.w1(32'h3b76bc16),
	.w2(32'h3b82b4ec),
	.w3(32'h3c35b564),
	.w4(32'h3aca1261),
	.w5(32'h39adda8b),
	.w6(32'h39dc8f57),
	.w7(32'h3b123b30),
	.w8(32'h3b4cfe3f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bdf53),
	.w1(32'h3b59832c),
	.w2(32'h3b5f9816),
	.w3(32'h3b42cbf4),
	.w4(32'h3b218fe9),
	.w5(32'h3aadbf1f),
	.w6(32'h3b8f854c),
	.w7(32'hbb265fd2),
	.w8(32'hbb8cebd4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07a0c9),
	.w1(32'hbcc6c244),
	.w2(32'hbc7a7175),
	.w3(32'hba60eb7f),
	.w4(32'hbc8caef6),
	.w5(32'hbb976d23),
	.w6(32'h3b853ccd),
	.w7(32'h39736c2e),
	.w8(32'hbb8a2a7f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf2bd5),
	.w1(32'hba4dff1d),
	.w2(32'hbae06afc),
	.w3(32'h3b546006),
	.w4(32'hbbca93b2),
	.w5(32'hbbb2c8d9),
	.w6(32'hbb581245),
	.w7(32'h3baa162f),
	.w8(32'h3bad1a8d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa332d7),
	.w1(32'hbc594304),
	.w2(32'hbc0c4884),
	.w3(32'h39dbb154),
	.w4(32'hbb8c2efc),
	.w5(32'hba0ca49c),
	.w6(32'h39af406f),
	.w7(32'hbacaf7c6),
	.w8(32'h3b65c850),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b981d6e),
	.w1(32'h3bb82026),
	.w2(32'h3b6076c0),
	.w3(32'h3b22bfff),
	.w4(32'hba42f216),
	.w5(32'h3adf1e80),
	.w6(32'h3bd6068b),
	.w7(32'hbae9690d),
	.w8(32'hbb46406d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c57c7a),
	.w1(32'hb798aaf6),
	.w2(32'h3846e238),
	.w3(32'hb8d58149),
	.w4(32'h36f8ba6f),
	.w5(32'h37c32a78),
	.w6(32'hb8eeacba),
	.w7(32'h3709d523),
	.w8(32'h37860f78),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380e0eb4),
	.w1(32'hb89b3722),
	.w2(32'hb75b1b46),
	.w3(32'h37dece09),
	.w4(32'hb7b25a3f),
	.w5(32'h38095159),
	.w6(32'hb5a8907b),
	.w7(32'hb8d729cb),
	.w8(32'hb89c576c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942e4c9),
	.w1(32'hb908454e),
	.w2(32'h37467c8f),
	.w3(32'hb88bc053),
	.w4(32'hb9164504),
	.w5(32'hb74e183b),
	.w6(32'hb844dcde),
	.w7(32'hb90dc933),
	.w8(32'hb8926f23),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1da496),
	.w1(32'hbb04bcf4),
	.w2(32'hba6d93f7),
	.w3(32'hba678596),
	.w4(32'hb955cbac),
	.w5(32'hba094027),
	.w6(32'h3aa84e12),
	.w7(32'h3ad3fb2f),
	.w8(32'h39b78459),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f0b80),
	.w1(32'hb7eabb19),
	.w2(32'hb8af20a8),
	.w3(32'h38f53922),
	.w4(32'h38d80a4d),
	.w5(32'hb6740f60),
	.w6(32'h390767ee),
	.w7(32'h391c00bb),
	.w8(32'hb78f0379),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac3ede),
	.w1(32'hbbb0d172),
	.w2(32'hbb0a9bcd),
	.w3(32'hbb38651d),
	.w4(32'h3adf609c),
	.w5(32'h3b336ad5),
	.w6(32'h3abb89ad),
	.w7(32'h3bbae4d0),
	.w8(32'h3b94bb83),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0cc7b),
	.w1(32'hbbe5b58b),
	.w2(32'hbb827e6f),
	.w3(32'hbbac2061),
	.w4(32'hba1ab507),
	.w5(32'hba9d4518),
	.w6(32'hb88d81dd),
	.w7(32'h3beacfa2),
	.w8(32'h3c03c766),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b60dc),
	.w1(32'h3a77a68b),
	.w2(32'h3a8efb36),
	.w3(32'h3b5167a4),
	.w4(32'hbab99f03),
	.w5(32'h3a830b9a),
	.w6(32'h3bb6f2fd),
	.w7(32'h3abc0527),
	.w8(32'h3a90af90),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89de134),
	.w1(32'hbb64115b),
	.w2(32'hbb77a777),
	.w3(32'h3b551bce),
	.w4(32'hbab363e6),
	.w5(32'hbb9cc1a5),
	.w6(32'h3ba1f376),
	.w7(32'h3b20bffe),
	.w8(32'hba998160),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb689b53),
	.w1(32'hbbf8890f),
	.w2(32'hbb46519b),
	.w3(32'h39b31bf8),
	.w4(32'hba33df89),
	.w5(32'hbb1f091c),
	.w6(32'h3ba5be42),
	.w7(32'h3b65b62d),
	.w8(32'hbaca0430),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4f516),
	.w1(32'hba88255b),
	.w2(32'h3a1cbaa4),
	.w3(32'h39f5a4d4),
	.w4(32'hb9ec36d2),
	.w5(32'hb8fa5f04),
	.w6(32'h39e8f611),
	.w7(32'h3a33f660),
	.w8(32'hb9d9b83b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46e029),
	.w1(32'hbace6b18),
	.w2(32'hb981cb23),
	.w3(32'hb973cf64),
	.w4(32'h3ad0307e),
	.w5(32'h3aac0218),
	.w6(32'h3b27f6a1),
	.w7(32'h3baf7b61),
	.w8(32'h3b892c3f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9cbc7),
	.w1(32'hb7fdb66d),
	.w2(32'hb734babb),
	.w3(32'hb89aa7a1),
	.w4(32'hb454e514),
	.w5(32'h3700c28a),
	.w6(32'hb87a0fa9),
	.w7(32'h36839268),
	.w8(32'hb747c940),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3858e478),
	.w1(32'hb66a7d01),
	.w2(32'h3819f109),
	.w3(32'h389c8b4c),
	.w4(32'hb7cce9ec),
	.w5(32'hb7093eba),
	.w6(32'h3808493d),
	.w7(32'h360b76da),
	.w8(32'hb7976f01),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381a1191),
	.w1(32'hb7814d93),
	.w2(32'h37398a5f),
	.w3(32'h37d9fa7f),
	.w4(32'hb63f963b),
	.w5(32'h36d0bce6),
	.w6(32'h38603338),
	.w7(32'hb7e2acca),
	.w8(32'h36eccd2a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa083f7),
	.w1(32'h3a899b7a),
	.w2(32'h3a2ad3ee),
	.w3(32'h3a835e76),
	.w4(32'h3a2a4fd2),
	.w5(32'h39264dc5),
	.w6(32'h3a426a2a),
	.w7(32'h39875126),
	.w8(32'hb948c499),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391249b9),
	.w1(32'h3b142e69),
	.w2(32'h39d223f3),
	.w3(32'h3b039ec0),
	.w4(32'hb9a6ad2a),
	.w5(32'hb94d5641),
	.w6(32'h3b5a42da),
	.w7(32'hba9cd7f6),
	.w8(32'hbadb8a70),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a82db1),
	.w1(32'h3a2b7239),
	.w2(32'h3a4a3cc0),
	.w3(32'hb90bd0e6),
	.w4(32'h395638ac),
	.w5(32'h3907cea5),
	.w6(32'h37876446),
	.w7(32'h38c203f6),
	.w8(32'h3912273a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25ce7a),
	.w1(32'hbac23afc),
	.w2(32'hba3fadf2),
	.w3(32'hbac89930),
	.w4(32'hba3a4c32),
	.w5(32'hbb0573b2),
	.w6(32'h3a9a9eb4),
	.w7(32'h3a9c5dbf),
	.w8(32'h3a85ef56),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b4331),
	.w1(32'hbb717c61),
	.w2(32'hbab2be4c),
	.w3(32'hb9409b7c),
	.w4(32'h3a8d3236),
	.w5(32'hbb2597f0),
	.w6(32'h3ba229ce),
	.w7(32'h3c0e609e),
	.w8(32'h3bb7a726),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be09ed5),
	.w1(32'h3bb41011),
	.w2(32'h3b830df6),
	.w3(32'h3b82d352),
	.w4(32'h3b0e4e7c),
	.w5(32'h3b046fd3),
	.w6(32'h3b32931f),
	.w7(32'hba8175b8),
	.w8(32'hbad0a7a7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb38787),
	.w1(32'hbc4db95a),
	.w2(32'hbb6591c6),
	.w3(32'hbc40c421),
	.w4(32'hbb028013),
	.w5(32'h3bc1f9e4),
	.w6(32'hbb86dec7),
	.w7(32'h3be8c1b2),
	.w8(32'h3b8e4035),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb3d52),
	.w1(32'h3bebaafd),
	.w2(32'h3b505b2a),
	.w3(32'h3bdcb688),
	.w4(32'h3bb02361),
	.w5(32'hb9984334),
	.w6(32'h3bb5083d),
	.w7(32'h3afe841b),
	.w8(32'h3aed4117),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f17d6),
	.w1(32'hbc3d0954),
	.w2(32'hbc116699),
	.w3(32'h3ab2939d),
	.w4(32'hbba37074),
	.w5(32'hbbe0c1fc),
	.w6(32'h3be8bbae),
	.w7(32'h3bb525b1),
	.w8(32'hb9299bdd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4021a),
	.w1(32'h3946e895),
	.w2(32'h39d9a044),
	.w3(32'h3afe94d7),
	.w4(32'hb8304fd2),
	.w5(32'hbafcc3fe),
	.w6(32'h3bed5ae0),
	.w7(32'h3b67ac44),
	.w8(32'hba91e377),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02a93c),
	.w1(32'h3b5fa00d),
	.w2(32'h394668b2),
	.w3(32'h3b0992bc),
	.w4(32'hbb5a6596),
	.w5(32'hbb127478),
	.w6(32'h3b9826ae),
	.w7(32'hbab60fd1),
	.w8(32'hbb252c09),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bab3b),
	.w1(32'h3b316041),
	.w2(32'h3a8028e2),
	.w3(32'h3b07070a),
	.w4(32'h3af1ea22),
	.w5(32'h3989bc41),
	.w6(32'h3ad6daed),
	.w7(32'h3aac1bad),
	.w8(32'h37e7a2b0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96c4d6),
	.w1(32'hbbb683b8),
	.w2(32'hbb776296),
	.w3(32'hba861fbc),
	.w4(32'hb9c40893),
	.w5(32'hbb4bc7dd),
	.w6(32'h3b37a0ab),
	.w7(32'h3bd83aae),
	.w8(32'h3b0f6c34),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53c91b),
	.w1(32'hbbf0549b),
	.w2(32'h3a8bd749),
	.w3(32'hbb248a4e),
	.w4(32'h3a9c22f5),
	.w5(32'h3bcd13e5),
	.w6(32'h3b0c78e1),
	.w7(32'h3bae924d),
	.w8(32'h3bba1952),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56e16b),
	.w1(32'hba764cd2),
	.w2(32'hbc1b60e1),
	.w3(32'hbb7da792),
	.w4(32'h3b873db6),
	.w5(32'h3bcc2f9d),
	.w6(32'hbc65ecb9),
	.w7(32'hbad1b70d),
	.w8(32'h3c19f5b8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc081ae),
	.w1(32'h3b80ffc4),
	.w2(32'hbba624ba),
	.w3(32'h3a3b78ae),
	.w4(32'hbb401306),
	.w5(32'hbbafe3e3),
	.w6(32'hbb854feb),
	.w7(32'hbc1a2ae1),
	.w8(32'hbc259e8a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61aa7d),
	.w1(32'h3b02cc52),
	.w2(32'h3a82fea4),
	.w3(32'h3b4d938c),
	.w4(32'hba744bcb),
	.w5(32'hbadca629),
	.w6(32'h3b323a72),
	.w7(32'h398bf260),
	.w8(32'hba7ffc92),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a7378),
	.w1(32'hbbb5b3d6),
	.w2(32'hba847f7e),
	.w3(32'hbb835b6f),
	.w4(32'h3c1325cc),
	.w5(32'h3bf750aa),
	.w6(32'h39d40924),
	.w7(32'h3bfe62ec),
	.w8(32'h3c21d147),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b426280),
	.w1(32'h3b73319a),
	.w2(32'h3b416a49),
	.w3(32'h3a8f476a),
	.w4(32'h3bab45ee),
	.w5(32'h3b5f9752),
	.w6(32'h3aae6cc0),
	.w7(32'h3b895c73),
	.w8(32'h3b5e28a8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce5d793),
	.w1(32'hbc1d03a5),
	.w2(32'hbc644e71),
	.w3(32'hbc3232b9),
	.w4(32'h3b642ad6),
	.w5(32'h3bcfd268),
	.w6(32'hba3db945),
	.w7(32'h3bd072ce),
	.w8(32'h3bfaede3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf49d9),
	.w1(32'h3b7a5ca2),
	.w2(32'h399439d3),
	.w3(32'hbb6b2f30),
	.w4(32'h3b400af0),
	.w5(32'h3b2bf4aa),
	.w6(32'hbb9472c2),
	.w7(32'h3a7d45d9),
	.w8(32'h3bb1a5f2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d8f0c),
	.w1(32'h39b80019),
	.w2(32'h392ce15c),
	.w3(32'h3a7f00d3),
	.w4(32'h39863c71),
	.w5(32'h37f497ab),
	.w6(32'h3a5a59d4),
	.w7(32'h38bc2589),
	.w8(32'hb91b9d16),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea3bb4),
	.w1(32'hba11396a),
	.w2(32'hbac436e5),
	.w3(32'h3ada7c63),
	.w4(32'hbaa910cb),
	.w5(32'hb9b48071),
	.w6(32'hb986465c),
	.w7(32'hba45c920),
	.w8(32'hbace862b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba101e86),
	.w1(32'h399c92f3),
	.w2(32'h3a8b0d06),
	.w3(32'h39085c9e),
	.w4(32'hb8296a19),
	.w5(32'hbaf15e22),
	.w6(32'h3b4c40d6),
	.w7(32'h3baa384a),
	.w8(32'h3b300cfc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fc305),
	.w1(32'h3af02675),
	.w2(32'hba3c288a),
	.w3(32'h3b236cba),
	.w4(32'hba41fbd1),
	.w5(32'hbb056046),
	.w6(32'h3b63c38f),
	.w7(32'hb88bcc59),
	.w8(32'hba5495e6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14881b),
	.w1(32'hbab32ac2),
	.w2(32'h395101f7),
	.w3(32'h3b198589),
	.w4(32'hbaa6301a),
	.w5(32'h3b2f5859),
	.w6(32'h39ee09cd),
	.w7(32'hbb49c789),
	.w8(32'hbac31226),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a8b40),
	.w1(32'hb9643219),
	.w2(32'h3a2f027f),
	.w3(32'h3a6a8bab),
	.w4(32'hb98b83f7),
	.w5(32'h3a78cfca),
	.w6(32'h3a41262f),
	.w7(32'hba3ed54d),
	.w8(32'hbac8c7f0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d4866),
	.w1(32'h3a694880),
	.w2(32'h3b8c3690),
	.w3(32'hbbc05c0c),
	.w4(32'hb942a2a9),
	.w5(32'h3b30347e),
	.w6(32'h3ab6beb2),
	.w7(32'h3b821030),
	.w8(32'h3c164f01),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81d6f0),
	.w1(32'hbbc84c3c),
	.w2(32'hbb97e77e),
	.w3(32'hbb20276a),
	.w4(32'hbc0442c5),
	.w5(32'hbc07b18a),
	.w6(32'h3aaf5964),
	.w7(32'hbb7eded5),
	.w8(32'hbbf8a91a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc8d2d),
	.w1(32'h3904a67c),
	.w2(32'h3a2bc53e),
	.w3(32'h38cd35e3),
	.w4(32'hb9aa475e),
	.w5(32'hb993b8f2),
	.w6(32'h3b055a12),
	.w7(32'h3ac49a66),
	.w8(32'h3aca150a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c049a4),
	.w1(32'hb980fd10),
	.w2(32'hb95d1c89),
	.w3(32'hb9c43eec),
	.w4(32'hb9e5aed0),
	.w5(32'hb95776f6),
	.w6(32'hb99f9542),
	.w7(32'hb991894e),
	.w8(32'hb93719af),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993521a),
	.w1(32'hba5a3276),
	.w2(32'hb948fe5a),
	.w3(32'hb791a5b2),
	.w4(32'hb94de8b9),
	.w5(32'hb9b7cbd4),
	.w6(32'h3a32eb2a),
	.w7(32'hb943d30e),
	.w8(32'hba3e7c0e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38037c62),
	.w1(32'h370f8257),
	.w2(32'h378bae5d),
	.w3(32'h382726e3),
	.w4(32'h37f7eb81),
	.w5(32'h3701fb7f),
	.w6(32'h37575853),
	.w7(32'hb7240df9),
	.w8(32'hb6a2ff23),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5f251),
	.w1(32'h3a318984),
	.w2(32'h3a645a16),
	.w3(32'h3a072d3c),
	.w4(32'h3a29efac),
	.w5(32'h3a2135e5),
	.w6(32'h3a161b7a),
	.w7(32'h398c98da),
	.w8(32'h39d52535),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d5dae),
	.w1(32'hb7655642),
	.w2(32'h3adaffe1),
	.w3(32'h38b20396),
	.w4(32'h3aba0701),
	.w5(32'h3b186c4b),
	.w6(32'h3b5d6f6f),
	.w7(32'h3b890387),
	.w8(32'h3b8ced66),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c3f0b),
	.w1(32'h39b3c5b5),
	.w2(32'h39d57a9d),
	.w3(32'h38c112e5),
	.w4(32'h3970e0f3),
	.w5(32'h39ee9d6c),
	.w6(32'h399d6b40),
	.w7(32'h39b5c5b5),
	.w8(32'h39152cba),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8043bc),
	.w1(32'hbb343e25),
	.w2(32'h392a86bd),
	.w3(32'hbb4c6ad6),
	.w4(32'h3a68e62a),
	.w5(32'h3b0ce7d2),
	.w6(32'hb97fb7a9),
	.w7(32'h3b3f38be),
	.w8(32'h3b984679),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b0b7),
	.w1(32'h3b4032fd),
	.w2(32'h3ace4317),
	.w3(32'h3bd2e88f),
	.w4(32'hbb1233f5),
	.w5(32'hbb057f73),
	.w6(32'h3ba7d134),
	.w7(32'hbb764190),
	.w8(32'hbbbfdf0c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39071838),
	.w1(32'h3789a73c),
	.w2(32'hb880b774),
	.w3(32'h38ba2ed9),
	.w4(32'h37bfe8f5),
	.w5(32'hb9111d80),
	.w6(32'h38fea50c),
	.w7(32'h3888442c),
	.w8(32'hb87eb760),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d7330),
	.w1(32'h399a6e4a),
	.w2(32'h3942db66),
	.w3(32'h397f57b0),
	.w4(32'h3954fa0a),
	.w5(32'h38ac7a96),
	.w6(32'h38c525de),
	.w7(32'h38ae2e7a),
	.w8(32'hb7bf19a9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782a4c0),
	.w1(32'hb745427a),
	.w2(32'h38bfb90e),
	.w3(32'h38a39d6e),
	.w4(32'h38108982),
	.w5(32'h381434cf),
	.w6(32'h385d9f4a),
	.w7(32'hb6404ea4),
	.w8(32'h382c58d8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d16716),
	.w1(32'h398f95ed),
	.w2(32'h3889ac81),
	.w3(32'h39f979f5),
	.w4(32'h39be132e),
	.w5(32'hb8f6862b),
	.w6(32'h39ca20b6),
	.w7(32'h39868019),
	.w8(32'h37c8885b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30a51e),
	.w1(32'hba3986e6),
	.w2(32'hba599381),
	.w3(32'h3ac5fb19),
	.w4(32'hbacdb322),
	.w5(32'hbba7f9f4),
	.w6(32'h3ab53600),
	.w7(32'h3b9fe207),
	.w8(32'h3c030c7f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb51b6c),
	.w1(32'hbbce50e5),
	.w2(32'hbabd46fb),
	.w3(32'hbb279942),
	.w4(32'hbb5da797),
	.w5(32'hbb0e2090),
	.w6(32'h3ae0ab58),
	.w7(32'h3b9be0da),
	.w8(32'h3b350ae6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad69a83),
	.w1(32'hba1126c6),
	.w2(32'h382c64b6),
	.w3(32'hba278f3b),
	.w4(32'h39ec8f4c),
	.w5(32'h39eaaee1),
	.w6(32'h3a5a7401),
	.w7(32'h3ab4b8dc),
	.w8(32'h3a63125b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecaef5),
	.w1(32'hbb845b46),
	.w2(32'hbb4f3a08),
	.w3(32'hb8bf06fc),
	.w4(32'hba61bfac),
	.w5(32'hbadfe295),
	.w6(32'hba2a8ab6),
	.w7(32'h3ae2def5),
	.w8(32'h3aeacf1c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b5973),
	.w1(32'hb8ed5fb5),
	.w2(32'h39af34b6),
	.w3(32'h3a3bc111),
	.w4(32'hb8be9d24),
	.w5(32'h3a4c3dc7),
	.w6(32'h3ac60a2c),
	.w7(32'h39b8476d),
	.w8(32'h3a0fd44d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919b17e),
	.w1(32'hbb67bfd2),
	.w2(32'hbb1743fd),
	.w3(32'h3ada68ac),
	.w4(32'hbb0ded29),
	.w5(32'hbb510aa0),
	.w6(32'h3b5a5314),
	.w7(32'h3af84e66),
	.w8(32'h399804a2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af45af9),
	.w1(32'hbb497b8e),
	.w2(32'hb9f19885),
	.w3(32'h3b98a063),
	.w4(32'hbb7294ce),
	.w5(32'hbaad0047),
	.w6(32'h3be5fe44),
	.w7(32'hba8f92f2),
	.w8(32'hbada70bc),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c069c),
	.w1(32'hbc032eb8),
	.w2(32'hbae39076),
	.w3(32'hbb3e6329),
	.w4(32'h390de295),
	.w5(32'h3aaf35df),
	.w6(32'h3ac095bc),
	.w7(32'h3be96b3f),
	.w8(32'h3bbabad6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40deed),
	.w1(32'h3acf9740),
	.w2(32'h399dd90c),
	.w3(32'h3a6ee23d),
	.w4(32'hbafd9d18),
	.w5(32'hbafbc05b),
	.w6(32'h3ac502cf),
	.w7(32'hbaed6c71),
	.w8(32'hbb66829a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0b49b),
	.w1(32'hbb9d0f77),
	.w2(32'hbb06a13b),
	.w3(32'hbb50e4e9),
	.w4(32'hbace0397),
	.w5(32'h390217d6),
	.w6(32'hba51012e),
	.w7(32'h3ae5db81),
	.w8(32'h3b085c87),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc66990),
	.w1(32'hbb8cd02d),
	.w2(32'hba9229a4),
	.w3(32'hbb8b618e),
	.w4(32'h3b91b683),
	.w5(32'h3b69b7ee),
	.w6(32'h3b65029f),
	.w7(32'h3bf983b4),
	.w8(32'h3be8185e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46c6f3),
	.w1(32'hba594a2e),
	.w2(32'hbb04f391),
	.w3(32'h36991108),
	.w4(32'hb9df8905),
	.w5(32'h3a40c14b),
	.w6(32'h3a679b87),
	.w7(32'h39b963c0),
	.w8(32'h3b01b193),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac2fa6),
	.w1(32'hbbdce06a),
	.w2(32'hbaf70015),
	.w3(32'hbb316d11),
	.w4(32'hbb242028),
	.w5(32'hbaee11ee),
	.w6(32'h3b265d83),
	.w7(32'h3b7f3b51),
	.w8(32'hb926b352),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c941f),
	.w1(32'hb7090ba7),
	.w2(32'h389ab0fd),
	.w3(32'hb8943cb4),
	.w4(32'hb71bbae6),
	.w5(32'h37e93168),
	.w6(32'h3a53e079),
	.w7(32'h3a56e6fc),
	.w8(32'h3a16fe94),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c524ee1),
	.w1(32'h3b3deea4),
	.w2(32'h3b402a63),
	.w3(32'h3bd8a422),
	.w4(32'hbb96bf00),
	.w5(32'hbb130934),
	.w6(32'h3ba436dc),
	.w7(32'hbbb0395a),
	.w8(32'hbbb02a60),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad45a7e),
	.w1(32'hba56e34d),
	.w2(32'hba166e1b),
	.w3(32'hba426c19),
	.w4(32'hba5880c7),
	.w5(32'hb6ce2b7f),
	.w6(32'h3a2ae3d8),
	.w7(32'h3acb40bc),
	.w8(32'h3adfeb0d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78795e8),
	.w1(32'hb82f3673),
	.w2(32'h38568082),
	.w3(32'hb8b9de7e),
	.w4(32'hb8af05aa),
	.w5(32'hb894b59a),
	.w6(32'h387877d6),
	.w7(32'h3865193f),
	.w8(32'h394c8a96),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d201ce),
	.w1(32'hb8c445c4),
	.w2(32'h388f9f92),
	.w3(32'hb893ddac),
	.w4(32'hb824df0b),
	.w5(32'hb7a31b03),
	.w6(32'hb75d34c1),
	.w7(32'hb85a4583),
	.w8(32'h392f3bf2),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e992e),
	.w1(32'hba519000),
	.w2(32'hb9ae44a0),
	.w3(32'hbb1a9d75),
	.w4(32'hba600327),
	.w5(32'hba29c783),
	.w6(32'h39a4ea53),
	.w7(32'h3a1b4d96),
	.w8(32'h3ad396c9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2a3cd),
	.w1(32'h3a4cc0f2),
	.w2(32'hbb13d215),
	.w3(32'hbadfc38e),
	.w4(32'hba51e25a),
	.w5(32'hba27bef1),
	.w6(32'h3981f756),
	.w7(32'hbaa30bec),
	.w8(32'hba11ee86),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa42801),
	.w1(32'hba4ae1ed),
	.w2(32'h3a3e7792),
	.w3(32'hb9ccd3ad),
	.w4(32'hba0e8893),
	.w5(32'hba40abaf),
	.w6(32'h3b86d565),
	.w7(32'h3b725d91),
	.w8(32'h3b79b42f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382bec22),
	.w1(32'hb8eee5e0),
	.w2(32'hb922b96e),
	.w3(32'h388969ec),
	.w4(32'hb80512bc),
	.w5(32'hb955e58c),
	.w6(32'h38b5d8a9),
	.w7(32'hb897dcdf),
	.w8(32'hb95b5d0a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b64d2),
	.w1(32'hbba4812c),
	.w2(32'hba91d280),
	.w3(32'hbb19b7de),
	.w4(32'hbb4918b8),
	.w5(32'hbb4807fa),
	.w6(32'h3b5504e2),
	.w7(32'h3b4c059a),
	.w8(32'hb8316c88),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81841d),
	.w1(32'hbac916b2),
	.w2(32'hbaba988d),
	.w3(32'h394619d8),
	.w4(32'hbb162c2a),
	.w5(32'hbb5f4f71),
	.w6(32'h3ad1bb7f),
	.w7(32'hb98f27bf),
	.w8(32'hbb253a80),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf53d3c),
	.w1(32'hbc067b89),
	.w2(32'hbbd8960c),
	.w3(32'hbad7cab2),
	.w4(32'h389a4a97),
	.w5(32'h3b65d040),
	.w6(32'h3aaeba51),
	.w7(32'h3bec12fb),
	.w8(32'h3be8762b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98def0),
	.w1(32'hbb215242),
	.w2(32'h3bda588e),
	.w3(32'h3bb91d79),
	.w4(32'hbb8fb623),
	.w5(32'h3b862478),
	.w6(32'h3bc199b1),
	.w7(32'hbb38dcfb),
	.w8(32'hbaf6f697),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43c410),
	.w1(32'h3af2d269),
	.w2(32'h3a2a6734),
	.w3(32'h3ac6913c),
	.w4(32'h398bbe68),
	.w5(32'hba23879c),
	.w6(32'h3abc6d62),
	.w7(32'hba677723),
	.w8(32'hbb22977a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b989d),
	.w1(32'h3b2a836f),
	.w2(32'h3ae768c1),
	.w3(32'h3b8f1113),
	.w4(32'h3b3f3fae),
	.w5(32'h3b61249a),
	.w6(32'h3b887c20),
	.w7(32'h3b4c7d34),
	.w8(32'h3b16d3ad),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109cdc),
	.w1(32'hbaea96c9),
	.w2(32'h3a88bb7d),
	.w3(32'hbb1836f9),
	.w4(32'hba8d2d38),
	.w5(32'h3a30e2dd),
	.w6(32'hb9147baf),
	.w7(32'h3aa07eae),
	.w8(32'h3b245f1d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba864d43),
	.w1(32'hba89001b),
	.w2(32'hba8379af),
	.w3(32'h3afb881d),
	.w4(32'hb9eb599d),
	.w5(32'h39fe9ba7),
	.w6(32'h3b2a6c37),
	.w7(32'hbac9d00b),
	.w8(32'hbad839db),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb11d6f),
	.w1(32'h3b7179d8),
	.w2(32'h3b253877),
	.w3(32'h3b630e1d),
	.w4(32'h3a925346),
	.w5(32'h3a8022c1),
	.w6(32'h3b526c54),
	.w7(32'h37d583d6),
	.w8(32'hba6d376f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaede62f),
	.w1(32'hbaabefa5),
	.w2(32'h39349ac3),
	.w3(32'hba404061),
	.w4(32'h3a284d5d),
	.w5(32'h3a8c9ca6),
	.w6(32'h39eddba5),
	.w7(32'h3b11dc7f),
	.w8(32'h3affea36),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ba29c),
	.w1(32'h395e5ca2),
	.w2(32'hb8e9c703),
	.w3(32'h39e8abb1),
	.w4(32'h39fda060),
	.w5(32'h39c20fb4),
	.w6(32'h39a44e85),
	.w7(32'h39ccaefd),
	.w8(32'h38f3b095),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa5561),
	.w1(32'hbbd1c549),
	.w2(32'hbb143522),
	.w3(32'hbb9514a5),
	.w4(32'hbafe8716),
	.w5(32'hb9ce3312),
	.w6(32'h3aaf3943),
	.w7(32'h3b6dc60e),
	.w8(32'h3b4fbe7c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba891fb1),
	.w1(32'h39a0ddb9),
	.w2(32'h39c6bca3),
	.w3(32'hb84ddb32),
	.w4(32'h3a869c09),
	.w5(32'h3a8b4d5d),
	.w6(32'h394c7cab),
	.w7(32'h39f41c8a),
	.w8(32'h3ac34adc),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c0e6b),
	.w1(32'hba97597d),
	.w2(32'h3b0d7712),
	.w3(32'h39c68ec8),
	.w4(32'hbab87391),
	.w5(32'hb7680c8a),
	.w6(32'h3b0c283c),
	.w7(32'h3aa030df),
	.w8(32'h3ac9709b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee8915),
	.w1(32'h399b2238),
	.w2(32'hb89a54f0),
	.w3(32'h372c43fb),
	.w4(32'h3951698f),
	.w5(32'h377ed38d),
	.w6(32'hb99fb607),
	.w7(32'h39122d24),
	.w8(32'h395c6c04),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be07762),
	.w1(32'h3b75d9aa),
	.w2(32'h3b2587a0),
	.w3(32'h3ba014aa),
	.w4(32'h3a42e08a),
	.w5(32'hba53be04),
	.w6(32'h3ba2954a),
	.w7(32'h3b1e2368),
	.w8(32'h381a31d4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39528751),
	.w1(32'h3992e5f5),
	.w2(32'h39b0d08f),
	.w3(32'h398fe92d),
	.w4(32'h39676c27),
	.w5(32'h39c2beea),
	.w6(32'h395096fb),
	.w7(32'h399ab615),
	.w8(32'h39a6f329),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928f356),
	.w1(32'hb9d3454f),
	.w2(32'hb9dd4a69),
	.w3(32'h398d91e0),
	.w4(32'hb9850511),
	.w5(32'hb9a69625),
	.w6(32'h39c826df),
	.w7(32'hb9bd3dcf),
	.w8(32'hb938ec52),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3eafb),
	.w1(32'hb9dd0fff),
	.w2(32'hb834cbbd),
	.w3(32'hb84922da),
	.w4(32'hbaccead6),
	.w5(32'h39a5b9dc),
	.w6(32'h39d72b00),
	.w7(32'h3a083035),
	.w8(32'h3a71f423),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb55f1),
	.w1(32'hbb1cb8d8),
	.w2(32'h3883d8cc),
	.w3(32'hbbdaac4b),
	.w4(32'hb9ba654d),
	.w5(32'hb95eafe5),
	.w6(32'hbb9af715),
	.w7(32'h3b83e45d),
	.w8(32'h3bf1c054),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b138dd2),
	.w1(32'h3b0e5863),
	.w2(32'h3ac00a7d),
	.w3(32'h3b0c60e1),
	.w4(32'h3acd38a1),
	.w5(32'h3a8505fd),
	.w6(32'h3aefe99b),
	.w7(32'h3aba32f4),
	.w8(32'h3a9c2808),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86384c),
	.w1(32'h3affeecd),
	.w2(32'h3a411015),
	.w3(32'h3abcd16f),
	.w4(32'hbab21e5b),
	.w5(32'hbb21c0c8),
	.w6(32'h3b77de53),
	.w7(32'h39e7f21d),
	.w8(32'hba921bf4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2290c),
	.w1(32'hbaa309a4),
	.w2(32'h3b14172d),
	.w3(32'h3afbf21d),
	.w4(32'hbb287ba6),
	.w5(32'hba320c16),
	.w6(32'h3ab56033),
	.w7(32'hbaca2c63),
	.w8(32'hbaa19312),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71e44),
	.w1(32'hbb9dd295),
	.w2(32'hbaa1b5f3),
	.w3(32'h3ae7c720),
	.w4(32'hba6e06b8),
	.w5(32'hb7751bcb),
	.w6(32'h3b8b58af),
	.w7(32'h3b38dd3c),
	.w8(32'h3b182aa5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba886ed4),
	.w1(32'hbb4fd293),
	.w2(32'hbb821b6a),
	.w3(32'h395929ed),
	.w4(32'hb9f48afc),
	.w5(32'hbad8beeb),
	.w6(32'h3b76fd13),
	.w7(32'h3b2f542b),
	.w8(32'h3b0d4be6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed4031),
	.w1(32'hbb95bd2c),
	.w2(32'hba6932af),
	.w3(32'hbb15ed9e),
	.w4(32'h39fcea8b),
	.w5(32'hba151b47),
	.w6(32'h3b2caf9b),
	.w7(32'h3bfa39c2),
	.w8(32'h3b61eab6),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2e18c),
	.w1(32'h3a77e776),
	.w2(32'h3a59e873),
	.w3(32'h3a2d92e8),
	.w4(32'h3ab6dea8),
	.w5(32'h3ab1aa1f),
	.w6(32'h39e6958e),
	.w7(32'h3ac632c0),
	.w8(32'h3af6a66a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00a825),
	.w1(32'hbb6e6dd1),
	.w2(32'hba549ad0),
	.w3(32'h3a45504f),
	.w4(32'hbb1f30a1),
	.w5(32'hbada9dd4),
	.w6(32'h3b62fdcf),
	.w7(32'h3acf4bea),
	.w8(32'hbaa71175),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65794ca),
	.w1(32'h37f77089),
	.w2(32'h37ece763),
	.w3(32'h38178689),
	.w4(32'h383219ca),
	.w5(32'h37e2fb12),
	.w6(32'h3791696a),
	.w7(32'hb6465562),
	.w8(32'hb7037466),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f3091),
	.w1(32'hba162ac5),
	.w2(32'h39e0e2d2),
	.w3(32'hb8b1712b),
	.w4(32'h3a0fe497),
	.w5(32'h3a9820a2),
	.w6(32'h39f1ab92),
	.w7(32'h3a893082),
	.w8(32'h3a8ef3bb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9698d9),
	.w1(32'hb913df6e),
	.w2(32'h39e653ee),
	.w3(32'h3a2a25db),
	.w4(32'hb9daa81f),
	.w5(32'h39467b69),
	.w6(32'h3946af82),
	.w7(32'hb9790fa2),
	.w8(32'hb9834296),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fdb19),
	.w1(32'hbb4bd560),
	.w2(32'hbb0d05ac),
	.w3(32'h39372d17),
	.w4(32'hbba759cf),
	.w5(32'hbb922cb7),
	.w6(32'h3b838d9e),
	.w7(32'h3986c1c9),
	.w8(32'hbb2af2b6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb606f6a0),
	.w1(32'h380ee211),
	.w2(32'h37ef212e),
	.w3(32'hb79fc7c3),
	.w4(32'hb856ef2b),
	.w5(32'hb7a02279),
	.w6(32'hb746a9b8),
	.w7(32'hb830b4b7),
	.w8(32'h364c6b15),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c84e43),
	.w1(32'hb99b627d),
	.w2(32'hb99daef6),
	.w3(32'hb9a9ca3e),
	.w4(32'hb955a901),
	.w5(32'hb95145f3),
	.w6(32'hb9031676),
	.w7(32'hb9013419),
	.w8(32'hb92ac857),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c6a3c),
	.w1(32'h39b015d5),
	.w2(32'h3b2f585c),
	.w3(32'h3b0fad10),
	.w4(32'h3a9a8e0a),
	.w5(32'h3b06bfa3),
	.w6(32'h3b12eb34),
	.w7(32'h3a924eaf),
	.w8(32'h3aa9ea23),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ef929),
	.w1(32'h38a8128c),
	.w2(32'h398cc8d8),
	.w3(32'h3b876fcf),
	.w4(32'h3b86d7e1),
	.w5(32'h3b6b2945),
	.w6(32'h3b2c04f7),
	.w7(32'h3b464aa5),
	.w8(32'h3b8c7e40),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8817ca),
	.w1(32'h3b25fb7a),
	.w2(32'hb88de4c2),
	.w3(32'hbb74786b),
	.w4(32'h3b8230fe),
	.w5(32'h3b1ac3d2),
	.w6(32'h391ff937),
	.w7(32'h3b210bbc),
	.w8(32'h3b629542),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b0413),
	.w1(32'hb91892c9),
	.w2(32'hb9aecc23),
	.w3(32'h3a0c8db3),
	.w4(32'hb9557d63),
	.w5(32'hb98d222c),
	.w6(32'h3a55461f),
	.w7(32'hb9272b39),
	.w8(32'h3860c185),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62684e),
	.w1(32'hbc004b81),
	.w2(32'hbb638301),
	.w3(32'hbb6120db),
	.w4(32'hb97494e5),
	.w5(32'hbb575e8b),
	.w6(32'h3b619a62),
	.w7(32'h3c2c2ecd),
	.w8(32'h3bc1a356),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d3991),
	.w1(32'hbc010edf),
	.w2(32'h3ab7bcf1),
	.w3(32'h3abf2feb),
	.w4(32'hbbe0ac8f),
	.w5(32'h3a9beb75),
	.w6(32'h3c1160a6),
	.w7(32'hba03d885),
	.w8(32'hbbd91a1e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8373c1),
	.w1(32'h37828d4a),
	.w2(32'h3aea7826),
	.w3(32'hba8abf3c),
	.w4(32'h3b055516),
	.w5(32'h3af455db),
	.w6(32'h3aa8ffd7),
	.w7(32'h3b311710),
	.w8(32'h3b00b0a0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a7dac5),
	.w1(32'hb8821341),
	.w2(32'hb8189c1c),
	.w3(32'hb8452c38),
	.w4(32'hb89166d2),
	.w5(32'hb8a0f07e),
	.w6(32'hb885b975),
	.w7(32'hb8b14e37),
	.w8(32'hb8ebd059),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba048761),
	.w1(32'hba044a4e),
	.w2(32'hba076644),
	.w3(32'hba204422),
	.w4(32'hb99af4d2),
	.w5(32'hba134cfb),
	.w6(32'hba2c7bcd),
	.w7(32'hb881f9ef),
	.w8(32'hb9e5ef00),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387e34fd),
	.w1(32'h37e402e7),
	.w2(32'h370203e8),
	.w3(32'h382dcd60),
	.w4(32'hb75ae025),
	.w5(32'hb5d2c85b),
	.w6(32'hb7ee13b3),
	.w7(32'hb80f69dc),
	.w8(32'hb78f2e2d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34440080),
	.w1(32'h3b36631b),
	.w2(32'h3b2bb8a8),
	.w3(32'hba8f58c7),
	.w4(32'h3af293d6),
	.w5(32'h3b20921d),
	.w6(32'hba0f189a),
	.w7(32'h3b22ed22),
	.w8(32'h3b195f33),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeca045),
	.w1(32'hbabde119),
	.w2(32'hb9e41510),
	.w3(32'hba9ca55d),
	.w4(32'h39aaad24),
	.w5(32'h3a96dfb6),
	.w6(32'h3ac8ba6e),
	.w7(32'h3adc3b89),
	.w8(32'h3afb600a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f57bc),
	.w1(32'h3ae67e43),
	.w2(32'h39490fc4),
	.w3(32'h3aec7394),
	.w4(32'hbad6f05f),
	.w5(32'hb9c58557),
	.w6(32'h3b7acf63),
	.w7(32'hb9ddc029),
	.w8(32'hbaacf6e8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923bd43),
	.w1(32'hb8957922),
	.w2(32'h3a1eebc0),
	.w3(32'h3a57cea9),
	.w4(32'hb93ec934),
	.w5(32'h3a3b0407),
	.w6(32'h3a54e5e8),
	.w7(32'hb829e9a0),
	.w8(32'h3a79ccf0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868fd5),
	.w1(32'hbab60e4d),
	.w2(32'hbbf5823e),
	.w3(32'hbb40714f),
	.w4(32'hbb4ac6b1),
	.w5(32'hbbd1e5b4),
	.w6(32'h3b384dbc),
	.w7(32'h3b3dd596),
	.w8(32'hbaa41137),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b4a57),
	.w1(32'hbbf08e78),
	.w2(32'hbbd890c8),
	.w3(32'hbc13054d),
	.w4(32'hbb8185e3),
	.w5(32'hbbeabbf1),
	.w6(32'hbbaa0dcc),
	.w7(32'h39d02563),
	.w8(32'h3b9fb521),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf07ecb),
	.w1(32'hbc0c2175),
	.w2(32'hbc1d582b),
	.w3(32'h3a9c4966),
	.w4(32'hbc1ae63b),
	.w5(32'hbc213f14),
	.w6(32'hba815a8d),
	.w7(32'hba900d09),
	.w8(32'hbbca0d20),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac45323),
	.w1(32'h3b87f93a),
	.w2(32'h3ad3424f),
	.w3(32'hbb184a83),
	.w4(32'h3b657d81),
	.w5(32'h3ad726bd),
	.w6(32'h3aac33b5),
	.w7(32'h3b02697c),
	.w8(32'h391b4aff),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28927d),
	.w1(32'h3a715687),
	.w2(32'h3b0d96a3),
	.w3(32'h3b6bfc5e),
	.w4(32'h3b805427),
	.w5(32'hbb424207),
	.w6(32'h3ac004a8),
	.w7(32'h3900d83e),
	.w8(32'hbaebf2be),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcba155),
	.w1(32'hbbcae1bd),
	.w2(32'hb9f7bc3c),
	.w3(32'h3b370fd1),
	.w4(32'hbbe52a0d),
	.w5(32'hbbe062eb),
	.w6(32'h3af53752),
	.w7(32'h3a329a28),
	.w8(32'hb9adbfa4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9be51),
	.w1(32'hbb34e792),
	.w2(32'hbb09cf7a),
	.w3(32'hbbc7e3b4),
	.w4(32'h3b9d5300),
	.w5(32'h3a9a6f16),
	.w6(32'hbb16fbb4),
	.w7(32'h3b928929),
	.w8(32'h3c19e0bd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbf016),
	.w1(32'h3b3e0acc),
	.w2(32'hbb785654),
	.w3(32'hb98bb517),
	.w4(32'h3a19c9b2),
	.w5(32'hba446db5),
	.w6(32'h3bdb2514),
	.w7(32'h3b6b67a9),
	.w8(32'h39264cbf),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11f1d2),
	.w1(32'h3c1d4f01),
	.w2(32'h3a5a3fc2),
	.w3(32'hbb04bc0e),
	.w4(32'h3c1b6de3),
	.w5(32'h3c00e302),
	.w6(32'hbae2bcc1),
	.w7(32'hbb25f067),
	.w8(32'h3bcdde79),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4e804),
	.w1(32'hbaaca575),
	.w2(32'hbb886a39),
	.w3(32'h3b167503),
	.w4(32'h3b6f4350),
	.w5(32'h3b71f9ae),
	.w6(32'h3a16ec44),
	.w7(32'h3bba28cc),
	.w8(32'h3bb46114),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb687a21),
	.w1(32'hbbc11316),
	.w2(32'hbbbafdb5),
	.w3(32'hbb90a9cd),
	.w4(32'hbbe7ec9f),
	.w5(32'hbb03c0b4),
	.w6(32'hbb5f59ae),
	.w7(32'hbaeaf0ad),
	.w8(32'h3992418f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbba3a1),
	.w1(32'h3b050d40),
	.w2(32'h394c4e9c),
	.w3(32'hbb961b47),
	.w4(32'h3b0fbddf),
	.w5(32'h3b2a4334),
	.w6(32'h3a85e378),
	.w7(32'h3aa3eda8),
	.w8(32'h3b581fa7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ec422),
	.w1(32'h3a96207f),
	.w2(32'hb93b8f82),
	.w3(32'hbb4c92ae),
	.w4(32'hbb11226e),
	.w5(32'hba1aabb9),
	.w6(32'hbb480508),
	.w7(32'h379d0f26),
	.w8(32'hba5be75a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb599bac),
	.w1(32'h39f690eb),
	.w2(32'h3b0278b2),
	.w3(32'hba76c645),
	.w4(32'hbab2253e),
	.w5(32'h3bd3039d),
	.w6(32'hbaa48d23),
	.w7(32'h3b706880),
	.w8(32'h3bd52e55),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a95e3),
	.w1(32'hbc0e68d9),
	.w2(32'hbbd55531),
	.w3(32'hbabd39a3),
	.w4(32'h3b4d565a),
	.w5(32'hbbe45580),
	.w6(32'h3b8bd43b),
	.w7(32'h3c176b00),
	.w8(32'h3c1addcf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22dd37),
	.w1(32'hbbbbcb37),
	.w2(32'h3be110c6),
	.w3(32'hbb9534e3),
	.w4(32'hba246c1e),
	.w5(32'h3af8f1f4),
	.w6(32'hbb0b99a5),
	.w7(32'h3bead3cc),
	.w8(32'h3b9c3814),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b623228),
	.w1(32'hbbb72c30),
	.w2(32'hbaa822c1),
	.w3(32'h3b98f3aa),
	.w4(32'hbae0386e),
	.w5(32'hbb23c443),
	.w6(32'h3c1cad62),
	.w7(32'h3b4dbde1),
	.w8(32'hbb1cc147),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc541bbf),
	.w1(32'hbbdf6602),
	.w2(32'hbb15b124),
	.w3(32'hbbd322a8),
	.w4(32'h3b891863),
	.w5(32'h3bac1b13),
	.w6(32'h3b446837),
	.w7(32'h3b68fb2a),
	.w8(32'h3b250e85),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0382f),
	.w1(32'h3aa4c6fa),
	.w2(32'hbb8a61e4),
	.w3(32'h3ae1b8ea),
	.w4(32'h3b8e7253),
	.w5(32'hbc0254e7),
	.w6(32'hbbae15f2),
	.w7(32'h3a3ce5e0),
	.w8(32'h3b071752),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a070359),
	.w1(32'hbb8fb2f4),
	.w2(32'hbc041585),
	.w3(32'hb95b5ea8),
	.w4(32'hbb4d3012),
	.w5(32'hbc14c859),
	.w6(32'hbba6ea1e),
	.w7(32'h3aaa07ec),
	.w8(32'hbb7e37ad),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1da59b),
	.w1(32'h3bfdbdb5),
	.w2(32'hbb702181),
	.w3(32'hbc815765),
	.w4(32'h3c29b58e),
	.w5(32'h3c234c97),
	.w6(32'hbc4b3f28),
	.w7(32'h3bc3a81a),
	.w8(32'h3c26bef6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eefce),
	.w1(32'hbb6f19e5),
	.w2(32'hbb83efba),
	.w3(32'hbb50900b),
	.w4(32'h3b510bf2),
	.w5(32'hbb6f2865),
	.w6(32'hba5e3308),
	.w7(32'h3bd5a656),
	.w8(32'h3b9f7ce5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fab7e),
	.w1(32'hbb855b98),
	.w2(32'hbab190de),
	.w3(32'hbc110acd),
	.w4(32'h3b8dadbe),
	.w5(32'h3b3b71fc),
	.w6(32'hba88a1f3),
	.w7(32'h3c6cf23c),
	.w8(32'h3c02d400),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842c25),
	.w1(32'hba98289a),
	.w2(32'h3b6062c0),
	.w3(32'h3b67e756),
	.w4(32'h3965e238),
	.w5(32'h3bfc3ace),
	.w6(32'h3b90513a),
	.w7(32'h3af6cf3e),
	.w8(32'hbb29c926),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fa1bb),
	.w1(32'h3b911cf9),
	.w2(32'h38de6e86),
	.w3(32'h3c1321a1),
	.w4(32'h3bbda485),
	.w5(32'h3abadab9),
	.w6(32'h3c443031),
	.w7(32'h3ad6d581),
	.w8(32'hba344a4e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb4375),
	.w1(32'hba290929),
	.w2(32'h3bc2dff9),
	.w3(32'h39c1d203),
	.w4(32'hbb92fb4d),
	.w5(32'hbbc4c804),
	.w6(32'h3aa6be0d),
	.w7(32'hbb3cb6f0),
	.w8(32'hbb5ab286),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba981145),
	.w1(32'h3b3f7e89),
	.w2(32'h3bb9b1e1),
	.w3(32'hb91b6287),
	.w4(32'hba868390),
	.w5(32'h3a8587a4),
	.w6(32'hbb0b0be0),
	.w7(32'hbab9da57),
	.w8(32'hbb09b445),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b936cb6),
	.w1(32'hb9dd884d),
	.w2(32'h3b1fd26a),
	.w3(32'h3b17a246),
	.w4(32'hbb2b141b),
	.w5(32'hbc168455),
	.w6(32'h3a8eb8b9),
	.w7(32'h3aa29f0e),
	.w8(32'hbb1246d3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf42d2),
	.w1(32'hbad21ddf),
	.w2(32'hbbae1b11),
	.w3(32'h3ba134e3),
	.w4(32'hbb31a0a6),
	.w5(32'h3b145e6f),
	.w6(32'hbac0bb55),
	.w7(32'hbaa69f30),
	.w8(32'h3b55247d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a2439),
	.w1(32'h3bc62d87),
	.w2(32'h3b37df8b),
	.w3(32'hbb79fb2b),
	.w4(32'h3b226e50),
	.w5(32'hbaed9ce2),
	.w6(32'hbae7913f),
	.w7(32'h3b4a3c7e),
	.w8(32'h3acb7238),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4248c6),
	.w1(32'hbc093183),
	.w2(32'hbad41deb),
	.w3(32'h39e7ab36),
	.w4(32'h3b14451e),
	.w5(32'hbbfa1820),
	.w6(32'hba7bdc94),
	.w7(32'h3af7b490),
	.w8(32'hbb8c9d9a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa92e1),
	.w1(32'h3a837cf8),
	.w2(32'hbad1d824),
	.w3(32'h3b3cfa4d),
	.w4(32'h3b1a0a0e),
	.w5(32'hbc048dcc),
	.w6(32'hbb892d83),
	.w7(32'h3b0f3d82),
	.w8(32'h39fad924),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06bf4d),
	.w1(32'hbbd14939),
	.w2(32'h3bc85788),
	.w3(32'h3a0f44c2),
	.w4(32'hbb76a36e),
	.w5(32'h3bb9ce4f),
	.w6(32'h39aaf2db),
	.w7(32'hbb11cd17),
	.w8(32'h382e0f8e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94d57f),
	.w1(32'hbb85e20f),
	.w2(32'hba7791fd),
	.w3(32'hbb3a6aa4),
	.w4(32'h3b76af08),
	.w5(32'hbbb81338),
	.w6(32'h3b576816),
	.w7(32'h3c16703f),
	.w8(32'h3bfcf891),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b92c),
	.w1(32'hbbe4b9cb),
	.w2(32'h3b915ec4),
	.w3(32'hbb5dca00),
	.w4(32'h3ae4a934),
	.w5(32'hbb2d102f),
	.w6(32'hba4dd68c),
	.w7(32'h3c0e528c),
	.w8(32'h39922fb4),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b2107),
	.w1(32'hbbe5477b),
	.w2(32'hbb10e535),
	.w3(32'h3bc88b29),
	.w4(32'hbb7b0362),
	.w5(32'hbbfe35b2),
	.w6(32'h3b325111),
	.w7(32'h3b92d99c),
	.w8(32'h3b923229),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d6bbb),
	.w1(32'hbb89ac21),
	.w2(32'hbaa25ab7),
	.w3(32'hb938f168),
	.w4(32'hbad44c0e),
	.w5(32'hb9a533a2),
	.w6(32'h3c234084),
	.w7(32'hbaa3b118),
	.w8(32'h3a9b7942),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb149609),
	.w1(32'h3c0a9f54),
	.w2(32'hbb5b0378),
	.w3(32'hba045f6a),
	.w4(32'h3bf9f4b0),
	.w5(32'hb9cee702),
	.w6(32'hba7d9db3),
	.w7(32'h3ba5c08b),
	.w8(32'h3b9dccdc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ccc0d),
	.w1(32'hbb30fd26),
	.w2(32'h3b958a24),
	.w3(32'hba3c8ab3),
	.w4(32'hba812cee),
	.w5(32'h3b960313),
	.w6(32'hba98a3b3),
	.w7(32'h3aab9442),
	.w8(32'hba871b2d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391cf2ae),
	.w1(32'hbbaba982),
	.w2(32'hba20b60d),
	.w3(32'hba9747c4),
	.w4(32'hbb312742),
	.w5(32'hbb14ddd6),
	.w6(32'h3b866a6f),
	.w7(32'h3bb624a9),
	.w8(32'h3b3bbc3c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c8c9b),
	.w1(32'hbb83e1cc),
	.w2(32'h3b0eb665),
	.w3(32'h3ad2e592),
	.w4(32'hbb8f32dd),
	.w5(32'h3c14f2d8),
	.w6(32'h3acbd3d1),
	.w7(32'h3aceeb6f),
	.w8(32'h3b92eb41),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc7058),
	.w1(32'h3b649709),
	.w2(32'hb9c89fa1),
	.w3(32'h3a95b008),
	.w4(32'hb97e0819),
	.w5(32'h39baf961),
	.w6(32'h3c53aefe),
	.w7(32'h3b8ce501),
	.w8(32'hba4403af),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf18de5),
	.w1(32'hbbc2ee59),
	.w2(32'hbae6472e),
	.w3(32'hbb0a3e86),
	.w4(32'hbbee98ae),
	.w5(32'hbb55f91b),
	.w6(32'h3b899b2b),
	.w7(32'h398b71b3),
	.w8(32'hbbb55ba7),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc122bf9),
	.w1(32'hbbd8c170),
	.w2(32'h3b877b20),
	.w3(32'hbb78ed88),
	.w4(32'h3a440a2d),
	.w5(32'hbbaf3787),
	.w6(32'hb8d68533),
	.w7(32'h3ba12194),
	.w8(32'h3b09d889),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a5183),
	.w1(32'hbc2e6b6a),
	.w2(32'hbba338f4),
	.w3(32'hba3f4177),
	.w4(32'hbafd4769),
	.w5(32'hbb2be375),
	.w6(32'h3a883587),
	.w7(32'h3b91808e),
	.w8(32'h3be87c53),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbf0d5),
	.w1(32'h39b21a35),
	.w2(32'hbaeeb1f6),
	.w3(32'hbb26530f),
	.w4(32'h3aff0741),
	.w5(32'hb89b899d),
	.w6(32'hbb293a84),
	.w7(32'hba41c916),
	.w8(32'h3ae530a3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e3a6),
	.w1(32'hbb47306d),
	.w2(32'hbb0842a4),
	.w3(32'h3b714e29),
	.w4(32'hbb98e5ef),
	.w5(32'hbb9583e0),
	.w6(32'hbaadbaf3),
	.w7(32'hba7c1062),
	.w8(32'hb95d558b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba07cec),
	.w1(32'hb923bf11),
	.w2(32'h3b826968),
	.w3(32'hbbbc2aa1),
	.w4(32'hba1c9843),
	.w5(32'h3b9e21f3),
	.w6(32'hbb3c0999),
	.w7(32'hba05e57d),
	.w8(32'h3ab05ea6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae48d53),
	.w1(32'hbb86b42d),
	.w2(32'hbb000ee0),
	.w3(32'h3c0c98f1),
	.w4(32'h3a51e360),
	.w5(32'h3bf5d7c1),
	.w6(32'h3c2c87ad),
	.w7(32'h3b88a117),
	.w8(32'h3bd22c02),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bdc24),
	.w1(32'hbaaaa7be),
	.w2(32'hbbcb603c),
	.w3(32'h3ab5cfc0),
	.w4(32'hbaf3c74d),
	.w5(32'hbc35c6d2),
	.w6(32'h3c6b77a6),
	.w7(32'h3a1ec5c2),
	.w8(32'hbb3de237),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c19f9),
	.w1(32'h3ab62a35),
	.w2(32'hbaaafeb1),
	.w3(32'hba9fc37a),
	.w4(32'h3b6fd368),
	.w5(32'h39728785),
	.w6(32'hbc131485),
	.w7(32'hbb01dbe9),
	.w8(32'hb9d051af),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5498bc),
	.w1(32'h3b92f623),
	.w2(32'hbacad012),
	.w3(32'hb7c2f2b2),
	.w4(32'h3b9154e5),
	.w5(32'h3b5ede1d),
	.w6(32'hbb5016c4),
	.w7(32'h3af6bcb6),
	.w8(32'h3b3391e1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c89d67),
	.w1(32'hbba321ec),
	.w2(32'hb952f466),
	.w3(32'h3a62ea6b),
	.w4(32'h3a4a09ec),
	.w5(32'hbc17bfe8),
	.w6(32'h3b44d923),
	.w7(32'hbb2bad83),
	.w8(32'hbb358f88),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fd6ca),
	.w1(32'hb8aa8751),
	.w2(32'h3aaece0f),
	.w3(32'h38a1f59b),
	.w4(32'hba390744),
	.w5(32'hbc264604),
	.w6(32'hbb2c113f),
	.w7(32'hba77a296),
	.w8(32'hbae88ab2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72a0d4),
	.w1(32'hbbef4f0a),
	.w2(32'h3bc2fb0f),
	.w3(32'h3b828e9f),
	.w4(32'hbbb6393e),
	.w5(32'h3af67d29),
	.w6(32'h3ae25b6e),
	.w7(32'hbb29178e),
	.w8(32'hbbe0ea7e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd0e4),
	.w1(32'hbc2ef5ef),
	.w2(32'hbad6fd49),
	.w3(32'h3c025dd4),
	.w4(32'hba66e2e1),
	.w5(32'hbb481d45),
	.w6(32'h3b2f72de),
	.w7(32'h3bc19b77),
	.w8(32'hb9ef288d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc443f0e),
	.w1(32'hbcb97166),
	.w2(32'hbc522969),
	.w3(32'h3b8b5d36),
	.w4(32'hbc94d872),
	.w5(32'hbc865156),
	.w6(32'h3c750219),
	.w7(32'h3aba627a),
	.w8(32'hba23d11e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbc63b),
	.w1(32'hbb098a25),
	.w2(32'hbad05309),
	.w3(32'hbb91bb03),
	.w4(32'hbbc244b1),
	.w5(32'hbb2812e2),
	.w6(32'hbaea39c8),
	.w7(32'hbb9317b7),
	.w8(32'hbbb55602),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3531c),
	.w1(32'hbbab4636),
	.w2(32'hbab458e1),
	.w3(32'hbac10083),
	.w4(32'hbb30c410),
	.w5(32'hbb8f35b3),
	.w6(32'hbb3770da),
	.w7(32'h3bcd4b6f),
	.w8(32'h3b8fed04),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule