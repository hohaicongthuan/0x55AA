module layer_10_featuremap_64(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf03a4d),
	.w1(32'h3b1ed842),
	.w2(32'hbad0252d),
	.w3(32'h3bf51748),
	.w4(32'h3b0ca740),
	.w5(32'hbba30e24),
	.w6(32'h3b9dcfd3),
	.w7(32'h3bf85c3c),
	.w8(32'h3c8d63ae),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52b5e7),
	.w1(32'hbb0afc37),
	.w2(32'h3bb51a85),
	.w3(32'h398a9278),
	.w4(32'hbc091859),
	.w5(32'hbbb6cee6),
	.w6(32'h3cb970bf),
	.w7(32'h3b26c788),
	.w8(32'h3b16f87e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc089e27),
	.w1(32'h3b8b62c8),
	.w2(32'hbc8ae7b8),
	.w3(32'hbc070035),
	.w4(32'h38521b5a),
	.w5(32'hbc627cca),
	.w6(32'h3a53d7bd),
	.w7(32'hba7d570d),
	.w8(32'hbbd44b64),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b81df),
	.w1(32'hbbb7069c),
	.w2(32'hbb3512a2),
	.w3(32'hbc28f303),
	.w4(32'h3b13431d),
	.w5(32'h3c86cbfc),
	.w6(32'h3c0b58d2),
	.w7(32'h3c92de0e),
	.w8(32'h3b435ede),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fd937),
	.w1(32'hbbbda320),
	.w2(32'h3ca899a8),
	.w3(32'h3c995fdd),
	.w4(32'h3c1dcbf9),
	.w5(32'h3b60bc27),
	.w6(32'hbc00311f),
	.w7(32'hbb962906),
	.w8(32'hbd04f7f1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cacad),
	.w1(32'h3a2512ec),
	.w2(32'h3b51e7d9),
	.w3(32'hb9b8e94a),
	.w4(32'hbbe00dbf),
	.w5(32'hbb8d44e8),
	.w6(32'hbd083eff),
	.w7(32'hbbdb5d8d),
	.w8(32'hbbad20b4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97842f),
	.w1(32'h3a70f853),
	.w2(32'h3af1ca40),
	.w3(32'hb9f53ae5),
	.w4(32'hbb481e15),
	.w5(32'h3a88ed96),
	.w6(32'hbae9db22),
	.w7(32'hbb9dd390),
	.w8(32'h3b6df545),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc040c7c),
	.w1(32'hbb930438),
	.w2(32'h3b0de323),
	.w3(32'hba8ed708),
	.w4(32'hbb97e866),
	.w5(32'h3b83db62),
	.w6(32'h3a171211),
	.w7(32'hbaef71b8),
	.w8(32'h3b907d55),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a835f2e),
	.w1(32'hbb1cfe19),
	.w2(32'hbbf0ef8f),
	.w3(32'h3aef31c7),
	.w4(32'h390cb5d1),
	.w5(32'hbc022839),
	.w6(32'h3bcd0459),
	.w7(32'h3ac1eb0c),
	.w8(32'hbb63a541),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc176050),
	.w1(32'hbbad1457),
	.w2(32'h3b1234ea),
	.w3(32'hbc6a9850),
	.w4(32'hbc0907db),
	.w5(32'h39c99081),
	.w6(32'hbbbe18f4),
	.w7(32'h3b14143f),
	.w8(32'hbb00231e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa62dbb),
	.w1(32'h3ac2d851),
	.w2(32'hbbcc42ed),
	.w3(32'h3adb6e98),
	.w4(32'h3a842605),
	.w5(32'hbc5e523a),
	.w6(32'h39a561f8),
	.w7(32'h3a459343),
	.w8(32'hbbe48597),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78cb30),
	.w1(32'hbaa38d5e),
	.w2(32'hbb677b3e),
	.w3(32'hbc8612b7),
	.w4(32'h3b074243),
	.w5(32'hbb9ca3e3),
	.w6(32'h3bc77d08),
	.w7(32'h3c9f56a5),
	.w8(32'hbb6c3df5),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c8e76),
	.w1(32'hbb3c1530),
	.w2(32'hbb46fb38),
	.w3(32'hbb84f483),
	.w4(32'hbaad811d),
	.w5(32'hbb9585f6),
	.w6(32'hbb5869f1),
	.w7(32'hbb2e0ee3),
	.w8(32'hbbac0641),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3975f8a5),
	.w1(32'hbb9401fd),
	.w2(32'h3be52ea1),
	.w3(32'hbb1ba6c4),
	.w4(32'h3b955b78),
	.w5(32'h3c8cb7ce),
	.w6(32'h3c544243),
	.w7(32'h3b9a745d),
	.w8(32'h3ba40485),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9573d7),
	.w1(32'h3c65845f),
	.w2(32'hbadf626f),
	.w3(32'h3d090584),
	.w4(32'h3c4a006a),
	.w5(32'hba2caaf0),
	.w6(32'hb9f8cde8),
	.w7(32'hbc4e4087),
	.w8(32'hbbb4d8f2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc7efb),
	.w1(32'hbb715d51),
	.w2(32'h3b747a1c),
	.w3(32'hbb657f60),
	.w4(32'hbb343442),
	.w5(32'h3ae3abf1),
	.w6(32'h3bcfcc84),
	.w7(32'h3be765bd),
	.w8(32'hba725b24),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b870fe3),
	.w1(32'h3b5fcaad),
	.w2(32'hba7fea4f),
	.w3(32'h3b49b244),
	.w4(32'h3a2c5305),
	.w5(32'hbba381d6),
	.w6(32'h3a0ee593),
	.w7(32'h399461ba),
	.w8(32'hbb8ca7e1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ce570),
	.w1(32'hbaee73d8),
	.w2(32'h3b73bf8f),
	.w3(32'h3a066ce3),
	.w4(32'hbb15bad6),
	.w5(32'h3b983346),
	.w6(32'h38564051),
	.w7(32'hba5bcb97),
	.w8(32'h396a51b2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59e4a1),
	.w1(32'hbb4afa77),
	.w2(32'hbb15207d),
	.w3(32'h3b3fe9e0),
	.w4(32'h3b172f59),
	.w5(32'hbac0648d),
	.w6(32'h3b8f6d02),
	.w7(32'h3bf5e109),
	.w8(32'hb9e6df97),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6beac9),
	.w1(32'h3b03bf46),
	.w2(32'h3b8aa9f1),
	.w3(32'h3b985998),
	.w4(32'h3c4d17b3),
	.w5(32'h3aee8e32),
	.w6(32'h3c83d946),
	.w7(32'h3c3d9bf5),
	.w8(32'h39c96791),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f549c),
	.w1(32'h3b89b4d9),
	.w2(32'hbb9b6644),
	.w3(32'h3ba221c2),
	.w4(32'h3b2c3cc9),
	.w5(32'hba0ef9b7),
	.w6(32'hba8b853d),
	.w7(32'h3b19f886),
	.w8(32'h3ab69839),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53c75a),
	.w1(32'hbc4e0fc0),
	.w2(32'hbb9f33fa),
	.w3(32'h3bb05586),
	.w4(32'hbbda98e8),
	.w5(32'h391f3ca6),
	.w6(32'h3cb0a703),
	.w7(32'h3c9f73db),
	.w8(32'hba8e6077),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb300),
	.w1(32'hbb89d045),
	.w2(32'hbb938941),
	.w3(32'h3ba29297),
	.w4(32'h3acde430),
	.w5(32'hbbe16399),
	.w6(32'hbc3b4c6e),
	.w7(32'hb9b36fb5),
	.w8(32'hbbf8b198),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba243d2),
	.w1(32'hbbc098b0),
	.w2(32'hbb7a5449),
	.w3(32'hbbe7e3d8),
	.w4(32'hbbf7bdf1),
	.w5(32'hba3656cd),
	.w6(32'hbc05ee77),
	.w7(32'hbbf0a408),
	.w8(32'hbb533a79),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d4bae),
	.w1(32'hbc1de4a7),
	.w2(32'hbbc203d8),
	.w3(32'h3b7592b5),
	.w4(32'hbada2c84),
	.w5(32'hbb9d8caa),
	.w6(32'h3b95ab76),
	.w7(32'h39a1b316),
	.w8(32'h3b59dc5d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada9596),
	.w1(32'h3b75b19d),
	.w2(32'hbc031a47),
	.w3(32'h3caa74ef),
	.w4(32'h3c836e5d),
	.w5(32'h3c4a2af0),
	.w6(32'h3c744779),
	.w7(32'h3c6e1b69),
	.w8(32'h3c74529e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc8c7c5),
	.w1(32'hbcd53baf),
	.w2(32'h39828254),
	.w3(32'hbb47b383),
	.w4(32'hbc72e0f8),
	.w5(32'hba138c8d),
	.w6(32'h3c2129c5),
	.w7(32'hbbabb567),
	.w8(32'h3a00f273),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f531da),
	.w1(32'h38c156fc),
	.w2(32'h3b5dd037),
	.w3(32'hba9d6910),
	.w4(32'hbaad10da),
	.w5(32'h390a584e),
	.w6(32'h36aa7e21),
	.w7(32'hb9b4d7a9),
	.w8(32'hbbdbfbef),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903ca6b),
	.w1(32'h3b1edf7c),
	.w2(32'hb9f537f6),
	.w3(32'hbb93a985),
	.w4(32'h3ae5e7d0),
	.w5(32'hbb57e0c8),
	.w6(32'hbbb3c826),
	.w7(32'h3a181e22),
	.w8(32'h3b72032e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08613c),
	.w1(32'hbbcd767d),
	.w2(32'h3abc01c0),
	.w3(32'h39b2cdab),
	.w4(32'h3ab52eb5),
	.w5(32'h3aa00ba9),
	.w6(32'h3b7183ee),
	.w7(32'h3c0d439d),
	.w8(32'hb80f5546),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205113),
	.w1(32'hbb84d51e),
	.w2(32'hbb36b74a),
	.w3(32'hbb6f152e),
	.w4(32'hbb36643e),
	.w5(32'hbb94a0ad),
	.w6(32'hbb6a796d),
	.w7(32'hbae84219),
	.w8(32'hbbc89641),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c56f8),
	.w1(32'hbc132cb2),
	.w2(32'hbc2d5f9d),
	.w3(32'h3aa0aa51),
	.w4(32'h3adc7007),
	.w5(32'hbc434b1a),
	.w6(32'hbb12e4a3),
	.w7(32'hbb074fe4),
	.w8(32'hbbf3310e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a7f15),
	.w1(32'hbc2fbd6a),
	.w2(32'h3b603ca3),
	.w3(32'hbbc86719),
	.w4(32'hbba3336f),
	.w5(32'hbb186c40),
	.w6(32'hbbf4846e),
	.w7(32'hbc0298fa),
	.w8(32'hbbc8fd65),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42623c),
	.w1(32'h3bc72dc0),
	.w2(32'h3b5dcd07),
	.w3(32'hb92081e6),
	.w4(32'h3b152ff9),
	.w5(32'h3bc35bc5),
	.w6(32'hbc00ab22),
	.w7(32'hbad1b561),
	.w8(32'h3c5860b3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25c198),
	.w1(32'hbba2f1e8),
	.w2(32'hbb1126e7),
	.w3(32'hbb82c4b0),
	.w4(32'hbad028de),
	.w5(32'hbb62d219),
	.w6(32'h3c297948),
	.w7(32'h3a9c5017),
	.w8(32'hbb88305d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa62688),
	.w1(32'h3af74abb),
	.w2(32'hbb82ec97),
	.w3(32'hba6f1509),
	.w4(32'h3a1ff357),
	.w5(32'hbad516d1),
	.w6(32'hbb1f0f83),
	.w7(32'hb9deea48),
	.w8(32'hba134c08),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c8e2b),
	.w1(32'hba2e3fdf),
	.w2(32'h3b396273),
	.w3(32'hbb70cb56),
	.w4(32'hbbe9eeab),
	.w5(32'h38442891),
	.w6(32'h3baa511a),
	.w7(32'hba82b1c4),
	.w8(32'hbb97786b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0b2e2),
	.w1(32'h3bdb2e23),
	.w2(32'hb99ea6c6),
	.w3(32'h3b0184a9),
	.w4(32'h3be1a62a),
	.w5(32'h3c610056),
	.w6(32'hbad9349d),
	.w7(32'h3b745536),
	.w8(32'h3c2d99be),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abbe40),
	.w1(32'h3ac85994),
	.w2(32'h3c899d03),
	.w3(32'h3bbf3f68),
	.w4(32'h3c0e157a),
	.w5(32'h3c31b57b),
	.w6(32'h3c4a40b2),
	.w7(32'h3c0c7e48),
	.w8(32'h3be59f6b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c920d25),
	.w1(32'h3b715fb2),
	.w2(32'h3b6005d7),
	.w3(32'h3c493a77),
	.w4(32'h3c3961ee),
	.w5(32'h3b6cc7f2),
	.w6(32'h3bf29595),
	.w7(32'h3c396665),
	.w8(32'h3c4f2875),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc373f),
	.w1(32'hbb153641),
	.w2(32'hbc1f6551),
	.w3(32'hbad702e4),
	.w4(32'hbbb6d999),
	.w5(32'hbbcfba5f),
	.w6(32'h3c38ae0f),
	.w7(32'h3c193162),
	.w8(32'h3ab3f1bb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70d6bd),
	.w1(32'hbc95b57a),
	.w2(32'hbb46ce7f),
	.w3(32'hbc12ec7d),
	.w4(32'hbc20d079),
	.w5(32'hbbd4a3f2),
	.w6(32'h3b0f81a4),
	.w7(32'hba96c4b4),
	.w8(32'hbc03d2b3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b646eb7),
	.w1(32'h3a90497f),
	.w2(32'hbbf23f0f),
	.w3(32'hba849d73),
	.w4(32'h39b1b928),
	.w5(32'hbb80da7a),
	.w6(32'hba4e563f),
	.w7(32'h3acb9e04),
	.w8(32'hbbe2093c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb888356),
	.w1(32'hba0a35dd),
	.w2(32'hbbb11354),
	.w3(32'hbacd876f),
	.w4(32'hb9fa7b17),
	.w5(32'hb78fd02c),
	.w6(32'hbaa59945),
	.w7(32'hbae73c29),
	.w8(32'h3b11e565),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17d93a),
	.w1(32'hbb8f15e2),
	.w2(32'hb9cf0d9a),
	.w3(32'hbaafeda8),
	.w4(32'hbc00f08b),
	.w5(32'hba5712c0),
	.w6(32'h3a09af3f),
	.w7(32'hbb4da4ad),
	.w8(32'h3afd8549),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09a424),
	.w1(32'hbc1e28cc),
	.w2(32'hba1f01f3),
	.w3(32'hbbd8b55d),
	.w4(32'hbb0aa6b7),
	.w5(32'hbb6325d8),
	.w6(32'h3b790046),
	.w7(32'h3b6189ec),
	.w8(32'hbbc9f636),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b572b0e),
	.w1(32'hbb749798),
	.w2(32'h3b57494d),
	.w3(32'h397d9def),
	.w4(32'h3b004218),
	.w5(32'hbb87be28),
	.w6(32'hbc1f30ad),
	.w7(32'h3b80702a),
	.w8(32'hbb8dae93),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d1361),
	.w1(32'h3a14469c),
	.w2(32'h3ad2fa51),
	.w3(32'hbb4f475b),
	.w4(32'hba9118f2),
	.w5(32'h3b031615),
	.w6(32'hbc17bf71),
	.w7(32'hbc1368f0),
	.w8(32'hbb5898df),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92019d),
	.w1(32'h3b23044c),
	.w2(32'h3a131aec),
	.w3(32'h3ba969cd),
	.w4(32'h3b6ad70d),
	.w5(32'h3b85bca2),
	.w6(32'h3a8ddfa5),
	.w7(32'hba0e2016),
	.w8(32'h3c4f5694),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d3d0a),
	.w1(32'hbb909db3),
	.w2(32'hbb9bff81),
	.w3(32'hba968198),
	.w4(32'hba400e2c),
	.w5(32'hbb76dea8),
	.w6(32'h3c7b702b),
	.w7(32'h3baab469),
	.w8(32'h3b9ce608),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a3a86),
	.w1(32'hbad5881f),
	.w2(32'hb9c7343b),
	.w3(32'hba36fdbc),
	.w4(32'h3b96ac49),
	.w5(32'h3b1c2c70),
	.w6(32'h399178d6),
	.w7(32'h37dd4bf1),
	.w8(32'hbc7914bd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babb236),
	.w1(32'h3b647e79),
	.w2(32'hbc05fcf4),
	.w3(32'h3ba64bcf),
	.w4(32'h3b038137),
	.w5(32'hbc1a3c3a),
	.w6(32'hbab84e19),
	.w7(32'hbbf59e31),
	.w8(32'hba7065bd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f4e80),
	.w1(32'hbbeedd0f),
	.w2(32'hbc85a963),
	.w3(32'hbbd1a856),
	.w4(32'hbb040524),
	.w5(32'hbc9d36d2),
	.w6(32'hbbe58b96),
	.w7(32'hbbde3b74),
	.w8(32'hbca94673),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc724a3d),
	.w1(32'hbc596a36),
	.w2(32'hba479357),
	.w3(32'hbca05af7),
	.w4(32'hbcb16f4d),
	.w5(32'hbc8fd382),
	.w6(32'hbc3939e9),
	.w7(32'hbc7c5ca1),
	.w8(32'hbc1abcc4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2dbfb),
	.w1(32'hbb74820b),
	.w2(32'hbb319c60),
	.w3(32'hbc50616c),
	.w4(32'hbbd3e22c),
	.w5(32'h3bcc365a),
	.w6(32'hbc345b46),
	.w7(32'h3b312168),
	.w8(32'h3c0e5716),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6bdf1),
	.w1(32'hbbd52f2f),
	.w2(32'hbc026343),
	.w3(32'h3b214046),
	.w4(32'h3b9248eb),
	.w5(32'hbb3bad6b),
	.w6(32'h3c51ea1e),
	.w7(32'h3c088a6b),
	.w8(32'hbbb542dd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a50a0),
	.w1(32'hbbe540bd),
	.w2(32'hbb267066),
	.w3(32'hbaf8ccc3),
	.w4(32'h37c0edda),
	.w5(32'hbb195d64),
	.w6(32'hbb6a3915),
	.w7(32'h3b7444f0),
	.w8(32'hbbbb31c0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba146eac),
	.w1(32'h3b517e95),
	.w2(32'hbaf7b7d3),
	.w3(32'hba602799),
	.w4(32'h3b15d222),
	.w5(32'hbb124ccd),
	.w6(32'hba495fc2),
	.w7(32'h3b4b7bcb),
	.w8(32'hbb17af68),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1e34c),
	.w1(32'h3926317a),
	.w2(32'h3b9bd356),
	.w3(32'hbb6d46b7),
	.w4(32'hbb172d78),
	.w5(32'h3bf57e12),
	.w6(32'hbbeb446e),
	.w7(32'hbb99938a),
	.w8(32'h3ca4b439),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aa2b2),
	.w1(32'h3c9d04e7),
	.w2(32'hbafc1abd),
	.w3(32'h3c497d54),
	.w4(32'h3c41df81),
	.w5(32'hbb09ad54),
	.w6(32'h3cbd03f6),
	.w7(32'h3c7b8432),
	.w8(32'hbb8ae293),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a082675),
	.w1(32'h3b20a7f8),
	.w2(32'h3ba0125e),
	.w3(32'h3b4db927),
	.w4(32'h38f4eb4f),
	.w5(32'h3c8e33b5),
	.w6(32'hbb15ceab),
	.w7(32'hbbdde4ee),
	.w8(32'h3c51687f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba991fd9),
	.w1(32'hbb239534),
	.w2(32'hbb34f891),
	.w3(32'h3c23d4cb),
	.w4(32'hbb4ff68c),
	.w5(32'hbbba68a6),
	.w6(32'h3caaab1e),
	.w7(32'h3c25dbac),
	.w8(32'hbaeb4631),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92c784),
	.w1(32'h3a5f88a8),
	.w2(32'hbb32680a),
	.w3(32'hbbbacba0),
	.w4(32'hba41a5f2),
	.w5(32'h3b10c91b),
	.w6(32'hbbce9134),
	.w7(32'h38a905a3),
	.w8(32'hba37ddac),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e3e18),
	.w1(32'hbb00d869),
	.w2(32'hbb448d83),
	.w3(32'h3b9e4951),
	.w4(32'h3b761131),
	.w5(32'h3b838331),
	.w6(32'hbb0736ad),
	.w7(32'h3ac42d3c),
	.w8(32'hbba9eee6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a51732),
	.w1(32'hbc12eb08),
	.w2(32'hbc152ab2),
	.w3(32'h3c1d6b3d),
	.w4(32'h3b9b9573),
	.w5(32'hbc0ad8ac),
	.w6(32'h3a629f20),
	.w7(32'h39b2a8b6),
	.w8(32'hbc6d3e23),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71aa77),
	.w1(32'hbc90676d),
	.w2(32'hbb2c3be6),
	.w3(32'hbc676c53),
	.w4(32'hbc6d76f3),
	.w5(32'h3b8c41f5),
	.w6(32'hbc5bc6f4),
	.w7(32'hbc424c28),
	.w8(32'h3bad572d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d67a9f),
	.w1(32'h3b63ab8f),
	.w2(32'hbb494680),
	.w3(32'h3b762dda),
	.w4(32'h3b9b4fd3),
	.w5(32'hbac5abd1),
	.w6(32'h3c10d748),
	.w7(32'h3bed02a4),
	.w8(32'hb9ce3723),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45378c),
	.w1(32'hbb3fafed),
	.w2(32'hbb85c8ca),
	.w3(32'h399f26f9),
	.w4(32'h38393da0),
	.w5(32'hbb983bf3),
	.w6(32'hb90f4172),
	.w7(32'h3bb785b5),
	.w8(32'hbc05c188),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22e889),
	.w1(32'hbb6bd367),
	.w2(32'h3c26c93f),
	.w3(32'hbc26050d),
	.w4(32'hbbb71fc0),
	.w5(32'h3bd4615e),
	.w6(32'hbbff0365),
	.w7(32'hbb8ef2b9),
	.w8(32'h3c24e4cb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28e7ab),
	.w1(32'h3bc9ac93),
	.w2(32'h3c6274ee),
	.w3(32'h3be6a8c4),
	.w4(32'h3b718183),
	.w5(32'h3c601f0e),
	.w6(32'h3c222e2e),
	.w7(32'h3be4ca90),
	.w8(32'h3c82258d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21f179),
	.w1(32'h38f08f18),
	.w2(32'hbb3570c2),
	.w3(32'h3c264ee2),
	.w4(32'h3bda28cd),
	.w5(32'hbb0895c5),
	.w6(32'h3c758d1f),
	.w7(32'h3c1943fe),
	.w8(32'hbbac0167),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae5280),
	.w1(32'hbbf7edf5),
	.w2(32'hbbac0a48),
	.w3(32'hbbaa34b4),
	.w4(32'hbbae3289),
	.w5(32'h39a92a68),
	.w6(32'hbbf7a6cd),
	.w7(32'hbaead65e),
	.w8(32'hba64e41e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53b0b1),
	.w1(32'hbbe0fc54),
	.w2(32'h3b9a2195),
	.w3(32'hbb4e4434),
	.w4(32'hbb584ca5),
	.w5(32'h3bd7afe7),
	.w6(32'hbb113221),
	.w7(32'hbb257cd1),
	.w8(32'h3bd0361d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bafad),
	.w1(32'hbbb8eceb),
	.w2(32'h3be5de6f),
	.w3(32'h3b3f8538),
	.w4(32'hbb7c25b4),
	.w5(32'h3bcf6aa8),
	.w6(32'h3ba5cab4),
	.w7(32'hbb160d8c),
	.w8(32'h3b11deb0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1dc4a),
	.w1(32'h3a02b04f),
	.w2(32'h39c9eeab),
	.w3(32'h3b213b82),
	.w4(32'h3b6ca6f6),
	.w5(32'hbb912099),
	.w6(32'hbb1eba97),
	.w7(32'hb9b8b628),
	.w8(32'hbc4ff53d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95251a),
	.w1(32'hb9951a84),
	.w2(32'hbbdd9645),
	.w3(32'hbb6bd4cf),
	.w4(32'hb9f2e40a),
	.w5(32'hbb8c15ce),
	.w6(32'hbc4a1ee6),
	.w7(32'hbbc00e74),
	.w8(32'hbb842ee5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00a279),
	.w1(32'h39fbd58d),
	.w2(32'h3b0a016d),
	.w3(32'hbc20018e),
	.w4(32'hbba6f447),
	.w5(32'hbbb227f4),
	.w6(32'hbbcf000f),
	.w7(32'hbc08c9d5),
	.w8(32'hbc15a69b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7262b3),
	.w1(32'hbc053a7e),
	.w2(32'h3b92459c),
	.w3(32'h3bc35fad),
	.w4(32'hbad9c430),
	.w5(32'hbbf54e12),
	.w6(32'hbb0f9236),
	.w7(32'hbc674bca),
	.w8(32'hbc162149),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0436aa),
	.w1(32'hbc560002),
	.w2(32'h38b5e797),
	.w3(32'hbb8d7230),
	.w4(32'hbc3c7911),
	.w5(32'hbbae3c33),
	.w6(32'hbc8174b1),
	.w7(32'hbb953576),
	.w8(32'h3a62b18e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65694e),
	.w1(32'h3a9c97fe),
	.w2(32'h3b22eb8a),
	.w3(32'hbb60f94c),
	.w4(32'hbc030e90),
	.w5(32'h3b969865),
	.w6(32'h3bbf3e41),
	.w7(32'h39eb5b1c),
	.w8(32'h3b6f301e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81e3c0),
	.w1(32'hbb8886ed),
	.w2(32'h3881aca1),
	.w3(32'h3bf15cb0),
	.w4(32'h3ac38b9d),
	.w5(32'h39af5cec),
	.w6(32'h3b8bce54),
	.w7(32'h3b4506c7),
	.w8(32'hbb65b6d7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac50f17),
	.w1(32'h3aba1879),
	.w2(32'h3b7e1211),
	.w3(32'hbb161303),
	.w4(32'hba8bb0d5),
	.w5(32'h3c05b973),
	.w6(32'hbbcb6fec),
	.w7(32'hbb23887b),
	.w8(32'hbb0ba316),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd73e75),
	.w1(32'hbc3575e2),
	.w2(32'h3ac3f846),
	.w3(32'h3b0e51b1),
	.w4(32'hbbf7f9ce),
	.w5(32'h3c5c5c95),
	.w6(32'hbb8c06fc),
	.w7(32'hbc0cfbdb),
	.w8(32'h3b708c8e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1328cb),
	.w1(32'h3a5f778e),
	.w2(32'h3a954f4e),
	.w3(32'h3c52d6d5),
	.w4(32'h3bb9919c),
	.w5(32'h3b7bf2ea),
	.w6(32'h3c1d8f18),
	.w7(32'h3c78576f),
	.w8(32'hbb9a7cf4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95682e),
	.w1(32'h3b047e3e),
	.w2(32'hba187899),
	.w3(32'hba50cf06),
	.w4(32'h3b0d3d0c),
	.w5(32'hbb96f852),
	.w6(32'hbbe42794),
	.w7(32'hbb17e2f9),
	.w8(32'hbbbc56a7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef4645),
	.w1(32'hba80455a),
	.w2(32'hbc18344c),
	.w3(32'hbbe620cc),
	.w4(32'hb93c62d1),
	.w5(32'hbbc076a4),
	.w6(32'h3b511d19),
	.w7(32'h38cb7413),
	.w8(32'hbc8ff892),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61a567),
	.w1(32'hbc8c3dbc),
	.w2(32'h3b556b24),
	.w3(32'hbc338227),
	.w4(32'hbc1b5422),
	.w5(32'h3b8a6324),
	.w6(32'hbc6fc9a5),
	.w7(32'hbbc534ad),
	.w8(32'h3ba25e64),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05f7b2),
	.w1(32'hbb400914),
	.w2(32'hb96d5baf),
	.w3(32'h3b900937),
	.w4(32'h3a9acb9a),
	.w5(32'hbae98c9a),
	.w6(32'h3baaa94c),
	.w7(32'h3b213277),
	.w8(32'hbc0e143c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8f73),
	.w1(32'h3a475d14),
	.w2(32'hbbb747c1),
	.w3(32'hbbb16b3a),
	.w4(32'hbb49d9cb),
	.w5(32'hbae080ff),
	.w6(32'h39013f27),
	.w7(32'h3bc5d207),
	.w8(32'hbad2c891),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2beff8),
	.w1(32'hbc16191b),
	.w2(32'hbc29e1a1),
	.w3(32'h3b00c004),
	.w4(32'hbb82e54a),
	.w5(32'hbc14e37b),
	.w6(32'h3c4cd679),
	.w7(32'h3c0875d3),
	.w8(32'hbc9a23d1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc944a5c),
	.w1(32'hbc984561),
	.w2(32'h3a620297),
	.w3(32'hbc432d22),
	.w4(32'hbc751529),
	.w5(32'h3bd528bd),
	.w6(32'hbc90a088),
	.w7(32'hbc6f70aa),
	.w8(32'h3c3fae65),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22b8ff),
	.w1(32'h3b960f4a),
	.w2(32'h3bf61db1),
	.w3(32'h3b57f2ea),
	.w4(32'h3c181f7d),
	.w5(32'h3ac389db),
	.w6(32'h3b48fe85),
	.w7(32'h3b2bd9bb),
	.w8(32'h3b8b7595),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c009f98),
	.w1(32'h3bab5dfc),
	.w2(32'hba8fc0e7),
	.w3(32'h3ac60acf),
	.w4(32'h39e99009),
	.w5(32'h3a2b11ab),
	.w6(32'h3bbf0f63),
	.w7(32'h3b65f203),
	.w8(32'h3b7fd1c0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b76e0a),
	.w1(32'hba8d94ae),
	.w2(32'hbb90994a),
	.w3(32'hba8b4729),
	.w4(32'hbb646a1c),
	.w5(32'hbb82e258),
	.w6(32'h3b69edb4),
	.w7(32'hba75d7d9),
	.w8(32'h395deb08),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad68c6d),
	.w1(32'hba8743d4),
	.w2(32'hbb1349ea),
	.w3(32'hbc0442e3),
	.w4(32'hbbc81e7c),
	.w5(32'hbaa9113c),
	.w6(32'hbb1ce110),
	.w7(32'hbba78779),
	.w8(32'hbb25d3a0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afba4bd),
	.w1(32'h3b371e4e),
	.w2(32'hbb7e6024),
	.w3(32'hbb0bc63e),
	.w4(32'h3b33e62f),
	.w5(32'h3a6261b5),
	.w6(32'h3bc30bb9),
	.w7(32'h3ba7d06e),
	.w8(32'hbc4b0bed),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4445),
	.w1(32'hbc39e169),
	.w2(32'hbaa915b6),
	.w3(32'h39373e7a),
	.w4(32'hba0326c4),
	.w5(32'hbaf8d0b2),
	.w6(32'h3b4d05f3),
	.w7(32'hbab58415),
	.w8(32'hbc3234d4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c4721),
	.w1(32'h39ad8a9b),
	.w2(32'hbaecf042),
	.w3(32'hb9cd3e64),
	.w4(32'hbacc0ecf),
	.w5(32'hbb511af4),
	.w6(32'hbb45040c),
	.w7(32'hbb861b91),
	.w8(32'hbb855ddd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4ed8b),
	.w1(32'hbb3be84d),
	.w2(32'h3bbffcfc),
	.w3(32'hbb888365),
	.w4(32'hbb68c39b),
	.w5(32'h3c2b7267),
	.w6(32'h3b0d1dc2),
	.w7(32'h3aa03f01),
	.w8(32'h3c44e042),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c975ee3),
	.w1(32'h3c87a84d),
	.w2(32'hbbc1ffe9),
	.w3(32'h3c7532a3),
	.w4(32'h3c82e676),
	.w5(32'hbb5962eb),
	.w6(32'h3c93c56b),
	.w7(32'h3c85e35c),
	.w8(32'hbc106cc4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd31476),
	.w1(32'hbb31fc1c),
	.w2(32'hbbcc674c),
	.w3(32'h3a92ffa2),
	.w4(32'hbb44edd2),
	.w5(32'hbc132f65),
	.w6(32'hbbdbb22a),
	.w7(32'hbbbb69f9),
	.w8(32'hbb816da5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffdd40),
	.w1(32'hbbe4814d),
	.w2(32'hba7b83d0),
	.w3(32'hbbfabfc8),
	.w4(32'hbb4d7ecd),
	.w5(32'hba86006c),
	.w6(32'hbb8a7cb9),
	.w7(32'hbba1db3d),
	.w8(32'hbb6b2d7d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba955c8),
	.w1(32'hba4be4be),
	.w2(32'hbc08eee7),
	.w3(32'hb913a1dc),
	.w4(32'hba128ef5),
	.w5(32'hbc2799c5),
	.w6(32'h3b519b52),
	.w7(32'h3be4c81d),
	.w8(32'hbc84d798),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46d95a),
	.w1(32'hbc348598),
	.w2(32'hbbaf09fa),
	.w3(32'hbc0794c4),
	.w4(32'hbbd3bf20),
	.w5(32'hbb804248),
	.w6(32'hbc82e7ed),
	.w7(32'hbc0daa5b),
	.w8(32'hbc065518),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f2b9e),
	.w1(32'hbb08fc54),
	.w2(32'hbac39d91),
	.w3(32'hbb0147ae),
	.w4(32'h39fb5924),
	.w5(32'hbb885c79),
	.w6(32'hbac9482e),
	.w7(32'hbc28528f),
	.w8(32'hbc247902),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ba09c),
	.w1(32'hbb20ba26),
	.w2(32'hbb34bf9d),
	.w3(32'hbb2c4f6b),
	.w4(32'hbb7e2266),
	.w5(32'hbb2cf344),
	.w6(32'hbbc43502),
	.w7(32'hba8d6995),
	.w8(32'hbc6d6446),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5eb0f),
	.w1(32'hbc21fd9e),
	.w2(32'h3bd6be45),
	.w3(32'hbbd74841),
	.w4(32'hbbe970a3),
	.w5(32'hb95a73b7),
	.w6(32'hbc1e48bc),
	.w7(32'hbbf87bc1),
	.w8(32'hbbb91bc9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24940d),
	.w1(32'h3b9c1f28),
	.w2(32'hba40d8c4),
	.w3(32'h3c611999),
	.w4(32'h3b3d2b9c),
	.w5(32'h3b3534a9),
	.w6(32'h3c80c0ac),
	.w7(32'h3c1abd40),
	.w8(32'hbb3c5060),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c260c23),
	.w1(32'h3b0bb344),
	.w2(32'hbbebc005),
	.w3(32'h3c046837),
	.w4(32'h3ba410ba),
	.w5(32'h3bac29ea),
	.w6(32'hba9f18a4),
	.w7(32'h3c04f69f),
	.w8(32'h3abf481a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca732c),
	.w1(32'hbc0f7857),
	.w2(32'h3b31c0cb),
	.w3(32'h3afc00cf),
	.w4(32'hbb44852a),
	.w5(32'h3aa4225f),
	.w6(32'h3bbf94c5),
	.w7(32'h3bcb932f),
	.w8(32'hbac6c2c6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1a89b),
	.w1(32'h3ba8b44f),
	.w2(32'hbab29599),
	.w3(32'h3b2a6c1c),
	.w4(32'hbb1a3331),
	.w5(32'h3b54630b),
	.w6(32'hbc12ba59),
	.w7(32'hbaa4a0a9),
	.w8(32'h3bd77ab1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d3637),
	.w1(32'hbbc77992),
	.w2(32'hbbb0d24f),
	.w3(32'h3ab953e4),
	.w4(32'hba179987),
	.w5(32'hbb7d3ffc),
	.w6(32'h3b7eb096),
	.w7(32'hbc20df97),
	.w8(32'hbb5fab00),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c2257),
	.w1(32'h3ac21adb),
	.w2(32'h3af50dde),
	.w3(32'h3c0f7091),
	.w4(32'hbaecb4de),
	.w5(32'h3b631cb9),
	.w6(32'h3c140235),
	.w7(32'h3b1185fb),
	.w8(32'h3c09eeb0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad74898),
	.w1(32'h3b25f4a2),
	.w2(32'hbb8febff),
	.w3(32'hbaafc9bd),
	.w4(32'hbad611b8),
	.w5(32'h3a3baaee),
	.w6(32'h3c379af3),
	.w7(32'h3ba24ed3),
	.w8(32'h3ae6b172),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5d099),
	.w1(32'h3b6adcfb),
	.w2(32'h3c5be39d),
	.w3(32'h3c215adb),
	.w4(32'h3c4e9b21),
	.w5(32'h3cb6e348),
	.w6(32'h3ba8d844),
	.w7(32'h3c0edc55),
	.w8(32'h3cca98d3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c957fcd),
	.w1(32'h3c6de01b),
	.w2(32'hbc8caa7e),
	.w3(32'h3cb8d84a),
	.w4(32'h3c83309a),
	.w5(32'hbc6d9236),
	.w6(32'h3cfbedbe),
	.w7(32'h3cc31a1a),
	.w8(32'hbd062464),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc01ba9),
	.w1(32'hbcd9bb4d),
	.w2(32'h3a9d963b),
	.w3(32'hbc84d35b),
	.w4(32'hbc57707c),
	.w5(32'h3c093898),
	.w6(32'hbcf09836),
	.w7(32'hbcca5e90),
	.w8(32'h3cb15e72),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03538a),
	.w1(32'h3c42e8f7),
	.w2(32'hbb9a68e0),
	.w3(32'h3c41ea55),
	.w4(32'h3c40d2e1),
	.w5(32'hbb47da87),
	.w6(32'h3cc64487),
	.w7(32'h3c8849f9),
	.w8(32'hbba4dd36),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc79ea6),
	.w1(32'hbb8b3fe9),
	.w2(32'hbb7669cd),
	.w3(32'h3ab133ee),
	.w4(32'h3b84ba34),
	.w5(32'hbc0b9beb),
	.w6(32'hbb3b9d1a),
	.w7(32'hba4c7b3a),
	.w8(32'hbbf7856f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc07b09),
	.w1(32'hbb9201d3),
	.w2(32'hba281837),
	.w3(32'h39109d87),
	.w4(32'hbb895349),
	.w5(32'hbad18d5b),
	.w6(32'hbb69fda7),
	.w7(32'hbb9d06bf),
	.w8(32'hbbfcfc5c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85ce3a),
	.w1(32'hbb12095d),
	.w2(32'h3b02b324),
	.w3(32'h3b8d27a3),
	.w4(32'h3b2c76b1),
	.w5(32'h3b701574),
	.w6(32'hbaf3faa6),
	.w7(32'hbbb14be8),
	.w8(32'h3b7a4c0b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d4285),
	.w1(32'hbb535b5a),
	.w2(32'hbb086e31),
	.w3(32'h3819dc6e),
	.w4(32'hba2db5c6),
	.w5(32'h3aa56049),
	.w6(32'h3acdd82b),
	.w7(32'hba8e3694),
	.w8(32'h3a89d5f6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc07dde),
	.w1(32'hbbf92549),
	.w2(32'hbb312116),
	.w3(32'hbb81262b),
	.w4(32'hbbe9ca6e),
	.w5(32'hbb8b2b51),
	.w6(32'hbb674b03),
	.w7(32'hbb2db27a),
	.w8(32'hbc7d099e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a2f06),
	.w1(32'hbc2307c9),
	.w2(32'hba38934b),
	.w3(32'h3b9f3ad5),
	.w4(32'hbb816a93),
	.w5(32'hbb026b2e),
	.w6(32'hbc189210),
	.w7(32'hbb1141d2),
	.w8(32'hbb17f649),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba603f43),
	.w1(32'h3b8436dc),
	.w2(32'hbb435827),
	.w3(32'h395efab9),
	.w4(32'h3b012da1),
	.w5(32'h3b742a59),
	.w6(32'h3ac81c8f),
	.w7(32'h3bc075fa),
	.w8(32'h3a34cc8f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf90bb1),
	.w1(32'h3af1a061),
	.w2(32'hbc1cbde4),
	.w3(32'h3b4b84bc),
	.w4(32'hb88cd2f2),
	.w5(32'hba9e16b2),
	.w6(32'h3c030536),
	.w7(32'h3b574e12),
	.w8(32'hbacb2232),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b28b6),
	.w1(32'h3b817a13),
	.w2(32'hbbbe27f1),
	.w3(32'h3b5448c8),
	.w4(32'hbb079c6b),
	.w5(32'hbb4440bd),
	.w6(32'h3b32f8f4),
	.w7(32'h3b9b0250),
	.w8(32'hbb76669a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a629749),
	.w1(32'hbbb39d9c),
	.w2(32'h39da2332),
	.w3(32'hb917610d),
	.w4(32'h3b7b36a8),
	.w5(32'h3c003e23),
	.w6(32'hbb624df8),
	.w7(32'hbb27cf77),
	.w8(32'h3ba01aa9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba1867),
	.w1(32'h39b10299),
	.w2(32'h3b1b444f),
	.w3(32'h3bcc6bee),
	.w4(32'hbb01c639),
	.w5(32'h3bfd02f6),
	.w6(32'h3c1e5e34),
	.w7(32'h3c696143),
	.w8(32'h3c4ac805),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9880593),
	.w1(32'hbb656013),
	.w2(32'hbbdaf6af),
	.w3(32'h3c3b528c),
	.w4(32'h3ba0f06c),
	.w5(32'hba8d0429),
	.w6(32'h3c482e29),
	.w7(32'h3bfe5de5),
	.w8(32'h3a90bcc3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd7517),
	.w1(32'hbbf9b12e),
	.w2(32'hbb8b6717),
	.w3(32'h3b28e56b),
	.w4(32'h3b28f64d),
	.w5(32'hbb883d89),
	.w6(32'h3bd729e4),
	.w7(32'hbb279d9b),
	.w8(32'hbc384b5c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0614b4),
	.w1(32'hbbba8e01),
	.w2(32'hbaac63ac),
	.w3(32'h3b04ace8),
	.w4(32'h3b28086b),
	.w5(32'h3bc885c7),
	.w6(32'hbc0d6103),
	.w7(32'hbc0599b8),
	.w8(32'h3c1304cf),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc125642),
	.w1(32'hbb9bfccb),
	.w2(32'hbb801135),
	.w3(32'h3b9924ce),
	.w4(32'h3b3d37c5),
	.w5(32'hbb67ac7b),
	.w6(32'h3c1bd3d3),
	.w7(32'h3c291cb0),
	.w8(32'hb95d78c5),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ee68b),
	.w1(32'hb9363ead),
	.w2(32'h3b369c55),
	.w3(32'h3b977d60),
	.w4(32'hbb0864e3),
	.w5(32'h3b830ff1),
	.w6(32'h3bfa2a6f),
	.w7(32'h3b3d415d),
	.w8(32'h3adf3ccd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff8d4e),
	.w1(32'hb9e42329),
	.w2(32'h3b26b4ad),
	.w3(32'h3b35b54c),
	.w4(32'h3a9ee5a2),
	.w5(32'h3bb5bf2e),
	.w6(32'h3a8f5d1a),
	.w7(32'h3aa4735b),
	.w8(32'h3b87ec09),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb077e2),
	.w1(32'h3c1ebe8c),
	.w2(32'hbc06a9b5),
	.w3(32'h3c20e002),
	.w4(32'h3b70d9a2),
	.w5(32'hbc04fa9b),
	.w6(32'h3c3099f6),
	.w7(32'h3b1c6a3d),
	.w8(32'hbc76f21a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fccca),
	.w1(32'hbbdad8d0),
	.w2(32'hbb2233fd),
	.w3(32'hbc962282),
	.w4(32'hbc7104d3),
	.w5(32'hbb7ab779),
	.w6(32'hbc803339),
	.w7(32'hbc818220),
	.w8(32'hbb72c4e5),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a1da0),
	.w1(32'h3a525c4b),
	.w2(32'hbaecd980),
	.w3(32'h3a4c970d),
	.w4(32'h3b53b0e7),
	.w5(32'h37b26966),
	.w6(32'hbb3619fa),
	.w7(32'h3b6270e8),
	.w8(32'h3b5e09d5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1761f6),
	.w1(32'hbb82e736),
	.w2(32'hb9b08517),
	.w3(32'hbae93778),
	.w4(32'hbb4d20d1),
	.w5(32'hba13903e),
	.w6(32'h3a058cef),
	.w7(32'hb9803e49),
	.w8(32'hbb998b64),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29d19c),
	.w1(32'hbaf2627e),
	.w2(32'hba537129),
	.w3(32'h39859d1b),
	.w4(32'h39fcc29d),
	.w5(32'hbb175a74),
	.w6(32'hbb302832),
	.w7(32'hbbb94f09),
	.w8(32'hbb8a5016),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab515ec),
	.w1(32'hbb83d6cc),
	.w2(32'hbbb5a329),
	.w3(32'hbb7bacb6),
	.w4(32'hbb82ae65),
	.w5(32'hbbc78e1b),
	.w6(32'hbb972b68),
	.w7(32'hbb937169),
	.w8(32'hb9b0560e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaec6f2),
	.w1(32'hbc31d9b5),
	.w2(32'hbc0c7d41),
	.w3(32'hbc04afea),
	.w4(32'hbb638b32),
	.w5(32'hbc318173),
	.w6(32'hbb728dcd),
	.w7(32'hbbabeb59),
	.w8(32'hbcc72d92),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c53c0),
	.w1(32'hbc11edc8),
	.w2(32'h3c27e326),
	.w3(32'hbc838fd7),
	.w4(32'hbc6a39ca),
	.w5(32'h3c245469),
	.w6(32'hbcaf81d1),
	.w7(32'hbc8c8c08),
	.w8(32'h3c70d6c2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c964ec1),
	.w1(32'h3c71b9b0),
	.w2(32'hba2bef61),
	.w3(32'h3c953352),
	.w4(32'h3c481c6f),
	.w5(32'h3b090ceb),
	.w6(32'h3cdb83e3),
	.w7(32'h3c759485),
	.w8(32'h3b99f283),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa59ba1),
	.w1(32'hbb00104a),
	.w2(32'h3b5ee675),
	.w3(32'hba58640e),
	.w4(32'hbb292081),
	.w5(32'h3b81acd3),
	.w6(32'h3ad0bdec),
	.w7(32'hba8ceaa7),
	.w8(32'hbc21459e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c9792),
	.w1(32'h3acbe3cb),
	.w2(32'h3ad78c3b),
	.w3(32'h3b78d82f),
	.w4(32'h3b6b34ef),
	.w5(32'h3a53e7c8),
	.w6(32'hbc227d58),
	.w7(32'hbbd9b438),
	.w8(32'hbb4384f8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba887d46),
	.w1(32'hba91e27e),
	.w2(32'hbb6b62f7),
	.w3(32'hbb88685e),
	.w4(32'h3a9a32fe),
	.w5(32'hbb7e52de),
	.w6(32'hbbc19af0),
	.w7(32'hbabc0319),
	.w8(32'hbc39bb9c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a50ed),
	.w1(32'hbcade1a0),
	.w2(32'hb979ff75),
	.w3(32'hbc4135e0),
	.w4(32'hbc61f022),
	.w5(32'h3b46a9bc),
	.w6(32'hbc0dd42d),
	.w7(32'hbc4a7e36),
	.w8(32'hbaaf4da4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e709),
	.w1(32'hbba39e8f),
	.w2(32'hbb899faf),
	.w3(32'h3b3c6d7b),
	.w4(32'hba51d0c3),
	.w5(32'hbb9acf6d),
	.w6(32'h3a25246a),
	.w7(32'hbb053633),
	.w8(32'hbc53f5c5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba122b4),
	.w1(32'h3b327eb8),
	.w2(32'h3c25b2fd),
	.w3(32'hbc3203ac),
	.w4(32'hbb07cd4c),
	.w5(32'h3b8a049f),
	.w6(32'hbc3aea04),
	.w7(32'h3b7fa2f1),
	.w8(32'h3b55cd2a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c339594),
	.w1(32'h3c111820),
	.w2(32'h3a935ebb),
	.w3(32'h3c212d95),
	.w4(32'h3b83e1bc),
	.w5(32'hba98e75d),
	.w6(32'h3c07d4a0),
	.w7(32'h3a9a9daf),
	.w8(32'hbb04aec3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b4ded),
	.w1(32'hbad628d5),
	.w2(32'hbb88284d),
	.w3(32'hbb36d021),
	.w4(32'hbb098bfb),
	.w5(32'hba6d64b9),
	.w6(32'hbbc098c1),
	.w7(32'hbaef1020),
	.w8(32'hbacddee4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926e0a),
	.w1(32'hbb3409db),
	.w2(32'hb9c38ddb),
	.w3(32'hbb2c103e),
	.w4(32'hbb777b0d),
	.w5(32'h3b43a4d2),
	.w6(32'hbb868d1b),
	.w7(32'hbbe9d005),
	.w8(32'hba312d0c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f1f47),
	.w1(32'h3b2c8ef4),
	.w2(32'hbace04df),
	.w3(32'hb982e4f4),
	.w4(32'h3c3711ec),
	.w5(32'hbb2bb544),
	.w6(32'hbacf5c20),
	.w7(32'h3b395c35),
	.w8(32'hb9f081d5),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a515a),
	.w1(32'hbb384aa5),
	.w2(32'hba4ad5d8),
	.w3(32'hbb2a5b34),
	.w4(32'hbb519316),
	.w5(32'h3b9e2276),
	.w6(32'hbbb8c059),
	.w7(32'hbafd8cce),
	.w8(32'hbab2d2d2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d0390),
	.w1(32'hbb1362f1),
	.w2(32'hbc120420),
	.w3(32'h3bf48719),
	.w4(32'h3b6cf01b),
	.w5(32'h3c16c5a9),
	.w6(32'h3bc1be74),
	.w7(32'hbb0334ee),
	.w8(32'h3c1c7bd7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc051e9a),
	.w1(32'h3abf9206),
	.w2(32'hb9a6ab3e),
	.w3(32'h3bc39bea),
	.w4(32'h3abe93a5),
	.w5(32'hbaa34f39),
	.w6(32'h3c75fc0d),
	.w7(32'h3c052761),
	.w8(32'h3b709bd0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d020b),
	.w1(32'hba0c1393),
	.w2(32'h3b3297fa),
	.w3(32'hbbb7b6f5),
	.w4(32'hbbcb76c8),
	.w5(32'h3b74655a),
	.w6(32'h3ba403fc),
	.w7(32'h3bcf6846),
	.w8(32'h3aca6e12),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b821e8c),
	.w1(32'hba4fd98c),
	.w2(32'hbc104362),
	.w3(32'h3b5fbe2b),
	.w4(32'h3a451f42),
	.w5(32'hbb99561e),
	.w6(32'h3b04002f),
	.w7(32'h3b97e8c5),
	.w8(32'hbbc19b16),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9cc6b),
	.w1(32'hbb85efa5),
	.w2(32'hbb5f6019),
	.w3(32'hbb3a027e),
	.w4(32'hbbadbbe5),
	.w5(32'hbc105e1d),
	.w6(32'hbc8ba5a0),
	.w7(32'hbc1910e6),
	.w8(32'hbc3bbfb8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c474da2),
	.w1(32'h3c65c33f),
	.w2(32'hba13539b),
	.w3(32'h3bbc21f0),
	.w4(32'h3cb7bd03),
	.w5(32'h3b6427c2),
	.w6(32'hbba7966f),
	.w7(32'h3c320705),
	.w8(32'h3c4a0033),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d61ba),
	.w1(32'h3b0ebbb0),
	.w2(32'hbab2bc06),
	.w3(32'hbbe59597),
	.w4(32'hbb381d7c),
	.w5(32'hbc037cf7),
	.w6(32'h3b960854),
	.w7(32'hbb04a9f5),
	.w8(32'hbb432bbf),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7366a3),
	.w1(32'h3b94f8bc),
	.w2(32'hbbd6262e),
	.w3(32'hbc904778),
	.w4(32'hbc128c8c),
	.w5(32'hbbb3c428),
	.w6(32'hbc32b467),
	.w7(32'hbc80e89e),
	.w8(32'h3b94ed27),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafe75c),
	.w1(32'h3bac7dcb),
	.w2(32'hbbda1998),
	.w3(32'hbc2afe42),
	.w4(32'hbb818b13),
	.w5(32'hbba39be1),
	.w6(32'hbacf6eb0),
	.w7(32'hbb687557),
	.w8(32'hbaf1a2b4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15b3e1),
	.w1(32'hbac4f738),
	.w2(32'hbc2cba16),
	.w3(32'hbbcaa8e9),
	.w4(32'h39452cd2),
	.w5(32'hbb0b764d),
	.w6(32'hbb257c1c),
	.w7(32'h3b9075ac),
	.w8(32'h3b9518c5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0f558),
	.w1(32'h39f00652),
	.w2(32'hbc3e7829),
	.w3(32'hbc2f79f1),
	.w4(32'hbbd74051),
	.w5(32'hbc8f63b4),
	.w6(32'h3b2a92fd),
	.w7(32'hbb9e2d82),
	.w8(32'h3b6dce5c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4541de),
	.w1(32'h3c371968),
	.w2(32'h3c512492),
	.w3(32'hbd1a90d2),
	.w4(32'hbb9f865e),
	.w5(32'h3bf5e8db),
	.w6(32'hbc9d880e),
	.w7(32'hbbb5f026),
	.w8(32'hbca2512f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc7a33e),
	.w1(32'hbc9f515a),
	.w2(32'hbbcba371),
	.w3(32'h3d62bf0f),
	.w4(32'h3c895442),
	.w5(32'hbb4c1ae7),
	.w6(32'h3cf43fe0),
	.w7(32'h3d11d7cd),
	.w8(32'hbbbdc5d6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a381b),
	.w1(32'hbc05aaa5),
	.w2(32'hbbd87905),
	.w3(32'hbb9117e0),
	.w4(32'hbc0021c7),
	.w5(32'hbcbd11c5),
	.w6(32'hbb7f14d4),
	.w7(32'h3ad51128),
	.w8(32'hbc84f95c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c900e14),
	.w1(32'h3ccba281),
	.w2(32'hbb57db8d),
	.w3(32'hbb97f042),
	.w4(32'h3d09c1bc),
	.w5(32'hbc22baf0),
	.w6(32'hbcfd207a),
	.w7(32'hbb782346),
	.w8(32'hbb83ae3b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43c3cd),
	.w1(32'hbc62fae3),
	.w2(32'hbbebdf4b),
	.w3(32'hbc04e3e4),
	.w4(32'h3ab17833),
	.w5(32'hbb2b5d98),
	.w6(32'hbc243a93),
	.w7(32'hbbae13ca),
	.w8(32'h3ad95efe),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb931209),
	.w1(32'h3b92cf5f),
	.w2(32'hbb8331a6),
	.w3(32'hbbac6d41),
	.w4(32'hbaa0522f),
	.w5(32'hbb43c20d),
	.w6(32'h3a8ee761),
	.w7(32'hbb5b8fe7),
	.w8(32'hbaecd01f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94efa9),
	.w1(32'hbbdd3fa9),
	.w2(32'hbc07e472),
	.w3(32'hbbe55b12),
	.w4(32'hbb9cb460),
	.w5(32'hbb137a39),
	.w6(32'hbb773e8e),
	.w7(32'hbc1f4de3),
	.w8(32'hbbbf56d0),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194b75),
	.w1(32'hbb4fe130),
	.w2(32'h398eb723),
	.w3(32'hbb751dbd),
	.w4(32'hbc4ab2e1),
	.w5(32'h3c34ec24),
	.w6(32'h3adb105f),
	.w7(32'hbc9c65ae),
	.w8(32'h3b62f6e3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ac60a),
	.w1(32'hbc8984de),
	.w2(32'hba8288ee),
	.w3(32'h3af988dd),
	.w4(32'hbbf9a6a0),
	.w5(32'hbcdd8953),
	.w6(32'h3bc287a4),
	.w7(32'hbb617238),
	.w8(32'hbcd78002),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42bbfc),
	.w1(32'h3c6822ec),
	.w2(32'h398482c7),
	.w3(32'hbb3fd044),
	.w4(32'h3c982d55),
	.w5(32'h3a0eec7d),
	.w6(32'hbcfb89d1),
	.w7(32'hbba33609),
	.w8(32'h3b372920),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf5dbf),
	.w1(32'h3bb79d89),
	.w2(32'hbc0101ee),
	.w3(32'h3a2e1d8f),
	.w4(32'h3b8db3ce),
	.w5(32'hbc3b2e70),
	.w6(32'h3bbd15af),
	.w7(32'h3b4590b5),
	.w8(32'hbbde1d22),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd092c5),
	.w1(32'hbc85f12f),
	.w2(32'hbb028257),
	.w3(32'hbc22dfb5),
	.w4(32'h3958d230),
	.w5(32'hbb90b113),
	.w6(32'hbc50f36a),
	.w7(32'hbb92aba8),
	.w8(32'hbb7b2258),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba53004),
	.w1(32'hbb9b07a2),
	.w2(32'hbc3b7b11),
	.w3(32'hbc3eb2df),
	.w4(32'hbbb535d0),
	.w5(32'hbb09aef1),
	.w6(32'hbb9df818),
	.w7(32'hbbd833bd),
	.w8(32'h3b3661e7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae19e30),
	.w1(32'h3c2141a9),
	.w2(32'hbb6b106f),
	.w3(32'hbc76f146),
	.w4(32'hbc173282),
	.w5(32'hbbf9dfbd),
	.w6(32'hbb125f65),
	.w7(32'hbb48cad7),
	.w8(32'hbc07539f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc8b21),
	.w1(32'hbba11026),
	.w2(32'h39d39459),
	.w3(32'hbc8662c1),
	.w4(32'hbbf4e0ae),
	.w5(32'h3c2d3e9e),
	.w6(32'hbc01fc07),
	.w7(32'hbb98e591),
	.w8(32'h3c245fa6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadabb3),
	.w1(32'hbc4a9d4c),
	.w2(32'h3b67f9f1),
	.w3(32'h3a71d326),
	.w4(32'hbc85866f),
	.w5(32'h3c315496),
	.w6(32'h3bb8a497),
	.w7(32'hbbecac56),
	.w8(32'h3af4ad16),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c475b),
	.w1(32'hbc0e48d5),
	.w2(32'h3bc3b178),
	.w3(32'h3c5e21ad),
	.w4(32'h3c133147),
	.w5(32'h3bdaad48),
	.w6(32'h3be6affb),
	.w7(32'h3c3c29d1),
	.w8(32'h3ab84c42),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30383f),
	.w1(32'hbc70e808),
	.w2(32'hbca985c6),
	.w3(32'hba8d7457),
	.w4(32'hbc1987df),
	.w5(32'hbc4eaa22),
	.w6(32'hbb978a50),
	.w7(32'hbae49e7c),
	.w8(32'h3bbeae4a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba078456),
	.w1(32'h3ccb5a33),
	.w2(32'h3b30605e),
	.w3(32'hbcaf31ae),
	.w4(32'h3ad2309f),
	.w5(32'h3c114824),
	.w6(32'hbc961e14),
	.w7(32'hbc4a220f),
	.w8(32'hbafdb36b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf18a4d),
	.w1(32'hbc09f8de),
	.w2(32'h3a4a55b2),
	.w3(32'h3c030b6e),
	.w4(32'h39e12953),
	.w5(32'hb7c382e4),
	.w6(32'h3c80dcba),
	.w7(32'h3c837037),
	.w8(32'h3c1835f1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba553edf),
	.w1(32'hbb1c2800),
	.w2(32'hbba3a2f7),
	.w3(32'hbb78d50d),
	.w4(32'hbbaf7963),
	.w5(32'hbc868245),
	.w6(32'h3c8bda87),
	.w7(32'h3c097801),
	.w8(32'hbc0127a1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97952d),
	.w1(32'h3c7456ee),
	.w2(32'hbb557b89),
	.w3(32'hbb187b51),
	.w4(32'h3c901e6d),
	.w5(32'hbc257762),
	.w6(32'hbc6f9a11),
	.w7(32'h3b4bdd6a),
	.w8(32'hbcda29c3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98f4e5),
	.w1(32'hba306035),
	.w2(32'h3b2ef6f2),
	.w3(32'h3cff48a3),
	.w4(32'h3cec86f6),
	.w5(32'h3c1d82a1),
	.w6(32'hbb2c804f),
	.w7(32'h3c9df8f0),
	.w8(32'h3b89ca5f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cdbdc),
	.w1(32'hbc79bcf1),
	.w2(32'h3bb0fc56),
	.w3(32'hbbaab5c7),
	.w4(32'hbca860db),
	.w5(32'hbb8f98c0),
	.w6(32'h3c9e88ed),
	.w7(32'h3b89b1d2),
	.w8(32'h3b114670),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be77b4b),
	.w1(32'h3a7ee34f),
	.w2(32'hbbf2321c),
	.w3(32'h3b7d1c16),
	.w4(32'h3b6b861b),
	.w5(32'h3b477a40),
	.w6(32'h3acb5017),
	.w7(32'h3b5fd09d),
	.w8(32'h39f0ddc4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e701f),
	.w1(32'h3bc93719),
	.w2(32'h3b958825),
	.w3(32'h39ae3b53),
	.w4(32'h3bd41c82),
	.w5(32'h3bfc644b),
	.w6(32'hba830172),
	.w7(32'h38ea859e),
	.w8(32'h3a3fee8e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba360ccc),
	.w1(32'h3b84fc10),
	.w2(32'hbb79c121),
	.w3(32'h3b6326c1),
	.w4(32'h3bf36e33),
	.w5(32'h3bf70d73),
	.w6(32'hbb1e81ee),
	.w7(32'h3b2bb9c2),
	.w8(32'h3bf6473c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75597b),
	.w1(32'hbcd192eb),
	.w2(32'hbc216aa5),
	.w3(32'h38cb535e),
	.w4(32'hbc948ed7),
	.w5(32'hba0a0770),
	.w6(32'h3c4c9b1f),
	.w7(32'hbb9d9cd2),
	.w8(32'h3bcde8bc),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8c91b),
	.w1(32'h3a11956d),
	.w2(32'hbc557b30),
	.w3(32'hbba479f7),
	.w4(32'hbb3cf81b),
	.w5(32'hbbbfa669),
	.w6(32'h3b1b2de2),
	.w7(32'hbbb3ac41),
	.w8(32'h3ada6649),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8e1e4),
	.w1(32'h3b9ccaeb),
	.w2(32'hbae78c30),
	.w3(32'hbc67b68f),
	.w4(32'hbb974bdf),
	.w5(32'h3af4e8b2),
	.w6(32'hbc146f22),
	.w7(32'h3a73af3e),
	.w8(32'h3ab0499f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4726a6),
	.w1(32'h3a57f57a),
	.w2(32'h3b8865d3),
	.w3(32'h3b4cf52c),
	.w4(32'h3a978e9a),
	.w5(32'h3b8d1212),
	.w6(32'hb8ecd595),
	.w7(32'hbaf38720),
	.w8(32'h3ab3350b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c515ce7),
	.w1(32'h3b678d9e),
	.w2(32'hbbd48864),
	.w3(32'h3c8e3b7f),
	.w4(32'h3c11ef85),
	.w5(32'hbca50929),
	.w6(32'h3c6b0421),
	.w7(32'h3c5c8c45),
	.w8(32'hbbe5982d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb6f743),
	.w1(32'h3c8640fd),
	.w2(32'h3c13b2b4),
	.w3(32'h3bd8c8fb),
	.w4(32'h3c82e693),
	.w5(32'h3c8b6faf),
	.w6(32'hbca454ef),
	.w7(32'hbac38a9e),
	.w8(32'h3bbfb905),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc854261),
	.w1(32'hbcccbdb7),
	.w2(32'hbc3582a7),
	.w3(32'h3c45ae13),
	.w4(32'hbca3f0d4),
	.w5(32'hbba3c6b9),
	.w6(32'h3c884756),
	.w7(32'h3be43dbe),
	.w8(32'hbac43057),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71f951),
	.w1(32'hbc94607b),
	.w2(32'hbc162c89),
	.w3(32'hbc444e35),
	.w4(32'hbc43973f),
	.w5(32'hbc1820bb),
	.w6(32'hbc5592f4),
	.w7(32'hbbeca6a8),
	.w8(32'hbb30c3d5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc239943),
	.w1(32'hbb8cd9ea),
	.w2(32'h3a854ecd),
	.w3(32'hbc925006),
	.w4(32'hba227cfa),
	.w5(32'h3a53149b),
	.w6(32'hbc72d690),
	.w7(32'hbc2297b3),
	.w8(32'h3b7b687e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29f301),
	.w1(32'h3b55fc5e),
	.w2(32'hbc13cfc6),
	.w3(32'hbb5fd0c2),
	.w4(32'hba00a127),
	.w5(32'hbc05d20f),
	.w6(32'h39f268fc),
	.w7(32'h3b03b2a9),
	.w8(32'hbc0cd0e0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b39d6),
	.w1(32'h391153ea),
	.w2(32'hbac47b79),
	.w3(32'hbc5ed98a),
	.w4(32'hb9fad7aa),
	.w5(32'hba567464),
	.w6(32'hbbf4b0fd),
	.w7(32'hbba35931),
	.w8(32'hbb0f5ba3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab19a69),
	.w1(32'h38faf54d),
	.w2(32'hbbc823ae),
	.w3(32'hbbcde6b4),
	.w4(32'hbb57514f),
	.w5(32'h3af844ae),
	.w6(32'hbbbf417e),
	.w7(32'h3a7b6269),
	.w8(32'hbb8e4e05),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb7a12),
	.w1(32'hbb525e54),
	.w2(32'h3c04e1fe),
	.w3(32'hbc589134),
	.w4(32'hbc4c33af),
	.w5(32'hbc2d6772),
	.w6(32'hbc648dbe),
	.w7(32'hbb7c190d),
	.w8(32'hbc43304b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09b16d),
	.w1(32'h3bffbc6b),
	.w2(32'h3aa7b436),
	.w3(32'h3c81eabc),
	.w4(32'h3c2867a3),
	.w5(32'h3be45109),
	.w6(32'hbbbcaf78),
	.w7(32'h3b5aae54),
	.w8(32'hba8e503d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd06dec),
	.w1(32'hba72aed0),
	.w2(32'h3b8841fa),
	.w3(32'h3c2ec359),
	.w4(32'h3bcb9fd6),
	.w5(32'hbc6cceab),
	.w6(32'h3b61e260),
	.w7(32'hba353133),
	.w8(32'hbc371d7a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca01bff),
	.w1(32'h3cb01470),
	.w2(32'hbb11d4cc),
	.w3(32'h3a97dd51),
	.w4(32'h3c4c862a),
	.w5(32'h3b3a5f31),
	.w6(32'hbc963865),
	.w7(32'hbb6d3518),
	.w8(32'hb9d9fafa),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce0282),
	.w1(32'hbb3eeecc),
	.w2(32'h3a572eb3),
	.w3(32'h3b6d7943),
	.w4(32'hbb2fad20),
	.w5(32'hbbe1a101),
	.w6(32'h3b1659c2),
	.w7(32'hbb906ff7),
	.w8(32'hbaf5b8de),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2d5a2),
	.w1(32'hbbd393f1),
	.w2(32'h3c40e834),
	.w3(32'hbc02498b),
	.w4(32'hbc1a9d7c),
	.w5(32'h3c6b313f),
	.w6(32'hbc6cb446),
	.w7(32'h3b893c79),
	.w8(32'h3ca25611),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b5a6f),
	.w1(32'hbcd9a8ba),
	.w2(32'h3b869697),
	.w3(32'h3c465f87),
	.w4(32'hbcc0532e),
	.w5(32'hbbccd780),
	.w6(32'h3cbd150a),
	.w7(32'h3b32f7cb),
	.w8(32'hbbf682d1),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83ebb5),
	.w1(32'hbb862b74),
	.w2(32'h3a89402c),
	.w3(32'hbc2f9fec),
	.w4(32'hbc29e59d),
	.w5(32'h3a60ceb1),
	.w6(32'hbbafe30f),
	.w7(32'hbc1419f5),
	.w8(32'hbb0f8f78),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd64dc6),
	.w1(32'hbba70864),
	.w2(32'h3b79792b),
	.w3(32'hbb4ef5ca),
	.w4(32'hbb9fe3e3),
	.w5(32'h3becb4af),
	.w6(32'h39cd3241),
	.w7(32'hb93f1351),
	.w8(32'h3bcb553a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24f913),
	.w1(32'hbcce1847),
	.w2(32'hbb4258e2),
	.w3(32'h3ba44521),
	.w4(32'hbca12f3a),
	.w5(32'hbbdc356b),
	.w6(32'h3cbbb2d0),
	.w7(32'hb931d41b),
	.w8(32'hbbe6a6c7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e201),
	.w1(32'hbb374b8a),
	.w2(32'h3b337ecb),
	.w3(32'hbbfe7238),
	.w4(32'hbb7c9535),
	.w5(32'h3a109c7a),
	.w6(32'hbc05658f),
	.w7(32'hbb1b8290),
	.w8(32'h3bb6ccaa),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad58ce5),
	.w1(32'hbbccbe03),
	.w2(32'hbaaf002e),
	.w3(32'hbbfeed95),
	.w4(32'hbb86433c),
	.w5(32'h3c579646),
	.w6(32'h3b88250d),
	.w7(32'hbbd19757),
	.w8(32'h3c48a517),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59cfcb),
	.w1(32'hbca16e69),
	.w2(32'h3afb82be),
	.w3(32'h3b4b004d),
	.w4(32'hbcadf313),
	.w5(32'h3c696af1),
	.w6(32'h3bc1e680),
	.w7(32'hbba40afb),
	.w8(32'h3c6bcf7f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd37724),
	.w1(32'hbc54230f),
	.w2(32'hbc249457),
	.w3(32'h3bf355d7),
	.w4(32'hbc4c1123),
	.w5(32'hbbec5070),
	.w6(32'h3cad0505),
	.w7(32'hbaf06841),
	.w8(32'hbc2b7473),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa8250),
	.w1(32'hbc2745f8),
	.w2(32'h3a7ac23d),
	.w3(32'h3b1ebad6),
	.w4(32'hbbc553f5),
	.w5(32'hba478adc),
	.w6(32'h3b9e5391),
	.w7(32'hba883cb0),
	.w8(32'hbaa8e146),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f8ac4),
	.w1(32'h3b217296),
	.w2(32'h3a3f6a0f),
	.w3(32'hbadac27b),
	.w4(32'hba128787),
	.w5(32'hbabd09cd),
	.w6(32'hba01ebb0),
	.w7(32'h3b9e1a1f),
	.w8(32'hbba43f1c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe9da2),
	.w1(32'h3b516d17),
	.w2(32'h3be0cc7b),
	.w3(32'h3bf1f13b),
	.w4(32'h3bd7af6d),
	.w5(32'h3b76b8f3),
	.w6(32'h39103118),
	.w7(32'h3b9f0b46),
	.w8(32'h3b716cab),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e11f),
	.w1(32'hbaaceabe),
	.w2(32'h3b638b18),
	.w3(32'h3bd513e8),
	.w4(32'hbb6123d5),
	.w5(32'h3bf1da03),
	.w6(32'h3c01732b),
	.w7(32'h3aba261a),
	.w8(32'hbb2f45ce),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcde97),
	.w1(32'h3a9a2325),
	.w2(32'hbc1bf9fe),
	.w3(32'h3bc0741b),
	.w4(32'h3c0bb9aa),
	.w5(32'hbb211397),
	.w6(32'hbb7f40a6),
	.w7(32'h3af88f24),
	.w8(32'hbb5ebdb6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa15697),
	.w1(32'hba9f45c0),
	.w2(32'hba56506c),
	.w3(32'hbc0c1661),
	.w4(32'h3c26d62f),
	.w5(32'hbc14880d),
	.w6(32'hbc0cbe8f),
	.w7(32'h398adf23),
	.w8(32'hb9eab672),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12c3db),
	.w1(32'hbc63fc70),
	.w2(32'hbb29a9be),
	.w3(32'h39dc5ceb),
	.w4(32'hbabdeb1d),
	.w5(32'h39d97609),
	.w6(32'hbbac310d),
	.w7(32'h3b3b16ad),
	.w8(32'h3c29f49c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15059b),
	.w1(32'h3c250ab3),
	.w2(32'hbc31c7fc),
	.w3(32'hbc34e44a),
	.w4(32'h3b590691),
	.w5(32'hbc4888db),
	.w6(32'hbacb06db),
	.w7(32'hbb58b9cd),
	.w8(32'hbba33def),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35249b),
	.w1(32'h3ca3cf2d),
	.w2(32'hbc43d246),
	.w3(32'hbc4121a7),
	.w4(32'h3c61fc66),
	.w5(32'hbc1eaf1c),
	.w6(32'hbc9f709c),
	.w7(32'hbbe7eaab),
	.w8(32'h3b33d8d9),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a937a),
	.w1(32'h391929c0),
	.w2(32'hbc0eec61),
	.w3(32'hbcb0d4d0),
	.w4(32'hbbbd1cb7),
	.w5(32'hbc504de8),
	.w6(32'hbc11d839),
	.w7(32'hbbc19edd),
	.w8(32'hba32a188),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd1957),
	.w1(32'h3857e3f7),
	.w2(32'hbbe79207),
	.w3(32'hbc85471b),
	.w4(32'hbc1a1f7f),
	.w5(32'hbba184ba),
	.w6(32'hbc42b32f),
	.w7(32'hbc205871),
	.w8(32'h3c0b556d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3007c4),
	.w1(32'h3a7e65d6),
	.w2(32'h3bde8270),
	.w3(32'hbb4f2a49),
	.w4(32'h3ba692e7),
	.w5(32'h3ad192f0),
	.w6(32'h3c7f0290),
	.w7(32'h3c25376e),
	.w8(32'h3b51035f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bc292),
	.w1(32'h3b83a01e),
	.w2(32'h39b7d478),
	.w3(32'hbc210235),
	.w4(32'hbc51f2c7),
	.w5(32'hbbda6129),
	.w6(32'hbc6ca549),
	.w7(32'hbca1a567),
	.w8(32'hbb8fc4e9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf36217),
	.w1(32'h3c14b1f0),
	.w2(32'hbb56e924),
	.w3(32'hba985405),
	.w4(32'h3c22614c),
	.w5(32'h3b49661f),
	.w6(32'hbc5c3c32),
	.w7(32'hbbb94784),
	.w8(32'h3be1f79a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ae678),
	.w1(32'hbc4985cd),
	.w2(32'h3c0f9081),
	.w3(32'hbb508780),
	.w4(32'hbc11594a),
	.w5(32'h3c3a49ef),
	.w6(32'h3bc370c3),
	.w7(32'h3bbca8c0),
	.w8(32'h3b7d48c5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd9f97),
	.w1(32'hbb79efa1),
	.w2(32'h3abe843e),
	.w3(32'h3b918731),
	.w4(32'hbbe42096),
	.w5(32'hbc762c5d),
	.w6(32'h3b83d668),
	.w7(32'hbabe23ab),
	.w8(32'hbc255102),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b922332),
	.w1(32'h3c0ced9f),
	.w2(32'h3b118a4b),
	.w3(32'h3bbf6de2),
	.w4(32'h3c1018cb),
	.w5(32'h3bb82779),
	.w6(32'hbc6c1654),
	.w7(32'h3b9fd0fd),
	.w8(32'h3bea4c3d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18568e),
	.w1(32'hbb4554f7),
	.w2(32'hbc1e0dce),
	.w3(32'h3bcbcc49),
	.w4(32'h3b01db99),
	.w5(32'hbb254f2d),
	.w6(32'h39c2947e),
	.w7(32'h3c85a1c0),
	.w8(32'hb9f2d9f8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e5d2e),
	.w1(32'hbab2548f),
	.w2(32'hba105aa6),
	.w3(32'hbb55d0f5),
	.w4(32'hbb9e6ec8),
	.w5(32'hbbcfe46b),
	.w6(32'h3a91c6de),
	.w7(32'h3b35fd80),
	.w8(32'hbc41ae62),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64f6e1),
	.w1(32'hbc056514),
	.w2(32'hbc033f88),
	.w3(32'hba0327ce),
	.w4(32'hbc7ee7e1),
	.w5(32'hbc9280ef),
	.w6(32'hbb762c43),
	.w7(32'h3b06176b),
	.w8(32'hbc0542c0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b947af8),
	.w1(32'h3bc22393),
	.w2(32'hbc189302),
	.w3(32'hbc101301),
	.w4(32'h3bda4a72),
	.w5(32'hbb9fc577),
	.w6(32'hbca6252c),
	.w7(32'h3a80dbbe),
	.w8(32'hbc0c4eca),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c701),
	.w1(32'h3bd6cc0f),
	.w2(32'h3c136833),
	.w3(32'hbc1d533f),
	.w4(32'hbaa20a53),
	.w5(32'h3b20b9d6),
	.w6(32'hbc7cb4c9),
	.w7(32'hbbc92b91),
	.w8(32'h3c06dc08),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c015a7c),
	.w1(32'hbbd07f14),
	.w2(32'hbc1261d4),
	.w3(32'h3cacb977),
	.w4(32'h3c17c8ad),
	.w5(32'hbc5ddc09),
	.w6(32'h3c27a5dd),
	.w7(32'h3c955d73),
	.w8(32'h3bc03345),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d23d1),
	.w1(32'h3c03b968),
	.w2(32'hbba1a900),
	.w3(32'hbcac36e8),
	.w4(32'hbb7758bf),
	.w5(32'hbc5730ac),
	.w6(32'hbc970bae),
	.w7(32'hbc0802f3),
	.w8(32'hbc40754e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29db52),
	.w1(32'h3ca29723),
	.w2(32'hba6c0d56),
	.w3(32'h388f517f),
	.w4(32'h3c6727c0),
	.w5(32'h3c543621),
	.w6(32'hbc23a5bc),
	.w7(32'h3b201779),
	.w8(32'h3a9d854d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc270c94),
	.w1(32'hbc99024f),
	.w2(32'hbc0f99fb),
	.w3(32'h3c5e9056),
	.w4(32'hbc691100),
	.w5(32'hbbd096d5),
	.w6(32'h3c8cde13),
	.w7(32'h3b7c55af),
	.w8(32'hbb999f0b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03a314),
	.w1(32'h3c2ddeb5),
	.w2(32'hbb6d589e),
	.w3(32'hb7730cc4),
	.w4(32'h3c44cbe2),
	.w5(32'hbc181825),
	.w6(32'hbae5c510),
	.w7(32'h3c60aba7),
	.w8(32'hbc0b89f6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9acfa0),
	.w1(32'h3c3d84d3),
	.w2(32'hbb342df9),
	.w3(32'hbc4052b7),
	.w4(32'h3c2bf5a6),
	.w5(32'hbb1808f7),
	.w6(32'hbc18dc98),
	.w7(32'h39b47ebe),
	.w8(32'h3b84127a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9d35f),
	.w1(32'h3bf84260),
	.w2(32'h3b20c766),
	.w3(32'hbbdcf8d1),
	.w4(32'h3682406b),
	.w5(32'h3bf6a03d),
	.w6(32'hbc21273a),
	.w7(32'hbc27dc7f),
	.w8(32'h3c11afd4),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b853c7f),
	.w1(32'h3aaf5827),
	.w2(32'h3b5fc805),
	.w3(32'h3bf89d85),
	.w4(32'h3bc2b094),
	.w5(32'h3a853331),
	.w6(32'hbada2780),
	.w7(32'hba935f97),
	.w8(32'h3831607a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18e850),
	.w1(32'h3b17bbb1),
	.w2(32'hba246352),
	.w3(32'hbab04ce5),
	.w4(32'h39fc806d),
	.w5(32'hbb0197e9),
	.w6(32'h3a3160ba),
	.w7(32'h3b234cb5),
	.w8(32'hbaff6f6d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba656f3d),
	.w1(32'hba8441c4),
	.w2(32'h3c09a0dc),
	.w3(32'hbb2e88f8),
	.w4(32'hba46ffd9),
	.w5(32'h3d0fa05c),
	.w6(32'hbb96995e),
	.w7(32'h392c959c),
	.w8(32'h3c8a3bf1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3ab7e),
	.w1(32'hbd18d79a),
	.w2(32'hba36f49b),
	.w3(32'h3caef38d),
	.w4(32'hbc6ca365),
	.w5(32'h3bda3b9c),
	.w6(32'h3d228060),
	.w7(32'h3cacc589),
	.w8(32'h3bf7e105),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae04fd0),
	.w1(32'hbb9c4be2),
	.w2(32'h3badf96e),
	.w3(32'h3c2d5709),
	.w4(32'h3a70e686),
	.w5(32'h3bb3b16f),
	.w6(32'h3c769178),
	.w7(32'h3c176595),
	.w8(32'h3b94d291),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68c80d),
	.w1(32'hba113eb9),
	.w2(32'hbae88f2a),
	.w3(32'h3b9261c5),
	.w4(32'hbaa22ad4),
	.w5(32'hbb7a1853),
	.w6(32'h3ac5d548),
	.w7(32'hbb802d5c),
	.w8(32'hbb964e89),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc977af7),
	.w1(32'hbbd86dc4),
	.w2(32'hbc40ca1d),
	.w3(32'hbcc4580f),
	.w4(32'hbc88569e),
	.w5(32'hbc94b66d),
	.w6(32'hbc9135b2),
	.w7(32'hbcc78edd),
	.w8(32'hbc241b75),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc891a9a),
	.w1(32'hbbe172f2),
	.w2(32'h3b9ff88d),
	.w3(32'hbcc01ce7),
	.w4(32'hbc66b41b),
	.w5(32'h3c4f3fb7),
	.w6(32'hbca37fba),
	.w7(32'hbc4a36ab),
	.w8(32'h3c61401d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule