module layer_10_featuremap_287(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c06b2),
	.w1(32'h3a82d98d),
	.w2(32'h3a8a1968),
	.w3(32'h398e23ed),
	.w4(32'h39c5b367),
	.w5(32'h3915723d),
	.w6(32'h3a198e0b),
	.w7(32'h3a3c8bdd),
	.w8(32'h3736bbe8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6da0550),
	.w1(32'h39780414),
	.w2(32'h38ecd8be),
	.w3(32'h389b6772),
	.w4(32'h388b85ed),
	.w5(32'hb86588a7),
	.w6(32'h360c56d2),
	.w7(32'h3944cc71),
	.w8(32'hb8e8b8aa),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9483402),
	.w1(32'hba575426),
	.w2(32'hba845db0),
	.w3(32'hb9c5c64b),
	.w4(32'hb99a836a),
	.w5(32'h39566e38),
	.w6(32'hba2032a2),
	.w7(32'hba6d6922),
	.w8(32'h3900b0c9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a3c25),
	.w1(32'h38c8bd1a),
	.w2(32'h38b0b1e6),
	.w3(32'h399d18f4),
	.w4(32'h39b26bb2),
	.w5(32'hbacb0b2e),
	.w6(32'h37108964),
	.w7(32'h38ee2858),
	.w8(32'hbacdfa94),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74274c),
	.w1(32'hba1d38e1),
	.w2(32'hb90a34bf),
	.w3(32'hbaa7fa56),
	.w4(32'hba4cf3b6),
	.w5(32'hb9705246),
	.w6(32'hbab34647),
	.w7(32'hba6dbaec),
	.w8(32'h388bbd7b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c7b98),
	.w1(32'h39adac93),
	.w2(32'h3a0bda4f),
	.w3(32'hb8d657c2),
	.w4(32'h379b9120),
	.w5(32'hb9ea09d3),
	.w6(32'h38a107bc),
	.w7(32'h39968a83),
	.w8(32'hb9cc8c69),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2ea2f),
	.w1(32'hb944ead7),
	.w2(32'hb91d5246),
	.w3(32'hb9ab3e97),
	.w4(32'hb9aabf67),
	.w5(32'hba23d8dd),
	.w6(32'hb9ceccb4),
	.w7(32'h38748f9a),
	.w8(32'hba11a182),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9925479),
	.w1(32'hba051ddc),
	.w2(32'hba7c264c),
	.w3(32'hba86c34b),
	.w4(32'hba3a28be),
	.w5(32'h3a1e6fd3),
	.w6(32'hba623eb2),
	.w7(32'hba7c60de),
	.w8(32'h3a29481c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20cfb2),
	.w1(32'h3a1dcd9f),
	.w2(32'h3a3063f0),
	.w3(32'h39adb8b3),
	.w4(32'h39e27d1f),
	.w5(32'hb82bae85),
	.w6(32'h398eb5c6),
	.w7(32'h3a04b690),
	.w8(32'h393f58a3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996ca72),
	.w1(32'h3a1a74f6),
	.w2(32'h3a41f8c9),
	.w3(32'h374859ba),
	.w4(32'h39fd929d),
	.w5(32'hba03674b),
	.w6(32'h3925c5c8),
	.w7(32'h3a2b2394),
	.w8(32'hb97587f1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf12db),
	.w1(32'hb8a1e09e),
	.w2(32'h38c5803a),
	.w3(32'hb917b84d),
	.w4(32'hb887c4f0),
	.w5(32'hba3366fb),
	.w6(32'h387f0497),
	.w7(32'h392196bf),
	.w8(32'hb892b307),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe4e4b),
	.w1(32'hb94de2b3),
	.w2(32'hb9120769),
	.w3(32'hb97fcf8a),
	.w4(32'hb9af770e),
	.w5(32'h391f1403),
	.w6(32'h3762218b),
	.w7(32'hb8314b16),
	.w8(32'h38f38bcb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cd17d),
	.w1(32'h39732adb),
	.w2(32'h39b82e2a),
	.w3(32'h390d95d4),
	.w4(32'h3a043ffd),
	.w5(32'hba3e5dde),
	.w6(32'h39609af5),
	.w7(32'h39c835a6),
	.w8(32'hba83daae),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bcda1),
	.w1(32'hba87d7b6),
	.w2(32'hb9b08061),
	.w3(32'hba6db9fa),
	.w4(32'hb9e520cf),
	.w5(32'h3a0b0781),
	.w6(32'hbaf119a6),
	.w7(32'hba95c665),
	.w8(32'h3a03ee88),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c18543),
	.w1(32'h39620eb1),
	.w2(32'hb6a4442a),
	.w3(32'h3a1e3eaa),
	.w4(32'h39f60538),
	.w5(32'h39dfc727),
	.w6(32'h39a87a07),
	.w7(32'h39eb403f),
	.w8(32'h38870e8c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392791ab),
	.w1(32'h3a11fb40),
	.w2(32'h3aabee28),
	.w3(32'h3a66ee82),
	.w4(32'h3af4bcf2),
	.w5(32'h39ef9f66),
	.w6(32'h398de198),
	.w7(32'h3ad0424c),
	.w8(32'h3a26e43e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a530365),
	.w1(32'h3a1d98f4),
	.w2(32'h39da12d4),
	.w3(32'h3856821c),
	.w4(32'h3962c6d7),
	.w5(32'hba070df5),
	.w6(32'hb6e8c7c6),
	.w7(32'h39749a6a),
	.w8(32'hba103e9e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37f35f),
	.w1(32'hb98d2ad9),
	.w2(32'h3904a8cf),
	.w3(32'hb9ae2d9b),
	.w4(32'h380bd02c),
	.w5(32'hb97da101),
	.w6(32'h37b237e3),
	.w7(32'h39b956eb),
	.w8(32'hb9f412d4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66c1cd),
	.w1(32'hba9f6a46),
	.w2(32'hba1c6184),
	.w3(32'hb9b72ed7),
	.w4(32'hb9a75fca),
	.w5(32'h3a637c6e),
	.w6(32'hba8ced17),
	.w7(32'hba023881),
	.w8(32'h3ac19594),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af92061),
	.w1(32'h3acbbf70),
	.w2(32'h3a9d6b3b),
	.w3(32'h398622cc),
	.w4(32'h39edf2c0),
	.w5(32'h3a0c17ad),
	.w6(32'h3a85a8f5),
	.w7(32'h3a4ab441),
	.w8(32'h39e5a9a9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39817f31),
	.w1(32'hb9caed59),
	.w2(32'h39e68e22),
	.w3(32'h39100998),
	.w4(32'h3a562be2),
	.w5(32'h3a405c5a),
	.w6(32'hb9582bbb),
	.w7(32'h3a20b8f4),
	.w8(32'h3a4076ce),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b7d07),
	.w1(32'h39df0b92),
	.w2(32'h384e9356),
	.w3(32'h39d8ec82),
	.w4(32'h3887dcf4),
	.w5(32'h3a0d0216),
	.w6(32'h39cbeccd),
	.w7(32'hb7719777),
	.w8(32'h3a828f06),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ef56),
	.w1(32'h3b070544),
	.w2(32'h3b160ca9),
	.w3(32'h3a9743e9),
	.w4(32'h3a989fef),
	.w5(32'hba82e3e5),
	.w6(32'h3a1d9f40),
	.w7(32'h3b1cb521),
	.w8(32'hbae874ae),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba198c4b),
	.w1(32'h3a211362),
	.w2(32'h3a1a8918),
	.w3(32'h39319c1d),
	.w4(32'h3a934b27),
	.w5(32'h3ad1672b),
	.w6(32'h391ed848),
	.w7(32'h3a8819e1),
	.w8(32'h3a7da848),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c0d3f),
	.w1(32'h3a8a92fe),
	.w2(32'h3a057bf0),
	.w3(32'h3b0c5cfa),
	.w4(32'h3b0de73e),
	.w5(32'h36a56b59),
	.w6(32'h3aabd1b4),
	.w7(32'h3aa714bb),
	.w8(32'hb85ce305),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a08a0e),
	.w1(32'hb77ffe3c),
	.w2(32'h393480d2),
	.w3(32'hb7d92c09),
	.w4(32'h3938a419),
	.w5(32'h3a07acfc),
	.w6(32'hb9c0009f),
	.w7(32'h38aeeece),
	.w8(32'h39b8e6b5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b3ba6),
	.w1(32'h383fb208),
	.w2(32'h39aeed4a),
	.w3(32'h39ef6d05),
	.w4(32'h3a2e291c),
	.w5(32'h388a9b11),
	.w6(32'hb8cca77c),
	.w7(32'h39acc389),
	.w8(32'h39853355),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27bf1c),
	.w1(32'h39e96db1),
	.w2(32'h3a52ff9a),
	.w3(32'hb73cb9ee),
	.w4(32'h39d55205),
	.w5(32'hba258041),
	.w6(32'h37fc32f4),
	.w7(32'h3a0bc1bb),
	.w8(32'hba0d1406),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ae3fb),
	.w1(32'h39b9ca35),
	.w2(32'h39f0c87c),
	.w3(32'h38ececd0),
	.w4(32'h3a024e59),
	.w5(32'hb8c6b497),
	.w6(32'hb8a7d93e),
	.w7(32'h392eda9f),
	.w8(32'hb98d73ad),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3887ffb5),
	.w1(32'h3995aace),
	.w2(32'h392e6b8c),
	.w3(32'h39d47bd3),
	.w4(32'h3a51d374),
	.w5(32'hb9e7569e),
	.w6(32'h39d5f561),
	.w7(32'h39ea0a0c),
	.w8(32'hb9c450a9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8811214),
	.w1(32'hb953676a),
	.w2(32'hb6e33438),
	.w3(32'hba288cf9),
	.w4(32'hba3d0cf9),
	.w5(32'hba933af5),
	.w6(32'hb8b54051),
	.w7(32'hb973cb58),
	.w8(32'hba225cb1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b09860),
	.w1(32'hba10effc),
	.w2(32'hba4afc90),
	.w3(32'hba814157),
	.w4(32'hba6eb9fc),
	.w5(32'h39f16100),
	.w6(32'hb9df2e89),
	.w7(32'hba85b5d4),
	.w8(32'h39016488),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95179cf),
	.w1(32'hb9d3d0a9),
	.w2(32'hbaba1daa),
	.w3(32'hb8fe3e6b),
	.w4(32'hba5577e9),
	.w5(32'hba3d4113),
	.w6(32'h38d99344),
	.w7(32'hba6c5423),
	.w8(32'hba5aa5e1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97e8d8),
	.w1(32'hb9ede714),
	.w2(32'hb996a959),
	.w3(32'hb9901be7),
	.w4(32'hb996e9f3),
	.w5(32'h385c6d59),
	.w6(32'h37d943d9),
	.w7(32'hb8b7f950),
	.w8(32'h392d4e8f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9795c06),
	.w1(32'hb8af75ee),
	.w2(32'h394a5d8b),
	.w3(32'h3a7282d3),
	.w4(32'h3aa420ea),
	.w5(32'h3aa40374),
	.w6(32'h39eef2b1),
	.w7(32'h3a945982),
	.w8(32'h3a3a558a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920fe43),
	.w1(32'hba4a6045),
	.w2(32'hbaa4eef9),
	.w3(32'h39e24641),
	.w4(32'hb8c8f502),
	.w5(32'hba000172),
	.w6(32'hb9c6e1b9),
	.w7(32'hba1f6fa1),
	.w8(32'hb9f92325),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9165c8),
	.w1(32'hba8041a3),
	.w2(32'hba6c41b6),
	.w3(32'hba374399),
	.w4(32'hba57edec),
	.w5(32'h3982bd0d),
	.w6(32'hba0b87e3),
	.w7(32'hb9c5d6cc),
	.w8(32'h39c08938),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987109c),
	.w1(32'h399526e1),
	.w2(32'hb943b5c2),
	.w3(32'h3a313e7b),
	.w4(32'h38fd8ba1),
	.w5(32'hba874a88),
	.w6(32'h39b7df92),
	.w7(32'h395d43d6),
	.w8(32'hb84e5457),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b4d8a),
	.w1(32'h3a7571c7),
	.w2(32'h39ad811e),
	.w3(32'hba269090),
	.w4(32'hba22b8ff),
	.w5(32'hbb24c53b),
	.w6(32'h39f64791),
	.w7(32'h39bc1c37),
	.w8(32'hbb10c598),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac32b87),
	.w1(32'hba9945a0),
	.w2(32'hba852289),
	.w3(32'hbaa21b22),
	.w4(32'hba67757c),
	.w5(32'hb9b80df1),
	.w6(32'hba7c7a46),
	.w7(32'hba731c9e),
	.w8(32'hb99e4293),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a63ebf),
	.w1(32'h3a1b84e0),
	.w2(32'h3a38ba15),
	.w3(32'h39fc2c83),
	.w4(32'h3933a26e),
	.w5(32'hb9acc23c),
	.w6(32'h397cc282),
	.w7(32'h3928e839),
	.w8(32'hb943ca16),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb871c064),
	.w1(32'hb9a5f16e),
	.w2(32'hb967d2f0),
	.w3(32'hba2d9a9c),
	.w4(32'hb9f709a7),
	.w5(32'h380c193a),
	.w6(32'hba2bee39),
	.w7(32'hb9d0236e),
	.w8(32'h381f47b3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a33479),
	.w1(32'hb9847874),
	.w2(32'hb8d062df),
	.w3(32'hb925c8dd),
	.w4(32'hb8676cb3),
	.w5(32'hb84a8a83),
	.w6(32'hb93a331d),
	.w7(32'hb91284a8),
	.w8(32'hb915dfd3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968e4d4),
	.w1(32'h38515afa),
	.w2(32'h397e0d66),
	.w3(32'hb982cec0),
	.w4(32'h39b880de),
	.w5(32'hba1e418b),
	.w6(32'hba0b0e87),
	.w7(32'h3a03ef9d),
	.w8(32'hba54a98e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f48667),
	.w1(32'hba7dd7fa),
	.w2(32'hbaa456a9),
	.w3(32'hba6c78db),
	.w4(32'hba622c38),
	.w5(32'h3922efe1),
	.w6(32'hba8d03fc),
	.w7(32'hba987c29),
	.w8(32'h3a0cb6c9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11515b),
	.w1(32'h39ff7256),
	.w2(32'h3934148c),
	.w3(32'h3793c7e0),
	.w4(32'h39947658),
	.w5(32'hb8589bac),
	.w6(32'h398dc4e7),
	.w7(32'h3a0e7912),
	.w8(32'h38d3ab05),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ca3b9),
	.w1(32'hb7004902),
	.w2(32'hb8e85f8e),
	.w3(32'h379a57eb),
	.w4(32'h39d713c7),
	.w5(32'h3adfdc19),
	.w6(32'hb8a8efaa),
	.w7(32'h3907ee2c),
	.w8(32'h3ad4674e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed3968),
	.w1(32'h3ad4a4eb),
	.w2(32'h3ae267f6),
	.w3(32'h3abeb658),
	.w4(32'h3ae300f3),
	.w5(32'h39dda5af),
	.w6(32'h3ac4e7b1),
	.w7(32'h3ad5c2ac),
	.w8(32'h39bb4833),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h352dfb5e),
	.w1(32'h39087529),
	.w2(32'h39ba6a82),
	.w3(32'hb88ad482),
	.w4(32'h390da905),
	.w5(32'h397c7faa),
	.w6(32'h39b32cf9),
	.w7(32'h3a0d4413),
	.w8(32'h3972b837),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0dff7),
	.w1(32'hb8a50270),
	.w2(32'hb98cf645),
	.w3(32'h3910cb9e),
	.w4(32'hb9023449),
	.w5(32'h3a218768),
	.w6(32'hb90997e3),
	.w7(32'hb9686113),
	.w8(32'h3a873fb8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77c226),
	.w1(32'h3aab6458),
	.w2(32'h39e42e89),
	.w3(32'h3a8b07ec),
	.w4(32'h3978b76b),
	.w5(32'hba0304fb),
	.w6(32'h3b123489),
	.w7(32'h397185f4),
	.w8(32'hb9a895a1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fcc2e8),
	.w1(32'h39878af6),
	.w2(32'h393c503e),
	.w3(32'hba3dea9f),
	.w4(32'hba2c6159),
	.w5(32'hba8ea128),
	.w6(32'hba2b3aa6),
	.w7(32'hb98f7da1),
	.w8(32'hba508ffa),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ae241),
	.w1(32'hba02f169),
	.w2(32'h39144b16),
	.w3(32'hba0dc867),
	.w4(32'hb9c9380b),
	.w5(32'hba362ec4),
	.w6(32'hb90e5fe9),
	.w7(32'hba2f6a96),
	.w8(32'hba4208e3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24fbeb),
	.w1(32'hb96fa1d5),
	.w2(32'hb7c0763d),
	.w3(32'hb9b195e4),
	.w4(32'hb9aa2593),
	.w5(32'h3a13b5bb),
	.w6(32'hb9db2e0d),
	.w7(32'hb5e4b8bb),
	.w8(32'h3a9c7af9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0ae98),
	.w1(32'h3a4da910),
	.w2(32'h3a04aa0a),
	.w3(32'hb9808c74),
	.w4(32'hb9ccf73e),
	.w5(32'hba5b2fac),
	.w6(32'h3a7e0f84),
	.w7(32'h39d6fa33),
	.w8(32'hba9b18fa),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92452e),
	.w1(32'hba756832),
	.w2(32'hb9b1d532),
	.w3(32'hb75b4fe9),
	.w4(32'h3a20f6d3),
	.w5(32'h38f51416),
	.w6(32'hba8f048a),
	.w7(32'h3722283d),
	.w8(32'hb7f6b1b9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39571cf4),
	.w1(32'h399ccedb),
	.w2(32'h393f9f38),
	.w3(32'h392a7ae6),
	.w4(32'h3907beff),
	.w5(32'hb9826280),
	.w6(32'hb904ede3),
	.w7(32'h38dfff71),
	.w8(32'hb9a6a32b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7da26),
	.w1(32'hba5c522c),
	.w2(32'hba3463d8),
	.w3(32'hb9e9b568),
	.w4(32'hb9d9f74c),
	.w5(32'hb77cf55c),
	.w6(32'hba077bfb),
	.w7(32'hba373b0d),
	.w8(32'hb7ffebf3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a0b7be),
	.w1(32'hb8748a95),
	.w2(32'hb9b50698),
	.w3(32'hb82436fc),
	.w4(32'hb901bf66),
	.w5(32'hba9456e0),
	.w6(32'hb9b60690),
	.w7(32'hb9949281),
	.w8(32'hba7937ec),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74f7dc),
	.w1(32'hba282f68),
	.w2(32'hba9a1c17),
	.w3(32'hba4866eb),
	.w4(32'hbaacb6d6),
	.w5(32'h391fe7e3),
	.w6(32'hb9ee8087),
	.w7(32'hbaa95c3a),
	.w8(32'h3a24ed19),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f4332),
	.w1(32'h3a60c308),
	.w2(32'h3a68e31d),
	.w3(32'hb9b92b2c),
	.w4(32'hb9eb9d79),
	.w5(32'h38a4a693),
	.w6(32'h39bf5310),
	.w7(32'h39fb7cdd),
	.w8(32'hb95e61a7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907378f),
	.w1(32'h390ceb29),
	.w2(32'h3a01b34d),
	.w3(32'h3921627a),
	.w4(32'h3a0eff4d),
	.w5(32'h391ab0ab),
	.w6(32'hb9fc5f8c),
	.w7(32'h39fdd120),
	.w8(32'hb8affeba),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973941e),
	.w1(32'hb9d75a2f),
	.w2(32'hb8bbae2f),
	.w3(32'h3997abd9),
	.w4(32'h391a91c8),
	.w5(32'hb8a24e99),
	.w6(32'hb4b13c6d),
	.w7(32'hb98b1408),
	.w8(32'hb94edfbd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3fdc8),
	.w1(32'h3979e0d2),
	.w2(32'h3a984dc8),
	.w3(32'h3a1f1eb6),
	.w4(32'h3a9724ee),
	.w5(32'hb8d7a22a),
	.w6(32'h380b7203),
	.w7(32'h3aeefa80),
	.w8(32'hb72100aa),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02996c),
	.w1(32'h38ce3665),
	.w2(32'h39aa3a71),
	.w3(32'hb99d8c43),
	.w4(32'hb83864dc),
	.w5(32'hb9827da3),
	.w6(32'h381058a5),
	.w7(32'h3a064e22),
	.w8(32'h39dd20d2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d62188),
	.w1(32'h3a05e3b2),
	.w2(32'h3a548e56),
	.w3(32'hb95b0dda),
	.w4(32'hb9cbfe8a),
	.w5(32'h38e6e42b),
	.w6(32'h3a7801d6),
	.w7(32'h3a156d4a),
	.w8(32'h38b60cc8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38155718),
	.w1(32'hb995ff67),
	.w2(32'hb9fb9517),
	.w3(32'hb91540d7),
	.w4(32'h3961e9c6),
	.w5(32'h3ac59e7f),
	.w6(32'hb8e86d1c),
	.w7(32'h386e17a8),
	.w8(32'h3ab25d04),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa58ecd),
	.w1(32'h3abb61dd),
	.w2(32'h3a9da02e),
	.w3(32'h3aaa845b),
	.w4(32'h3ac811b8),
	.w5(32'hb99547c1),
	.w6(32'h3a9c82db),
	.w7(32'h3ac91dd7),
	.w8(32'hb98640cc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982901c),
	.w1(32'h3a09d836),
	.w2(32'h39f514ca),
	.w3(32'h387ab2a2),
	.w4(32'h39dd91e7),
	.w5(32'hb9874128),
	.w6(32'h39b9d9a8),
	.w7(32'h3a3e5296),
	.w8(32'hb9c91909),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82bb947),
	.w1(32'h3927022a),
	.w2(32'hb9e9d863),
	.w3(32'hb86859ce),
	.w4(32'h39983934),
	.w5(32'hb9fbde10),
	.w6(32'hb9ff7200),
	.w7(32'hb6b99fb8),
	.w8(32'hba0b378d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9783423),
	.w1(32'hba14b582),
	.w2(32'hb8da5f10),
	.w3(32'hb90565ca),
	.w4(32'h395a4e31),
	.w5(32'h3a39dc0d),
	.w6(32'hba309220),
	.w7(32'hb851e6fc),
	.w8(32'h39cf412a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983367f),
	.w1(32'h380a5e63),
	.w2(32'h3a451d7a),
	.w3(32'hb99d12c6),
	.w4(32'h39c4056b),
	.w5(32'h38ee2a4c),
	.w6(32'hb9e9e375),
	.w7(32'h3a0bf7d7),
	.w8(32'hba21f166),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfffe7),
	.w1(32'h3a8f0f89),
	.w2(32'h3a62abbf),
	.w3(32'h398b9bdf),
	.w4(32'h392af4d9),
	.w5(32'hb83b62b0),
	.w6(32'hba149ee7),
	.w7(32'hb9a03d3f),
	.w8(32'hb9cff0f4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c3d4a),
	.w1(32'hb8502048),
	.w2(32'h39e46588),
	.w3(32'h39a0cf79),
	.w4(32'h3a19210d),
	.w5(32'h39e7ed6d),
	.w6(32'h3a111e7c),
	.w7(32'h3a2d766e),
	.w8(32'h39f4ea9c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3974f2fa),
	.w1(32'h3a060653),
	.w2(32'h39d500ee),
	.w3(32'h3a54f3f2),
	.w4(32'h3a016cd3),
	.w5(32'h3943d621),
	.w6(32'h3a67f60b),
	.w7(32'h3a044c1a),
	.w8(32'h39ccc57b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a44fee),
	.w1(32'h3a3188f5),
	.w2(32'h3a70d237),
	.w3(32'h397742a5),
	.w4(32'h399f181d),
	.w5(32'hb937ce18),
	.w6(32'h39ba438a),
	.w7(32'h3a241d09),
	.w8(32'h392b66bc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a1ce95),
	.w1(32'h3a7c2baa),
	.w2(32'h3aa5f3be),
	.w3(32'h3994dd9f),
	.w4(32'hb8206745),
	.w5(32'h3810343c),
	.w6(32'h39185b10),
	.w7(32'h3a71a9ad),
	.w8(32'h39b694e6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1eb4d3),
	.w1(32'h38f33876),
	.w2(32'hb9ebdaee),
	.w3(32'hba45377c),
	.w4(32'hba5a4984),
	.w5(32'h388a2b83),
	.w6(32'hb9ffefa1),
	.w7(32'hba07b6f3),
	.w8(32'hb8afb6b0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97634d7),
	.w1(32'h38572f26),
	.w2(32'h3978f751),
	.w3(32'h39020fb7),
	.w4(32'h39eb57ef),
	.w5(32'h3a2850a6),
	.w6(32'hb949c38d),
	.w7(32'h39b3f0a0),
	.w8(32'h3a41c678),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a8af7),
	.w1(32'h3a6cc26e),
	.w2(32'h3a86a9d5),
	.w3(32'h39b93677),
	.w4(32'h39d83386),
	.w5(32'h38fd31dd),
	.w6(32'h39a0318f),
	.w7(32'h3a69c0ec),
	.w8(32'h399f5880),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f7878),
	.w1(32'hb9d2a0b6),
	.w2(32'hb98c5951),
	.w3(32'hb8ad4527),
	.w4(32'hb98b6bc2),
	.w5(32'h39953ac2),
	.w6(32'hb939bc2b),
	.w7(32'hb9dd1faa),
	.w8(32'h38c4c69e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b64a09),
	.w1(32'hb95506f7),
	.w2(32'hb96153ac),
	.w3(32'hb8778c33),
	.w4(32'hb90afe22),
	.w5(32'h390ce8b2),
	.w6(32'h38873a8f),
	.w7(32'h37a24865),
	.w8(32'h3932c997),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b395c5),
	.w1(32'hb899cb02),
	.w2(32'hb90fc5cb),
	.w3(32'h38494b00),
	.w4(32'hb9accc4d),
	.w5(32'h3a920447),
	.w6(32'hba5b6284),
	.w7(32'hb993d32a),
	.w8(32'h3a95b8f0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7beba7),
	.w1(32'h3aa3c74b),
	.w2(32'h3ade3fb8),
	.w3(32'h3ae7d937),
	.w4(32'h3af9d001),
	.w5(32'h3a205e7e),
	.w6(32'h3ae78506),
	.w7(32'h3aeb1841),
	.w8(32'h3a43fefa),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e875d),
	.w1(32'h3a8ffc28),
	.w2(32'h3a8d5bb0),
	.w3(32'h399c3ae7),
	.w4(32'h39a4c6bb),
	.w5(32'hb9f4b470),
	.w6(32'hb9826a66),
	.w7(32'h3a34d56b),
	.w8(32'hb87411f4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922ec56),
	.w1(32'hb8a87583),
	.w2(32'h3987428a),
	.w3(32'hb9df7b10),
	.w4(32'hb967189a),
	.w5(32'hb9ca3235),
	.w6(32'hb91e568c),
	.w7(32'h39ad78c1),
	.w8(32'hb9809065),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bccff8),
	.w1(32'hba9251b1),
	.w2(32'hbaa399a3),
	.w3(32'hba07f1a8),
	.w4(32'hb9999a79),
	.w5(32'h39806217),
	.w6(32'hba4f7b94),
	.w7(32'hba3bdc49),
	.w8(32'hb90df9f4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa49a3),
	.w1(32'h3a870f27),
	.w2(32'h39e32b8b),
	.w3(32'hb991c86f),
	.w4(32'hb9cbd0df),
	.w5(32'hb810ba36),
	.w6(32'hb9c58d9e),
	.w7(32'hb9dd5faa),
	.w8(32'hb6c9fd5f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938bf76),
	.w1(32'h39053507),
	.w2(32'h38e46958),
	.w3(32'hb89b50f0),
	.w4(32'h37ad5428),
	.w5(32'h37ee3a3e),
	.w6(32'hb956c6ce),
	.w7(32'h3957518f),
	.w8(32'h3979ebe5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bd538),
	.w1(32'h38ff1cd0),
	.w2(32'hb88b7c3f),
	.w3(32'hb9599c9b),
	.w4(32'hb9d1fad8),
	.w5(32'h38e343ba),
	.w6(32'hb9bb47d4),
	.w7(32'hb9f0b263),
	.w8(32'h37a9e436),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3863ddd2),
	.w1(32'h3aae0adc),
	.w2(32'h39ee9cb9),
	.w3(32'h3ab7a8ea),
	.w4(32'h3a17b99e),
	.w5(32'hba811b3d),
	.w6(32'h3af0b2c0),
	.w7(32'h3a52c6bf),
	.w8(32'hbac71aac),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86479e),
	.w1(32'hb98d7897),
	.w2(32'h3a670c6b),
	.w3(32'hb82a46b2),
	.w4(32'h3a71440d),
	.w5(32'hba692534),
	.w6(32'hba6b4e24),
	.w7(32'h3a8aa30e),
	.w8(32'hba76d1f1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10e3c7),
	.w1(32'hb9e67dd9),
	.w2(32'hba43bdfc),
	.w3(32'hba545cb5),
	.w4(32'hba530302),
	.w5(32'hb95b9d11),
	.w6(32'hba7698e6),
	.w7(32'hba40a252),
	.w8(32'hb9e98fb3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9603ba4),
	.w1(32'hb848b886),
	.w2(32'hb9a70bf6),
	.w3(32'h3a1edda1),
	.w4(32'h39d9abf5),
	.w5(32'h3a1d53d6),
	.w6(32'h388fc6ab),
	.w7(32'h39965780),
	.w8(32'h3a4290f2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06ca84),
	.w1(32'h3a0f5fe4),
	.w2(32'h3a8cf88c),
	.w3(32'h3980d4b7),
	.w4(32'h3a06be37),
	.w5(32'hb931f6ef),
	.w6(32'h38b9ec9f),
	.w7(32'h3a6a40b4),
	.w8(32'h39276fbf),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cc045),
	.w1(32'h39308875),
	.w2(32'h38eb4a6f),
	.w3(32'hb9e4fc14),
	.w4(32'hb9fa1036),
	.w5(32'hbaa55005),
	.w6(32'hb9fc9ac2),
	.w7(32'hb9737ae6),
	.w8(32'hba9adb5b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d90ed),
	.w1(32'hb9b583aa),
	.w2(32'hb926670a),
	.w3(32'hba46017c),
	.w4(32'hb9c1b34c),
	.w5(32'hba10703b),
	.w6(32'hba2fdddc),
	.w7(32'hba149e2b),
	.w8(32'hba26a875),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7c144),
	.w1(32'hba8eb30e),
	.w2(32'hbaa18327),
	.w3(32'hba9f69e1),
	.w4(32'hbab91f38),
	.w5(32'h3ba9b996),
	.w6(32'hbaff58ff),
	.w7(32'hbac33920),
	.w8(32'hbb0f6dec),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfaf39),
	.w1(32'hbb0bc567),
	.w2(32'hbbb02894),
	.w3(32'hbb6a0ef3),
	.w4(32'hbb77cc95),
	.w5(32'hbc2359e8),
	.w6(32'hbad17adc),
	.w7(32'hbaa7064e),
	.w8(32'hbcba3a64),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d3622),
	.w1(32'hbc3f0a02),
	.w2(32'hbb99f106),
	.w3(32'hbcf87d2d),
	.w4(32'h3a65035a),
	.w5(32'hbb0addfd),
	.w6(32'hbd1aa006),
	.w7(32'hba39976c),
	.w8(32'h3ae32055),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9273bb),
	.w1(32'h3c0c88ed),
	.w2(32'h3b927678),
	.w3(32'h3ac8f13f),
	.w4(32'hbb490a2e),
	.w5(32'h3c57b8b7),
	.w6(32'h3c64a2d6),
	.w7(32'hbbcdc3cd),
	.w8(32'h3ab8a5b4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cd16d),
	.w1(32'hbb6b60e6),
	.w2(32'hbb838cf7),
	.w3(32'h3b6e76f8),
	.w4(32'h3b6e58bd),
	.w5(32'hb9ad942a),
	.w6(32'hbb8108a1),
	.w7(32'hb8853f65),
	.w8(32'hbb88d3f2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ed30),
	.w1(32'hbc170d1a),
	.w2(32'hba07dcd5),
	.w3(32'hbc055c8c),
	.w4(32'h3aaa35e9),
	.w5(32'hbccbdcf5),
	.w6(32'hbc08c649),
	.w7(32'hbc222150),
	.w8(32'hbd7bbeff),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd11be0c),
	.w1(32'hbbc69926),
	.w2(32'h3cc5b0f9),
	.w3(32'hbcd03a8a),
	.w4(32'h3c73aad1),
	.w5(32'hbaafe59c),
	.w6(32'hb9058dbd),
	.w7(32'h3d5c25be),
	.w8(32'h3c8aa224),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53faa9),
	.w1(32'h3b9a5914),
	.w2(32'hbc6eea31),
	.w3(32'h3c078d39),
	.w4(32'hbc15cb7c),
	.w5(32'hbcd8174b),
	.w6(32'hbad27ea5),
	.w7(32'hbc95e32c),
	.w8(32'hbcf49d90),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4a1f5),
	.w1(32'h3b7d0c6d),
	.w2(32'h3ce19251),
	.w3(32'hbc168cab),
	.w4(32'h3bcf525f),
	.w5(32'hbc841e36),
	.w6(32'hbc2b4674),
	.w7(32'h3cfd4a4c),
	.w8(32'hbc845244),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc732c7b),
	.w1(32'hbb7923a2),
	.w2(32'h3c97981b),
	.w3(32'hbc861b7a),
	.w4(32'hbbb3bd0a),
	.w5(32'h3c4752f7),
	.w6(32'hbbd4de2a),
	.w7(32'h3cadf665),
	.w8(32'h3c8a9485),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37fd82),
	.w1(32'hbbc11d7e),
	.w2(32'hbc247476),
	.w3(32'hba62b7b6),
	.w4(32'hbbe1ea3b),
	.w5(32'h3c05ef51),
	.w6(32'hbbbd4b6c),
	.w7(32'hbc8cb8ed),
	.w8(32'hbaee2a29),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b1369),
	.w1(32'hbb0f5e7c),
	.w2(32'hbc0897b2),
	.w3(32'hbb7bf921),
	.w4(32'hbbe0d5fd),
	.w5(32'h3cd9d363),
	.w6(32'hbb9d2b5a),
	.w7(32'hbbf64d1b),
	.w8(32'h3cc9e838),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d9803),
	.w1(32'hbc0e89cd),
	.w2(32'hbcc2fb43),
	.w3(32'h3c4ad6f5),
	.w4(32'hbae78da1),
	.w5(32'hbb07d719),
	.w6(32'hbb48ed79),
	.w7(32'hbcb7f9ca),
	.w8(32'h3bd54b05),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c7390),
	.w1(32'h3b118f66),
	.w2(32'h3c5a1a9c),
	.w3(32'h3b856f05),
	.w4(32'hba8b6276),
	.w5(32'h3a6ebeee),
	.w6(32'h3a9f4b2d),
	.w7(32'hbbac60b4),
	.w8(32'hbbf9db50),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27311c),
	.w1(32'h3b343174),
	.w2(32'hbb1a6a1f),
	.w3(32'h3a92fe23),
	.w4(32'hbb281a76),
	.w5(32'h3bfc017f),
	.w6(32'hba1ef676),
	.w7(32'hbb8f1a27),
	.w8(32'h3c84eaa9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a57b5),
	.w1(32'hbc1eba05),
	.w2(32'hbc00df28),
	.w3(32'h3af23c04),
	.w4(32'hbc27a215),
	.w5(32'hba9e46ab),
	.w6(32'hbc6001c0),
	.w7(32'hbcba32e4),
	.w8(32'hbc240dd7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9abb0),
	.w1(32'hba49dac8),
	.w2(32'h39d29034),
	.w3(32'h3b0f8f6e),
	.w4(32'h3a84a25a),
	.w5(32'hbc92371b),
	.w6(32'hbac452e8),
	.w7(32'hbb0823ad),
	.w8(32'hbcabe7d3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc6afb),
	.w1(32'h3ae74e25),
	.w2(32'h3bddb3c6),
	.w3(32'hbc9bb179),
	.w4(32'h3c1a563b),
	.w5(32'hbaec9e8b),
	.w6(32'hbccd2bfe),
	.w7(32'h3ad291aa),
	.w8(32'hbbeb8091),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73277f),
	.w1(32'hbad6a389),
	.w2(32'h39f7ae11),
	.w3(32'hbba5d7b0),
	.w4(32'h39b3c2ad),
	.w5(32'h3cbf37df),
	.w6(32'hbc46a522),
	.w7(32'hb9906b9e),
	.w8(32'h3d09eed0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca55471),
	.w1(32'h3a0ac327),
	.w2(32'hbccda434),
	.w3(32'h3c39a4e8),
	.w4(32'hbc422450),
	.w5(32'hbb025459),
	.w6(32'h3c3c7e4a),
	.w7(32'hbcbf1ed2),
	.w8(32'hbc13946e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ba1b6),
	.w1(32'hbbb56b3c),
	.w2(32'hbc44d721),
	.w3(32'h3af6197d),
	.w4(32'h3ad7a7f3),
	.w5(32'hbae4940d),
	.w6(32'h3bcd2703),
	.w7(32'h3c817687),
	.w8(32'hbab1d1f6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad5c3c),
	.w1(32'hbb272366),
	.w2(32'hbae4da5d),
	.w3(32'hbbedf164),
	.w4(32'hbbce8acd),
	.w5(32'hbc4a2847),
	.w6(32'hbb768cad),
	.w7(32'hbbbecfa6),
	.w8(32'hbcfe05b0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc704cc9),
	.w1(32'h3c579a6f),
	.w2(32'h3d0183b9),
	.w3(32'hbc9de04e),
	.w4(32'h3c44cba0),
	.w5(32'h3acc3442),
	.w6(32'h3c0ee490),
	.w7(32'h3d2d76f9),
	.w8(32'hbbb56069),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1abbcb),
	.w1(32'h3bd4a800),
	.w2(32'h3b9139ea),
	.w3(32'hbc2c0332),
	.w4(32'hb9dea8bb),
	.w5(32'h3bf2fd26),
	.w6(32'hbb545f63),
	.w7(32'h3b4249a8),
	.w8(32'h3c3437d7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2616c6),
	.w1(32'hbbacd3cd),
	.w2(32'hbae0efbc),
	.w3(32'h3bcadd4f),
	.w4(32'h3be4ad99),
	.w5(32'h3b90ff58),
	.w6(32'h3b09b88d),
	.w7(32'h3b81ef26),
	.w8(32'h3b444fe8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b240f49),
	.w1(32'h3a41f9b2),
	.w2(32'h3c1e589c),
	.w3(32'h3c002287),
	.w4(32'h3ac05667),
	.w5(32'hbb6c19a7),
	.w6(32'hbb28e003),
	.w7(32'h3bf83d1a),
	.w8(32'h3c40e69f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4bb92),
	.w1(32'hbc16e16a),
	.w2(32'h3af90899),
	.w3(32'h3c2a3108),
	.w4(32'h3c5e9df5),
	.w5(32'h3bc125b5),
	.w6(32'h3b435276),
	.w7(32'h3c067a57),
	.w8(32'h3b99f472),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07acb8),
	.w1(32'hba75421b),
	.w2(32'hb97a707e),
	.w3(32'h3bb2fc26),
	.w4(32'h3c18476a),
	.w5(32'h3b479e70),
	.w6(32'hb9d082f8),
	.w7(32'h3b2338ef),
	.w8(32'hbbf79e13),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb457457),
	.w1(32'hbb1e379e),
	.w2(32'hbbf8267e),
	.w3(32'hb9574983),
	.w4(32'hba35206d),
	.w5(32'h3c99537d),
	.w6(32'h3ba6b3c7),
	.w7(32'hbbaebb1d),
	.w8(32'h3cff360d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91dc92),
	.w1(32'hbb892fc6),
	.w2(32'hbcce3a44),
	.w3(32'h3c3279c1),
	.w4(32'hbbb73e1b),
	.w5(32'hbbfaa39c),
	.w6(32'h3bdc567b),
	.w7(32'hbcb6b2bc),
	.w8(32'hbcc41265),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe757f5),
	.w1(32'hbb79ca0c),
	.w2(32'h3c79e49f),
	.w3(32'hbc177ed7),
	.w4(32'h3bc658df),
	.w5(32'h3c8008a3),
	.w6(32'hbc0a4419),
	.w7(32'h3c4763c0),
	.w8(32'h3998fd91),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ad545),
	.w1(32'hbbb4f19a),
	.w2(32'hbb21f099),
	.w3(32'h39ac22ee),
	.w4(32'hb9579b06),
	.w5(32'hbbccf943),
	.w6(32'hbbac0778),
	.w7(32'hbbe780ca),
	.w8(32'h3b8f0421),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba470934),
	.w1(32'h3a5249bf),
	.w2(32'hbb0c7b8b),
	.w3(32'h3b4dacb1),
	.w4(32'h3b9cbd6a),
	.w5(32'hbbacee97),
	.w6(32'hbb5dcc31),
	.w7(32'hb8351164),
	.w8(32'hbb68ca7a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44813d),
	.w1(32'hbb39309f),
	.w2(32'h3b2bdf4e),
	.w3(32'hbc289aa4),
	.w4(32'hbc546129),
	.w5(32'h3c1f1b0c),
	.w6(32'hba6f8a42),
	.w7(32'h3a504fd7),
	.w8(32'h3cc023a4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56a9c3),
	.w1(32'hba15c082),
	.w2(32'hbb9a7ecc),
	.w3(32'h3c207146),
	.w4(32'h3b0d0cde),
	.w5(32'h3c7963e0),
	.w6(32'h3bb2bdbf),
	.w7(32'hbc0e1cee),
	.w8(32'h3c230390),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c503367),
	.w1(32'hbc784c19),
	.w2(32'h3b0695c4),
	.w3(32'hbbf5f450),
	.w4(32'h3c15529b),
	.w5(32'h3cecf758),
	.w6(32'hbab41c3b),
	.w7(32'h3be81ca5),
	.w8(32'h3ceede28),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37c211),
	.w1(32'hbc11e612),
	.w2(32'hbcaaba0a),
	.w3(32'h3c8e4e35),
	.w4(32'hbb47a0fe),
	.w5(32'h3c92b27b),
	.w6(32'hba5e927a),
	.w7(32'hbce8d65d),
	.w8(32'h3d007f18),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c772410),
	.w1(32'h3b2e4624),
	.w2(32'hbc732d06),
	.w3(32'h3c7fdc44),
	.w4(32'hbb2d64e0),
	.w5(32'h3cab4423),
	.w6(32'h3c2104fa),
	.w7(32'hbc887194),
	.w8(32'h3cdab292),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa7d64),
	.w1(32'hbc331089),
	.w2(32'hbbc88ed4),
	.w3(32'h3c466972),
	.w4(32'hbc066b32),
	.w5(32'h3ca22275),
	.w6(32'h394e3036),
	.w7(32'hbcbb68e6),
	.w8(32'h3cf77638),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67a6e9),
	.w1(32'hbae582dd),
	.w2(32'hbc9f6f1c),
	.w3(32'h3c6641ed),
	.w4(32'hbc03f9a7),
	.w5(32'h3cd21058),
	.w6(32'h3bde4d69),
	.w7(32'hbcbf16be),
	.w8(32'h3ce5abc8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fbfc2),
	.w1(32'hbc37cc73),
	.w2(32'hbcc839d1),
	.w3(32'h3c709626),
	.w4(32'hbb49421f),
	.w5(32'h3c918c5b),
	.w6(32'hb9a0a7b9),
	.w7(32'hbce01d2a),
	.w8(32'h3c9cfa2e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c366339),
	.w1(32'hbc13de7a),
	.w2(32'hba9ef645),
	.w3(32'h3c0029d4),
	.w4(32'h3a3e9d0e),
	.w5(32'hbc0a6254),
	.w6(32'hbc254018),
	.w7(32'hbc8d11ce),
	.w8(32'hbbad4900),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc58ae3),
	.w1(32'hbaeea70f),
	.w2(32'h3b853205),
	.w3(32'hbc079fba),
	.w4(32'hbc5907a4),
	.w5(32'hbce66ffd),
	.w6(32'h3b873431),
	.w7(32'hbba56fd8),
	.w8(32'hbc80d0b0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc923541),
	.w1(32'h3a9f8130),
	.w2(32'h3d03cfce),
	.w3(32'hbbe0fc97),
	.w4(32'h3c6faf11),
	.w5(32'h3c03fd5f),
	.w6(32'hbb5b0f6c),
	.w7(32'h3d0a8d05),
	.w8(32'hbc19deb5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb592c80),
	.w1(32'hbc60f3d2),
	.w2(32'h3a95576e),
	.w3(32'hbc921f94),
	.w4(32'hb81cf9de),
	.w5(32'hbb307f7b),
	.w6(32'hbc5377c6),
	.w7(32'h3c0943fd),
	.w8(32'h3c3800e3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9ed5c),
	.w1(32'h3a857d7f),
	.w2(32'h3c10edc4),
	.w3(32'h3bbfe4fc),
	.w4(32'hbaf93fab),
	.w5(32'h3bb751ae),
	.w6(32'hbb846cc7),
	.w7(32'hbc5ab2b2),
	.w8(32'h3bc52dab),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8930e3),
	.w1(32'hbc5b26c3),
	.w2(32'hbc5a00e3),
	.w3(32'h3b8f3071),
	.w4(32'h3b93ec07),
	.w5(32'h3cb4b094),
	.w6(32'hbc5f9a72),
	.w7(32'hbc455d96),
	.w8(32'h3d0102d3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ffacc),
	.w1(32'h3ac90460),
	.w2(32'hbc4c34f8),
	.w3(32'h3c4ed41f),
	.w4(32'hbbcf0983),
	.w5(32'hbc709412),
	.w6(32'hbb448a5d),
	.w7(32'hbce45765),
	.w8(32'hbc9ff676),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0911d6),
	.w1(32'h3ba611ce),
	.w2(32'h3ce27186),
	.w3(32'hbb8ba949),
	.w4(32'h3c3066fb),
	.w5(32'hbb32af45),
	.w6(32'hbc0f4d3c),
	.w7(32'h3ceeb83f),
	.w8(32'hbcd1ac8a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31f96c),
	.w1(32'h3c2f6710),
	.w2(32'h3c30c301),
	.w3(32'h3b81f3a5),
	.w4(32'h3c04553d),
	.w5(32'h3a08733a),
	.w6(32'h3acef4d7),
	.w7(32'h3cc61802),
	.w8(32'hba515bc9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02d73e),
	.w1(32'hbc3285bb),
	.w2(32'h3b388a57),
	.w3(32'h3a4dfc97),
	.w4(32'h3b061752),
	.w5(32'h3b8a0b93),
	.w6(32'hba8c2cc0),
	.w7(32'hbb2b9441),
	.w8(32'h3afbb5ad),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad556c6),
	.w1(32'hbb8c92a1),
	.w2(32'hbbc7698f),
	.w3(32'h3c2d875c),
	.w4(32'h3c62c2e0),
	.w5(32'h3d0830b3),
	.w6(32'h3b095bb9),
	.w7(32'h3b57d16d),
	.w8(32'h3d1edfc7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb1d39),
	.w1(32'hbac637c6),
	.w2(32'hbd0a75a9),
	.w3(32'h3c335355),
	.w4(32'hbc934ae2),
	.w5(32'hba4156bc),
	.w6(32'h3c294caa),
	.w7(32'hbcfa7c2a),
	.w8(32'hba9ced2b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aebe0),
	.w1(32'h3aca815a),
	.w2(32'h3b5dfe89),
	.w3(32'hbabd02de),
	.w4(32'hbab9f91b),
	.w5(32'h3b5a7a1b),
	.w6(32'h3b1878f8),
	.w7(32'hbb408ba7),
	.w8(32'h3befa311),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f35a9a),
	.w1(32'hbbc37566),
	.w2(32'h3c4efd89),
	.w3(32'h3b14de03),
	.w4(32'h3bf0688b),
	.w5(32'h3b81a26d),
	.w6(32'hbb3c7027),
	.w7(32'h3bbffc6a),
	.w8(32'hbc3dca09),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc90253),
	.w1(32'h3b37a2d3),
	.w2(32'h3be0ebed),
	.w3(32'hbbd269e1),
	.w4(32'hbb522676),
	.w5(32'h3ba3f7dc),
	.w6(32'hbb802c7d),
	.w7(32'h3c05ee58),
	.w8(32'h3ca872a4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3b05d),
	.w1(32'hbabc6c16),
	.w2(32'hbb054547),
	.w3(32'h3c48e875),
	.w4(32'hbb736473),
	.w5(32'h3bdd81e3),
	.w6(32'hbaa0703f),
	.w7(32'hbcc1369e),
	.w8(32'h3c4fecbc),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1962fb),
	.w1(32'hbb83b21c),
	.w2(32'hbbf38c14),
	.w3(32'h39986a45),
	.w4(32'hbc10455e),
	.w5(32'h3cb16c5b),
	.w6(32'hbb066ac1),
	.w7(32'hbc9e483b),
	.w8(32'h3ca6a1bd),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c191d88),
	.w1(32'hbb535072),
	.w2(32'hbc543d80),
	.w3(32'h3bf93e75),
	.w4(32'h3af62cbc),
	.w5(32'h3c31b4d1),
	.w6(32'h3ac90e00),
	.w7(32'hbc1efa7c),
	.w8(32'h3b1ceebc),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb784dd),
	.w1(32'hbc224c2e),
	.w2(32'hbbc56a1d),
	.w3(32'h3bd6415d),
	.w4(32'h3ba27aa1),
	.w5(32'h3b6330fa),
	.w6(32'h3bb40fb2),
	.w7(32'h3b420bfa),
	.w8(32'h3992a2e3),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18b0b5),
	.w1(32'hbc02e22a),
	.w2(32'hbb4d8d67),
	.w3(32'h3aea6d80),
	.w4(32'h3ac791a1),
	.w5(32'hbc0754ba),
	.w6(32'hba8cf45b),
	.w7(32'h3b538112),
	.w8(32'hbc593131),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5bbfa),
	.w1(32'hbb4dd16b),
	.w2(32'h38b4d60a),
	.w3(32'hbbeaf8f5),
	.w4(32'h3a250074),
	.w5(32'hbb006d13),
	.w6(32'hbc809bdb),
	.w7(32'hba57a542),
	.w8(32'hbc0fc80c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f9b8),
	.w1(32'hbb846b42),
	.w2(32'h3c191470),
	.w3(32'hbc07d137),
	.w4(32'hbba15cff),
	.w5(32'hbc2e8c45),
	.w6(32'hbbd6030c),
	.w7(32'h3c5eb91a),
	.w8(32'hbcd00781),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93b0ae),
	.w1(32'h3c4f506d),
	.w2(32'h3c6786ae),
	.w3(32'hbc98d9c1),
	.w4(32'h3b3a6d8c),
	.w5(32'hbc4b0b6d),
	.w6(32'hbc96f817),
	.w7(32'h3c4e9349),
	.w8(32'hbca092cb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9baa87),
	.w1(32'hbbe3ae07),
	.w2(32'h3cd33497),
	.w3(32'hbc1933a4),
	.w4(32'h3c63a088),
	.w5(32'h3c16c9cd),
	.w6(32'hbc4b4dc2),
	.w7(32'h3cab32ba),
	.w8(32'h3c1ef640),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c326fb7),
	.w1(32'h3b3ec336),
	.w2(32'hbbe24e0c),
	.w3(32'h3b893003),
	.w4(32'h398ad354),
	.w5(32'hbc66c968),
	.w6(32'h3c05baf2),
	.w7(32'h38a92849),
	.w8(32'hbc4790a7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5d467),
	.w1(32'h3c014d87),
	.w2(32'h3c4d6300),
	.w3(32'hbc6f42ef),
	.w4(32'h3c570cf0),
	.w5(32'hbc2edffb),
	.w6(32'hbc8894e7),
	.w7(32'h3c9bd016),
	.w8(32'hbc226d28),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac06bd1),
	.w1(32'hbb362d03),
	.w2(32'hbc9436e6),
	.w3(32'hbc449557),
	.w4(32'h3b434ea4),
	.w5(32'h3c45f24e),
	.w6(32'h3bf2820b),
	.w7(32'h3ca1dd2d),
	.w8(32'h3c05a612),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3e0a2),
	.w1(32'hbafd90f6),
	.w2(32'hbc4bcbc0),
	.w3(32'h3c176f95),
	.w4(32'hbb3f919a),
	.w5(32'h39675691),
	.w6(32'hbb925017),
	.w7(32'hbca0298d),
	.w8(32'h3b5371b0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2da81),
	.w1(32'hb9b49c41),
	.w2(32'hbaead938),
	.w3(32'h3b97e852),
	.w4(32'h3b4e1f36),
	.w5(32'h3cbb6e8f),
	.w6(32'h3c0b0c90),
	.w7(32'h381d0283),
	.w8(32'h3c3f1d62),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c3ff9),
	.w1(32'hbc599c70),
	.w2(32'hbd23e32e),
	.w3(32'h3adefa1d),
	.w4(32'hbb87a965),
	.w5(32'hbabe34dd),
	.w6(32'h3c73bb80),
	.w7(32'hbc92d524),
	.w8(32'hbc044a8c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7b293),
	.w1(32'h3baf287d),
	.w2(32'h3c220eb1),
	.w3(32'hbaa0b5a0),
	.w4(32'hba6bf860),
	.w5(32'h3c9e21a0),
	.w6(32'hbb70df67),
	.w7(32'h3b4c576d),
	.w8(32'h3d166aa3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91e9dc),
	.w1(32'hbb38d480),
	.w2(32'hbca23fe8),
	.w3(32'h3c02b60a),
	.w4(32'hbc3f2a60),
	.w5(32'hbc9f9ad7),
	.w6(32'h3ba35f35),
	.w7(32'hbcd2ed61),
	.w8(32'hbcd9f777),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2e4bb),
	.w1(32'h3c49d41e),
	.w2(32'h3cccfac5),
	.w3(32'hbbe290ff),
	.w4(32'h3aef8269),
	.w5(32'h3c5fe9f5),
	.w6(32'h3b820277),
	.w7(32'h3d08bb3d),
	.w8(32'h3c9f414d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5db01),
	.w1(32'h3a9ca2c3),
	.w2(32'h3a8c1a37),
	.w3(32'h3c43713f),
	.w4(32'h3c345f24),
	.w5(32'hbbaabe27),
	.w6(32'hbcb3a93c),
	.w7(32'hbc914e21),
	.w8(32'hbc2e8294),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29f042),
	.w1(32'h3c3b5990),
	.w2(32'h3c36237e),
	.w3(32'hbb15d31c),
	.w4(32'h3c38ce49),
	.w5(32'h3bc5284a),
	.w6(32'h3c1e1528),
	.w7(32'h3c594a58),
	.w8(32'hba054943),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3353a0),
	.w1(32'h3c27b054),
	.w2(32'h3b58cc33),
	.w3(32'h3bd5a304),
	.w4(32'hbbce5d6d),
	.w5(32'hbb5398de),
	.w6(32'h3c46f7e0),
	.w7(32'hbb115bf7),
	.w8(32'hbc141933),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc36e75),
	.w1(32'hbb3f784d),
	.w2(32'hbc101ffd),
	.w3(32'hbc1c9533),
	.w4(32'hbb4b66b2),
	.w5(32'h3cc89332),
	.w6(32'hb9f56e86),
	.w7(32'hbc058782),
	.w8(32'h3d28c09f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5685f),
	.w1(32'hbb9ada77),
	.w2(32'hbce0cf51),
	.w3(32'h3c20cf7c),
	.w4(32'hbcb939fb),
	.w5(32'hbc38a2d5),
	.w6(32'h3b8f4ee1),
	.w7(32'hbd0e292c),
	.w8(32'hba797b25),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd06786),
	.w1(32'h3bf2b74b),
	.w2(32'h3cdeaba6),
	.w3(32'h3b0e00fb),
	.w4(32'h3c0a0b5f),
	.w5(32'h3cf40b5c),
	.w6(32'h3b5e6413),
	.w7(32'h3ce63f4c),
	.w8(32'h3d1d32ca),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe0347),
	.w1(32'hbc2b0e96),
	.w2(32'hbd1feb85),
	.w3(32'h3bac5d16),
	.w4(32'hbcbdd0de),
	.w5(32'hbb7eb00f),
	.w6(32'h3a3b548d),
	.w7(32'hbd28dc3a),
	.w8(32'hbc1c55fe),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cda55),
	.w1(32'hbcec0fe3),
	.w2(32'hbc431bc1),
	.w3(32'hbd002d5f),
	.w4(32'h3b5ab5e9),
	.w5(32'hbc0de982),
	.w6(32'hbcef86db),
	.w7(32'h3b85b885),
	.w8(32'hbc59c648),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cd405),
	.w1(32'h3c483379),
	.w2(32'h3c9b2360),
	.w3(32'h3a9b71af),
	.w4(32'h3c10d14c),
	.w5(32'h3b8d6163),
	.w6(32'h3b8beef8),
	.w7(32'h3cd4810e),
	.w8(32'h3a924600),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8992ca),
	.w1(32'h3b227475),
	.w2(32'h3c08ed62),
	.w3(32'hbc4a8e2a),
	.w4(32'hbb5fa846),
	.w5(32'hbc2bfdfd),
	.w6(32'hbc05ce91),
	.w7(32'hbb7dec08),
	.w8(32'hbc2f95ec),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e3bb4),
	.w1(32'hbc8d1c6a),
	.w2(32'hbb8396cd),
	.w3(32'hbc3bcc0f),
	.w4(32'h3b13d25a),
	.w5(32'hbb37fe2c),
	.w6(32'hbc2b35ed),
	.w7(32'h3ac2b93a),
	.w8(32'hbb2bf813),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb10d73),
	.w1(32'hbab252e4),
	.w2(32'h3c39d1f0),
	.w3(32'h3b262d68),
	.w4(32'h3b6fac25),
	.w5(32'h3c19fd41),
	.w6(32'h3b8aa365),
	.w7(32'h3bb93fcb),
	.w8(32'hbbe2662c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fcccd),
	.w1(32'hbbe14f4e),
	.w2(32'h3b809027),
	.w3(32'hba7198ac),
	.w4(32'h3be300f8),
	.w5(32'hbaf441f6),
	.w6(32'hbb8ad87d),
	.w7(32'h3a2e509a),
	.w8(32'hbae4608a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7ea38),
	.w1(32'h3bbc17f6),
	.w2(32'h3bd9b091),
	.w3(32'hba74deaf),
	.w4(32'h3b75bd7a),
	.w5(32'hbb35a32c),
	.w6(32'h3b071bd8),
	.w7(32'h3befb89e),
	.w8(32'hbc241246),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e4d67),
	.w1(32'hbc2895bc),
	.w2(32'h3bddbcc5),
	.w3(32'hbbbd8b4d),
	.w4(32'hbb056a24),
	.w5(32'h3ce7eb77),
	.w6(32'hbc6acbe7),
	.w7(32'h3be8debc),
	.w8(32'h3d351063),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbfe1da),
	.w1(32'hbb9d65ee),
	.w2(32'hbcec02f7),
	.w3(32'h3c05abc2),
	.w4(32'hbc960550),
	.w5(32'h3c19d4ec),
	.w6(32'h3bf62814),
	.w7(32'hbd01ef42),
	.w8(32'h3b88f8cb),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b169287),
	.w1(32'h3caeb455),
	.w2(32'hbbd1daff),
	.w3(32'h3b4e0256),
	.w4(32'hbb94dbdc),
	.w5(32'h3c011d52),
	.w6(32'h3cf54f26),
	.w7(32'h3b5dd64c),
	.w8(32'h3b5a2063),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b615213),
	.w1(32'hbc0fe034),
	.w2(32'hbc04c432),
	.w3(32'h3b999de4),
	.w4(32'hba3adcb6),
	.w5(32'h3bb6c336),
	.w6(32'hb91216dc),
	.w7(32'hbc0ce93d),
	.w8(32'h3ca65282),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3234ca),
	.w1(32'hbbb009d2),
	.w2(32'hbc2f9172),
	.w3(32'h3be405c8),
	.w4(32'hbb6ac904),
	.w5(32'h3c18a901),
	.w6(32'hbb734f89),
	.w7(32'hbcb2f4a7),
	.w8(32'hbbbad251),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b037887),
	.w1(32'h3b13ce14),
	.w2(32'h3b80257e),
	.w3(32'hba19c374),
	.w4(32'h3be33a28),
	.w5(32'hbbd00104),
	.w6(32'h3b902aef),
	.w7(32'h3c24804a),
	.w8(32'hbc5fd70d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbe515),
	.w1(32'hbbd5e208),
	.w2(32'h3b769fea),
	.w3(32'hbbac5369),
	.w4(32'h3bdcd3ea),
	.w5(32'hba18fb1a),
	.w6(32'hbbfd88a4),
	.w7(32'h3bf8f45a),
	.w8(32'hbac2e873),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae42d2),
	.w1(32'hbc180387),
	.w2(32'h3b4451b1),
	.w3(32'hbb602200),
	.w4(32'h3c25eca9),
	.w5(32'h3b31a700),
	.w6(32'hb9103b83),
	.w7(32'h3b5844dc),
	.w8(32'hbbac1012),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae19532),
	.w1(32'h3b967d41),
	.w2(32'h3bba7637),
	.w3(32'hbb91ce4f),
	.w4(32'hba8057e5),
	.w5(32'h3c4ba773),
	.w6(32'hbaa1d67f),
	.w7(32'h3b3ff236),
	.w8(32'h3c4e1087),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6372c),
	.w1(32'hbc3532d4),
	.w2(32'h3b0fdec7),
	.w3(32'h3a37d827),
	.w4(32'hbc117208),
	.w5(32'h3bbdf275),
	.w6(32'hbc83ffc1),
	.w7(32'hbc854014),
	.w8(32'h3ca3238a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac11dc8),
	.w1(32'h3b83cfd2),
	.w2(32'hbb221654),
	.w3(32'h3c9df4fd),
	.w4(32'hb89da678),
	.w5(32'hbba9c7de),
	.w6(32'h3b8112b4),
	.w7(32'hbbde1902),
	.w8(32'hbc474483),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b69c4),
	.w1(32'hbc619514),
	.w2(32'hbb4df303),
	.w3(32'hbc806343),
	.w4(32'hbadd62f8),
	.w5(32'hbab6b55b),
	.w6(32'hbca5559a),
	.w7(32'hbc2926e7),
	.w8(32'hbb4995cb),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58a4e4),
	.w1(32'h3bfd61e9),
	.w2(32'h3bea776b),
	.w3(32'hbaa3c037),
	.w4(32'h3b706f01),
	.w5(32'hbc021238),
	.w6(32'hbc9dec48),
	.w7(32'h3b7c6499),
	.w8(32'hbb320713),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c7595),
	.w1(32'h3bdff590),
	.w2(32'hbac6b9cd),
	.w3(32'hbb97fbe4),
	.w4(32'h39ca9d45),
	.w5(32'hba8a2738),
	.w6(32'h3b8bfd3d),
	.w7(32'hbafdfd43),
	.w8(32'h3be82220),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28c690),
	.w1(32'h3b65f3aa),
	.w2(32'hbc0069ce),
	.w3(32'h3b4472dd),
	.w4(32'hb9b2d9c6),
	.w5(32'hbb03b138),
	.w6(32'h3b3166c0),
	.w7(32'hbbcc93e3),
	.w8(32'h3b6033c6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee4cc8),
	.w1(32'h3b94d4f4),
	.w2(32'hbaf5d593),
	.w3(32'h3b8b0bf7),
	.w4(32'h3b875d49),
	.w5(32'hbd064a1d),
	.w6(32'h3bbf0055),
	.w7(32'h3b35ca35),
	.w8(32'hbcf560fa),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbcad57),
	.w1(32'hbb5c5c5e),
	.w2(32'h3c8c3070),
	.w3(32'hbc2ece04),
	.w4(32'h3bbcbd8e),
	.w5(32'h3c05cc68),
	.w6(32'hbb9e7353),
	.w7(32'h3c838e5a),
	.w8(32'h3bd58975),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5e4b9),
	.w1(32'hbbf37108),
	.w2(32'hba8593e6),
	.w3(32'hb92b6c0d),
	.w4(32'hbbf064d7),
	.w5(32'hbd286e41),
	.w6(32'hbcc1f5fa),
	.w7(32'hbcacfeaa),
	.w8(32'hbd4dd810),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce57135),
	.w1(32'h3c27c778),
	.w2(32'h3d4f309f),
	.w3(32'hbc785f25),
	.w4(32'h3cc440e9),
	.w5(32'hbada7f22),
	.w6(32'hbbdc8259),
	.w7(32'h3d705428),
	.w8(32'hbc1856ec),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aa006),
	.w1(32'h3a2729b0),
	.w2(32'h3c21583f),
	.w3(32'hbbd70adf),
	.w4(32'h3a93ada6),
	.w5(32'hbbf5cb28),
	.w6(32'hbc0bf10e),
	.w7(32'hbb25d872),
	.w8(32'hbc9dd025),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c5f04),
	.w1(32'hbab23757),
	.w2(32'h3c8a605e),
	.w3(32'hbca34fc4),
	.w4(32'h3b12630c),
	.w5(32'h39af79e1),
	.w6(32'hbcabd52f),
	.w7(32'h3c69d9df),
	.w8(32'hbc345f71),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b0cec),
	.w1(32'hbbdb54eb),
	.w2(32'hbaffec82),
	.w3(32'hbad68f54),
	.w4(32'h3a708ebd),
	.w5(32'h3ca56911),
	.w6(32'h3abc977a),
	.w7(32'h3b8ddf3c),
	.w8(32'h3cf5886d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8b485),
	.w1(32'hbbb6af53),
	.w2(32'hbc5815b1),
	.w3(32'h3cb9cb4d),
	.w4(32'h3ba0e30c),
	.w5(32'hbbf67d9c),
	.w6(32'h3ba3a2b3),
	.w7(32'hbc8cdb53),
	.w8(32'hbb50bb45),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7c2c6),
	.w1(32'hbb8f01e6),
	.w2(32'h39a807c6),
	.w3(32'hbb9829c0),
	.w4(32'hbb8fe64f),
	.w5(32'hbd03f443),
	.w6(32'h3c2ede4d),
	.w7(32'h3c2410dd),
	.w8(32'hbd255738),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5a269),
	.w1(32'h3c00d895),
	.w2(32'h3ce642a7),
	.w3(32'hbc4198fb),
	.w4(32'h3be93d62),
	.w5(32'h39d69ad3),
	.w6(32'hbbc0cf70),
	.w7(32'h3d0e6fce),
	.w8(32'hbc095cb5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe3ce6),
	.w1(32'hbc3eab8c),
	.w2(32'h3b8cdc71),
	.w3(32'hbc9c5aa9),
	.w4(32'h3b781a60),
	.w5(32'h3c63fd68),
	.w6(32'hbc6fdc27),
	.w7(32'h3b452120),
	.w8(32'h3c49b9c2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf469e),
	.w1(32'hbb78c912),
	.w2(32'hb96db751),
	.w3(32'h3b393747),
	.w4(32'h3b3fe5d6),
	.w5(32'hbb5ccda8),
	.w6(32'hbbb55143),
	.w7(32'hbc3b7bba),
	.w8(32'hbbf990a6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb589c34),
	.w1(32'h3a2de67f),
	.w2(32'h3bee6ffa),
	.w3(32'hbc00d248),
	.w4(32'hbb039323),
	.w5(32'h3c0e19d0),
	.w6(32'hbb9ab58d),
	.w7(32'h3806a25e),
	.w8(32'h3c6f0b72),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c354280),
	.w1(32'hbc1b2e2c),
	.w2(32'hbc49277c),
	.w3(32'h3bb6c6c5),
	.w4(32'h3b41e717),
	.w5(32'hbacefd4f),
	.w6(32'hbaa12905),
	.w7(32'hbbd4b404),
	.w8(32'h3c03e577),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca00d2),
	.w1(32'hbba562d1),
	.w2(32'hba4179a5),
	.w3(32'hbbad91b9),
	.w4(32'hbc7403c9),
	.w5(32'h3a7de4d2),
	.w6(32'hbb80f42f),
	.w7(32'hbc9c8003),
	.w8(32'hbac2890b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f6c29),
	.w1(32'hba8daa86),
	.w2(32'hba89bae9),
	.w3(32'h3b3338b1),
	.w4(32'h3b9cae48),
	.w5(32'h3cb7b1ff),
	.w6(32'h3bdcb5e7),
	.w7(32'h3bc5b4d6),
	.w8(32'h3d0ae403),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97b2ad),
	.w1(32'h3a8c3714),
	.w2(32'hbc945343),
	.w3(32'h3c7f1c4d),
	.w4(32'hbb99fc8a),
	.w5(32'h3c71ab77),
	.w6(32'h3bb00f87),
	.w7(32'hbcce5e92),
	.w8(32'h3c4f1801),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c549c),
	.w1(32'hbc4311cb),
	.w2(32'h3bb5660d),
	.w3(32'h3ae12a75),
	.w4(32'hb8a1cfa1),
	.w5(32'h3b1be2c5),
	.w6(32'hbb9eb30a),
	.w7(32'h3bc05792),
	.w8(32'h3c3d6d2b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39698da6),
	.w1(32'h3965ec4f),
	.w2(32'h3b417ca8),
	.w3(32'h3b900cd1),
	.w4(32'h3ba20c33),
	.w5(32'hbb05d09d),
	.w6(32'h3bfee31d),
	.w7(32'h3c12bf6e),
	.w8(32'hbc8cb30e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8ee38),
	.w1(32'hbc722396),
	.w2(32'h3b41bd1e),
	.w3(32'hbc9b4e79),
	.w4(32'hbaf0049e),
	.w5(32'hb9ff8c99),
	.w6(32'hbce5d269),
	.w7(32'hbb38f079),
	.w8(32'h3c063bd7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb309c7f),
	.w1(32'hbc22300e),
	.w2(32'hbb3bfe54),
	.w3(32'hbc6ed557),
	.w4(32'h3c3c8add),
	.w5(32'h3af6e3aa),
	.w6(32'hbc85bb40),
	.w7(32'hbc1b3d30),
	.w8(32'h3ba612a6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03adb9),
	.w1(32'hbb869dee),
	.w2(32'hbb6521d4),
	.w3(32'hbbee7ef7),
	.w4(32'hbc12aa17),
	.w5(32'h3ba43e0b),
	.w6(32'hbc1cf6a5),
	.w7(32'hbc177162),
	.w8(32'h3ab7b05b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b8053),
	.w1(32'hbbcc1d73),
	.w2(32'h3b126ea3),
	.w3(32'hbbdc0a2e),
	.w4(32'h3bd43844),
	.w5(32'h3c8449c6),
	.w6(32'hbc23b482),
	.w7(32'hbb70480f),
	.w8(32'hbc0f5fd0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e484b),
	.w1(32'h3b9b85d2),
	.w2(32'h3c4c393d),
	.w3(32'h3c1478c9),
	.w4(32'hbcdc7022),
	.w5(32'hbac64ae2),
	.w6(32'h3c312144),
	.w7(32'h3c7063d3),
	.w8(32'hbc92550b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36895b),
	.w1(32'hbc084762),
	.w2(32'hbc2af4dd),
	.w3(32'hbb729fcb),
	.w4(32'h3b0e799a),
	.w5(32'hbbd73181),
	.w6(32'h3c559ee3),
	.w7(32'h3c5074c5),
	.w8(32'hbc18bcbb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c3866),
	.w1(32'hbb46761d),
	.w2(32'h3bb692c7),
	.w3(32'hbc5f2f52),
	.w4(32'h3c469ace),
	.w5(32'hba010620),
	.w6(32'hbc878d74),
	.w7(32'h3a382f5d),
	.w8(32'hb9d78958),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b76e77),
	.w1(32'hba3c8f35),
	.w2(32'hba365de9),
	.w3(32'hba5697c6),
	.w4(32'hba0805ed),
	.w5(32'hba0f066d),
	.w6(32'hba4d0949),
	.w7(32'hba37eace),
	.w8(32'hba384064),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9917d20),
	.w1(32'h398b9fe1),
	.w2(32'h37592636),
	.w3(32'h3983572a),
	.w4(32'h39aca349),
	.w5(32'h3a915db8),
	.w6(32'h3a8b9262),
	.w7(32'h3a3c9e40),
	.w8(32'h3af77cb6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dedb3),
	.w1(32'h39d8fccf),
	.w2(32'h39ff3347),
	.w3(32'h3a866c50),
	.w4(32'h39bd8c9a),
	.w5(32'h39b5b3ca),
	.w6(32'h3abb25a6),
	.w7(32'h3a880354),
	.w8(32'hb9810f09),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385fb385),
	.w1(32'h3987d5a6),
	.w2(32'hb8a2fd13),
	.w3(32'h3867d6c3),
	.w4(32'h3a82844c),
	.w5(32'h3a05b787),
	.w6(32'h3afc7747),
	.w7(32'h3a68d7ac),
	.w8(32'h394baae9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad9558),
	.w1(32'h38f505e4),
	.w2(32'h39c38207),
	.w3(32'h398bc553),
	.w4(32'h39f600d6),
	.w5(32'h3a119e32),
	.w6(32'h390c4602),
	.w7(32'h399787ca),
	.w8(32'h3ae9cf88),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ef854),
	.w1(32'h373ab42f),
	.w2(32'h393f18b3),
	.w3(32'h3a93669e),
	.w4(32'hb7978e30),
	.w5(32'h39da6a69),
	.w6(32'h3a918ef8),
	.w7(32'h3a1e6369),
	.w8(32'h3a1cfa0a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e099a5),
	.w1(32'hb94d5127),
	.w2(32'hba36d0ae),
	.w3(32'hbaa2bce5),
	.w4(32'hbac74ded),
	.w5(32'hb82aa674),
	.w6(32'hb9e306ca),
	.w7(32'hb9738fba),
	.w8(32'hb7e1c7e3),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdbb61),
	.w1(32'hb88f2fc6),
	.w2(32'h3a877c01),
	.w3(32'h3867cf73),
	.w4(32'h3a39c720),
	.w5(32'h3a67103f),
	.w6(32'h38b3fe63),
	.w7(32'h3a618e33),
	.w8(32'hb9fe2151),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955c52b),
	.w1(32'h399df75c),
	.w2(32'h39c495bb),
	.w3(32'h3995f828),
	.w4(32'h3a39b571),
	.w5(32'hba424238),
	.w6(32'hb9ae4778),
	.w7(32'h395fe41c),
	.w8(32'hba2192e2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1de3dc),
	.w1(32'hb95cece1),
	.w2(32'hb734a52d),
	.w3(32'hba1222b6),
	.w4(32'hb996c9a3),
	.w5(32'hbaa8cf25),
	.w6(32'h393b842e),
	.w7(32'h39a52b75),
	.w8(32'hba963586),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48107c),
	.w1(32'hba8a5d0e),
	.w2(32'hba66ca9c),
	.w3(32'hbab9b6e8),
	.w4(32'hba8b7ab8),
	.w5(32'hb9f51d23),
	.w6(32'hba86a092),
	.w7(32'hba8efd8a),
	.w8(32'h382994af),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e20da),
	.w1(32'hba3b1419),
	.w2(32'hbaa6503c),
	.w3(32'hb995f199),
	.w4(32'hba87ccb7),
	.w5(32'hb92da7cd),
	.w6(32'hb9fcf765),
	.w7(32'hba5b5bde),
	.w8(32'hb9d4a4b3),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b00963),
	.w1(32'hb97b021b),
	.w2(32'hba95deeb),
	.w3(32'hba25dc79),
	.w4(32'h3980b3a2),
	.w5(32'h39ef8cf7),
	.w6(32'hba24a5d1),
	.w7(32'hba3be05c),
	.w8(32'hb8727dfc),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92168b),
	.w1(32'hb8e88cbd),
	.w2(32'hb95dbaa1),
	.w3(32'h3a459243),
	.w4(32'h3a2d6803),
	.w5(32'h3a9749d9),
	.w6(32'h3a0bdb79),
	.w7(32'h39e5eee6),
	.w8(32'h3a12d108),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2145cd),
	.w1(32'hb926dacb),
	.w2(32'hb7a01132),
	.w3(32'h3a2adac5),
	.w4(32'h3a7f0f2d),
	.w5(32'h398d245b),
	.w6(32'hb9930835),
	.w7(32'h39084ea9),
	.w8(32'hb7c1bbc3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38590d49),
	.w1(32'h3a3a84b7),
	.w2(32'h3a38e285),
	.w3(32'h3a119e17),
	.w4(32'h3a5ef1b9),
	.w5(32'hb9a95012),
	.w6(32'h3a823984),
	.w7(32'h393c66d0),
	.w8(32'hb9e66493),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba803ad7),
	.w1(32'h38a9cbd8),
	.w2(32'hb9bbd559),
	.w3(32'hb93aabad),
	.w4(32'h3a1ab1ad),
	.w5(32'h39b52e2d),
	.w6(32'hb996f95f),
	.w7(32'h39ad5174),
	.w8(32'hb89b1d04),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfc9c7),
	.w1(32'hb9880580),
	.w2(32'hb9b21ef9),
	.w3(32'hb9296099),
	.w4(32'h3926ef21),
	.w5(32'h3a767f8f),
	.w6(32'h3aabd50f),
	.w7(32'h38f3efc1),
	.w8(32'h3a489e94),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a408124),
	.w1(32'h397f0b4a),
	.w2(32'h38a16bc6),
	.w3(32'h39d37f18),
	.w4(32'h3a53ab7c),
	.w5(32'hb7c7e390),
	.w6(32'h3987f9dd),
	.w7(32'h3a1af229),
	.w8(32'h39e6d998),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390aa048),
	.w1(32'hb9934dea),
	.w2(32'hb936d7b1),
	.w3(32'hba13e765),
	.w4(32'hba476da6),
	.w5(32'hba4f9601),
	.w6(32'h3a01d87d),
	.w7(32'hba201f54),
	.w8(32'hb94542c8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba639cc4),
	.w1(32'hba3604f1),
	.w2(32'hba08e2fb),
	.w3(32'hba2216e3),
	.w4(32'hba11261f),
	.w5(32'hba50fda3),
	.w6(32'hb90e8399),
	.w7(32'h39b48a9c),
	.w8(32'hb91e1516),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca980f),
	.w1(32'hbae2e750),
	.w2(32'hbac4936d),
	.w3(32'hb9e0fba6),
	.w4(32'hba1ce8c8),
	.w5(32'hb74b3d07),
	.w6(32'hba0378fe),
	.w7(32'hba482501),
	.w8(32'h390b1bd6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf9619),
	.w1(32'hb9eb4a4f),
	.w2(32'hb974b913),
	.w3(32'hb8edf2e3),
	.w4(32'hb93d557c),
	.w5(32'hb8f97b0a),
	.w6(32'h3a7645cb),
	.w7(32'h39a1588c),
	.w8(32'h39e71e10),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60951c),
	.w1(32'hb9392f9a),
	.w2(32'hb9ce13a4),
	.w3(32'h3a012a9f),
	.w4(32'h3966b304),
	.w5(32'h3a820315),
	.w6(32'h39b12cb3),
	.w7(32'hb8b4154f),
	.w8(32'hb84c16d2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989637c),
	.w1(32'h39afee02),
	.w2(32'h3999e2c7),
	.w3(32'h3ae87edf),
	.w4(32'h3a6b5eb2),
	.w5(32'hba50d22b),
	.w6(32'h3a9d8eb7),
	.w7(32'hb9edc52a),
	.w8(32'hb9b4e772),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a093b74),
	.w1(32'hb89b1045),
	.w2(32'hb9bae76c),
	.w3(32'hb9101782),
	.w4(32'hb8b6b6c2),
	.w5(32'h390b49d4),
	.w6(32'hb9fe9d8d),
	.w7(32'hb9fb41d7),
	.w8(32'h3aac14cb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b6d6f9),
	.w1(32'h3a1231b9),
	.w2(32'hb7a1d975),
	.w3(32'h39921951),
	.w4(32'h3a1c0419),
	.w5(32'hb928bf74),
	.w6(32'h3b2aa2df),
	.w7(32'h3a7402dc),
	.w8(32'h389714bd),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bf3b45),
	.w1(32'h376bd5e6),
	.w2(32'h3800e39b),
	.w3(32'h3a28c27e),
	.w4(32'h3a9003bb),
	.w5(32'hba941792),
	.w6(32'h3a2b7549),
	.w7(32'h3a3a2b54),
	.w8(32'hba5d2598),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df7101),
	.w1(32'h37cdb8ea),
	.w2(32'hb95ebdfb),
	.w3(32'hba8d6a0c),
	.w4(32'hba131f14),
	.w5(32'h39ef00f8),
	.w6(32'hb9c96736),
	.w7(32'hb9cbcf10),
	.w8(32'h39b543a9),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39200531),
	.w1(32'hb7a5175d),
	.w2(32'hba4cb708),
	.w3(32'h39cc5570),
	.w4(32'hb7a2528c),
	.w5(32'hba28e3ca),
	.w6(32'h39a4fbea),
	.w7(32'hb9b59569),
	.w8(32'hb8db632f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule