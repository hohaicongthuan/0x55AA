module layer_6_featuremap_109(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09244b),
	.w1(32'hbb614e47),
	.w2(32'hbb6a1ed8),
	.w3(32'h35f26caf),
	.w4(32'h3a98f760),
	.w5(32'h3af792b8),
	.w6(32'hbad8147d),
	.w7(32'hba434d94),
	.w8(32'hb9e86bcd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac34823),
	.w1(32'hbbcaad39),
	.w2(32'hbbb892cc),
	.w3(32'h3ad63013),
	.w4(32'h3b06da6d),
	.w5(32'h3b7d0c37),
	.w6(32'h3c0474f7),
	.w7(32'h3c40a23a),
	.w8(32'h3c892a3a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b175),
	.w1(32'h3baffb9d),
	.w2(32'hb947f5e3),
	.w3(32'h3a93aa90),
	.w4(32'hbafc173c),
	.w5(32'hb9f41d42),
	.w6(32'h3c1aedb0),
	.w7(32'hbb282fd5),
	.w8(32'hbbd33ccc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd1c674),
	.w1(32'hbc32589c),
	.w2(32'hbc12490b),
	.w3(32'hbb9e6c6a),
	.w4(32'hba7626c1),
	.w5(32'hba2aaf1d),
	.w6(32'hba8cf542),
	.w7(32'h3be9a831),
	.w8(32'h3c129b6b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2595eb),
	.w1(32'hba9fb212),
	.w2(32'hbb8451bd),
	.w3(32'h3ad2957a),
	.w4(32'h3ba99ccd),
	.w5(32'h3c3e1185),
	.w6(32'hbb2336db),
	.w7(32'h3aac85e1),
	.w8(32'hba40a5b5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebc743),
	.w1(32'h3c0e28d4),
	.w2(32'h3ae8d201),
	.w3(32'h3bd35188),
	.w4(32'h3ab1440b),
	.w5(32'hb9ca7633),
	.w6(32'h3b5ba8d6),
	.w7(32'hbb7d2b3e),
	.w8(32'hbb88c535),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d229a),
	.w1(32'h39a0849a),
	.w2(32'h3c07cbcc),
	.w3(32'hbbd7d394),
	.w4(32'hba5803ea),
	.w5(32'h3b2bbc2d),
	.w6(32'hbb4d8618),
	.w7(32'h3c03b736),
	.w8(32'h3c304884),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05b350),
	.w1(32'h3c2c7ee9),
	.w2(32'h3c889521),
	.w3(32'h39367156),
	.w4(32'hb99bd9c0),
	.w5(32'h3b3eea55),
	.w6(32'h3ba4dabf),
	.w7(32'hbb265314),
	.w8(32'hbae1dbbb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc98764),
	.w1(32'h3b695b10),
	.w2(32'h39622a96),
	.w3(32'hbaec4aad),
	.w4(32'h3aa0a177),
	.w5(32'h3b4aedf1),
	.w6(32'hbb9c58ef),
	.w7(32'h3b458306),
	.w8(32'h3c8aa9bf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4e7ee),
	.w1(32'h3c3a8273),
	.w2(32'h3bfa81ea),
	.w3(32'hba3b660b),
	.w4(32'hbc239f63),
	.w5(32'hbc1a4017),
	.w6(32'h3b0f7700),
	.w7(32'hbbf2a601),
	.w8(32'hbbc3b230),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f095f),
	.w1(32'h3ca2eca1),
	.w2(32'h3bba1288),
	.w3(32'h3c428b6c),
	.w4(32'h3c24427a),
	.w5(32'h3c0e7b31),
	.w6(32'h3cc96137),
	.w7(32'h3c91a2a0),
	.w8(32'h3c62447b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2de74),
	.w1(32'hbaf30aa9),
	.w2(32'hbb595ef7),
	.w3(32'hbb44079a),
	.w4(32'hbb72e947),
	.w5(32'hbb39ffe9),
	.w6(32'hbb5e4172),
	.w7(32'hbb4b187d),
	.w8(32'hbb6ba845),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4de817),
	.w1(32'h3b0e116a),
	.w2(32'hba86014c),
	.w3(32'h3b3bcd86),
	.w4(32'h398af065),
	.w5(32'h3bd66c29),
	.w6(32'h3ae0338e),
	.w7(32'h3a27edb4),
	.w8(32'h3bfe803a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dfb74),
	.w1(32'hbaac3057),
	.w2(32'hba53a7b7),
	.w3(32'h3c540dab),
	.w4(32'h3c9d2bc8),
	.w5(32'h3ccf3a92),
	.w6(32'h3c0fa741),
	.w7(32'h3c4063ca),
	.w8(32'h3ca02a15),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fb750),
	.w1(32'hbc3e257b),
	.w2(32'hbaaf03dd),
	.w3(32'hbb968a5f),
	.w4(32'h3b772e7c),
	.w5(32'h3bcd0747),
	.w6(32'hbba570e8),
	.w7(32'h3c40e753),
	.w8(32'h3c466a39),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd37bf),
	.w1(32'h3a0b680b),
	.w2(32'hbb0d9688),
	.w3(32'h3ae1fa78),
	.w4(32'hba713ae7),
	.w5(32'hbb3bdb1d),
	.w6(32'h3baa1025),
	.w7(32'hb8bbbe69),
	.w8(32'hba073fe2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf0145),
	.w1(32'h3c5e0cfd),
	.w2(32'h3c39d653),
	.w3(32'h3c19d96c),
	.w4(32'h3cb39822),
	.w5(32'h3c44839d),
	.w6(32'h3c0d4bd0),
	.w7(32'h3c72de69),
	.w8(32'h3c51a94e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f39a8),
	.w1(32'h3b3ccf49),
	.w2(32'h3b12f579),
	.w3(32'hb928822a),
	.w4(32'hbb277deb),
	.w5(32'hbb2ccf8f),
	.w6(32'h3b3cc18f),
	.w7(32'h3ad8a717),
	.w8(32'h3a511339),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c0886),
	.w1(32'h39e7055f),
	.w2(32'h36e1276b),
	.w3(32'h39fafc9d),
	.w4(32'h3a70d5ce),
	.w5(32'hbb3eee97),
	.w6(32'hb9de275b),
	.w7(32'h39dccd4f),
	.w8(32'hbaf8aae0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaba50),
	.w1(32'hbab61b74),
	.w2(32'h3bd21abc),
	.w3(32'h3b70b1a4),
	.w4(32'h3882ebf4),
	.w5(32'h3bf1e998),
	.w6(32'h3be8a1e6),
	.w7(32'h3b818ac3),
	.w8(32'h3c5d1570),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d5bf1),
	.w1(32'hbb4c19c1),
	.w2(32'hba0918ba),
	.w3(32'h3ab6882b),
	.w4(32'h3bc991a5),
	.w5(32'h3bf96cde),
	.w6(32'h3b95c0c5),
	.w7(32'h3c0fab33),
	.w8(32'h3c39bfbf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81fdde),
	.w1(32'h3a55a836),
	.w2(32'h3b768717),
	.w3(32'h3c10da64),
	.w4(32'h3c9af179),
	.w5(32'h3c8f662e),
	.w6(32'h3ca7aa0c),
	.w7(32'h3cf026c9),
	.w8(32'h3d046b15),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca553b8),
	.w1(32'hbcaf07bb),
	.w2(32'hbc8bdad9),
	.w3(32'hbca7ac96),
	.w4(32'hbc4d1469),
	.w5(32'h3a40057f),
	.w6(32'hbcac148e),
	.w7(32'hbc8913cd),
	.w8(32'h3c0cc715),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b733c2e),
	.w1(32'hbaa20815),
	.w2(32'h3bbeecf2),
	.w3(32'h3c43611b),
	.w4(32'h3c7854d7),
	.w5(32'h3c911343),
	.w6(32'h3ce180eb),
	.w7(32'h3d157d21),
	.w8(32'h3cf6c464),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7dfe2),
	.w1(32'hbc032341),
	.w2(32'hbc98d771),
	.w3(32'hbcbe3185),
	.w4(32'hbb16f4db),
	.w5(32'hbb2b6441),
	.w6(32'hbc4b4115),
	.w7(32'hbac52d7b),
	.w8(32'h3aa8e5e4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850294),
	.w1(32'h3be571c6),
	.w2(32'h395a81ef),
	.w3(32'hbc1031f0),
	.w4(32'hbb73bc17),
	.w5(32'h3b2bda64),
	.w6(32'hbb8869b8),
	.w7(32'hbb8f52e9),
	.w8(32'h3b84d8f0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed44cf),
	.w1(32'h397b2644),
	.w2(32'h3b72dce7),
	.w3(32'h3c3e2502),
	.w4(32'h3b254949),
	.w5(32'h3c014fe3),
	.w6(32'h3c7df819),
	.w7(32'h3c7dc6b0),
	.w8(32'h3c916a41),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0626f),
	.w1(32'h3b53a56d),
	.w2(32'h3bb8d5be),
	.w3(32'h3b001ff1),
	.w4(32'h3b496245),
	.w5(32'h3ac472a0),
	.w6(32'h3b5600be),
	.w7(32'h3bedc992),
	.w8(32'h3b9eb70a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b18f6),
	.w1(32'hbbfb9b8f),
	.w2(32'h39b44970),
	.w3(32'hba28ebf6),
	.w4(32'h3b61cbd5),
	.w5(32'h3baa6377),
	.w6(32'hbb3ea7b2),
	.w7(32'h3b718419),
	.w8(32'h3bca77c4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab735ca),
	.w1(32'hb911ea4b),
	.w2(32'h3b0e4e5a),
	.w3(32'hbc87ee07),
	.w4(32'hbbc13e38),
	.w5(32'hbb05b287),
	.w6(32'hbbc44063),
	.w7(32'hb9330c8c),
	.w8(32'h3b8e6ee2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba763fe),
	.w1(32'hbc02fc0d),
	.w2(32'hbc9b7bc1),
	.w3(32'hba21ad0d),
	.w4(32'hb99badea),
	.w5(32'h3b7fc1d0),
	.w6(32'h3ba2cc70),
	.w7(32'h3a937468),
	.w8(32'h3b8c3cdc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc86717),
	.w1(32'h3c2ee475),
	.w2(32'hbb3c04be),
	.w3(32'h3c0559d9),
	.w4(32'h3c27b0ae),
	.w5(32'h3c0b8607),
	.w6(32'h3bc21b46),
	.w7(32'h3bdaa58f),
	.w8(32'hb9a19be7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53986a),
	.w1(32'hbb28d009),
	.w2(32'h3c0addd7),
	.w3(32'hbc182713),
	.w4(32'h39f59916),
	.w5(32'h3aecbab5),
	.w6(32'h3b6b0fe5),
	.w7(32'h3c769276),
	.w8(32'h3be64a58),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39be59),
	.w1(32'h3bb610e4),
	.w2(32'h3c5c478b),
	.w3(32'h3ba165b8),
	.w4(32'h3bcfaa0f),
	.w5(32'hbae76cdd),
	.w6(32'h3c05e712),
	.w7(32'h3beae699),
	.w8(32'h3c188ae2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28dc49),
	.w1(32'hba2b74e6),
	.w2(32'hbb5ff8c0),
	.w3(32'hba937182),
	.w4(32'hbb524b41),
	.w5(32'hbb57a320),
	.w6(32'hbb170b0a),
	.w7(32'hbb837c45),
	.w8(32'hbb6780f3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc20393),
	.w1(32'h3b68121b),
	.w2(32'hbc0ca61f),
	.w3(32'hbc1f1f68),
	.w4(32'hbbb8841b),
	.w5(32'hbc18d646),
	.w6(32'hb9fa38b5),
	.w7(32'hbbcea393),
	.w8(32'hbbb81ddb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd29967),
	.w1(32'h3b8b6198),
	.w2(32'h3ae38374),
	.w3(32'h3b718660),
	.w4(32'h3b878117),
	.w5(32'h3ba56655),
	.w6(32'h3abd7d2b),
	.w7(32'hba235f87),
	.w8(32'h3a47584f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb976d7),
	.w1(32'hba4c5983),
	.w2(32'h3b440651),
	.w3(32'h39280332),
	.w4(32'h3bd5d6c2),
	.w5(32'h3b87f477),
	.w6(32'h3b279fa3),
	.w7(32'h3be1c7ab),
	.w8(32'h3bb0dfdf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e3976),
	.w1(32'h3c0a37e8),
	.w2(32'h3b48846a),
	.w3(32'h3b06298e),
	.w4(32'hbb4c159d),
	.w5(32'h3b932bbf),
	.w6(32'h3abf5770),
	.w7(32'hbaad5911),
	.w8(32'h3b45d7e9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba35d5e),
	.w1(32'h3bbbfe7f),
	.w2(32'h3a3cf6c9),
	.w3(32'h3d00b26d),
	.w4(32'h3cc2bf2b),
	.w5(32'h3cf64097),
	.w6(32'h3d1322c6),
	.w7(32'h3d201b9b),
	.w8(32'h3d50bbfe),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2eba87),
	.w1(32'h3c386d7b),
	.w2(32'h3c20de5a),
	.w3(32'h3c55a759),
	.w4(32'h3c5e9a62),
	.w5(32'h3b8e1361),
	.w6(32'h3c2bd32e),
	.w7(32'h3c93499f),
	.w8(32'h3bb0cded),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf5d15),
	.w1(32'h3a932c13),
	.w2(32'h3ba621ac),
	.w3(32'h3b813048),
	.w4(32'h3bd0b421),
	.w5(32'h3c0072b2),
	.w6(32'h3b86d961),
	.w7(32'h3c2b3578),
	.w8(32'h3c51f1ad),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe6d77),
	.w1(32'hbb283067),
	.w2(32'hbba5b1dc),
	.w3(32'h3a44f150),
	.w4(32'h3ab8487c),
	.w5(32'h3bb1e09a),
	.w6(32'hbb162ef3),
	.w7(32'hbb314b93),
	.w8(32'h3b4e570e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d5a49),
	.w1(32'hbb050373),
	.w2(32'hbc2ecf27),
	.w3(32'hb9060927),
	.w4(32'h3afe6238),
	.w5(32'hbb49f961),
	.w6(32'h39b2313b),
	.w7(32'h3aa7c8f8),
	.w8(32'h3b7d6843),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc073936),
	.w1(32'hbc06e70e),
	.w2(32'hbbb8864e),
	.w3(32'h3bad20fc),
	.w4(32'h3bc76feb),
	.w5(32'h3bb6e6f4),
	.w6(32'h3c1255b9),
	.w7(32'h3bfbe394),
	.w8(32'h3c0b888b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cc20f),
	.w1(32'h3c0995b3),
	.w2(32'hbc02e17b),
	.w3(32'hbc0100ac),
	.w4(32'hbbad941c),
	.w5(32'hbc09c813),
	.w6(32'h3b178457),
	.w7(32'hbc27eeee),
	.w8(32'hbc2b602c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5ce2b),
	.w1(32'hbc5353fd),
	.w2(32'hbc830de4),
	.w3(32'h3a96b0c7),
	.w4(32'hbb5213c2),
	.w5(32'h3cbfc6b5),
	.w6(32'hbb0706ba),
	.w7(32'h3a9707a1),
	.w8(32'h3d062122),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8ca95),
	.w1(32'hb981a19b),
	.w2(32'h3b80d9fc),
	.w3(32'hbc00bd05),
	.w4(32'hba760523),
	.w5(32'hbb60587a),
	.w6(32'hbc014ccf),
	.w7(32'h37d27e2a),
	.w8(32'h3b263001),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02467f),
	.w1(32'hba03d8df),
	.w2(32'hbb9666c4),
	.w3(32'h3c49e28a),
	.w4(32'h3c4d174b),
	.w5(32'h3c3ac10a),
	.w6(32'h3c10afbd),
	.w7(32'h3c120904),
	.w8(32'h3bcad78c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394fe7ba),
	.w1(32'h3bd021e4),
	.w2(32'h3af232f4),
	.w3(32'hbb8ac24f),
	.w4(32'hbaeda07f),
	.w5(32'hbb34c784),
	.w6(32'h3b096494),
	.w7(32'hba810379),
	.w8(32'h39bf0ab5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1889b2),
	.w1(32'h3b9f4c81),
	.w2(32'h3ba2d6ff),
	.w3(32'h3a829994),
	.w4(32'h3ba46ab3),
	.w5(32'h3c6a228f),
	.w6(32'h3b49f219),
	.w7(32'h3c3a135c),
	.w8(32'h3cc7763a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca48a16),
	.w1(32'h3ac0beb3),
	.w2(32'h3bfac3cb),
	.w3(32'h3be4a444),
	.w4(32'h3c382198),
	.w5(32'h3c42ec1f),
	.w6(32'h3bdb9c0c),
	.w7(32'h3c52b122),
	.w8(32'h3c7686c7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d2038),
	.w1(32'hbb4c40f6),
	.w2(32'h3bcfe1ea),
	.w3(32'h3bc079c5),
	.w4(32'h3c23e1bc),
	.w5(32'h3c6e6d88),
	.w6(32'h3ac4c844),
	.w7(32'h3c17ab6a),
	.w8(32'h3c6d6960),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84ccca),
	.w1(32'hbc681c1a),
	.w2(32'hbbc2f348),
	.w3(32'h3ba8f5f3),
	.w4(32'h3c9d96de),
	.w5(32'h3ca34b8d),
	.w6(32'h3beab475),
	.w7(32'h3cb65f5d),
	.w8(32'h3cb552dd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c8b7c),
	.w1(32'hbadae057),
	.w2(32'h3aa501a1),
	.w3(32'h3b582a0e),
	.w4(32'h3c12d43a),
	.w5(32'h3c460b4e),
	.w6(32'h3b8f1be8),
	.w7(32'h3c8e7b4f),
	.w8(32'h3cc055ed),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9df97e),
	.w1(32'hba5b6321),
	.w2(32'hbcd2bfa7),
	.w3(32'hbc600614),
	.w4(32'hbb560237),
	.w5(32'hbc1f69a4),
	.w6(32'hbb9b7077),
	.w7(32'hbbb4b18d),
	.w8(32'hbcb252e5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc47152),
	.w1(32'h398708bf),
	.w2(32'h3c088fb3),
	.w3(32'h3c1cf59a),
	.w4(32'h3c621ce6),
	.w5(32'h3c751348),
	.w6(32'h3c01d58b),
	.w7(32'h3c755b13),
	.w8(32'h3c7de9f6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4da587),
	.w1(32'h3c74a391),
	.w2(32'hbc87ce81),
	.w3(32'h3ba6d52f),
	.w4(32'hbc1c5f2e),
	.w5(32'hba37ccd0),
	.w6(32'h3c661aa6),
	.w7(32'hbc9cbfde),
	.w8(32'h3b3d7ad4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc891365),
	.w1(32'hbbd424a0),
	.w2(32'hbc2cb7d7),
	.w3(32'hbba03990),
	.w4(32'hbb8fc54d),
	.w5(32'hbbd47448),
	.w6(32'h39b3211f),
	.w7(32'hbb2154b0),
	.w8(32'hbbb40796),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcef270a),
	.w1(32'hbc811cd6),
	.w2(32'hbd00fc52),
	.w3(32'hbca083df),
	.w4(32'hbb9c2d3a),
	.w5(32'h3aec8004),
	.w6(32'hbbd8ca2c),
	.w7(32'hbba09534),
	.w8(32'h3c54af87),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d59b8ea),
	.w1(32'h3ca338e6),
	.w2(32'h3c6a25d2),
	.w3(32'hbb19ee59),
	.w4(32'h3b5aa621),
	.w5(32'h3c506773),
	.w6(32'hbc4b8b60),
	.w7(32'hbc3823ce),
	.w8(32'hbbc1e65b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce88e4d),
	.w1(32'hbc946dca),
	.w2(32'hbd0983cb),
	.w3(32'hbc8e6960),
	.w4(32'hbcbbb7f6),
	.w5(32'h3aa8a57c),
	.w6(32'hbc0efbe3),
	.w7(32'hbce4c08c),
	.w8(32'h3d297c87),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1693db),
	.w1(32'h3c50889c),
	.w2(32'hbcb8d29e),
	.w3(32'hbcca9773),
	.w4(32'hbc27b762),
	.w5(32'h3bd2d2ef),
	.w6(32'hbced4789),
	.w7(32'hbd27c535),
	.w8(32'h3cb28f67),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d15e657),
	.w1(32'hbb95d93c),
	.w2(32'hba87793d),
	.w3(32'hbaa56fb4),
	.w4(32'hba530ee2),
	.w5(32'h3a79ac4b),
	.w6(32'h3aa305b5),
	.w7(32'hbb958d02),
	.w8(32'h3b3133f8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule