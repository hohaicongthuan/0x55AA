module layer_8_featuremap_121(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b65bf),
	.w1(32'hbcf2f420),
	.w2(32'hbc0982ce),
	.w3(32'h3af34035),
	.w4(32'hbc3a9343),
	.w5(32'h3c478e9f),
	.w6(32'hbc5dbba7),
	.w7(32'hbcbf7172),
	.w8(32'h3c6e1ba8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca14374),
	.w1(32'h3d082fc9),
	.w2(32'h3c4d7cc9),
	.w3(32'h3c81304e),
	.w4(32'h3c55bcc6),
	.w5(32'h3c0b37c0),
	.w6(32'h3d4d34b4),
	.w7(32'h3d101b83),
	.w8(32'hbca7fbdc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7b6d9),
	.w1(32'hbb04a125),
	.w2(32'h393bb582),
	.w3(32'h3b10b596),
	.w4(32'h3b7ebaee),
	.w5(32'h3bddd025),
	.w6(32'hbc227c5a),
	.w7(32'h3c17b30b),
	.w8(32'hbbbbc3d6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0d0ea),
	.w1(32'hbc410be0),
	.w2(32'hbca88af0),
	.w3(32'h3b4ceaee),
	.w4(32'hbc56e100),
	.w5(32'h3b9ee06b),
	.w6(32'h3bd80760),
	.w7(32'hbc294ad2),
	.w8(32'hbc1e1f2d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8df53e),
	.w1(32'h3c8daf74),
	.w2(32'hbc8f8fc3),
	.w3(32'h38b1f2df),
	.w4(32'h3b33d262),
	.w5(32'h3b667e1a),
	.w6(32'h3ca8d9bb),
	.w7(32'hbcc582c8),
	.w8(32'h3cdc25fd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfb3e32),
	.w1(32'h3c05cf9f),
	.w2(32'h3cd09479),
	.w3(32'h3b34c4f7),
	.w4(32'h3c61016d),
	.w5(32'h3bbfaaf0),
	.w6(32'h3ae404a7),
	.w7(32'h3d2086be),
	.w8(32'hbc2a1f6d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19c268),
	.w1(32'h3c59049b),
	.w2(32'hbc2730ba),
	.w3(32'hbc22a822),
	.w4(32'h3bcfcda0),
	.w5(32'h3c380603),
	.w6(32'hbbe3334a),
	.w7(32'h381c9843),
	.w8(32'h3c2a9537),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b5340),
	.w1(32'hbbf09530),
	.w2(32'hbc3386c5),
	.w3(32'h3bb81763),
	.w4(32'hbce9fe6f),
	.w5(32'h3c279640),
	.w6(32'h3b778189),
	.w7(32'hbc15da63),
	.w8(32'h3d399ba6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd67d62),
	.w1(32'hbc79bb5e),
	.w2(32'hbc941f00),
	.w3(32'hbb8b88ac),
	.w4(32'hbc6f3fba),
	.w5(32'h3bcfcf00),
	.w6(32'hbcb3cc48),
	.w7(32'hbcb8ad3f),
	.w8(32'h3c17c1a0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca2d60),
	.w1(32'hba2bbb8b),
	.w2(32'h3c9654b0),
	.w3(32'h3bdb3051),
	.w4(32'h3b0fa38d),
	.w5(32'h3ca69265),
	.w6(32'h3c923f0a),
	.w7(32'h3ce3ea15),
	.w8(32'hbb80435e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccfb33b),
	.w1(32'h3b082a62),
	.w2(32'hbc87d160),
	.w3(32'hbc934488),
	.w4(32'hba26c2da),
	.w5(32'hbbf00d65),
	.w6(32'hbc172f45),
	.w7(32'hbca9094a),
	.w8(32'h37de667c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbcf28),
	.w1(32'hbac93248),
	.w2(32'h3c685ec6),
	.w3(32'hba6846fc),
	.w4(32'h3b9774fa),
	.w5(32'hbc3d5fb6),
	.w6(32'h3af98d43),
	.w7(32'h3bad75c0),
	.w8(32'h3a83506b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63a056),
	.w1(32'h3c25fb51),
	.w2(32'h3b7ab76d),
	.w3(32'hbb908689),
	.w4(32'h3a670499),
	.w5(32'h3ae4c5c4),
	.w6(32'h3bd1e56e),
	.w7(32'hbba1a683),
	.w8(32'hbb91e9ac),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68a626),
	.w1(32'h3b41a340),
	.w2(32'h3bd4f43c),
	.w3(32'hbb4cd179),
	.w4(32'hbba8d8b8),
	.w5(32'hbad0096a),
	.w6(32'h3ae8ac3b),
	.w7(32'hbb40a322),
	.w8(32'hbc294801),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd0269),
	.w1(32'hbb1ba5a2),
	.w2(32'hbb26ab9e),
	.w3(32'hbba4834d),
	.w4(32'hbb73ed7e),
	.w5(32'h3ae3d85c),
	.w6(32'hbc23f0da),
	.w7(32'hbb81cae9),
	.w8(32'hbb9377e4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d638f),
	.w1(32'h3bc0335e),
	.w2(32'hbc00f643),
	.w3(32'h3a8dcc3e),
	.w4(32'hba93a52d),
	.w5(32'h3b938bd7),
	.w6(32'h3a927a8c),
	.w7(32'h3bbcd301),
	.w8(32'h3bdbc378),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0e76b),
	.w1(32'h3bd54e34),
	.w2(32'h3ca190a8),
	.w3(32'hbb35a297),
	.w4(32'hbcb87a6e),
	.w5(32'hbc8680ef),
	.w6(32'hbc124aca),
	.w7(32'h3c204660),
	.w8(32'hbc951c0a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3443f4),
	.w1(32'hbc519435),
	.w2(32'hbb627a05),
	.w3(32'hbb5f6a15),
	.w4(32'h3c834eac),
	.w5(32'h3a6abe8e),
	.w6(32'hbb3f32dc),
	.w7(32'hbb299809),
	.w8(32'hbc884876),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0cd13e),
	.w1(32'hbc474792),
	.w2(32'h3d00f0b6),
	.w3(32'hbba67632),
	.w4(32'h3c4ae909),
	.w5(32'hbb166bac),
	.w6(32'hb9cbe3e5),
	.w7(32'h3d1b6fc2),
	.w8(32'hbc15baaa),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd98ace),
	.w1(32'hbc65e4de),
	.w2(32'hbc9c4a0a),
	.w3(32'hbbecd168),
	.w4(32'h3c2b024a),
	.w5(32'h3c7c0d79),
	.w6(32'hbc43b3a6),
	.w7(32'hbb22ad42),
	.w8(32'hba3fd457),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb95743),
	.w1(32'h3cb840de),
	.w2(32'h3c8fda0f),
	.w3(32'h3c3a1a57),
	.w4(32'h3b005bab),
	.w5(32'hbc06d94f),
	.w6(32'h3ba0cd88),
	.w7(32'h3c3f284b),
	.w8(32'hbcebcac6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde72e2),
	.w1(32'hbc0427fe),
	.w2(32'h3c93b4fc),
	.w3(32'h3a074c69),
	.w4(32'hbc8fff90),
	.w5(32'h3c445e80),
	.w6(32'hbcc85b6f),
	.w7(32'hbc1414fa),
	.w8(32'h3ba0dda8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce04f09),
	.w1(32'hbbb6309b),
	.w2(32'hbca56b4d),
	.w3(32'h3bd64761),
	.w4(32'hbc5a8c47),
	.w5(32'h3d095543),
	.w6(32'h3ca1e301),
	.w7(32'hbca38d9c),
	.w8(32'h3d6b986d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca263a),
	.w1(32'hbb0c62b1),
	.w2(32'hbc9b424b),
	.w3(32'hbb847779),
	.w4(32'h3a71a456),
	.w5(32'hbbd2b650),
	.w6(32'h3c64091d),
	.w7(32'hbc3394c0),
	.w8(32'h3bf8520d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb663cfe),
	.w1(32'h3a29d912),
	.w2(32'h3b8e7fa4),
	.w3(32'hbb21cd3f),
	.w4(32'hb9ca531d),
	.w5(32'hbb65cee4),
	.w6(32'hba57fd69),
	.w7(32'h3c05737c),
	.w8(32'h3b3c9799),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfadc32),
	.w1(32'h3c162e18),
	.w2(32'h3c17a3d3),
	.w3(32'h3bc0785d),
	.w4(32'hbc3df029),
	.w5(32'h3c28b5a8),
	.w6(32'h3c1801dd),
	.w7(32'hbb63f21e),
	.w8(32'h3bbcd0cc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03a4ed),
	.w1(32'h39b4027c),
	.w2(32'h3c136dcc),
	.w3(32'h3938798b),
	.w4(32'hbbf0d761),
	.w5(32'hbc0c7ad6),
	.w6(32'hbc3ea515),
	.w7(32'h3c3aac88),
	.w8(32'hbca6cf80),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8553e1),
	.w1(32'hbcf1732e),
	.w2(32'hbbe1149a),
	.w3(32'h3bf45275),
	.w4(32'hbd34d1af),
	.w5(32'hbc729b1b),
	.w6(32'hbcc308ae),
	.w7(32'hbd02c524),
	.w8(32'hbca6d25c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fac55),
	.w1(32'hb9232da5),
	.w2(32'hbbe68fd8),
	.w3(32'h3be27a2d),
	.w4(32'hbc44aa5f),
	.w5(32'h3c6e3571),
	.w6(32'h3c1f7319),
	.w7(32'h3cd841f3),
	.w8(32'hbcb52176),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03e23c),
	.w1(32'hbc393fb8),
	.w2(32'h3bcca965),
	.w3(32'h3bc0a33a),
	.w4(32'h3bc71fe5),
	.w5(32'hbcea1b2d),
	.w6(32'h3ce22b16),
	.w7(32'h3c48d49a),
	.w8(32'hbc38631a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc0af9),
	.w1(32'hbc139990),
	.w2(32'hb92ba798),
	.w3(32'hbb31f41a),
	.w4(32'hba5e3503),
	.w5(32'h3aade3f3),
	.w6(32'hbc10eefb),
	.w7(32'hbb454d62),
	.w8(32'hbacf1e57),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d39b4),
	.w1(32'hba7f0ccc),
	.w2(32'h3c3b81aa),
	.w3(32'hba594bb5),
	.w4(32'hbc6b75b7),
	.w5(32'hbb942f40),
	.w6(32'hbac4f2af),
	.w7(32'h3c2e0a55),
	.w8(32'hbce178b9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87d445),
	.w1(32'hbc572244),
	.w2(32'hbbe7ca27),
	.w3(32'h3b80bf63),
	.w4(32'h3c9e210a),
	.w5(32'hbc75fa69),
	.w6(32'hbb747c4b),
	.w7(32'hbb8b2bfe),
	.w8(32'hbb443401),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce21871),
	.w1(32'hbbbe31fb),
	.w2(32'h3c9efcf2),
	.w3(32'hbc00c56d),
	.w4(32'hbc08d2be),
	.w5(32'hbc7c5d5e),
	.w6(32'hbbba9fa0),
	.w7(32'h3ca51277),
	.w8(32'hbcbbd3c9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb377aa1),
	.w1(32'h3b7a0ea1),
	.w2(32'h3ad9b256),
	.w3(32'h3ba191d5),
	.w4(32'h3c67daec),
	.w5(32'h3bf221e2),
	.w6(32'hbc59cce9),
	.w7(32'hba28936b),
	.w8(32'hbb8d6b02),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b8e48),
	.w1(32'h3bed64bc),
	.w2(32'hbd094475),
	.w3(32'h3b905945),
	.w4(32'h3b579ec6),
	.w5(32'h3c9bd4a2),
	.w6(32'h3b71e579),
	.w7(32'hbbe34e30),
	.w8(32'h3d7c0895),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa27757),
	.w1(32'hbb4e269b),
	.w2(32'h391331e8),
	.w3(32'hbc83b253),
	.w4(32'h3ae3f67e),
	.w5(32'h3990e93e),
	.w6(32'h3c9980c5),
	.w7(32'h3a8fbd1b),
	.w8(32'hbc576055),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ccc70),
	.w1(32'h3bb6427d),
	.w2(32'h3b336a1d),
	.w3(32'h3b13294d),
	.w4(32'h3a235b2d),
	.w5(32'hbc64954c),
	.w6(32'h3a9cf688),
	.w7(32'h3bd50c06),
	.w8(32'hba8eb3f6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbbe39),
	.w1(32'hbc955c44),
	.w2(32'h3c9b69e6),
	.w3(32'h3b9cb328),
	.w4(32'h3c10d5f5),
	.w5(32'hbc6592c2),
	.w6(32'hbb3caa66),
	.w7(32'h3d555aa3),
	.w8(32'hbd2bc25b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ef1df),
	.w1(32'hbc7bc30b),
	.w2(32'hbc05fcfa),
	.w3(32'h3b39ae45),
	.w4(32'hba8c4ba0),
	.w5(32'h3bc58ec2),
	.w6(32'h3c3cbc72),
	.w7(32'hbb41d2b4),
	.w8(32'h3bc97ae1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3ff4),
	.w1(32'h3a706961),
	.w2(32'h3b86f2b8),
	.w3(32'hbb6c33c8),
	.w4(32'hbc2c89f2),
	.w5(32'hbb4ffc3a),
	.w6(32'hbb3de363),
	.w7(32'h3ad9762f),
	.w8(32'hbc8594f0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5fe9b),
	.w1(32'h3bfbadb9),
	.w2(32'hbceba86b),
	.w3(32'hbc044b9d),
	.w4(32'hbb2958a6),
	.w5(32'h3c12f1f7),
	.w6(32'hbc562093),
	.w7(32'hbc3cce7b),
	.w8(32'h3d132a0e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9c1d2),
	.w1(32'h3bc7746a),
	.w2(32'hbc1c1325),
	.w3(32'hba229c47),
	.w4(32'hbbfa9097),
	.w5(32'hbc4be662),
	.w6(32'hbc2e149a),
	.w7(32'hbc283e6d),
	.w8(32'h3a210d45),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceed50c),
	.w1(32'hbba9faeb),
	.w2(32'h3a9e39ec),
	.w3(32'hbaa71054),
	.w4(32'hbb6290f9),
	.w5(32'h3b0f53c3),
	.w6(32'h3bbf9975),
	.w7(32'hbc12217f),
	.w8(32'h3b913963),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8fa2c),
	.w1(32'hbb2a6134),
	.w2(32'hbca367d0),
	.w3(32'hbbb29d29),
	.w4(32'hbc114b97),
	.w5(32'h3bf20b4f),
	.w6(32'h3b6faf87),
	.w7(32'h3c5efcb6),
	.w8(32'h3be19b95),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b6113),
	.w1(32'h3bd5453e),
	.w2(32'hbca73fc7),
	.w3(32'hbc1b512a),
	.w4(32'hbb1859d7),
	.w5(32'h3c4b367b),
	.w6(32'h3c517ab4),
	.w7(32'hbd084aac),
	.w8(32'h3d8d7aeb),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c445efd),
	.w1(32'h3c8efba6),
	.w2(32'hbbb9bca3),
	.w3(32'hbb037f38),
	.w4(32'hbc5ef861),
	.w5(32'hbc100b86),
	.w6(32'h3c814e7a),
	.w7(32'hbbbcff8f),
	.w8(32'hbc9c1728),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b613bae),
	.w1(32'hbc2cd49f),
	.w2(32'hbc2a619d),
	.w3(32'h3c6b9b9b),
	.w4(32'hbc6b588e),
	.w5(32'hbbba6a1b),
	.w6(32'hbbe74dd8),
	.w7(32'h3c8f03ae),
	.w8(32'h3ccdc29d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc410c1d),
	.w1(32'hba25be6b),
	.w2(32'h3c91a888),
	.w3(32'hbc50f705),
	.w4(32'h3b8ab968),
	.w5(32'hbc8376b3),
	.w6(32'h3cd5f8d2),
	.w7(32'h3c17360b),
	.w8(32'hbc762cfa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6f47f),
	.w1(32'h3aa630f2),
	.w2(32'h3bfa527b),
	.w3(32'hbc191ee5),
	.w4(32'hbcd6c3d4),
	.w5(32'hbcc0c18d),
	.w6(32'hba766c4f),
	.w7(32'h3c4c50ce),
	.w8(32'hbca27930),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066768),
	.w1(32'hbc231180),
	.w2(32'hbcf4d423),
	.w3(32'hbae8dae7),
	.w4(32'h3caf6437),
	.w5(32'h3cab4eea),
	.w6(32'h3be364fa),
	.w7(32'h3c14614e),
	.w8(32'h3d850d4d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2782d9),
	.w1(32'hbba4fa30),
	.w2(32'h3d2ec340),
	.w3(32'hbc997457),
	.w4(32'hbc5a96b6),
	.w5(32'hbca2818b),
	.w6(32'h3c24f508),
	.w7(32'h3c8e09d1),
	.w8(32'hbb0f053c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55e29d),
	.w1(32'hbc4323d0),
	.w2(32'hba967ecb),
	.w3(32'h3c29b403),
	.w4(32'hb9edb034),
	.w5(32'h3adecfed),
	.w6(32'hbc481248),
	.w7(32'hbba72204),
	.w8(32'hbc913c91),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc087413),
	.w1(32'hbc7e2bfb),
	.w2(32'h3ba37dcd),
	.w3(32'hbc0555ff),
	.w4(32'hbbc37fac),
	.w5(32'h3b85aa8e),
	.w6(32'hbc6829a5),
	.w7(32'hbba8e8ca),
	.w8(32'h3b5ea989),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9f7d6),
	.w1(32'hb8575587),
	.w2(32'h3b9316dc),
	.w3(32'hbba73e2e),
	.w4(32'hbbc29329),
	.w5(32'hbc0b23dd),
	.w6(32'hbb10e6ff),
	.w7(32'hbc0ef23f),
	.w8(32'h3c0feb0f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7bcc4),
	.w1(32'hbc7001bf),
	.w2(32'h3a699754),
	.w3(32'h3c27f267),
	.w4(32'hbc4099a0),
	.w5(32'h3c94791b),
	.w6(32'hbc93d7cb),
	.w7(32'hbc9c215e),
	.w8(32'h3d01fe3a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46d431),
	.w1(32'hbbace43d),
	.w2(32'h3b6855e3),
	.w3(32'hbc8adbda),
	.w4(32'h3c67a131),
	.w5(32'h3c759be0),
	.w6(32'h3b7830e5),
	.w7(32'h3bf9eff6),
	.w8(32'h3b75c748),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60e330),
	.w1(32'h3bc70599),
	.w2(32'hbb259a5f),
	.w3(32'h3b6e5c4f),
	.w4(32'hbc6ca954),
	.w5(32'h3cef5522),
	.w6(32'h3b5a19b2),
	.w7(32'hbcd785b6),
	.w8(32'h3d37a79c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c881eb2),
	.w1(32'hbca9e33e),
	.w2(32'h3966a8ca),
	.w3(32'h3bcfd595),
	.w4(32'hbbbd2c63),
	.w5(32'h3b075042),
	.w6(32'h3c6f677d),
	.w7(32'hbc160bdf),
	.w8(32'h3bd7384f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381fdeeb),
	.w1(32'h3b0fcaf5),
	.w2(32'h3b7d7338),
	.w3(32'hbbd93795),
	.w4(32'hbc277af4),
	.w5(32'h3b1b8ea9),
	.w6(32'h38adc2e4),
	.w7(32'hbc3726dd),
	.w8(32'h3c5f72e8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91b471),
	.w1(32'h3bd217da),
	.w2(32'hbb6752df),
	.w3(32'h3b9b5521),
	.w4(32'h3baa194f),
	.w5(32'h3b8fc2ff),
	.w6(32'hbb2633cb),
	.w7(32'h3c8525a5),
	.w8(32'h3d68f269),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf79684),
	.w1(32'h3b773f4e),
	.w2(32'hbc822b71),
	.w3(32'hbcfb3434),
	.w4(32'hbc610bf0),
	.w5(32'hbb05df2c),
	.w6(32'hbbe8f1ea),
	.w7(32'hbc214762),
	.w8(32'h3a53ccb4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bfaff),
	.w1(32'h3b286af7),
	.w2(32'h3b334d67),
	.w3(32'h3b29d7bc),
	.w4(32'hbbac38f9),
	.w5(32'hbc54e149),
	.w6(32'h3bbf8bc9),
	.w7(32'h3b7f923c),
	.w8(32'hbd2be0dc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce83d26),
	.w1(32'hba3c95ea),
	.w2(32'h3c5acee3),
	.w3(32'h3c08348b),
	.w4(32'hbb065855),
	.w5(32'hbaa06d11),
	.w6(32'h3ae4b4f5),
	.w7(32'h3a76b5b3),
	.w8(32'hbca44432),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f2496),
	.w1(32'h3abf4a39),
	.w2(32'hbb002bc2),
	.w3(32'hba97a9a3),
	.w4(32'hbc30c53c),
	.w5(32'h3af953a2),
	.w6(32'hbad35b80),
	.w7(32'hbc64cc81),
	.w8(32'hbc05de7f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8851ed),
	.w1(32'hbc6e556b),
	.w2(32'h3adb6607),
	.w3(32'h3b3edb3f),
	.w4(32'hbca1b110),
	.w5(32'hbcca709d),
	.w6(32'hbc041801),
	.w7(32'hbbb7512d),
	.w8(32'hbc5120cb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86aba3),
	.w1(32'hbbc755ae),
	.w2(32'hbd1275f0),
	.w3(32'hb903f3c2),
	.w4(32'h3ce81c95),
	.w5(32'hbc91adcd),
	.w6(32'h3b356513),
	.w7(32'h3c0c137e),
	.w8(32'h3cf6ccf3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d62edc5),
	.w1(32'hbb8f514c),
	.w2(32'h3c80d18b),
	.w3(32'h3ba75873),
	.w4(32'h3b69a822),
	.w5(32'hbc60d0a5),
	.w6(32'hbb6bff04),
	.w7(32'h3b840c9d),
	.w8(32'hbaa81de2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd72848),
	.w1(32'h3b0b6611),
	.w2(32'h3c4dc27a),
	.w3(32'hbbca6707),
	.w4(32'hbb2dc6c3),
	.w5(32'h3b6c7ead),
	.w6(32'hbcc5ef69),
	.w7(32'hba85bd88),
	.w8(32'hbc7f2682),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc401ccf),
	.w1(32'hbc173751),
	.w2(32'h3c77df85),
	.w3(32'h3b693c21),
	.w4(32'h3b52d279),
	.w5(32'hbc4ca990),
	.w6(32'h3b1f8e2b),
	.w7(32'h3c15834a),
	.w8(32'hbc151a71),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb08715),
	.w1(32'h3ba2b1af),
	.w2(32'hbc25d4aa),
	.w3(32'h3bd7c876),
	.w4(32'h3b3e9d4e),
	.w5(32'h3b93e883),
	.w6(32'h3b09825b),
	.w7(32'h3b7112ce),
	.w8(32'h3cb3010f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b312351),
	.w1(32'h3ba67987),
	.w2(32'h3b76db12),
	.w3(32'hbb64e0d0),
	.w4(32'hbc5a9511),
	.w5(32'hbbb6f110),
	.w6(32'h3abbcb74),
	.w7(32'h3c166998),
	.w8(32'hbce24529),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbddd6b),
	.w1(32'h3ca30d97),
	.w2(32'h3b2d7080),
	.w3(32'h3c3a9a01),
	.w4(32'hbc28ef2f),
	.w5(32'h3c39d868),
	.w6(32'h3c8da50a),
	.w7(32'hbc329c40),
	.w8(32'h3bfbe4fa),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88d400),
	.w1(32'h3a50abd2),
	.w2(32'hbce1295b),
	.w3(32'h3c4702c0),
	.w4(32'hbc699829),
	.w5(32'h3c479511),
	.w6(32'h3b555d42),
	.w7(32'hbd3216a9),
	.w8(32'h3bf522dd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd10f26d),
	.w1(32'h3c5046ff),
	.w2(32'hbbdb9004),
	.w3(32'h3cac4509),
	.w4(32'hbb257f3c),
	.w5(32'hbc9df491),
	.w6(32'h3c8a700c),
	.w7(32'h3bccc97d),
	.w8(32'h3bc36bf5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb233d3),
	.w1(32'hbcae48ce),
	.w2(32'h3cf01cc8),
	.w3(32'hbc2a1451),
	.w4(32'h3be7b617),
	.w5(32'h3c9d13ce),
	.w6(32'hbca11c40),
	.w7(32'h3c957a38),
	.w8(32'h3c131420),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09a5b9),
	.w1(32'h3c8a5525),
	.w2(32'hba9c2752),
	.w3(32'h3b845e19),
	.w4(32'h3b004562),
	.w5(32'h3b09faa1),
	.w6(32'h3c940713),
	.w7(32'h3b09ae63),
	.w8(32'h3bccb37e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a4fa1),
	.w1(32'hbb99abea),
	.w2(32'hb9877920),
	.w3(32'h3b18556f),
	.w4(32'h3be86340),
	.w5(32'h3c023c66),
	.w6(32'hba8cb749),
	.w7(32'h3b696b60),
	.w8(32'h3bf19f88),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee441b),
	.w1(32'hb8207c60),
	.w2(32'h3bb736fa),
	.w3(32'h3b391290),
	.w4(32'h3b95d6d4),
	.w5(32'h3c301c7e),
	.w6(32'hbb413968),
	.w7(32'h3a76771d),
	.w8(32'h3c0de067),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb7161),
	.w1(32'h3a333e2a),
	.w2(32'h3b53cbc6),
	.w3(32'h3b6676f9),
	.w4(32'h3ac865c1),
	.w5(32'hbb01cecf),
	.w6(32'hb9d4b314),
	.w7(32'h3bdc0016),
	.w8(32'hbbf83d7d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c60bc),
	.w1(32'h3b579089),
	.w2(32'hbbf9a746),
	.w3(32'h3b202d00),
	.w4(32'hbb10a19b),
	.w5(32'hbb868479),
	.w6(32'h3b01868d),
	.w7(32'hbc7b0caa),
	.w8(32'h3d371c52),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9040a3),
	.w1(32'hbb8cae3f),
	.w2(32'hba4c68d7),
	.w3(32'hbc93e3bc),
	.w4(32'hbc09941b),
	.w5(32'hbbc423db),
	.w6(32'h3aa2b893),
	.w7(32'h3b747729),
	.w8(32'h3aab7db0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fe28a),
	.w1(32'hbc8764ec),
	.w2(32'h3cbc06e3),
	.w3(32'h3a89b862),
	.w4(32'hbc106b3b),
	.w5(32'h3b78dd3e),
	.w6(32'hbc0e1668),
	.w7(32'h3b907862),
	.w8(32'h3c898de6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc074df6),
	.w1(32'h3b844a77),
	.w2(32'hbb62ad54),
	.w3(32'hbbc32919),
	.w4(32'h3c2ac67e),
	.w5(32'hbc611404),
	.w6(32'h3c9e2670),
	.w7(32'h3c27105e),
	.w8(32'hbb3d615a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98c405),
	.w1(32'hbacd911a),
	.w2(32'h3c4af864),
	.w3(32'hbc0e4bbe),
	.w4(32'hbcaee217),
	.w5(32'h3ced0838),
	.w6(32'hbab88bbd),
	.w7(32'h3bfb65bf),
	.w8(32'h3cdc3926),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1c873f),
	.w1(32'h3c5cbd6d),
	.w2(32'hbc7067b2),
	.w3(32'hbc35d271),
	.w4(32'h39d35489),
	.w5(32'hbc4b4b55),
	.w6(32'hbc6248ce),
	.w7(32'h3baf5e4d),
	.w8(32'hbbc22d62),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc560260),
	.w1(32'hbbead608),
	.w2(32'h3c071411),
	.w3(32'h3b6d1245),
	.w4(32'hbb01fef0),
	.w5(32'hbb55e67e),
	.w6(32'hbbcb3efb),
	.w7(32'h3acd660c),
	.w8(32'hbb1d02d8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc146793),
	.w1(32'hbbae0154),
	.w2(32'h3b74515b),
	.w3(32'h3be0cbb8),
	.w4(32'h3b66fa91),
	.w5(32'h3a69b512),
	.w6(32'hbb846cd3),
	.w7(32'h3c1a47d2),
	.w8(32'hbbd70576),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af257cc),
	.w1(32'h38fe8b9a),
	.w2(32'h3b211fbb),
	.w3(32'hbb234723),
	.w4(32'hbb216926),
	.w5(32'hbaf6ff7d),
	.w6(32'h3b7fb787),
	.w7(32'hbb8b7f7b),
	.w8(32'hbbc85b5d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f07c8),
	.w1(32'hbb4a9323),
	.w2(32'h3c33907c),
	.w3(32'hbbd726f6),
	.w4(32'hbc1b6f6a),
	.w5(32'hbb262b37),
	.w6(32'hbc147b8c),
	.w7(32'h3a14add8),
	.w8(32'h3cf882f8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd43002),
	.w1(32'hba4f9f5e),
	.w2(32'hbbf1e538),
	.w3(32'h3bbb6b1a),
	.w4(32'h3b9a7788),
	.w5(32'hbaae366d),
	.w6(32'h3b4715c4),
	.w7(32'hb96b3d81),
	.w8(32'hbc1b9eaa),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10d487),
	.w1(32'hbb94f532),
	.w2(32'h3c28c073),
	.w3(32'hbbaad3b7),
	.w4(32'h3c755f05),
	.w5(32'hbc5a605c),
	.w6(32'hbbf5def1),
	.w7(32'h3ae4e7bb),
	.w8(32'h3ba86333),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd22ea),
	.w1(32'hbbcc74bf),
	.w2(32'h3bd92204),
	.w3(32'hbbb1fbe6),
	.w4(32'hb99b8640),
	.w5(32'hbd0ac860),
	.w6(32'h3bc5ee55),
	.w7(32'hbc1a0023),
	.w8(32'h3c4dba07),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7baea),
	.w1(32'hbba58024),
	.w2(32'h3bcc5d25),
	.w3(32'h3c600b8b),
	.w4(32'h39d5dac1),
	.w5(32'h3cbdc6e0),
	.w6(32'hbc4a6d32),
	.w7(32'h3d278eab),
	.w8(32'hbc7ee285),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0798c5),
	.w1(32'h3c20a6ec),
	.w2(32'h3bcc4fad),
	.w3(32'hbc186cb6),
	.w4(32'h3c4fc1aa),
	.w5(32'h3bd6ef11),
	.w6(32'hbc310adf),
	.w7(32'h3b94ccf1),
	.w8(32'h3b67f7d9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbba55),
	.w1(32'h3b37ff69),
	.w2(32'hbb7bca3c),
	.w3(32'h3bed7bb3),
	.w4(32'h39e39363),
	.w5(32'hbc8a69c7),
	.w6(32'h3b8ff35e),
	.w7(32'hbb5b67ec),
	.w8(32'hbaede8f1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb129a9),
	.w1(32'hbbce53e4),
	.w2(32'hbbce1ee6),
	.w3(32'hbbda1938),
	.w4(32'hbc480e3c),
	.w5(32'h3c7a0c2a),
	.w6(32'hbb32e03b),
	.w7(32'hba8b9ad4),
	.w8(32'h3c8be002),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbcb57f),
	.w1(32'hbbbaecfe),
	.w2(32'h3ab16f20),
	.w3(32'h3ad26aba),
	.w4(32'hbc1e5a8c),
	.w5(32'h3d1ed32a),
	.w6(32'h3c2f3774),
	.w7(32'h3c206e51),
	.w8(32'h3cb926bc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd006f06),
	.w1(32'h3c0eda30),
	.w2(32'hbb4eb966),
	.w3(32'hbc18a984),
	.w4(32'hbb05ebc9),
	.w5(32'hbb1192d1),
	.w6(32'hbc99f5fa),
	.w7(32'hbb697308),
	.w8(32'hbbdb56d6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4a610),
	.w1(32'h3b6f9972),
	.w2(32'h3b9d79ab),
	.w3(32'hbb87e3fb),
	.w4(32'hbacecc76),
	.w5(32'hbc1e6f13),
	.w6(32'hbb75bf18),
	.w7(32'h3cf83936),
	.w8(32'hbcbc61c7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38baf6),
	.w1(32'h3c04632a),
	.w2(32'h3ba666a6),
	.w3(32'h3c9bebd1),
	.w4(32'h3c0f7d14),
	.w5(32'h39825781),
	.w6(32'h3c671eb9),
	.w7(32'h3bcde7ef),
	.w8(32'hbb1a0d26),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b368ca1),
	.w1(32'hbc315e28),
	.w2(32'h3bcdc356),
	.w3(32'h3bed7636),
	.w4(32'h3b58660d),
	.w5(32'hbc7f5933),
	.w6(32'hbc8f9dca),
	.w7(32'hbb95ad0e),
	.w8(32'hbc197d1f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc703a7),
	.w1(32'h3b20262a),
	.w2(32'hba1515ae),
	.w3(32'hbbebcb7f),
	.w4(32'hbc42ea3d),
	.w5(32'hbb3c30b4),
	.w6(32'hbc39d27a),
	.w7(32'h3c0b013f),
	.w8(32'h3d43fe1e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e89c5),
	.w1(32'hbc692b1a),
	.w2(32'hbbc1568d),
	.w3(32'h3b65641f),
	.w4(32'hbbb3982e),
	.w5(32'hbb1cbbeb),
	.w6(32'hbce1bdb1),
	.w7(32'hbb2d6f15),
	.w8(32'hba815501),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4d492),
	.w1(32'hb8e48214),
	.w2(32'h3ba1e46d),
	.w3(32'hbaff0d47),
	.w4(32'hbb1b14a5),
	.w5(32'hbc1d85d7),
	.w6(32'h3b961993),
	.w7(32'h3c11fa6e),
	.w8(32'hbc7348c2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e9845),
	.w1(32'hbb9ffde0),
	.w2(32'hbba26632),
	.w3(32'h3b9f5d49),
	.w4(32'h3b56fd9c),
	.w5(32'h3be49958),
	.w6(32'h3b9061b7),
	.w7(32'h3cd94211),
	.w8(32'hbcf1f05e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e554),
	.w1(32'h3c725bcb),
	.w2(32'h3c23a190),
	.w3(32'h3c38943d),
	.w4(32'hbc911588),
	.w5(32'h3c46cb63),
	.w6(32'h3ce3f343),
	.w7(32'hbc401099),
	.w8(32'h3ca6515a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75675d),
	.w1(32'hbbfaf5cc),
	.w2(32'hbb37818b),
	.w3(32'h3bfcbcbf),
	.w4(32'h3ae2ad46),
	.w5(32'hb9a1906e),
	.w6(32'h3c0490f1),
	.w7(32'h3adadfca),
	.w8(32'h3b33c8a6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bafe8),
	.w1(32'h3a9e4732),
	.w2(32'h3b9ef109),
	.w3(32'h3b646660),
	.w4(32'h3b524528),
	.w5(32'hbc2d4423),
	.w6(32'h3a37e626),
	.w7(32'hbbaecc8a),
	.w8(32'h3cf6025d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b883792),
	.w1(32'hbb8c01aa),
	.w2(32'hbc80e33c),
	.w3(32'h3b9c31d2),
	.w4(32'h3c58778f),
	.w5(32'hbcdbe0e0),
	.w6(32'h3baf0523),
	.w7(32'h3c793d91),
	.w8(32'hbd6c5fc0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd2047),
	.w1(32'hba4634fb),
	.w2(32'h3a2420eb),
	.w3(32'h3bb87d56),
	.w4(32'hbb5bf3e2),
	.w5(32'h3c1ee080),
	.w6(32'h3d0144dc),
	.w7(32'h3b055243),
	.w8(32'hbca15e95),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb672722),
	.w1(32'hbba09790),
	.w2(32'h3c3143d0),
	.w3(32'hbb8cf50a),
	.w4(32'hbc38f21f),
	.w5(32'hbc1a5e6c),
	.w6(32'h3b5a4504),
	.w7(32'hbd1a3ce1),
	.w8(32'h3cbbf5b9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41f511),
	.w1(32'hbbd5edec),
	.w2(32'hbb96b0ff),
	.w3(32'hbc2e9368),
	.w4(32'h3aaff6cb),
	.w5(32'hbc57b4da),
	.w6(32'h3c3bcd36),
	.w7(32'h3c0c66c9),
	.w8(32'hbc86a43f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb203e21),
	.w1(32'hbca8746f),
	.w2(32'hbca4ff2c),
	.w3(32'hbc13f891),
	.w4(32'hbc2cb9b7),
	.w5(32'hbc8af468),
	.w6(32'hbc4b0c44),
	.w7(32'hbbe81061),
	.w8(32'hbc6717a4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78a334),
	.w1(32'hbccbb513),
	.w2(32'h3bae38ce),
	.w3(32'hbcb1dd88),
	.w4(32'h3c92201d),
	.w5(32'hbd152bcd),
	.w6(32'hbcb4d6a8),
	.w7(32'h3a0c2c2a),
	.w8(32'hbd146cfe),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c72b2),
	.w1(32'h3ae4e6d2),
	.w2(32'hbcafaae4),
	.w3(32'hbb118c5f),
	.w4(32'hbc2cfa40),
	.w5(32'h3c59fc2f),
	.w6(32'h3c8779ac),
	.w7(32'hbc3b0370),
	.w8(32'h3b8110b2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba06d66),
	.w1(32'h3c60bc12),
	.w2(32'hbc12bd55),
	.w3(32'hbc4a748f),
	.w4(32'hbbdcb3f2),
	.w5(32'hbbe1e5b6),
	.w6(32'h3c7a8c9c),
	.w7(32'hbc9cf32b),
	.w8(32'hbc6aad77),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf13eb1),
	.w1(32'h3a72ee88),
	.w2(32'hbb9110a2),
	.w3(32'hbbc3a6f5),
	.w4(32'h3af26f09),
	.w5(32'hba29c355),
	.w6(32'h393a9722),
	.w7(32'h3a8589c5),
	.w8(32'h3b505e2c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba91601),
	.w1(32'h39db9bf6),
	.w2(32'h3bfc1764),
	.w3(32'h39d00b91),
	.w4(32'hbc0576b0),
	.w5(32'h3b939dc5),
	.w6(32'hbad6be1c),
	.w7(32'hbcdc01a3),
	.w8(32'hbaf79300),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44de6f),
	.w1(32'h3b16d158),
	.w2(32'h3b72254d),
	.w3(32'hbc063ac9),
	.w4(32'hbbe92dcf),
	.w5(32'hbcad8bbe),
	.w6(32'hbc0e99e5),
	.w7(32'hbca00f23),
	.w8(32'hbb71ecc1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d007f),
	.w1(32'h3b93b1d7),
	.w2(32'h3b8aef3c),
	.w3(32'hbbe8e5a9),
	.w4(32'h3b31403a),
	.w5(32'hbab42325),
	.w6(32'h3c9a4179),
	.w7(32'h3bd4d8a2),
	.w8(32'h3c18cf41),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8277b1),
	.w1(32'hbb8e27a7),
	.w2(32'h3c8c1935),
	.w3(32'h3a6aecdf),
	.w4(32'h3b4f2ff0),
	.w5(32'hbc8c5dc1),
	.w6(32'h3abe3fc4),
	.w7(32'h3ca862a2),
	.w8(32'hbb3b89ae),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc1271),
	.w1(32'hbc50d434),
	.w2(32'hbaeed81b),
	.w3(32'h3b84858c),
	.w4(32'h3b78be40),
	.w5(32'h3a87cbea),
	.w6(32'hbb8ee0bf),
	.w7(32'h3a82bd0d),
	.w8(32'h3b37b0db),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc787c),
	.w1(32'h3a2d5c7e),
	.w2(32'hbb774c31),
	.w3(32'h3ad667d3),
	.w4(32'hbbd4ac85),
	.w5(32'hbce30a28),
	.w6(32'hb99623e3),
	.w7(32'hbc246c06),
	.w8(32'h3c914541),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e6fef),
	.w1(32'hbcd2fa06),
	.w2(32'hbbd0f90a),
	.w3(32'h3c2b3d51),
	.w4(32'h3c37be85),
	.w5(32'hbac69b56),
	.w6(32'h3c8cbaf1),
	.w7(32'h3d18aa09),
	.w8(32'hbda0c8b1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4a211),
	.w1(32'h3c96bc58),
	.w2(32'hbb1ea548),
	.w3(32'h3bb2ab55),
	.w4(32'hbbaa799b),
	.w5(32'h3b9c6147),
	.w6(32'h3cb827d1),
	.w7(32'hbb8feec1),
	.w8(32'h3c31161a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94fda6),
	.w1(32'h3b472c5f),
	.w2(32'hbc63da3a),
	.w3(32'hbab1eb17),
	.w4(32'hba20c4a5),
	.w5(32'hbc156940),
	.w6(32'h3b89edac),
	.w7(32'hbcd0ea36),
	.w8(32'hbc4bf503),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d2610),
	.w1(32'hbc0ac45f),
	.w2(32'hbb87dc43),
	.w3(32'hbc868985),
	.w4(32'hbc02b442),
	.w5(32'h39efcf2c),
	.w6(32'hbc87fc46),
	.w7(32'hbc36312c),
	.w8(32'h3aa94ea3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule