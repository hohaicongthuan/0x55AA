module layer_8_featuremap_6(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce7aad8),
	.w1(32'h3a01e924),
	.w2(32'h3b85b787),
	.w3(32'h3cbf449f),
	.w4(32'hbb9f76c7),
	.w5(32'h3c232fb0),
	.w6(32'hbc21f1d3),
	.w7(32'h3b53954d),
	.w8(32'h3c5876d2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52c42d),
	.w1(32'hbbea729b),
	.w2(32'hbc0b53b5),
	.w3(32'hbb86fb5b),
	.w4(32'hbb27f228),
	.w5(32'hbbe70da7),
	.w6(32'hbaab0300),
	.w7(32'h3b257434),
	.w8(32'h3a752e20),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21fdef),
	.w1(32'h3abf08ee),
	.w2(32'hba86c35c),
	.w3(32'hbb25d9b7),
	.w4(32'h3a69b598),
	.w5(32'hbb32d4fc),
	.w6(32'h3bab3a30),
	.w7(32'h3a324254),
	.w8(32'h38aa8feb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfc505),
	.w1(32'h3c265f32),
	.w2(32'h3c5b213b),
	.w3(32'hbb60357c),
	.w4(32'h3c97d628),
	.w5(32'h3c9ba073),
	.w6(32'h3b8a9cf2),
	.w7(32'h3cac93fc),
	.w8(32'h3c62696e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c9baf),
	.w1(32'hbb4d0277),
	.w2(32'hbb5f84bb),
	.w3(32'h3b4e601b),
	.w4(32'h3ac48176),
	.w5(32'hbaad2b89),
	.w6(32'h3b267009),
	.w7(32'h3b121680),
	.w8(32'hb9597344),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51de3c),
	.w1(32'h3c096f6b),
	.w2(32'h3a1769f2),
	.w3(32'h3aa94fa3),
	.w4(32'h3c4ed82e),
	.w5(32'hbc5144a8),
	.w6(32'h3c2a62d4),
	.w7(32'hbbf30d14),
	.w8(32'hbcbdc991),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ca031),
	.w1(32'hbb9ab661),
	.w2(32'hbb106250),
	.w3(32'h38f1fd50),
	.w4(32'hbb2de80b),
	.w5(32'hb9dce67e),
	.w6(32'hbb1b1cfc),
	.w7(32'hb983097b),
	.w8(32'h3a6fd5e7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16aa72),
	.w1(32'h3af7cbe8),
	.w2(32'h3c8de00c),
	.w3(32'hbae6f947),
	.w4(32'h3bf10ec5),
	.w5(32'h3bf7e81d),
	.w6(32'h3b63939b),
	.w7(32'h39392d0c),
	.w8(32'h3a5884ec),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f6dfc),
	.w1(32'hbccb683a),
	.w2(32'hbcca4f66),
	.w3(32'h3bed8299),
	.w4(32'hbcbc0142),
	.w5(32'hbcb489a6),
	.w6(32'h39f91db6),
	.w7(32'hbcc3d040),
	.w8(32'hbcbe2e76),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4575fd),
	.w1(32'h3a7b53d8),
	.w2(32'h3c1b47a1),
	.w3(32'hbce5a7f8),
	.w4(32'h3b921eb6),
	.w5(32'h3bd05b3b),
	.w6(32'hbcf06d2e),
	.w7(32'h3b319920),
	.w8(32'h3bb7c08f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8b662),
	.w1(32'h3bb513e6),
	.w2(32'h3c48332e),
	.w3(32'hbc04e512),
	.w4(32'hbb769f03),
	.w5(32'h3be6655e),
	.w6(32'hbbd68be8),
	.w7(32'hbc059236),
	.w8(32'h3c108389),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcda7f0),
	.w1(32'h3b9d7682),
	.w2(32'h3ba604f0),
	.w3(32'hbb03ccbb),
	.w4(32'h3be06298),
	.w5(32'h3c546fd6),
	.w6(32'h3b35bd11),
	.w7(32'h3c54eab5),
	.w8(32'h3c042eea),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac0121),
	.w1(32'hbbf46d27),
	.w2(32'hbc664dad),
	.w3(32'h3b07ed06),
	.w4(32'hb9fd34af),
	.w5(32'hbc3a67d3),
	.w6(32'h3b84ba11),
	.w7(32'h3bce6b89),
	.w8(32'hbb198aa6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc035fe5),
	.w1(32'hbc7c06dd),
	.w2(32'hbccb97fe),
	.w3(32'hbb0ec3d3),
	.w4(32'hbcfc337c),
	.w5(32'hbd458fee),
	.w6(32'hb982756e),
	.w7(32'hbcbb25fd),
	.w8(32'hbd17d395),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f975b),
	.w1(32'h3c7e6101),
	.w2(32'h3cdf29f2),
	.w3(32'hbd0cdee4),
	.w4(32'h3cf95ff7),
	.w5(32'h3d3ce436),
	.w6(32'hbcdabafb),
	.w7(32'h3cdcf051),
	.w8(32'h3d211e9d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc40805),
	.w1(32'hb9b28109),
	.w2(32'h3b18d8bd),
	.w3(32'h3d2421f6),
	.w4(32'h3af23535),
	.w5(32'hb916a872),
	.w6(32'h3d0f66aa),
	.w7(32'hbb1492ba),
	.w8(32'hbafa90a4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a861cf7),
	.w1(32'hbbd2da3e),
	.w2(32'h3a8ca7f9),
	.w3(32'hbbaf6bb7),
	.w4(32'hbc4c54c0),
	.w5(32'h3bd974d2),
	.w6(32'hbb98e838),
	.w7(32'hbbf973d2),
	.w8(32'h3c2f6485),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda693e),
	.w1(32'h3becbf06),
	.w2(32'h3c03cd9e),
	.w3(32'h3c38ee7d),
	.w4(32'h3c31ee64),
	.w5(32'h3ad5e126),
	.w6(32'h3bbd0014),
	.w7(32'h3c3eb0b2),
	.w8(32'h3b90495d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cd879),
	.w1(32'h3b84c0b0),
	.w2(32'h3cdea339),
	.w3(32'hbd0ec56b),
	.w4(32'hbcfe1ba5),
	.w5(32'h3cb90966),
	.w6(32'hbbbb6e62),
	.w7(32'h3c335418),
	.w8(32'h3d10e8cb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ca273),
	.w1(32'h3c86d548),
	.w2(32'h3cbe3119),
	.w3(32'h3c8c5d8c),
	.w4(32'h3d2a90b0),
	.w5(32'h3d484549),
	.w6(32'h3b8767e3),
	.w7(32'h3cb862a0),
	.w8(32'h3cf967d8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cff15e5),
	.w1(32'hb9fc2be5),
	.w2(32'hbcde7c34),
	.w3(32'h3d340933),
	.w4(32'hbce1688f),
	.w5(32'hbd593f2b),
	.w6(32'h3cf23139),
	.w7(32'hbceb983a),
	.w8(32'hbd229bb9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33e113),
	.w1(32'h3ae99bf2),
	.w2(32'hbb94986b),
	.w3(32'hbce07cc5),
	.w4(32'hbbb436f1),
	.w5(32'hbc69cc9f),
	.w6(32'hbc94f3f8),
	.w7(32'hbb8c87d9),
	.w8(32'hbc3d94bb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8f484),
	.w1(32'hbc203491),
	.w2(32'h3cc3d6c2),
	.w3(32'hbc20b198),
	.w4(32'hbbd839cb),
	.w5(32'h3c23da74),
	.w6(32'hbc8ee288),
	.w7(32'hbc5aec46),
	.w8(32'h3c5c7aba),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4adc02),
	.w1(32'h3b5eac26),
	.w2(32'h3ad88f27),
	.w3(32'h3ba1eae0),
	.w4(32'hbafbc707),
	.w5(32'hbbb25953),
	.w6(32'h3b23efc9),
	.w7(32'hbbcec982),
	.w8(32'hbc44c04d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd25bac),
	.w1(32'h3b2b1575),
	.w2(32'hba1d958c),
	.w3(32'hba139370),
	.w4(32'h3bc31d06),
	.w5(32'h3ba37b20),
	.w6(32'hbb86575f),
	.w7(32'h3b8fd8ac),
	.w8(32'h3b7c03ff),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb948296),
	.w1(32'h3c0a333b),
	.w2(32'h3c456556),
	.w3(32'h3a90cc6a),
	.w4(32'h3c4f4794),
	.w5(32'h3c6e5a85),
	.w6(32'h3b249c61),
	.w7(32'h3c399581),
	.w8(32'h3c535524),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58958e),
	.w1(32'h3bfe464d),
	.w2(32'h3c8b8028),
	.w3(32'h3c8abe10),
	.w4(32'h3c50bdd7),
	.w5(32'h3c9cd2b5),
	.w6(32'h3c4606cb),
	.w7(32'h3bd0d803),
	.w8(32'h3c653853),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd41265a),
	.w1(32'h3cea4a61),
	.w2(32'hbd0f3175),
	.w3(32'hbc6d0750),
	.w4(32'hbcf05259),
	.w5(32'hbdcb98e8),
	.w6(32'hbd1cd04b),
	.w7(32'hbd0dc4d5),
	.w8(32'hbd682dad),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8169c),
	.w1(32'h3ba1dd5f),
	.w2(32'h3c565f80),
	.w3(32'hbbc6ffb6),
	.w4(32'h3c25973f),
	.w5(32'h3c6575ce),
	.w6(32'h3a0ea91b),
	.w7(32'h3ba65283),
	.w8(32'h3c188f17),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fe311),
	.w1(32'h3b5b071e),
	.w2(32'h3c3a4598),
	.w3(32'h3bef4935),
	.w4(32'h3c0fafd0),
	.w5(32'h3c957760),
	.w6(32'hba9f8000),
	.w7(32'h3c2332ca),
	.w8(32'h3cb0cd2b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c129dea),
	.w1(32'hbbdb62ea),
	.w2(32'hbadbe41f),
	.w3(32'h3c913615),
	.w4(32'hbbf42fe1),
	.w5(32'hbb15dc18),
	.w6(32'h3cc11096),
	.w7(32'hbb97ff89),
	.w8(32'h3ac6580e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886dfe),
	.w1(32'hbcb0c218),
	.w2(32'hbca5b567),
	.w3(32'hbbe1fe9a),
	.w4(32'hbce16139),
	.w5(32'hbcdaeca6),
	.w6(32'hbb1375e6),
	.w7(32'hbcc36bdf),
	.w8(32'hbcb48e6c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62b558),
	.w1(32'hb9576574),
	.w2(32'h395b29b7),
	.w3(32'hbc8d6b28),
	.w4(32'hba7f5770),
	.w5(32'hbacdf8f2),
	.w6(32'hbc6d88dd),
	.w7(32'h3a51c073),
	.w8(32'hba200a31),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68223f),
	.w1(32'hbbcd0d78),
	.w2(32'hbb15c0ec),
	.w3(32'h3b13e702),
	.w4(32'hbb075268),
	.w5(32'h3b3a5f93),
	.w6(32'h3b3e2c94),
	.w7(32'hbbac932d),
	.w8(32'h39998b29),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4da696),
	.w1(32'hbb6dbe57),
	.w2(32'hbbf0248f),
	.w3(32'hbbc9721f),
	.w4(32'h3a21f7eb),
	.w5(32'hbbc962e7),
	.w6(32'hbc592d1a),
	.w7(32'hbb98236b),
	.w8(32'hbc33480a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3874f3),
	.w1(32'hbaabfe8f),
	.w2(32'h3aa9c4e4),
	.w3(32'hbc6de84f),
	.w4(32'hbbda5500),
	.w5(32'hbb547450),
	.w6(32'hbbf43436),
	.w7(32'h3aeee1b6),
	.w8(32'h3accab5e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc7fb9),
	.w1(32'hbb05cdb7),
	.w2(32'hba9d26f6),
	.w3(32'h3b7a880f),
	.w4(32'h3abe0180),
	.w5(32'hbb818bde),
	.w6(32'h3b55d07c),
	.w7(32'hba47baea),
	.w8(32'hbbd7ae6f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16856d),
	.w1(32'h3a5630ee),
	.w2(32'h3a95cfbc),
	.w3(32'hbc49e769),
	.w4(32'h3c0dad10),
	.w5(32'hbb3d7dcb),
	.w6(32'hbc49da68),
	.w7(32'h3be59f7f),
	.w8(32'h3bcf0826),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc087eea),
	.w1(32'h3a8e3a09),
	.w2(32'hbb59e43e),
	.w3(32'hbbddc8df),
	.w4(32'hba9f9c91),
	.w5(32'h3b83bc23),
	.w6(32'hbba07f16),
	.w7(32'hbbff1b1b),
	.w8(32'hbbc0db1b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae81531),
	.w1(32'h3bd19f67),
	.w2(32'h3bc5f97e),
	.w3(32'hba6223fa),
	.w4(32'h3b69d4e1),
	.w5(32'h3c330d60),
	.w6(32'hbbd3e9bc),
	.w7(32'h3ba29eac),
	.w8(32'h3c24f84e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c87f5),
	.w1(32'h3d29cc18),
	.w2(32'h3d2ec601),
	.w3(32'h3ca28454),
	.w4(32'h3d6a11ba),
	.w5(32'h3d2fc230),
	.w6(32'h3cc8b86c),
	.w7(32'h3d3c78e3),
	.w8(32'h3d057b2e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a584b),
	.w1(32'hbca8a39a),
	.w2(32'hbc979f2e),
	.w3(32'h3c7cd950),
	.w4(32'hbcec9f12),
	.w5(32'hbcf06ac5),
	.w6(32'h3c5f718f),
	.w7(32'hbcc891a6),
	.w8(32'hbcb79c62),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2543b6),
	.w1(32'hbb93af07),
	.w2(32'hbb81730a),
	.w3(32'hbca45612),
	.w4(32'hbb831414),
	.w5(32'hbb1a5865),
	.w6(32'hbc8c85e4),
	.w7(32'hbb89df36),
	.w8(32'hbb439dbf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06c2bb),
	.w1(32'h3b1794a9),
	.w2(32'h3b963a10),
	.w3(32'hbb08fab1),
	.w4(32'hb9cc231c),
	.w5(32'hba653430),
	.w6(32'hbb035374),
	.w7(32'hbb0838a6),
	.w8(32'h3a8ac9e3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad66f7),
	.w1(32'hbca80768),
	.w2(32'h3abd9057),
	.w3(32'hbbb479ee),
	.w4(32'hbc922036),
	.w5(32'h3b87dedf),
	.w6(32'hbb75f0d3),
	.w7(32'hbbaeaf63),
	.w8(32'h3c43c85a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc8de76),
	.w1(32'hbc68f471),
	.w2(32'h3c12828b),
	.w3(32'hbc805d6c),
	.w4(32'hbb7a255e),
	.w5(32'h3bf9c828),
	.w6(32'hbbc0a699),
	.w7(32'hbb8e103f),
	.w8(32'h3c4a3136),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf9e75),
	.w1(32'hbc054982),
	.w2(32'hbc0351a1),
	.w3(32'h3b1bbee6),
	.w4(32'hbc004a7f),
	.w5(32'hbbd9e903),
	.w6(32'h390c6c09),
	.w7(32'hbc0307dd),
	.w8(32'hbb74a3ec),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1b8e4),
	.w1(32'hbc0e354f),
	.w2(32'h3b4fdbc5),
	.w3(32'hbce21ec6),
	.w4(32'hbccc5656),
	.w5(32'hbc05b436),
	.w6(32'hbc67e493),
	.w7(32'hbc098fbf),
	.w8(32'h3c1ec2bf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d380e),
	.w1(32'h3c8dbc3f),
	.w2(32'h3cae39ca),
	.w3(32'h3a375de9),
	.w4(32'h3cb19437),
	.w5(32'h3cc51e88),
	.w6(32'h3b76e377),
	.w7(32'h3c86925c),
	.w8(32'h3ca2bfc8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc69dc7),
	.w1(32'h3c3665df),
	.w2(32'h3c8912c4),
	.w3(32'h3c9fae4c),
	.w4(32'h3c6081a0),
	.w5(32'h3c88a194),
	.w6(32'h3cca4b04),
	.w7(32'h3c41544c),
	.w8(32'h3b6b339f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5efeed),
	.w1(32'hbc71566c),
	.w2(32'hbc8f91c3),
	.w3(32'hba812562),
	.w4(32'hbc5b5ae2),
	.w5(32'hbc7de29c),
	.w6(32'h3b672142),
	.w7(32'hbc402a29),
	.w8(32'hbcb135ec),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa526d),
	.w1(32'hbbb9db56),
	.w2(32'h3b56730b),
	.w3(32'hbc00187e),
	.w4(32'hbc329278),
	.w5(32'hba6b9880),
	.w6(32'hbb45faf1),
	.w7(32'h39d50f59),
	.w8(32'h3ab30352),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ba492),
	.w1(32'hbb0fe11e),
	.w2(32'h3b361733),
	.w3(32'h3aa05fea),
	.w4(32'hba1876ef),
	.w5(32'h3b1baf9b),
	.w6(32'hbb13e040),
	.w7(32'h3b9b9c34),
	.w8(32'h390b4adc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc469747),
	.w1(32'hbc15c026),
	.w2(32'h3b831e42),
	.w3(32'hba51908c),
	.w4(32'h3c60eacc),
	.w5(32'h3cb31901),
	.w6(32'hbc3548ca),
	.w7(32'h3ae7c9e3),
	.w8(32'h3c800396),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb772533),
	.w1(32'hba30a053),
	.w2(32'hbb93d81d),
	.w3(32'h3bb139e0),
	.w4(32'h3b164be5),
	.w5(32'hba092251),
	.w6(32'h3aace800),
	.w7(32'h3bff000d),
	.w8(32'h3aaa0924),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca23729),
	.w1(32'hbc8b725f),
	.w2(32'h3a72e8ec),
	.w3(32'hbd0ce651),
	.w4(32'hbcc22e15),
	.w5(32'hbb75a7d0),
	.w6(32'hbc33a725),
	.w7(32'h3ab4d651),
	.w8(32'h3c02a875),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b69f0),
	.w1(32'hbc0b04a6),
	.w2(32'hbbbad89a),
	.w3(32'hba435cba),
	.w4(32'hbb3c6647),
	.w5(32'h3b6cd4f1),
	.w6(32'hbb4a4713),
	.w7(32'hbc0da8b1),
	.w8(32'hbb605fca),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba82617),
	.w1(32'hbba73efc),
	.w2(32'h3ae5028c),
	.w3(32'hbb81b7c4),
	.w4(32'hbb4bad00),
	.w5(32'h3b1eee10),
	.w6(32'hbba81edf),
	.w7(32'hbbfbeed2),
	.w8(32'hbb4fc832),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95f3a6),
	.w1(32'hbb302403),
	.w2(32'h3ad7c3fe),
	.w3(32'h3792a313),
	.w4(32'hbbe09b9d),
	.w5(32'hbb01bcff),
	.w6(32'hbae8a050),
	.w7(32'hbc19c37b),
	.w8(32'hbb89610c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb098a27),
	.w1(32'h3bb6c1cf),
	.w2(32'h3ba65fba),
	.w3(32'hbb0fd3ae),
	.w4(32'h3c1f14f3),
	.w5(32'h3c217cdf),
	.w6(32'hbc148983),
	.w7(32'h3a01647c),
	.w8(32'h3b30e8e9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01a0d6),
	.w1(32'hb9c274cd),
	.w2(32'h3babf797),
	.w3(32'h3a0b23b2),
	.w4(32'h3b746515),
	.w5(32'hba77796b),
	.w6(32'hbb0e04d1),
	.w7(32'hbb87b412),
	.w8(32'hbbbb2772),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7e703),
	.w1(32'hbaf8597e),
	.w2(32'h3818d93f),
	.w3(32'hbc305b69),
	.w4(32'hba17fa0d),
	.w5(32'h3b87c879),
	.w6(32'hbc67642a),
	.w7(32'hbc0ea648),
	.w8(32'h3a90beff),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97f81c),
	.w1(32'hbc502b5a),
	.w2(32'hbbc0fe53),
	.w3(32'h39888220),
	.w4(32'h3b6a9e89),
	.w5(32'h3c4d4721),
	.w6(32'h3c010b5e),
	.w7(32'h3c81aa5e),
	.w8(32'h3c73dfa3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabd28e),
	.w1(32'hbba914fe),
	.w2(32'h3b8ad526),
	.w3(32'hbbfc6992),
	.w4(32'h3a8ee6d3),
	.w5(32'h3b70aade),
	.w6(32'hbbb8692a),
	.w7(32'hbb15a27d),
	.w8(32'hbb161611),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fb0b13),
	.w1(32'hba7f8957),
	.w2(32'hb92562d9),
	.w3(32'hba413dee),
	.w4(32'hbb400b23),
	.w5(32'hbbd3d06b),
	.w6(32'hbbfe663a),
	.w7(32'hbb1dddee),
	.w8(32'hbb3c9e98),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba576226),
	.w1(32'h3c16237c),
	.w2(32'h3bb1c959),
	.w3(32'hbbebd60f),
	.w4(32'h3b8a8daa),
	.w5(32'hba35c9de),
	.w6(32'hbb0798e7),
	.w7(32'h3ba0e283),
	.w8(32'hb92e572c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f51f8),
	.w1(32'h3bfccd48),
	.w2(32'h3b3786b3),
	.w3(32'h3bd9941a),
	.w4(32'h3c104cd2),
	.w5(32'h3b8e8f21),
	.w6(32'h3b959a88),
	.w7(32'h3bb47cb4),
	.w8(32'h3ad37146),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8c326),
	.w1(32'h3ba6fb6f),
	.w2(32'h3bbc236a),
	.w3(32'hbc11c55d),
	.w4(32'h3c9005f4),
	.w5(32'h3cb8fae6),
	.w6(32'h3ae6813a),
	.w7(32'h3cab1b26),
	.w8(32'h3c9983f6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb73140),
	.w1(32'h3a2bab5d),
	.w2(32'h3b108f0b),
	.w3(32'h3c7d8768),
	.w4(32'h3b1b92fb),
	.w5(32'h3a17f27e),
	.w6(32'h3c403dda),
	.w7(32'h3ac663be),
	.w8(32'h3b0610cb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d063e8f),
	.w1(32'h3cb71e7a),
	.w2(32'h3c6976f5),
	.w3(32'hbbb224db),
	.w4(32'hbce25ce3),
	.w5(32'hbd0920c8),
	.w6(32'hbc0bb8ce),
	.w7(32'hbcdf16da),
	.w8(32'hb98a843c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e04ea),
	.w1(32'hbc83591f),
	.w2(32'h3c0913eb),
	.w3(32'hba88d340),
	.w4(32'hbc0d95c7),
	.w5(32'h3c8ca381),
	.w6(32'hbb1db62c),
	.w7(32'hbc7684f4),
	.w8(32'h3c3d573f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1db3f0),
	.w1(32'hbbb8b664),
	.w2(32'h3bdcf7b3),
	.w3(32'h3ba37195),
	.w4(32'hb9717d80),
	.w5(32'h3c0234c2),
	.w6(32'hbb466d86),
	.w7(32'hbc44641a),
	.w8(32'h3bd08aef),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c74006),
	.w1(32'hbb0d7a9b),
	.w2(32'hbc173842),
	.w3(32'h3c364b2c),
	.w4(32'hbbaf70ca),
	.w5(32'hbc1ce08a),
	.w6(32'hbc227916),
	.w7(32'hbbb36222),
	.w8(32'hbc2adaa8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa2e28),
	.w1(32'hbc1ad7ea),
	.w2(32'h3ba7c255),
	.w3(32'hbc16a68a),
	.w4(32'h3cb88fc0),
	.w5(32'hba95a0cd),
	.w6(32'hbb938852),
	.w7(32'h3b16b3fe),
	.w8(32'h3b24911b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc78422),
	.w1(32'hbcbc4381),
	.w2(32'hbc0a51bb),
	.w3(32'h3c0167c0),
	.w4(32'hbcc78e6f),
	.w5(32'h3c3f64ca),
	.w6(32'hbbd1eb5e),
	.w7(32'hbca8ed23),
	.w8(32'h3baaab34),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87861f),
	.w1(32'h3a583ca2),
	.w2(32'h3c085a95),
	.w3(32'h3c647307),
	.w4(32'h3b8b72dc),
	.w5(32'hbb147e9a),
	.w6(32'hbc01d473),
	.w7(32'hbb0602ec),
	.w8(32'h3c9637b0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e3a2),
	.w1(32'hbc6f9efb),
	.w2(32'hbb97be4f),
	.w3(32'h3c4473b3),
	.w4(32'hbcbb8109),
	.w5(32'h3bb8907a),
	.w6(32'h3c324ebc),
	.w7(32'hbd179360),
	.w8(32'h3cc1aa50),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86828e),
	.w1(32'h3a4a6971),
	.w2(32'h3b3d399a),
	.w3(32'h3c974685),
	.w4(32'hbc7ed06a),
	.w5(32'hbb733bd8),
	.w6(32'h3bbf2ab6),
	.w7(32'hbbcfb68b),
	.w8(32'h3c332d9d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8658a),
	.w1(32'hbcedc544),
	.w2(32'h3c443c3a),
	.w3(32'hbc0395a2),
	.w4(32'hbc558c3f),
	.w5(32'h3ca3ccda),
	.w6(32'hbb176c37),
	.w7(32'hbc4224fc),
	.w8(32'h3c867871),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164a13),
	.w1(32'hbb80ecce),
	.w2(32'hbc2902e0),
	.w3(32'h3befc764),
	.w4(32'h3c84e1d5),
	.w5(32'h3c3ed7e4),
	.w6(32'h3a3f6921),
	.w7(32'hbaa21b11),
	.w8(32'hbbb71447),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe094a7),
	.w1(32'h3c4f3304),
	.w2(32'hbcc87445),
	.w3(32'h3c975b03),
	.w4(32'hbc7597df),
	.w5(32'hbbaaa6b2),
	.w6(32'hbc134601),
	.w7(32'hbb0a7768),
	.w8(32'hbbff983a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bb0f4),
	.w1(32'h3c22f79e),
	.w2(32'h3a31337c),
	.w3(32'h3c75a55c),
	.w4(32'h3bf82b0b),
	.w5(32'h3ab999cd),
	.w6(32'hbc8ef7bf),
	.w7(32'hbc279122),
	.w8(32'hbc2f1cc4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb741fc),
	.w1(32'h394a842f),
	.w2(32'h3b03c8ae),
	.w3(32'hbb6d68a7),
	.w4(32'hbd16e7fb),
	.w5(32'h3c28f81f),
	.w6(32'hbab1dcd3),
	.w7(32'hbcd43e82),
	.w8(32'h3c751876),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb922c),
	.w1(32'hbc8d8509),
	.w2(32'hbc2b6595),
	.w3(32'h3d2f5b80),
	.w4(32'h3c57c433),
	.w5(32'h3c6fa4a6),
	.w6(32'h3d3304d4),
	.w7(32'h3c5809c6),
	.w8(32'h388688a4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a7b3e),
	.w1(32'hbd29f350),
	.w2(32'h3c634a09),
	.w3(32'h3b910c1a),
	.w4(32'hbcfff9f8),
	.w5(32'h3cb90d97),
	.w6(32'h3ca7bdda),
	.w7(32'hbcea1cf2),
	.w8(32'h3cc3d52a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15af60),
	.w1(32'hbc4ab3aa),
	.w2(32'h3c637720),
	.w3(32'h3c8f1b03),
	.w4(32'h3cd91b74),
	.w5(32'h3c9d971d),
	.w6(32'hba722a59),
	.w7(32'h3c5963a2),
	.w8(32'h3c123609),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc269038),
	.w1(32'hbcb3d416),
	.w2(32'hbbc2e15e),
	.w3(32'h3c4b325e),
	.w4(32'hbd2d0df5),
	.w5(32'h3cd3ac5c),
	.w6(32'h3b9cd15a),
	.w7(32'hbc6487b7),
	.w8(32'h3c4d7d5b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c131588),
	.w1(32'hbd070ea1),
	.w2(32'h392dfa6b),
	.w3(32'h3c1de90e),
	.w4(32'hbcc48e1a),
	.w5(32'h3c47c333),
	.w6(32'h3cb14bcf),
	.w7(32'hbcdd1e03),
	.w8(32'h3c4671ca),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8da75),
	.w1(32'h3bbf5c27),
	.w2(32'h3c01bd3c),
	.w3(32'h3c312495),
	.w4(32'hba7c2f54),
	.w5(32'h3d1f3599),
	.w6(32'h3ba2cd1a),
	.w7(32'h3b1499af),
	.w8(32'h3c67ed84),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17f756),
	.w1(32'h3b4d9f26),
	.w2(32'hba5f7814),
	.w3(32'h3b644b25),
	.w4(32'hbc116da1),
	.w5(32'hbb92d7f9),
	.w6(32'h3c3144d6),
	.w7(32'h39f3eab5),
	.w8(32'hbaadd49e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96db15),
	.w1(32'hbc6a767c),
	.w2(32'h3cd6a639),
	.w3(32'hbb45f2a8),
	.w4(32'hbad7053b),
	.w5(32'h3d3fd223),
	.w6(32'h3b5512ae),
	.w7(32'hbc89b6a6),
	.w8(32'h3ce27548),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c2797),
	.w1(32'hbb4b378d),
	.w2(32'hbcf84895),
	.w3(32'h3abf86f0),
	.w4(32'hbd1d5a22),
	.w5(32'hbd02e3f4),
	.w6(32'hbc2ad25c),
	.w7(32'hbc5600c4),
	.w8(32'hbcc3e976),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb285451),
	.w1(32'h3bdc4c07),
	.w2(32'hbc4a6d78),
	.w3(32'h3ae5b149),
	.w4(32'h3ae1f755),
	.w5(32'hbc0cbed9),
	.w6(32'hbc1d7640),
	.w7(32'hbc0cae0b),
	.w8(32'hbc6d19e7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaae5b),
	.w1(32'hbad5ec1b),
	.w2(32'hbab1c6d8),
	.w3(32'hbc198851),
	.w4(32'h3a603a93),
	.w5(32'h3a8c82af),
	.w6(32'hbbdd4193),
	.w7(32'hbb926758),
	.w8(32'h3a8f9e67),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc931f0),
	.w1(32'hbc6cc844),
	.w2(32'hbc89dce0),
	.w3(32'h3a941885),
	.w4(32'hbccb9ee0),
	.w5(32'hbd5b4ca7),
	.w6(32'hbb7ca3e0),
	.w7(32'hbc798c13),
	.w8(32'hbcca6ae1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd34082f),
	.w1(32'hbcd53f04),
	.w2(32'hbaa1a179),
	.w3(32'hbd0139c9),
	.w4(32'hbc85897e),
	.w5(32'h3c9061aa),
	.w6(32'hbc6cd45f),
	.w7(32'hbc94bd65),
	.w8(32'h3c797725),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf84a6c),
	.w1(32'hbaf41d88),
	.w2(32'hbb77eb4b),
	.w3(32'h3baf8eab),
	.w4(32'hbb42fc4f),
	.w5(32'hb9f99446),
	.w6(32'hbbab40b6),
	.w7(32'hbb06e031),
	.w8(32'hbad4b861),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed8ff3),
	.w1(32'h3c244445),
	.w2(32'h3c1b0813),
	.w3(32'hbb91b32f),
	.w4(32'h3ae08854),
	.w5(32'h3bc479a8),
	.w6(32'hbb033ec7),
	.w7(32'hbc73c883),
	.w8(32'h3c24a8df),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefe6e3),
	.w1(32'h3c0d3880),
	.w2(32'hbb72a4d1),
	.w3(32'h3cac4ae3),
	.w4(32'h3b450763),
	.w5(32'hb9450791),
	.w6(32'h3c214661),
	.w7(32'h3b2917d4),
	.w8(32'hba9872d1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36cada),
	.w1(32'h3be055f2),
	.w2(32'hbbdb29f8),
	.w3(32'hbba9ccf2),
	.w4(32'h3a4ab468),
	.w5(32'hbc4e165b),
	.w6(32'hbb950bdb),
	.w7(32'h3b8388fd),
	.w8(32'hbb33e418),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba950b74),
	.w1(32'hbcf7a6d3),
	.w2(32'h3ba278e9),
	.w3(32'h3c5372c4),
	.w4(32'hbc9279f6),
	.w5(32'h3c9c8545),
	.w6(32'h3bfd4319),
	.w7(32'hbc32781f),
	.w8(32'h3cd652f8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3ccb1),
	.w1(32'h3c07b4f2),
	.w2(32'hbba426eb),
	.w3(32'h3c227b99),
	.w4(32'hba0824a1),
	.w5(32'hbc4fd6e8),
	.w6(32'hbc486a69),
	.w7(32'hbb988d4c),
	.w8(32'h3c4956b8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f6471),
	.w1(32'h3ac67403),
	.w2(32'hbc6d2340),
	.w3(32'h3b70bf40),
	.w4(32'hbb70c81e),
	.w5(32'hbc96b92f),
	.w6(32'hbb11ea7a),
	.w7(32'hbc5eb963),
	.w8(32'hbcd0b724),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab6771),
	.w1(32'h3d136569),
	.w2(32'h3c4d0d65),
	.w3(32'hbb0cd4d2),
	.w4(32'h3d04ccb5),
	.w5(32'h3bbbd15c),
	.w6(32'hbc08e1c8),
	.w7(32'h3cbc5897),
	.w8(32'hbac8ab71),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcbc44),
	.w1(32'hbc777bd9),
	.w2(32'hbab92ec3),
	.w3(32'hb9d44cfd),
	.w4(32'hbbdfa56f),
	.w5(32'h3d0d5cb1),
	.w6(32'h3c24626f),
	.w7(32'hbbcf1330),
	.w8(32'h3cb70651),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf42706),
	.w1(32'hbc0c4c2c),
	.w2(32'h3ba10dd3),
	.w3(32'h3c430cf5),
	.w4(32'hbc7949f9),
	.w5(32'h3b335f90),
	.w6(32'hbd218577),
	.w7(32'hbc86c42f),
	.w8(32'h3b7221c5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11ae2e),
	.w1(32'h3c571bb0),
	.w2(32'h3ab8e507),
	.w3(32'h3b8e802c),
	.w4(32'h3c087945),
	.w5(32'hbb6a661a),
	.w6(32'h3bf19b75),
	.w7(32'h3c1aa9e5),
	.w8(32'hbb8b6c9d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9079a7),
	.w1(32'hbc95dcab),
	.w2(32'hbc1aacf9),
	.w3(32'hbb972f17),
	.w4(32'hbc82c487),
	.w5(32'hbc047831),
	.w6(32'hbb23d93f),
	.w7(32'hbccf8bfb),
	.w8(32'hbca43064),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe4da8),
	.w1(32'hbcb79de4),
	.w2(32'h3b2cf9a4),
	.w3(32'hbc25a6bf),
	.w4(32'hbcb06aff),
	.w5(32'hbc1cef58),
	.w6(32'hbbf6692c),
	.w7(32'h39af599a),
	.w8(32'h3c8b347c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c469655),
	.w1(32'hbca20e72),
	.w2(32'h3bf52de8),
	.w3(32'h3cae4d0c),
	.w4(32'h39c23b41),
	.w5(32'h3ca0d1a7),
	.w6(32'h3c20a35c),
	.w7(32'hbc113a4d),
	.w8(32'h3c0eec88),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91d640),
	.w1(32'hbd11001b),
	.w2(32'hbca18c89),
	.w3(32'hbb738d03),
	.w4(32'hbc03cb5b),
	.w5(32'hbcfc71b4),
	.w6(32'hbb376547),
	.w7(32'hbced2951),
	.w8(32'hbbf9ac13),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9225fe),
	.w1(32'hbb4c2fc2),
	.w2(32'h3cc1da72),
	.w3(32'h3c53a631),
	.w4(32'hbb135e71),
	.w5(32'h3c25bae3),
	.w6(32'h38c6fe8e),
	.w7(32'hbba1a0f1),
	.w8(32'h3b874a7d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f1ef7),
	.w1(32'hb992146b),
	.w2(32'hbb54efc5),
	.w3(32'hbc0f9395),
	.w4(32'hbaa48835),
	.w5(32'hbbfbc351),
	.w6(32'h3c17974c),
	.w7(32'h39d2a55d),
	.w8(32'hbb94d19c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45ddaa),
	.w1(32'h3db5af51),
	.w2(32'hbe400d32),
	.w3(32'hbaab5398),
	.w4(32'hbe584171),
	.w5(32'h3eaf3ff7),
	.w6(32'h3bcb991a),
	.w7(32'h3db8fc18),
	.w8(32'hbe1157cf),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3de50fd7),
	.w1(32'hbc1be7d8),
	.w2(32'h3c86404b),
	.w3(32'hbe2cf8d4),
	.w4(32'h3a515558),
	.w5(32'h3c83e044),
	.w6(32'h3d8887c8),
	.w7(32'hbc187657),
	.w8(32'h3c123c37),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ebbae),
	.w1(32'h3b655b57),
	.w2(32'hbba0d333),
	.w3(32'hbc191e07),
	.w4(32'hb975882a),
	.w5(32'hbc08b4d9),
	.w6(32'hbbde6e06),
	.w7(32'hb9fc0ac1),
	.w8(32'hbbe082a9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4990fe),
	.w1(32'hbc8ac12a),
	.w2(32'h3c874b27),
	.w3(32'hbbfcf920),
	.w4(32'hbc0cd1fe),
	.w5(32'hbc533521),
	.w6(32'hbbf1d3cb),
	.w7(32'hbc7b62aa),
	.w8(32'hba4cf38d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d687a),
	.w1(32'hbc725ae0),
	.w2(32'h3b68e326),
	.w3(32'hbaa19cd9),
	.w4(32'hbc99c407),
	.w5(32'h3d332543),
	.w6(32'hbc0edfa2),
	.w7(32'hbbbaa01e),
	.w8(32'hbbc583d0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ea5a1),
	.w1(32'hbce877f9),
	.w2(32'hbc30abb5),
	.w3(32'hbc9825e5),
	.w4(32'hbae6066d),
	.w5(32'h3c900615),
	.w6(32'h3d0d7a9f),
	.w7(32'hbb9be416),
	.w8(32'hbc7ae884),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c6d48),
	.w1(32'hbb857b06),
	.w2(32'hbb1511ac),
	.w3(32'hbca1e805),
	.w4(32'hbb432e2b),
	.w5(32'hbb4f8413),
	.w6(32'h3aa1b73b),
	.w7(32'hbb3c79cd),
	.w8(32'hbb938e96),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01b3e9),
	.w1(32'hbc0ea987),
	.w2(32'hbb34c4ff),
	.w3(32'hb5095700),
	.w4(32'h3b04d3c1),
	.w5(32'h3c09b10b),
	.w6(32'hbc333f2e),
	.w7(32'h3ab31218),
	.w8(32'h3c00339b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9acccd),
	.w1(32'h3b4e05b5),
	.w2(32'hbb5b1923),
	.w3(32'h3c10282a),
	.w4(32'hbb9b74be),
	.w5(32'hbbbef20b),
	.w6(32'h3b4dd689),
	.w7(32'hbb838e97),
	.w8(32'hbbaff322),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a684018),
	.w1(32'h3b83a776),
	.w2(32'hbb3942f2),
	.w3(32'hbb991789),
	.w4(32'h3af3920b),
	.w5(32'hbc01f1ed),
	.w6(32'hbbf92cd1),
	.w7(32'hbb1b1001),
	.w8(32'hbc2314f3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5898f3),
	.w1(32'hbc03c8a2),
	.w2(32'hbcc1fd57),
	.w3(32'hbb89e176),
	.w4(32'hbd43bd9b),
	.w5(32'h3ca054c6),
	.w6(32'hbbb31393),
	.w7(32'hbc557f27),
	.w8(32'h3b0b67fe),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc368a3b),
	.w1(32'h3bcc3293),
	.w2(32'h3bdde5e4),
	.w3(32'hbb00aa4a),
	.w4(32'h3cd21e09),
	.w5(32'h3cda8d76),
	.w6(32'hbcd1cdcd),
	.w7(32'h3c21e90c),
	.w8(32'h3c36685e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc005504),
	.w1(32'hbb98c6fc),
	.w2(32'hbc17069f),
	.w3(32'h3c104e88),
	.w4(32'hbc0668ea),
	.w5(32'hbbe36e47),
	.w6(32'hbb3ed8e2),
	.w7(32'hbc54c33c),
	.w8(32'h3bc4bbcc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49a75d),
	.w1(32'hbb7c2193),
	.w2(32'hbb8b0548),
	.w3(32'hbb754fb1),
	.w4(32'hbb2a1795),
	.w5(32'hbbf6e887),
	.w6(32'hbc5657a8),
	.w7(32'h3921cfa4),
	.w8(32'hbbd84128),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb745aec),
	.w1(32'hbd39316a),
	.w2(32'h3c7cf66b),
	.w3(32'hbc818b90),
	.w4(32'hbd124a80),
	.w5(32'hbcbba1c9),
	.w6(32'hbc23e5bb),
	.w7(32'hbd3e3c5e),
	.w8(32'h3bfe2d34),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule