module layer_10_featuremap_340(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabca8c3),
	.w1(32'h3abb3a20),
	.w2(32'hbb2645fe),
	.w3(32'hbb3a780b),
	.w4(32'hbb1315e3),
	.w5(32'hba5bce65),
	.w6(32'hba968838),
	.w7(32'hbb3f1dbe),
	.w8(32'h3b595d0a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9866e4e),
	.w1(32'h3b2a1633),
	.w2(32'h3ac2e499),
	.w3(32'hbb1fa8f9),
	.w4(32'h3982bf95),
	.w5(32'h3b15d651),
	.w6(32'h3b24fd79),
	.w7(32'h3abe7229),
	.w8(32'h3ba08d9a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad99dd2),
	.w1(32'h3b051ccd),
	.w2(32'hba87b9ff),
	.w3(32'h3b02ffdf),
	.w4(32'h3b09a7ec),
	.w5(32'hba62dd43),
	.w6(32'h3b795615),
	.w7(32'h3b880f63),
	.w8(32'h3aeb8ed3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bb984),
	.w1(32'hba2304f7),
	.w2(32'hba451374),
	.w3(32'h391abb50),
	.w4(32'h39898e6c),
	.w5(32'h3a43acfb),
	.w6(32'h3b40ca2f),
	.w7(32'h39cb2f26),
	.w8(32'hbb752372),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b458b9c),
	.w1(32'hba9f1c9d),
	.w2(32'h3aeae99e),
	.w3(32'hbad30103),
	.w4(32'h3a9e0d73),
	.w5(32'hba8baf01),
	.w6(32'hbaf861b9),
	.w7(32'hbb35d0fe),
	.w8(32'h399097c6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9ab48),
	.w1(32'hbb580431),
	.w2(32'hbb1ec7cc),
	.w3(32'hb96efaa2),
	.w4(32'h3b035f8c),
	.w5(32'h3a8ec05c),
	.w6(32'h3a96209e),
	.w7(32'h376f7c60),
	.w8(32'h3af4a4f0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba959645),
	.w1(32'hb88bcea1),
	.w2(32'h3b3e49e2),
	.w3(32'h3ae000f4),
	.w4(32'h3b4af154),
	.w5(32'hbb9369fe),
	.w6(32'h3b93b896),
	.w7(32'h3ae59339),
	.w8(32'hbb7c7120),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb468333),
	.w1(32'hbb4a4229),
	.w2(32'hbb7cbc8e),
	.w3(32'hbb2a45fc),
	.w4(32'hbab00786),
	.w5(32'hba008320),
	.w6(32'hba2da3ee),
	.w7(32'hbb459784),
	.w8(32'hbb547e19),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ab0bd),
	.w1(32'hbb73ecb0),
	.w2(32'hbae84f8b),
	.w3(32'hb81f9fdb),
	.w4(32'h3a64645f),
	.w5(32'hbaa1331a),
	.w6(32'hbaddac32),
	.w7(32'hbab1adca),
	.w8(32'hb779ecea),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f9552),
	.w1(32'hbb0305a3),
	.w2(32'hbac4e407),
	.w3(32'h3a8487df),
	.w4(32'h3b0f1860),
	.w5(32'hba98bb99),
	.w6(32'h39f7d9e4),
	.w7(32'hb981ad52),
	.w8(32'hba91cb52),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94be20),
	.w1(32'hbac702d5),
	.w2(32'h3a36c3a0),
	.w3(32'hba9cdda3),
	.w4(32'h3b4245d7),
	.w5(32'hbaf68558),
	.w6(32'h3b8d3a2a),
	.w7(32'hba8d7c48),
	.w8(32'hba5a57b6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e7c1a),
	.w1(32'hba1f677d),
	.w2(32'h39ad4afc),
	.w3(32'hbb7189b1),
	.w4(32'hbae77850),
	.w5(32'hbab59c3d),
	.w6(32'h3b25864b),
	.w7(32'hb7c62e58),
	.w8(32'h3a9b0f05),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3c264),
	.w1(32'hbb999ce9),
	.w2(32'hba959a6d),
	.w3(32'hbb03a7cd),
	.w4(32'hbb029e3b),
	.w5(32'hbac451d1),
	.w6(32'h3b888d02),
	.w7(32'h3b7ef5a5),
	.w8(32'hbb091907),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10ee76),
	.w1(32'hbb2cb69a),
	.w2(32'hba1a5ee7),
	.w3(32'hba187d30),
	.w4(32'h3b0992cf),
	.w5(32'hbb30209c),
	.w6(32'hbb3ca0e8),
	.w7(32'hba138176),
	.w8(32'hba4458e0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bdf45),
	.w1(32'hbb2854a3),
	.w2(32'hba6b5f89),
	.w3(32'hbb0536a3),
	.w4(32'h394ebff7),
	.w5(32'hbb052165),
	.w6(32'h3a842b06),
	.w7(32'h3ae98890),
	.w8(32'hbb2f97e6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d32a3),
	.w1(32'hbb29254d),
	.w2(32'h3ac799fc),
	.w3(32'hbb3d0c49),
	.w4(32'hbbca20b0),
	.w5(32'h3a95c349),
	.w6(32'h3ad5f04d),
	.w7(32'hba59ff94),
	.w8(32'hb943dc44),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4181f4),
	.w1(32'hbb63d8cc),
	.w2(32'hbacfe99e),
	.w3(32'hbac4b4a6),
	.w4(32'h3ab6fde1),
	.w5(32'h3a884709),
	.w6(32'h3b4d0ac1),
	.w7(32'hba20ea70),
	.w8(32'h3b774cf0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a6b68),
	.w1(32'hbac3f7ea),
	.w2(32'hbb03674b),
	.w3(32'h3af99ab3),
	.w4(32'h3b6234f7),
	.w5(32'h3b82a843),
	.w6(32'h3af4c91f),
	.w7(32'hbb08767e),
	.w8(32'hba64e802),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06979e),
	.w1(32'h3a1d73a1),
	.w2(32'hb984a1df),
	.w3(32'h3bae2d45),
	.w4(32'h3b32fa33),
	.w5(32'hbba0dfbc),
	.w6(32'h3b65cba8),
	.w7(32'h3b3aeec3),
	.w8(32'hbaaac26d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63b370),
	.w1(32'hba1b2f7d),
	.w2(32'hba0035f2),
	.w3(32'h3a6cb795),
	.w4(32'h3b3a091d),
	.w5(32'hbb83f4a5),
	.w6(32'h3abc5014),
	.w7(32'h3984b1ff),
	.w8(32'hbba66831),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53b661),
	.w1(32'h3abed466),
	.w2(32'hb9f592a9),
	.w3(32'h3b189acc),
	.w4(32'hbb56e42c),
	.w5(32'h3a257fde),
	.w6(32'h38f46e94),
	.w7(32'hbacfa7cc),
	.w8(32'hba35de16),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04f04b),
	.w1(32'hba13005a),
	.w2(32'hba26c25a),
	.w3(32'h3abadeeb),
	.w4(32'h3a95f4c4),
	.w5(32'hba6270b0),
	.w6(32'hbb12548e),
	.w7(32'hba8093b8),
	.w8(32'h3a0f23a1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba800cf0),
	.w1(32'hbb2cc578),
	.w2(32'h397e4d25),
	.w3(32'h3a9bfb98),
	.w4(32'hbab3d7f6),
	.w5(32'h3916a5e1),
	.w6(32'hba1a5ea4),
	.w7(32'hbb8a1ffa),
	.w8(32'hbbb3f6b1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac26832),
	.w1(32'hbb62fc76),
	.w2(32'h3af4138f),
	.w3(32'hba8ccd84),
	.w4(32'hbbaf3b89),
	.w5(32'h3ae065ea),
	.w6(32'hba4d5cca),
	.w7(32'hbb748ae7),
	.w8(32'hb9e6011f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abce5cb),
	.w1(32'h3bda7fe6),
	.w2(32'h3b829b1c),
	.w3(32'hbacb49fc),
	.w4(32'hbab60cc5),
	.w5(32'hb8b97f31),
	.w6(32'h3c051269),
	.w7(32'hbaf5642e),
	.w8(32'hbaf86ec2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab7956),
	.w1(32'hbb6d5b76),
	.w2(32'hb9e1444a),
	.w3(32'hb920186a),
	.w4(32'h3aff39d6),
	.w5(32'hb8b939ef),
	.w6(32'hba0201b9),
	.w7(32'hba2049f0),
	.w8(32'h3b085691),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82165d),
	.w1(32'hbaf01254),
	.w2(32'h3a0867e9),
	.w3(32'hbb355446),
	.w4(32'hba37d361),
	.w5(32'hbae591c6),
	.w6(32'hbb5856fa),
	.w7(32'h3ac65a70),
	.w8(32'hba6aacab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20e5a5),
	.w1(32'hba7a419f),
	.w2(32'hbb333a6e),
	.w3(32'hba7962a2),
	.w4(32'hba895dff),
	.w5(32'h3a23669f),
	.w6(32'hbabce525),
	.w7(32'hbb2a55a5),
	.w8(32'hbb2d8e71),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb5334),
	.w1(32'hbb263ccb),
	.w2(32'hba85583d),
	.w3(32'hb947800f),
	.w4(32'h3b533c1a),
	.w5(32'hbb5788b5),
	.w6(32'h3a884bf1),
	.w7(32'hba408507),
	.w8(32'h3a2df191),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba437c7e),
	.w1(32'hbbe6c7da),
	.w2(32'hbb7c5774),
	.w3(32'hbba8b7b2),
	.w4(32'h3b27e51d),
	.w5(32'h3b255278),
	.w6(32'hbb74db5f),
	.w7(32'hbb139741),
	.w8(32'hbb160df6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a2c23),
	.w1(32'h3c2c2c4b),
	.w2(32'h3b96e845),
	.w3(32'h3bf5fc9b),
	.w4(32'h3a3840f8),
	.w5(32'hb93e81c7),
	.w6(32'hbb74a5a8),
	.w7(32'hbbd20ec6),
	.w8(32'h3acf28c0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63818b),
	.w1(32'h3c057455),
	.w2(32'h3b942f71),
	.w3(32'h3af17bd5),
	.w4(32'h3981cdee),
	.w5(32'hbb030db2),
	.w6(32'h3c115d23),
	.w7(32'h3abde60f),
	.w8(32'hbb6cf7e5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb211e50),
	.w1(32'h3b8bb342),
	.w2(32'h3a2d89e9),
	.w3(32'hbb8a607c),
	.w4(32'hba407028),
	.w5(32'hbb15a708),
	.w6(32'hbb883e87),
	.w7(32'hb9cc12c2),
	.w8(32'h3afec51b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba7873),
	.w1(32'hbb396cc8),
	.w2(32'hbb13912f),
	.w3(32'hbb3a4a4f),
	.w4(32'h3b36aca0),
	.w5(32'hbafecee0),
	.w6(32'h3ac7843b),
	.w7(32'hbb96ac61),
	.w8(32'hba419cd9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d6f44),
	.w1(32'hba08fa85),
	.w2(32'hba2a5e8c),
	.w3(32'h3a392b53),
	.w4(32'hbb0c047f),
	.w5(32'h3b4b90e9),
	.w6(32'h3bc66535),
	.w7(32'hb9f0ea5a),
	.w8(32'hbc13dda8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb088c2b),
	.w1(32'h3b65825f),
	.w2(32'hbb023a76),
	.w3(32'h3b8a0fd7),
	.w4(32'h3b52c903),
	.w5(32'h3915e1a5),
	.w6(32'hbc0cb200),
	.w7(32'hbc3bd26f),
	.w8(32'hbb3c6251),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b140afc),
	.w1(32'h3b5831de),
	.w2(32'h37bef088),
	.w3(32'hba419d54),
	.w4(32'hbb47201b),
	.w5(32'hba0e4b68),
	.w6(32'hba1976e7),
	.w7(32'hbbf2b72d),
	.w8(32'h3b179a2e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a920ad7),
	.w1(32'hbafb4cbe),
	.w2(32'h3aa25ecb),
	.w3(32'hba56f00d),
	.w4(32'h3b250b7b),
	.w5(32'hbb4bbf38),
	.w6(32'hb9fcb78f),
	.w7(32'h3ae75a75),
	.w8(32'hbbab6289),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a924c5c),
	.w1(32'h3c2f73c5),
	.w2(32'h3bc12803),
	.w3(32'hba9fdd69),
	.w4(32'h3a86f620),
	.w5(32'h3a8618ed),
	.w6(32'hbbc78f52),
	.w7(32'hbc0f78cc),
	.w8(32'hbb122797),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a5068),
	.w1(32'hbbdd4dd8),
	.w2(32'hbbea2bb5),
	.w3(32'h3b2f2a80),
	.w4(32'hbb212eac),
	.w5(32'hbad2478f),
	.w6(32'hbb505c64),
	.w7(32'hbb3607e9),
	.w8(32'hb90282c2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ad16d),
	.w1(32'hbb0245ba),
	.w2(32'h3acbb8c6),
	.w3(32'hbb83f19b),
	.w4(32'h3a343c14),
	.w5(32'hba036178),
	.w6(32'h39488fea),
	.w7(32'hbb03ad56),
	.w8(32'h3aa92372),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945a6f3),
	.w1(32'hba396a14),
	.w2(32'h3ab4b8bb),
	.w3(32'hb9a472f9),
	.w4(32'h3ab8341a),
	.w5(32'hb9cb126d),
	.w6(32'h39e200da),
	.w7(32'hb93fb272),
	.w8(32'h3ac68d2c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21fb45),
	.w1(32'h3afde52c),
	.w2(32'h38f6921b),
	.w3(32'h385f770e),
	.w4(32'hba84bb9e),
	.w5(32'hbb0e39fc),
	.w6(32'h3bd625c8),
	.w7(32'h3a4cefc7),
	.w8(32'hbabe9608),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43c9e1),
	.w1(32'h3acb99fe),
	.w2(32'h3b8a5eb1),
	.w3(32'hbb2b7e85),
	.w4(32'h3b4fdf7d),
	.w5(32'h3b2696b0),
	.w6(32'h3c3ea2d8),
	.w7(32'hbb7a30fa),
	.w8(32'hbb6ba172),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94e5bb),
	.w1(32'hbac8558b),
	.w2(32'hbb3888c8),
	.w3(32'h3bb62d8d),
	.w4(32'h3b378b9d),
	.w5(32'hbac5c7ab),
	.w6(32'hbb9cc41c),
	.w7(32'h3a440011),
	.w8(32'hba552c1f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43c7e5),
	.w1(32'hbabfe1d7),
	.w2(32'h39c5d24d),
	.w3(32'hbb1e268a),
	.w4(32'hbb28ca95),
	.w5(32'hb89c28ed),
	.w6(32'hba8c18a8),
	.w7(32'hbb4ff89e),
	.w8(32'hbba43b3c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae29310),
	.w1(32'hbb91de8f),
	.w2(32'hbb2c5074),
	.w3(32'h3ad3e059),
	.w4(32'h3aa8f4da),
	.w5(32'hba0b8543),
	.w6(32'hbbe81e7c),
	.w7(32'hb9801996),
	.w8(32'hbab60bb5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c9fcb),
	.w1(32'h3a94e20b),
	.w2(32'h3adfc358),
	.w3(32'hba66a69c),
	.w4(32'h3974802b),
	.w5(32'hbb59b3c7),
	.w6(32'h39bf867c),
	.w7(32'hb9882ad8),
	.w8(32'h3acb8566),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13ee68),
	.w1(32'h3acd02c3),
	.w2(32'h3ae56787),
	.w3(32'hb9b06ef4),
	.w4(32'hba51b983),
	.w5(32'hba61ac96),
	.w6(32'h3a988470),
	.w7(32'h3b131d93),
	.w8(32'hb9e66df8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa637be),
	.w1(32'hbae223f6),
	.w2(32'hb9d61641),
	.w3(32'hba960106),
	.w4(32'hb98842c2),
	.w5(32'h3b576096),
	.w6(32'hbb78b569),
	.w7(32'hbac243e2),
	.w8(32'h3ade039b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad209f5),
	.w1(32'hba7eb2a7),
	.w2(32'h3ad4c1fa),
	.w3(32'hbb684510),
	.w4(32'hbb014bf5),
	.w5(32'hbad1acb7),
	.w6(32'hbb814c55),
	.w7(32'hbbaca75b),
	.w8(32'h3b177edc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f3c5a),
	.w1(32'h3b004c04),
	.w2(32'hba32fb2e),
	.w3(32'h3af66770),
	.w4(32'h3b869ba4),
	.w5(32'hbadb5f37),
	.w6(32'h3ba9128c),
	.w7(32'hbb79fd62),
	.w8(32'hba00010f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1207c3),
	.w1(32'hbb95da2c),
	.w2(32'h3ad44dc9),
	.w3(32'hbb47b470),
	.w4(32'h39ab39e1),
	.w5(32'hba62a47d),
	.w6(32'hb99b740b),
	.w7(32'hbb20478a),
	.w8(32'h3af137e1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e5b7b),
	.w1(32'hbaaa685b),
	.w2(32'hbb3048a5),
	.w3(32'hbba921b6),
	.w4(32'h398c4c38),
	.w5(32'hbb2361d8),
	.w6(32'hbadc3539),
	.w7(32'hbb51eb56),
	.w8(32'h3afc97f9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae685f2),
	.w1(32'h37533b84),
	.w2(32'hbaad3c00),
	.w3(32'hb921ea8e),
	.w4(32'hbb179f28),
	.w5(32'h3b831e13),
	.w6(32'h3c0b546d),
	.w7(32'h3a76fb08),
	.w8(32'h3bce8ee1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa662d),
	.w1(32'h3acf6f21),
	.w2(32'h3be3d8b7),
	.w3(32'h3b4cf4f7),
	.w4(32'h3b077033),
	.w5(32'h39a6d53d),
	.w6(32'h3c728009),
	.w7(32'h3bc05d2d),
	.w8(32'hba1a00e9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58336a),
	.w1(32'h3b7e2942),
	.w2(32'h3b8befd5),
	.w3(32'h3aa3da41),
	.w4(32'h3aeb20c0),
	.w5(32'hbb802fec),
	.w6(32'h3b8cefdb),
	.w7(32'h397642ac),
	.w8(32'hbab36d99),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d32ea),
	.w1(32'hbbcd010e),
	.w2(32'hbb5c4332),
	.w3(32'hbb2ab407),
	.w4(32'h3992c251),
	.w5(32'hb9f9875a),
	.w6(32'hbb7de002),
	.w7(32'hbb68865a),
	.w8(32'hbaeed189),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb095cf4),
	.w1(32'hbb099b04),
	.w2(32'h391753d6),
	.w3(32'hbafe01a9),
	.w4(32'hb95a5e85),
	.w5(32'h3ab4efb6),
	.w6(32'hbb3db241),
	.w7(32'hbaff8191),
	.w8(32'h3b9dcd08),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35f8c3),
	.w1(32'h3af8b767),
	.w2(32'h3b6ff4b5),
	.w3(32'hbb002002),
	.w4(32'h3b13825d),
	.w5(32'hbb161cb0),
	.w6(32'h3ac79b2b),
	.w7(32'h3b7b87da),
	.w8(32'hbae8add2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2e5d2),
	.w1(32'h3a6ea0d9),
	.w2(32'h3ab7208b),
	.w3(32'hb9942f11),
	.w4(32'h3a548912),
	.w5(32'hbb1f5499),
	.w6(32'hb973fd1b),
	.w7(32'hbb59a6ca),
	.w8(32'hbb136f33),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9b221),
	.w1(32'hbb5c9e26),
	.w2(32'hbb25da9d),
	.w3(32'hbac3b1d1),
	.w4(32'hbaf573f3),
	.w5(32'hbb887edf),
	.w6(32'h3aec8953),
	.w7(32'hba52c0ea),
	.w8(32'hbb8d4bca),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c5e17),
	.w1(32'hbb44bbc4),
	.w2(32'hbb5fd982),
	.w3(32'hbb57238e),
	.w4(32'hbbb607d1),
	.w5(32'hbb3974ea),
	.w6(32'h3b445be6),
	.w7(32'hbb56e0f0),
	.w8(32'hbb09a390),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae17c1),
	.w1(32'hbac30da9),
	.w2(32'hbae7eaf9),
	.w3(32'hbaa5e783),
	.w4(32'hba10eec3),
	.w5(32'hbb306366),
	.w6(32'hba933891),
	.w7(32'hbb3fd6a1),
	.w8(32'hbbc7ab8c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87b35e),
	.w1(32'hbbba5fe4),
	.w2(32'hba6667cd),
	.w3(32'h3aba76be),
	.w4(32'h3985e8ba),
	.w5(32'h3ae200be),
	.w6(32'h3bac345b),
	.w7(32'hb968d6bd),
	.w8(32'h3bd38ee0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11ad09),
	.w1(32'h39b2c58d),
	.w2(32'h39a49f79),
	.w3(32'hba387660),
	.w4(32'h398e660d),
	.w5(32'hba988419),
	.w6(32'h3c515c93),
	.w7(32'h3b8de160),
	.w8(32'hbb08eaf7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fab508),
	.w1(32'hbaf6da0d),
	.w2(32'hbb3e9f6c),
	.w3(32'hbb28407d),
	.w4(32'hba114b6e),
	.w5(32'hbb134189),
	.w6(32'h39be436e),
	.w7(32'hbb727325),
	.w8(32'hb7a305fe),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff888d),
	.w1(32'hba339bfd),
	.w2(32'hba8b8558),
	.w3(32'hba589a6b),
	.w4(32'h39e5a52b),
	.w5(32'hba933aee),
	.w6(32'h3a8cbac6),
	.w7(32'hba60d150),
	.w8(32'hbb8ed200),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0d923),
	.w1(32'h3aa03469),
	.w2(32'h3bcaeef9),
	.w3(32'hbb268a0e),
	.w4(32'h399612c8),
	.w5(32'h3b08b7cd),
	.w6(32'hba98c9ff),
	.w7(32'h3aea35bc),
	.w8(32'h3acc5c1e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0f885),
	.w1(32'h3a2ab43f),
	.w2(32'hbb5754e3),
	.w3(32'h3be43d93),
	.w4(32'h3c165a02),
	.w5(32'hbb05b8db),
	.w6(32'h3af536bf),
	.w7(32'hbba19acd),
	.w8(32'hbb094a70),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae76009),
	.w1(32'h3a978701),
	.w2(32'hbae72a13),
	.w3(32'h39eca7ef),
	.w4(32'hbaf3ded6),
	.w5(32'hba5436b5),
	.w6(32'hbaea0f60),
	.w7(32'hba89a86c),
	.w8(32'hbb5d4deb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2d243),
	.w1(32'h393266a0),
	.w2(32'hbaeec3cf),
	.w3(32'h3b2b0800),
	.w4(32'hbb0e6441),
	.w5(32'h3ba948bf),
	.w6(32'hbb5f3a0f),
	.w7(32'hbb1c02f8),
	.w8(32'hbbec5abd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23ca59),
	.w1(32'h3a41ebd3),
	.w2(32'hbaaab36b),
	.w3(32'h3c219861),
	.w4(32'h3baf0d4c),
	.w5(32'h3ad1f405),
	.w6(32'hbbe456a9),
	.w7(32'hbbe533d4),
	.w8(32'h3b448bbd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68a02c),
	.w1(32'h3a27df15),
	.w2(32'hbb31afde),
	.w3(32'h39ef8c33),
	.w4(32'h3be194ff),
	.w5(32'hbac84129),
	.w6(32'hb8477728),
	.w7(32'hbb825448),
	.w8(32'hba965b84),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb272729),
	.w1(32'hbb27ff56),
	.w2(32'hbad7d2d5),
	.w3(32'hbb363cc5),
	.w4(32'hba350e7e),
	.w5(32'h39ff7c2f),
	.w6(32'h3b901d0b),
	.w7(32'hbac9bbd4),
	.w8(32'h3b33a4ef),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08aba8),
	.w1(32'hba025e04),
	.w2(32'hbab4b89c),
	.w3(32'h3a6996d5),
	.w4(32'h3acf0388),
	.w5(32'h3a29388a),
	.w6(32'h3ac3eb95),
	.w7(32'hba651c0f),
	.w8(32'hba48faea),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98532ed),
	.w1(32'hba636ede),
	.w2(32'h3b8eb9d0),
	.w3(32'hbb1814c2),
	.w4(32'hbac5cbd2),
	.w5(32'hbaa2c6f6),
	.w6(32'h3a3a39a4),
	.w7(32'hbb0c2a2b),
	.w8(32'hbb6679b2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5440c3),
	.w1(32'hbaab94d1),
	.w2(32'hbb4b9710),
	.w3(32'hb9fca358),
	.w4(32'h3b606542),
	.w5(32'h3a072f4e),
	.w6(32'hbb429c5d),
	.w7(32'hbb9d8949),
	.w8(32'hbb1ec546),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0986df),
	.w1(32'hbac7a6bd),
	.w2(32'hbb68bad8),
	.w3(32'h3b2df9b8),
	.w4(32'h3b22eb5c),
	.w5(32'hbb3042ac),
	.w6(32'hbb09c5f9),
	.w7(32'hbb350f24),
	.w8(32'h3a652692),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbeac1),
	.w1(32'hb9f23527),
	.w2(32'hb925e504),
	.w3(32'hbae26472),
	.w4(32'h3aa5aef0),
	.w5(32'hbb65c61a),
	.w6(32'h3aff2f05),
	.w7(32'hba4655d8),
	.w8(32'h38d4269c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e4118),
	.w1(32'hbaf0ba84),
	.w2(32'hbba07c31),
	.w3(32'hbb017bcb),
	.w4(32'hbb6722b5),
	.w5(32'h3b743e39),
	.w6(32'hbb6a79e5),
	.w7(32'hbb2f53c0),
	.w8(32'h3a74a28f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fd3dd),
	.w1(32'h3b3dbb6e),
	.w2(32'h3af203e9),
	.w3(32'h3b9f968d),
	.w4(32'h3b8799a3),
	.w5(32'hbb26c42e),
	.w6(32'hb83bd4bf),
	.w7(32'hbb613165),
	.w8(32'hbbb686e8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1517f3),
	.w1(32'hba87c356),
	.w2(32'h3b5e5551),
	.w3(32'hba452977),
	.w4(32'h3a9dfd4a),
	.w5(32'h3aff95fc),
	.w6(32'hbb6d2529),
	.w7(32'hbb70213c),
	.w8(32'h3b5677ef),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09f5df),
	.w1(32'h3b6bfd7e),
	.w2(32'h3b9f296e),
	.w3(32'h3a487fc6),
	.w4(32'h39cc107e),
	.w5(32'hbadbb8fb),
	.w6(32'h3bdc5f66),
	.w7(32'h3c3457d6),
	.w8(32'h3ad5b18b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993bf88),
	.w1(32'hba1d6809),
	.w2(32'hba842d4f),
	.w3(32'hb98fd385),
	.w4(32'h39962767),
	.w5(32'hbb9cf7d1),
	.w6(32'h39c90425),
	.w7(32'hbb04a2c1),
	.w8(32'hbae98ffd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab85bae),
	.w1(32'h388e24a1),
	.w2(32'h39f1de71),
	.w3(32'hbb2dd2c9),
	.w4(32'hb9920c92),
	.w5(32'hbb6a2cf9),
	.w6(32'h3b2e8576),
	.w7(32'hbb410e2f),
	.w8(32'hbaceca2f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4952fd),
	.w1(32'hbb56ad4e),
	.w2(32'hbb3c2759),
	.w3(32'hbb966cc7),
	.w4(32'hbaf7b35d),
	.w5(32'hbad45842),
	.w6(32'hbb831ef6),
	.w7(32'hb97c3a26),
	.w8(32'hbb89451b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0e819),
	.w1(32'h390ab9d5),
	.w2(32'hb9e645d7),
	.w3(32'hbb51b55d),
	.w4(32'hbac91044),
	.w5(32'h3a9538b6),
	.w6(32'hbb3b9321),
	.w7(32'hbb64f5dc),
	.w8(32'h3ab13943),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad05c1f),
	.w1(32'hbabc74e3),
	.w2(32'h3a838208),
	.w3(32'h3a810eef),
	.w4(32'h3b39af16),
	.w5(32'hbb01130d),
	.w6(32'h3b39f621),
	.w7(32'h3ac2f2d0),
	.w8(32'hba82cfa9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d08d4),
	.w1(32'hbc18cff3),
	.w2(32'hbbe67a65),
	.w3(32'hbb82ea05),
	.w4(32'h3a1c89b0),
	.w5(32'h3b533ac8),
	.w6(32'hbbb8adf1),
	.w7(32'hbba6b7df),
	.w8(32'h3b56ad7b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dd09c),
	.w1(32'hba90f17b),
	.w2(32'hbad95f9b),
	.w3(32'h3acc6c3b),
	.w4(32'hbb2be53f),
	.w5(32'h3a9cfa25),
	.w6(32'h3a20bd5a),
	.w7(32'hbb46bb91),
	.w8(32'hb9f813f7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f4c22),
	.w1(32'hbbeda13f),
	.w2(32'hba506521),
	.w3(32'h3ab54143),
	.w4(32'h3aa5e34f),
	.w5(32'h3bd8e724),
	.w6(32'h3aaf330a),
	.w7(32'hbadff70e),
	.w8(32'h3bcb9742),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05ccee),
	.w1(32'h3c545f09),
	.w2(32'h3c625725),
	.w3(32'hbbafa3c3),
	.w4(32'hbb90a45d),
	.w5(32'h3b18ec9b),
	.w6(32'h3c368f01),
	.w7(32'h3929f0a8),
	.w8(32'h3b9fe1f7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89516d),
	.w1(32'hbaee61f9),
	.w2(32'hbb918b58),
	.w3(32'hb92f410d),
	.w4(32'hb9c910a9),
	.w5(32'hbae2ccd4),
	.w6(32'h3bbdb9e1),
	.w7(32'hbabe9ea6),
	.w8(32'hbb29b889),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23152d),
	.w1(32'hbb4b5750),
	.w2(32'hbb0ea164),
	.w3(32'hbb1106a3),
	.w4(32'hbafd03e8),
	.w5(32'hbaa0ce87),
	.w6(32'hbb949af4),
	.w7(32'hbba44574),
	.w8(32'h3b1ff834),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc4bb5),
	.w1(32'hbaa8894a),
	.w2(32'h3b30b022),
	.w3(32'hbbaf22fd),
	.w4(32'hbb8bf02f),
	.w5(32'h3af7b3bf),
	.w6(32'h3c43e595),
	.w7(32'h3c095e1e),
	.w8(32'hbabd1889),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc7c7b),
	.w1(32'hba643872),
	.w2(32'hbb6c051f),
	.w3(32'h3bba15ac),
	.w4(32'h3b84b399),
	.w5(32'h381bc217),
	.w6(32'hbba3ade0),
	.w7(32'hbb27da2f),
	.w8(32'hbb91275c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc96d6),
	.w1(32'h3b552106),
	.w2(32'h3b5e4e38),
	.w3(32'hb794307c),
	.w4(32'hbaa68643),
	.w5(32'hb84ee602),
	.w6(32'hbbb64b39),
	.w7(32'hbb895afd),
	.w8(32'hbaba0559),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ecf1c),
	.w1(32'h3a004241),
	.w2(32'hba38bffe),
	.w3(32'hba181f23),
	.w4(32'hb9b92659),
	.w5(32'hb789a349),
	.w6(32'hbaaf2d5a),
	.w7(32'hba0d10af),
	.w8(32'hbb3edad1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62c397),
	.w1(32'h3abee4e7),
	.w2(32'h39aa172a),
	.w3(32'hbb5a6cfe),
	.w4(32'hbb79df25),
	.w5(32'h39b25b15),
	.w6(32'hba62d74a),
	.w7(32'hbb42fe5f),
	.w8(32'h39eb1e32),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f5934),
	.w1(32'h3b0eca2a),
	.w2(32'hb9f853d6),
	.w3(32'hbaaeeead),
	.w4(32'hbb3b0476),
	.w5(32'hbb5db147),
	.w6(32'h3adf7c02),
	.w7(32'hbaf30171),
	.w8(32'hbab636a3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb8807),
	.w1(32'hbb0cdbd3),
	.w2(32'hbb804398),
	.w3(32'hbb2be74a),
	.w4(32'hbaefb111),
	.w5(32'h3a44bd0f),
	.w6(32'hba95b00f),
	.w7(32'hbb2f5be4),
	.w8(32'hbabe3332),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15f9aa),
	.w1(32'h3934bdd9),
	.w2(32'h3b16aa27),
	.w3(32'hbab6653e),
	.w4(32'hba84a433),
	.w5(32'hbb719fd4),
	.w6(32'hbb1a3a2a),
	.w7(32'hbab8dfe4),
	.w8(32'hbb59480c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82c1b6),
	.w1(32'hbba18572),
	.w2(32'hbb93e152),
	.w3(32'hbb6782b4),
	.w4(32'hbb0916a4),
	.w5(32'hb9517ead),
	.w6(32'hbb5ac9e5),
	.w7(32'hbb2397a3),
	.w8(32'h3b09121b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54a8fe),
	.w1(32'hb7c902d7),
	.w2(32'h3aa01a59),
	.w3(32'hbae70620),
	.w4(32'hbb0c75de),
	.w5(32'h3a3c90ff),
	.w6(32'h3aac4354),
	.w7(32'h3b429d2f),
	.w8(32'hb994699b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eec4a),
	.w1(32'h3a98a10d),
	.w2(32'hb950e32f),
	.w3(32'hbaace12b),
	.w4(32'hba126a5f),
	.w5(32'hb9c2cb3b),
	.w6(32'hba23c294),
	.w7(32'h37d3708d),
	.w8(32'hbad4101d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4c093),
	.w1(32'h3a9bdc15),
	.w2(32'hbafdb2ef),
	.w3(32'hbb3617d2),
	.w4(32'h3ac22eee),
	.w5(32'hba6826e8),
	.w6(32'hbaaaf59b),
	.w7(32'h3ab49f4b),
	.w8(32'hbab32721),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35177f),
	.w1(32'h3b121741),
	.w2(32'h3b0462cc),
	.w3(32'hbb4868e6),
	.w4(32'hbb1444dc),
	.w5(32'h3b50b2f6),
	.w6(32'h3a7197d7),
	.w7(32'hb98e5023),
	.w8(32'h3b47695a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5921),
	.w1(32'h3b6168b1),
	.w2(32'h3a8ef299),
	.w3(32'h3ad8594c),
	.w4(32'h3a62cb09),
	.w5(32'hbaf740c3),
	.w6(32'h3b51a041),
	.w7(32'h3b15a345),
	.w8(32'hbb329b0e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e2739),
	.w1(32'hbac1e10b),
	.w2(32'hb9a51747),
	.w3(32'hbac8d9fd),
	.w4(32'hbb191ff9),
	.w5(32'hb9f2a02b),
	.w6(32'hba1738fb),
	.w7(32'h39ad3e3c),
	.w8(32'h3a7b0a10),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b292343),
	.w1(32'h3a94060a),
	.w2(32'h3a873315),
	.w3(32'hbadca140),
	.w4(32'hbb219457),
	.w5(32'h3a8ed290),
	.w6(32'hb9c4e44c),
	.w7(32'hbb0ae302),
	.w8(32'hb9097804),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0ae3c),
	.w1(32'h3b0b04ef),
	.w2(32'hb98e17ab),
	.w3(32'hb98e7199),
	.w4(32'hbb059814),
	.w5(32'h3b5e5411),
	.w6(32'hba84d35d),
	.w7(32'hba911f8f),
	.w8(32'h3a9b6d6f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd123e),
	.w1(32'hb932f3b5),
	.w2(32'h3abe837d),
	.w3(32'h3b55f0b5),
	.w4(32'h3b4f5251),
	.w5(32'hba87ea8c),
	.w6(32'h3b2a0f90),
	.w7(32'h3b76c667),
	.w8(32'hba693710),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae408b9),
	.w1(32'h39b3a1be),
	.w2(32'hbb2ef553),
	.w3(32'hba11e1b5),
	.w4(32'hb93abf15),
	.w5(32'h39f56eb4),
	.w6(32'h3acea6d9),
	.w7(32'hbb139934),
	.w8(32'h3a12e53c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a3d2a),
	.w1(32'h3a9f53c6),
	.w2(32'hba32b9e5),
	.w3(32'h3aafa15f),
	.w4(32'hb8ab5108),
	.w5(32'h3abd5a93),
	.w6(32'h3a3698e2),
	.w7(32'hba60916b),
	.w8(32'hba302115),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48d28b),
	.w1(32'h3a8ebb01),
	.w2(32'hba27ac84),
	.w3(32'h3981277b),
	.w4(32'hba9c4253),
	.w5(32'h3abdc21d),
	.w6(32'hb9d9f418),
	.w7(32'hba88709d),
	.w8(32'h39a8355c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5e8a3),
	.w1(32'hbab533cc),
	.w2(32'h3997911a),
	.w3(32'h3b108e24),
	.w4(32'h3ae01203),
	.w5(32'h3a3ee977),
	.w6(32'hbaf36317),
	.w7(32'h38fd00e8),
	.w8(32'h3ac58983),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4afa76),
	.w1(32'hba5c73e7),
	.w2(32'hb9c675e2),
	.w3(32'hbaa80f19),
	.w4(32'h3aed16cd),
	.w5(32'hbac4a23d),
	.w6(32'h3b4ebfbe),
	.w7(32'hba1cd3f1),
	.w8(32'hbadde265),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0726ed),
	.w1(32'hb9e64e42),
	.w2(32'h3ab3450d),
	.w3(32'hba515a4b),
	.w4(32'h3a487733),
	.w5(32'hba8499c5),
	.w6(32'hbade8436),
	.w7(32'hb8c8eef5),
	.w8(32'h3a97c8ef),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac43529),
	.w1(32'h3ab6944c),
	.w2(32'h38933f93),
	.w3(32'hbb3fa405),
	.w4(32'hbb0da124),
	.w5(32'h39a204cd),
	.w6(32'h3a8331b5),
	.w7(32'h39b339fb),
	.w8(32'h3ab3b65d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a2da6),
	.w1(32'hb94bb71f),
	.w2(32'h390f0566),
	.w3(32'hbad14a74),
	.w4(32'hbaaa628a),
	.w5(32'hba3acbf1),
	.w6(32'hba3b5ae7),
	.w7(32'h3a0dfa0c),
	.w8(32'hbaebf101),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9abf6d),
	.w1(32'h3a7e51a1),
	.w2(32'h3a5ce856),
	.w3(32'hb95b9abc),
	.w4(32'hba950fee),
	.w5(32'h3b80d434),
	.w6(32'h39ddd2de),
	.w7(32'h3a4a8d68),
	.w8(32'h3ade665a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf73513),
	.w1(32'hba5f6b3f),
	.w2(32'h3a2bc56b),
	.w3(32'h3b44b59a),
	.w4(32'h3b5a5ea9),
	.w5(32'hba5ee36b),
	.w6(32'h3b116b71),
	.w7(32'hba3bf3c1),
	.w8(32'hbb9a12eb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5310dd),
	.w1(32'hbb11d267),
	.w2(32'h3a30f104),
	.w3(32'h3b1dca8c),
	.w4(32'h3a3ae878),
	.w5(32'h3b3ee631),
	.w6(32'h3aa2b9ae),
	.w7(32'h3b5d161e),
	.w8(32'hb95c1591),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a2d09),
	.w1(32'h3a095577),
	.w2(32'hb9ef91f1),
	.w3(32'h3b717c9b),
	.w4(32'h3b179735),
	.w5(32'hbb4c347c),
	.w6(32'hba2e8a9b),
	.w7(32'hbb0555d0),
	.w8(32'hbafada4d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae7738),
	.w1(32'hbb7b4cb4),
	.w2(32'hbb8e613b),
	.w3(32'hba9399e6),
	.w4(32'h3b316249),
	.w5(32'hb9bc6d12),
	.w6(32'h3aca252a),
	.w7(32'hb9c8975b),
	.w8(32'hba3ff82d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d09b5b),
	.w1(32'h3b1506f7),
	.w2(32'h3b34ad0a),
	.w3(32'hbab4619f),
	.w4(32'hbaaa54d5),
	.w5(32'hba4c1c84),
	.w6(32'hb8bc2de1),
	.w7(32'hbae42cf3),
	.w8(32'hba8c09db),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91bcbd8),
	.w1(32'hbb12af2d),
	.w2(32'hbafea4cf),
	.w3(32'h3995d463),
	.w4(32'hb9779814),
	.w5(32'hbb41bcb6),
	.w6(32'h3b10c8f8),
	.w7(32'h3a45dcef),
	.w8(32'hbb016dfa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cab7b),
	.w1(32'hba7932d3),
	.w2(32'hb949e1a8),
	.w3(32'hbb8b458c),
	.w4(32'hbb42e95a),
	.w5(32'h3b2ca0b4),
	.w6(32'hb9e83c68),
	.w7(32'hb9980795),
	.w8(32'hbb926e47),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcac5c),
	.w1(32'hbb39bfee),
	.w2(32'h3a208ccf),
	.w3(32'h3aa1c982),
	.w4(32'h3aea06e8),
	.w5(32'h3a71900a),
	.w6(32'hba9089a5),
	.w7(32'hbab5a31e),
	.w8(32'hba1e7964),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991f6d2),
	.w1(32'h3a102c65),
	.w2(32'hb9f2f25c),
	.w3(32'h3a58a077),
	.w4(32'hb99abf54),
	.w5(32'h3b176bc5),
	.w6(32'h3995259b),
	.w7(32'hb97c74cd),
	.w8(32'h3b6bef1f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ed60f),
	.w1(32'h3b6dafc0),
	.w2(32'h3b39529e),
	.w3(32'h3b03b432),
	.w4(32'h3ac997be),
	.w5(32'hbb8d1d5f),
	.w6(32'h3abbb0d2),
	.w7(32'h389574a2),
	.w8(32'hbb80f179),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06aeba),
	.w1(32'hbb76e351),
	.w2(32'hbac8dc1a),
	.w3(32'hbb167f65),
	.w4(32'hbb56dd57),
	.w5(32'h38a205b5),
	.w6(32'hbab22aa7),
	.w7(32'h3b0a8fee),
	.w8(32'hba182843),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16e9b2),
	.w1(32'hba3db8fc),
	.w2(32'h38f5c611),
	.w3(32'hb9a6306f),
	.w4(32'hbab47467),
	.w5(32'h390e8432),
	.w6(32'hb8a9ccee),
	.w7(32'h38761437),
	.w8(32'hbadd35f3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389714e1),
	.w1(32'hb9da72c7),
	.w2(32'hba21baa4),
	.w3(32'hba80bf80),
	.w4(32'h39cc9c85),
	.w5(32'hbad9e46d),
	.w6(32'hbb4f627f),
	.w7(32'hbb25dfb3),
	.w8(32'h3979a31d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94306f),
	.w1(32'h3a8b803c),
	.w2(32'hb9b52ba6),
	.w3(32'hbb4e74e9),
	.w4(32'hbb876329),
	.w5(32'h3aa84152),
	.w6(32'hbb4b447f),
	.w7(32'hbb455bf0),
	.w8(32'h3a8bea1c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897bdc3),
	.w1(32'h3a20aa4a),
	.w2(32'h39ff30bd),
	.w3(32'h3af40cf9),
	.w4(32'h39f325b9),
	.w5(32'hb91d799f),
	.w6(32'h3ad5631a),
	.w7(32'h3a92d353),
	.w8(32'hba00f66d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac394ec),
	.w1(32'hbaafb2bf),
	.w2(32'h376fa937),
	.w3(32'hb9d2e85c),
	.w4(32'hbaa4b62f),
	.w5(32'h3a1520c5),
	.w6(32'hb81223d3),
	.w7(32'h3a2b3094),
	.w8(32'h39a24b12),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b3c8e),
	.w1(32'h3a3f4ab0),
	.w2(32'h3a8c4722),
	.w3(32'h3a298174),
	.w4(32'hb9d6ff94),
	.w5(32'hba88f039),
	.w6(32'h3a028d30),
	.w7(32'h3a1dd25d),
	.w8(32'hbae0e0a8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacb651),
	.w1(32'h39f1509b),
	.w2(32'hb9c11052),
	.w3(32'hbacd94e2),
	.w4(32'hbb68ff7b),
	.w5(32'h3b4d6815),
	.w6(32'h3974bd8f),
	.w7(32'hba6aec83),
	.w8(32'h3a2dbd73),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38eb7d),
	.w1(32'hbb3a315a),
	.w2(32'hbb395b77),
	.w3(32'h3a73f8c7),
	.w4(32'h3a866c52),
	.w5(32'hbbc3dc56),
	.w6(32'h3a5e728f),
	.w7(32'h3adb5e0d),
	.w8(32'hbb0a8718),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398efa8d),
	.w1(32'h3a841db2),
	.w2(32'hbb021b76),
	.w3(32'hbb8cdd8d),
	.w4(32'hba1d8a18),
	.w5(32'h3b73db12),
	.w6(32'hbab9d007),
	.w7(32'hba15ae86),
	.w8(32'h3b4b463e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64186c),
	.w1(32'h3b0c69e6),
	.w2(32'h3affe14c),
	.w3(32'h3adb114f),
	.w4(32'h3a18b669),
	.w5(32'h3a836080),
	.w6(32'h38b1efaa),
	.w7(32'h39392bf7),
	.w8(32'h3b144960),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95890bc),
	.w1(32'h3a1c6ab5),
	.w2(32'h39511106),
	.w3(32'hbb19c5f1),
	.w4(32'hbae9faa5),
	.w5(32'hba156e9a),
	.w6(32'h3afd11bc),
	.w7(32'hb880d49a),
	.w8(32'h385f42c4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39454ea2),
	.w1(32'h3b4960c5),
	.w2(32'h3b3c96c0),
	.w3(32'hbb486361),
	.w4(32'hbb471c17),
	.w5(32'h387e7c84),
	.w6(32'h3a843150),
	.w7(32'hb92bc410),
	.w8(32'hb870e80b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96d9a0),
	.w1(32'h399dc600),
	.w2(32'hb9353d89),
	.w3(32'h393824ff),
	.w4(32'hbaa64942),
	.w5(32'hbb71875d),
	.w6(32'hb959c954),
	.w7(32'hb947d3e5),
	.w8(32'h364677bc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75e7f1),
	.w1(32'hbab69539),
	.w2(32'hbaaa0909),
	.w3(32'hbb559fe2),
	.w4(32'hbb3c11d6),
	.w5(32'hbaf55890),
	.w6(32'hba4c374e),
	.w7(32'hbb3cb17a),
	.w8(32'hbb525261),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe0d98),
	.w1(32'hba9a5021),
	.w2(32'hbb0ab963),
	.w3(32'hba595dfa),
	.w4(32'h3a15e6ae),
	.w5(32'hb996bdd5),
	.w6(32'h3abbf4dc),
	.w7(32'h38961858),
	.w8(32'hb96d804a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e7b3e),
	.w1(32'hba270f1e),
	.w2(32'hb98caffc),
	.w3(32'hbb3615e3),
	.w4(32'hbb6818e6),
	.w5(32'h3b0616c2),
	.w6(32'hba752a87),
	.w7(32'hbb5e8000),
	.w8(32'h3ad13bb6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b359100),
	.w1(32'h3a775bb0),
	.w2(32'h3b304a0c),
	.w3(32'h3b152668),
	.w4(32'h3b02a59b),
	.w5(32'h3a027762),
	.w6(32'hba274f83),
	.w7(32'h3ac27013),
	.w8(32'hba57353e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9da6ea),
	.w1(32'hb946de26),
	.w2(32'h3912b1a8),
	.w3(32'hba9c5d26),
	.w4(32'hb8a38a22),
	.w5(32'hbb7bde30),
	.w6(32'hbad3dca5),
	.w7(32'hbad602f2),
	.w8(32'h3afb4d13),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8651730),
	.w1(32'hba007cba),
	.w2(32'hbb90707c),
	.w3(32'hbbc7b133),
	.w4(32'hbb9a595a),
	.w5(32'hb9c8757a),
	.w6(32'hbaaa191c),
	.w7(32'hbb12b0e3),
	.w8(32'hbb1681ed),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eacdc),
	.w1(32'hbb1aa4d8),
	.w2(32'hbb972ddd),
	.w3(32'h3ab232fb),
	.w4(32'hba9d26d8),
	.w5(32'hb965d539),
	.w6(32'h3aac60a1),
	.w7(32'hbb017692),
	.w8(32'h3b04ea50),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73c315),
	.w1(32'h3b33e74c),
	.w2(32'h3ae1c8ca),
	.w3(32'hbb269d95),
	.w4(32'hbb5c2c4b),
	.w5(32'hb99884a2),
	.w6(32'h3b19fd69),
	.w7(32'hb982b108),
	.w8(32'h3b3b3d90),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b010de3),
	.w1(32'h3aa93d80),
	.w2(32'h37f2cd2f),
	.w3(32'hbae36126),
	.w4(32'h3a5d905e),
	.w5(32'hbb1b9c89),
	.w6(32'h3a07f7c2),
	.w7(32'h3a8d978f),
	.w8(32'hbb662e20),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922d2e),
	.w1(32'hbad33cb5),
	.w2(32'hb9c01f32),
	.w3(32'hbae4949b),
	.w4(32'hbb204f3a),
	.w5(32'hbac2b5a1),
	.w6(32'hb9d3eff8),
	.w7(32'h3a0403fa),
	.w8(32'hbadf715e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef31fb),
	.w1(32'hbadb90ed),
	.w2(32'hbb0b020e),
	.w3(32'h3a173c08),
	.w4(32'h3af685b8),
	.w5(32'hbab26d90),
	.w6(32'h3a6225f8),
	.w7(32'h3a15b43c),
	.w8(32'hbb5670d5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03f3cb),
	.w1(32'h3a0cd297),
	.w2(32'h3a9037cb),
	.w3(32'hb95e4057),
	.w4(32'hba86a7cf),
	.w5(32'hbb558d32),
	.w6(32'h3ad0d7f1),
	.w7(32'h3a49c3c8),
	.w8(32'hbb0530a4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989b9d7),
	.w1(32'hbb229376),
	.w2(32'hbb818f9c),
	.w3(32'hba10decc),
	.w4(32'hbace90cd),
	.w5(32'hba40932f),
	.w6(32'h390b8c23),
	.w7(32'hbb055723),
	.w8(32'h3a287adc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadcce9),
	.w1(32'h3aa130ba),
	.w2(32'hbb4a924c),
	.w3(32'hba3cbdab),
	.w4(32'hbb1337c8),
	.w5(32'hbb31abd1),
	.w6(32'hba8d7d4a),
	.w7(32'hbb574603),
	.w8(32'hbacc5384),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2898fe),
	.w1(32'h3a71190c),
	.w2(32'hba21f014),
	.w3(32'hbb01ed66),
	.w4(32'hbb7c8a90),
	.w5(32'hb9ac4d4c),
	.w6(32'hba6cd7d6),
	.w7(32'hbb28b872),
	.w8(32'hba99730c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf6bd8),
	.w1(32'h3a8f48b3),
	.w2(32'h3a09353b),
	.w3(32'hba03ee76),
	.w4(32'hba986ddb),
	.w5(32'h3a6484ad),
	.w6(32'h39919d26),
	.w7(32'hba26a21c),
	.w8(32'hbb149c26),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8524b),
	.w1(32'hbb3cfd14),
	.w2(32'hbb246367),
	.w3(32'h3b880a27),
	.w4(32'hb9e539bd),
	.w5(32'hbadc4a21),
	.w6(32'h3b816007),
	.w7(32'h3b40c840),
	.w8(32'hbb3cae56),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1336a),
	.w1(32'hba7449f8),
	.w2(32'hba301426),
	.w3(32'hbb59321c),
	.w4(32'hbb68b02b),
	.w5(32'hbaa7a1bf),
	.w6(32'hbb1ac510),
	.w7(32'hbadccc29),
	.w8(32'h3b1af362),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4603e),
	.w1(32'hbb1496c2),
	.w2(32'hbbb2b016),
	.w3(32'hba9548a5),
	.w4(32'hbac49b2c),
	.w5(32'h3ae24ed1),
	.w6(32'h3b8439e2),
	.w7(32'h3b023ce7),
	.w8(32'h3b83d00d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5c199),
	.w1(32'h3a3c7f6c),
	.w2(32'h3ad7a4d9),
	.w3(32'h3ab2cd1c),
	.w4(32'h3b33ab74),
	.w5(32'hba9ad319),
	.w6(32'h3b9329be),
	.w7(32'h3b44f198),
	.w8(32'hbb8a778e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb443edc),
	.w1(32'hbb855267),
	.w2(32'hbade2f2f),
	.w3(32'h3b40352e),
	.w4(32'h3abe6090),
	.w5(32'hbb67cd4c),
	.w6(32'hba283ee2),
	.w7(32'h3af1519c),
	.w8(32'hbb3b6d77),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf36f24),
	.w1(32'h3b2c78ad),
	.w2(32'h3b77ada0),
	.w3(32'hbac968f7),
	.w4(32'hba0f0b84),
	.w5(32'hbaa056b9),
	.w6(32'h385bba33),
	.w7(32'h3a90806e),
	.w8(32'hbb02a5f9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada3c26),
	.w1(32'hb96d1902),
	.w2(32'h393674e0),
	.w3(32'hba58566c),
	.w4(32'hbabaf059),
	.w5(32'hba942ae0),
	.w6(32'hbb86033f),
	.w7(32'hbb0a24cf),
	.w8(32'hba702d5e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa160e1),
	.w1(32'h3aa7d17d),
	.w2(32'hb7ffa179),
	.w3(32'hbb159c85),
	.w4(32'hbb2fb7e0),
	.w5(32'hb9bde158),
	.w6(32'hba809625),
	.w7(32'hba33abde),
	.w8(32'h3adad279),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9debbf0),
	.w1(32'hba9f5898),
	.w2(32'h3a699f25),
	.w3(32'hbacbec94),
	.w4(32'h37afd117),
	.w5(32'h3b28d8de),
	.w6(32'h3aa2c34e),
	.w7(32'h3a5bb8fd),
	.w8(32'hbb1969ce),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba849f24),
	.w1(32'hb76d49c6),
	.w2(32'h3b0352af),
	.w3(32'hbaba7404),
	.w4(32'hbb34f0e7),
	.w5(32'hbb05f729),
	.w6(32'hb8f57227),
	.w7(32'hba00664f),
	.w8(32'h3974a760),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdb832),
	.w1(32'hb9f50754),
	.w2(32'hba581d73),
	.w3(32'hbb1869fd),
	.w4(32'hbb878454),
	.w5(32'hb9857bea),
	.w6(32'hbaa9415f),
	.w7(32'hbaa732db),
	.w8(32'hb7cfd57b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cbf4f),
	.w1(32'h3b0edd6a),
	.w2(32'h3b0d0f44),
	.w3(32'hba3a96cc),
	.w4(32'h391a645f),
	.w5(32'h3aa2beaa),
	.w6(32'h39673131),
	.w7(32'hba670bd0),
	.w8(32'h3ac2eeb3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab50879),
	.w1(32'h3b05dc3e),
	.w2(32'hb9d5e1ae),
	.w3(32'hbb0effee),
	.w4(32'hbb0a6d90),
	.w5(32'h3b877eea),
	.w6(32'h389dba59),
	.w7(32'hbb4dedc4),
	.w8(32'h3b416b37),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cde015),
	.w1(32'h39f5a78d),
	.w2(32'h3b14a8fd),
	.w3(32'h3ba3be73),
	.w4(32'h3b9d676c),
	.w5(32'h3abfb086),
	.w6(32'h3b4eabf7),
	.w7(32'h3b9a7dbf),
	.w8(32'h3a56de0a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfc0ee),
	.w1(32'hbaac6aec),
	.w2(32'hbaf6e85c),
	.w3(32'h3b0ef666),
	.w4(32'h3b074154),
	.w5(32'h3acb0e1d),
	.w6(32'h3a356c43),
	.w7(32'h3a9e5989),
	.w8(32'h3b1206a2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a80c8),
	.w1(32'h3a819ab7),
	.w2(32'h3b109e44),
	.w3(32'h3a4d8d91),
	.w4(32'h3aa5cecf),
	.w5(32'hbba922ee),
	.w6(32'hb9c3480d),
	.w7(32'h3ac8d9df),
	.w8(32'hbba95c5d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b96b3),
	.w1(32'hba101d2e),
	.w2(32'hba4500a3),
	.w3(32'hbad5187e),
	.w4(32'hbb7ba159),
	.w5(32'h3aa00e67),
	.w6(32'hba6c5b6f),
	.w7(32'hbb4e5eef),
	.w8(32'h3a1658f9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01eb8c),
	.w1(32'h39c74566),
	.w2(32'h3a73d786),
	.w3(32'h39e72440),
	.w4(32'h399351ee),
	.w5(32'hb8d72a33),
	.w6(32'h3910c96b),
	.w7(32'h3910bd21),
	.w8(32'hb88de9f9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa73e92),
	.w1(32'h39d9bd98),
	.w2(32'hba44772d),
	.w3(32'hbb193b42),
	.w4(32'hbae46827),
	.w5(32'hbb607375),
	.w6(32'hba8b30c1),
	.w7(32'hbb215940),
	.w8(32'hbb3d9c18),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d1715),
	.w1(32'h3b0c7584),
	.w2(32'h3b0bd0c6),
	.w3(32'hba25066a),
	.w4(32'h39909b05),
	.w5(32'h39c495ca),
	.w6(32'h3934da48),
	.w7(32'h3b0c09b9),
	.w8(32'hbb1716f1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa607f),
	.w1(32'hbb1c7960),
	.w2(32'hbaf51dc2),
	.w3(32'h3a9ba33f),
	.w4(32'hb8991de0),
	.w5(32'hbb5ea66c),
	.w6(32'h3aeb6270),
	.w7(32'h3ae65b70),
	.w8(32'hbb53bb0f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7881d2),
	.w1(32'hbade0fc1),
	.w2(32'hbb59fb4d),
	.w3(32'hba776ba7),
	.w4(32'hbb622c80),
	.w5(32'hbab9670c),
	.w6(32'h38c70832),
	.w7(32'hb8d81ac4),
	.w8(32'hba54b45c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924e866),
	.w1(32'h391b4488),
	.w2(32'h39c6bb9d),
	.w3(32'h3a879827),
	.w4(32'hb8fc3af3),
	.w5(32'h3a2bd700),
	.w6(32'hb774912b),
	.w7(32'h3b035360),
	.w8(32'hb992b389),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a960912),
	.w1(32'h3a8ccc56),
	.w2(32'hb9897369),
	.w3(32'h3a5085f9),
	.w4(32'h3b25908f),
	.w5(32'h3a2775ed),
	.w6(32'h3aa79ce0),
	.w7(32'h3b12f317),
	.w8(32'h3ac07eb7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b096940),
	.w1(32'h3a64cdc7),
	.w2(32'h3a9fe32a),
	.w3(32'hb989b99f),
	.w4(32'h3a01d627),
	.w5(32'h3b8cde46),
	.w6(32'hba0b9857),
	.w7(32'h3a8fe7af),
	.w8(32'h3b9270f8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdf45f),
	.w1(32'hbb986674),
	.w2(32'hbb775754),
	.w3(32'h3bd8abeb),
	.w4(32'h3b734dcb),
	.w5(32'hbae941c6),
	.w6(32'h3b67e779),
	.w7(32'hba6ba942),
	.w8(32'hbb1cda83),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3929021b),
	.w1(32'hbad903a8),
	.w2(32'hba55e2d4),
	.w3(32'h3abb2768),
	.w4(32'h3af9ef8f),
	.w5(32'h3a9a1eed),
	.w6(32'hba91f3ef),
	.w7(32'h3ac5dbb9),
	.w8(32'h3a81a1dc),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92811f),
	.w1(32'h3b263428),
	.w2(32'h3ad4c86f),
	.w3(32'hbb15acc3),
	.w4(32'hbb379d51),
	.w5(32'hbac60cc0),
	.w6(32'h3a98f894),
	.w7(32'hbaa9d3ef),
	.w8(32'hbb2a2496),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bd483),
	.w1(32'hbb56df45),
	.w2(32'hba8972a1),
	.w3(32'h3a343944),
	.w4(32'hbb0848ad),
	.w5(32'h390723d1),
	.w6(32'h3b921487),
	.w7(32'h3b76c7f6),
	.w8(32'hba982b5a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e0c07),
	.w1(32'h3a8ce420),
	.w2(32'h3b23bc76),
	.w3(32'h3ab05d6e),
	.w4(32'hb7ddfb01),
	.w5(32'h3b3b741a),
	.w6(32'h3add4898),
	.w7(32'h3b60ef30),
	.w8(32'hb814ff28),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43058d),
	.w1(32'hbb4cd30f),
	.w2(32'hbb1b36be),
	.w3(32'h3af923b3),
	.w4(32'hbb46378f),
	.w5(32'h3a4ab8d0),
	.w6(32'h3b41cbd8),
	.w7(32'h3abbda8b),
	.w8(32'hbb27cd56),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bf8d3),
	.w1(32'hbb863df3),
	.w2(32'hbb03676b),
	.w3(32'h3acf5128),
	.w4(32'hbabe1773),
	.w5(32'hbaf0e767),
	.w6(32'h3b1ca9c0),
	.w7(32'hb9d1feb6),
	.w8(32'hbadeab04),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a024e15),
	.w1(32'h3aae68fa),
	.w2(32'h3a6f5a51),
	.w3(32'h39030adb),
	.w4(32'hbaf3921e),
	.w5(32'h3be16c00),
	.w6(32'h395d1759),
	.w7(32'hba4984af),
	.w8(32'h3b460a19),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db278),
	.w1(32'h3991388a),
	.w2(32'h3b00ce4d),
	.w3(32'h3bfc5ba9),
	.w4(32'h3bbcc363),
	.w5(32'hbb568183),
	.w6(32'h3bb296db),
	.w7(32'h3bd75747),
	.w8(32'hbb831929),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99535b),
	.w1(32'hba53d4bf),
	.w2(32'hbb13c306),
	.w3(32'hbb012e58),
	.w4(32'hbb4c0cec),
	.w5(32'h3ae4e2b2),
	.w6(32'hbb154423),
	.w7(32'hbab4078a),
	.w8(32'h39e0784e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b371021),
	.w1(32'h3adcdf0d),
	.w2(32'h39fa090f),
	.w3(32'hbac90330),
	.w4(32'hbb0a6019),
	.w5(32'hba56c0a9),
	.w6(32'hbb304baa),
	.w7(32'hba9d2f4e),
	.w8(32'h3b374fd2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b020645),
	.w1(32'h3b21faca),
	.w2(32'h3aa120f1),
	.w3(32'hba3606f5),
	.w4(32'h3a450ea2),
	.w5(32'hba5d0749),
	.w6(32'h3b14a84f),
	.w7(32'h3a6fbf8d),
	.w8(32'h387d038c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a177ade),
	.w1(32'h3ad2af83),
	.w2(32'h3a42e374),
	.w3(32'hbafc5cca),
	.w4(32'hb9f7ec63),
	.w5(32'h370a273a),
	.w6(32'hb9c88115),
	.w7(32'hba8dcef1),
	.w8(32'hba850bc3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb486335),
	.w1(32'hbb7f24c8),
	.w2(32'hbb20df7f),
	.w3(32'h3a95ce2a),
	.w4(32'h3ae8ff80),
	.w5(32'h3a9caa2d),
	.w6(32'h3b724265),
	.w7(32'h3bc8dc7b),
	.w8(32'hbaacf4f1),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb183863),
	.w1(32'hba946a8e),
	.w2(32'h3a1bbd14),
	.w3(32'h39add317),
	.w4(32'h37e45e8d),
	.w5(32'h397d677d),
	.w6(32'h3ade74fe),
	.w7(32'h3aabf4bc),
	.w8(32'hba55ba11),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa27de2),
	.w1(32'h3a1314b8),
	.w2(32'h3acc0112),
	.w3(32'h3a47668d),
	.w4(32'hbab3c070),
	.w5(32'h3a45c5be),
	.w6(32'h3b07db0b),
	.w7(32'h3ae0d012),
	.w8(32'hbad98d74),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ff2a),
	.w1(32'hbb378421),
	.w2(32'hbb3efb39),
	.w3(32'h3b086922),
	.w4(32'h3b081d28),
	.w5(32'hba739355),
	.w6(32'hb9caefef),
	.w7(32'hba59fd6d),
	.w8(32'hba81bd37),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef5f86),
	.w1(32'h3a133c78),
	.w2(32'h3a465638),
	.w3(32'hba68163d),
	.w4(32'hbac3d93f),
	.w5(32'hba84f3e2),
	.w6(32'hbb427c44),
	.w7(32'hbb65a92a),
	.w8(32'hbb2a29d3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d83b1),
	.w1(32'hb8549509),
	.w2(32'hbaad9bf3),
	.w3(32'hbb1714af),
	.w4(32'hbad81695),
	.w5(32'h39ce6f6b),
	.w6(32'hbad0a972),
	.w7(32'hbb042c1f),
	.w8(32'h3b077663),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89c346),
	.w1(32'h39bc3c40),
	.w2(32'hb9e1a07a),
	.w3(32'hb9828402),
	.w4(32'hba698a37),
	.w5(32'hb900c326),
	.w6(32'h39ea4114),
	.w7(32'hba5e4d83),
	.w8(32'hba84e09e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12d3a7),
	.w1(32'h3af7460a),
	.w2(32'h3ab8c551),
	.w3(32'h39870e1c),
	.w4(32'hb9e17dd5),
	.w5(32'hbb6e7bda),
	.w6(32'hb98b13e1),
	.w7(32'h39f01578),
	.w8(32'h38a8223e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bf1711),
	.w1(32'h3a0caa38),
	.w2(32'h39ce5674),
	.w3(32'hbb2cdd3b),
	.w4(32'hbac7581f),
	.w5(32'hba99bfb9),
	.w6(32'hbab4797f),
	.w7(32'h38c89d10),
	.w8(32'hba22d1e2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a360464),
	.w1(32'hba177305),
	.w2(32'hbae748d1),
	.w3(32'hba9ac46c),
	.w4(32'hbacaec02),
	.w5(32'h3a2d033b),
	.w6(32'hba631c76),
	.w7(32'hbaad6773),
	.w8(32'hb9292226),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82746c),
	.w1(32'h39c43209),
	.w2(32'h39c3f953),
	.w3(32'hbaa88ced),
	.w4(32'hba9c3d96),
	.w5(32'h3badf2cc),
	.w6(32'hbadb0b9a),
	.w7(32'hba800c3c),
	.w8(32'h3bab8225),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a885c22),
	.w1(32'h3b41a985),
	.w2(32'h3b26b747),
	.w3(32'h3bce7e92),
	.w4(32'h3be10505),
	.w5(32'h3aa2909e),
	.w6(32'h3bbdec69),
	.w7(32'h3bb94e02),
	.w8(32'h361a788c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0dfb9),
	.w1(32'hbacb8ed2),
	.w2(32'hbab9a09f),
	.w3(32'h38c357f6),
	.w4(32'h3ab4c3f1),
	.w5(32'hba31c937),
	.w6(32'hba7d7819),
	.w7(32'hbab30673),
	.w8(32'hbabd0cb7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a621fb8),
	.w1(32'h3b03af31),
	.w2(32'h3a6726c3),
	.w3(32'hbad9bafb),
	.w4(32'hbb2a1eb4),
	.w5(32'hbb57a9f4),
	.w6(32'h38ca9e25),
	.w7(32'hba9ca14a),
	.w8(32'hba549ba1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21c107),
	.w1(32'h3b7511c2),
	.w2(32'h3a4e8b72),
	.w3(32'hbbc0f83e),
	.w4(32'hbb3d2892),
	.w5(32'hba3995d7),
	.w6(32'hbb45da1b),
	.w7(32'hbb306673),
	.w8(32'hbb2133a5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a439700),
	.w1(32'hbb243a0c),
	.w2(32'hbae11432),
	.w3(32'h39d612ef),
	.w4(32'h3ac23df9),
	.w5(32'h39ececf0),
	.w6(32'h3a40f15e),
	.w7(32'hb9a493e1),
	.w8(32'hb9e65b5c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40e32e),
	.w1(32'hb98ee531),
	.w2(32'hb98b00a5),
	.w3(32'hbaa3b9ee),
	.w4(32'hb9b6701e),
	.w5(32'hbb6cf55e),
	.w6(32'hbb12d425),
	.w7(32'hbb0ef1f3),
	.w8(32'hbb1c5342),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3de6fa),
	.w1(32'h3a7ebf79),
	.w2(32'h3a9a1a13),
	.w3(32'hbb4a99fc),
	.w4(32'hbab378a6),
	.w5(32'hbb5beb16),
	.w6(32'hbac5cbdf),
	.w7(32'hba2fd9ba),
	.w8(32'hbb76a3b0),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82a6af),
	.w1(32'hbabdb75f),
	.w2(32'hb9e43c96),
	.w3(32'hbb0d71a6),
	.w4(32'hbaf268ce),
	.w5(32'hba5ec1f8),
	.w6(32'hbb3dd376),
	.w7(32'hb9e43eda),
	.w8(32'hba0a444e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2794de),
	.w1(32'h3993a637),
	.w2(32'hb98361c8),
	.w3(32'h39c2c18f),
	.w4(32'hba476669),
	.w5(32'hbb1752ff),
	.w6(32'h37e1cde1),
	.w7(32'h380be04b),
	.w8(32'h3b17c3b5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13a8c3),
	.w1(32'h3ba3f91b),
	.w2(32'h39fd7830),
	.w3(32'hbb468b0a),
	.w4(32'hba5dad03),
	.w5(32'h379a3dd2),
	.w6(32'hb785a4f1),
	.w7(32'hbb68f3ae),
	.w8(32'h391bd778),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a2459),
	.w1(32'h3a3cff08),
	.w2(32'h3b2e2e12),
	.w3(32'h3ac82265),
	.w4(32'h3ad1e95e),
	.w5(32'hba3c5e14),
	.w6(32'hb9f37b37),
	.w7(32'h3ae4ea87),
	.w8(32'h3abd76ec),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba375151),
	.w1(32'h38a052b7),
	.w2(32'h3a537b38),
	.w3(32'hbb07ba4c),
	.w4(32'hba8ec194),
	.w5(32'h3b5c3c5c),
	.w6(32'h3a68f421),
	.w7(32'h3ad22744),
	.w8(32'h3b729c20),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b149d92),
	.w1(32'h3abfcb05),
	.w2(32'h3a6589d1),
	.w3(32'h3b577c28),
	.w4(32'h3ae0ab94),
	.w5(32'h391e3a0a),
	.w6(32'h3af9c699),
	.w7(32'h3b6d3558),
	.w8(32'hb982c6be),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfd021),
	.w1(32'hbbbcf17a),
	.w2(32'hbaa8c593),
	.w3(32'h3afb28f7),
	.w4(32'h380f5dc0),
	.w5(32'hbb97a191),
	.w6(32'h3a3da3d8),
	.w7(32'hb9fb6779),
	.w8(32'hbaab3253),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab0405),
	.w1(32'h3990d39c),
	.w2(32'hbab3944d),
	.w3(32'hba622b00),
	.w4(32'hbb6a386a),
	.w5(32'h3a7be954),
	.w6(32'hbb1cb861),
	.w7(32'hbb714658),
	.w8(32'h3a47a9ef),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a04a79),
	.w1(32'hba9b3331),
	.w2(32'hba2edda8),
	.w3(32'hb9faedc3),
	.w4(32'hb960f195),
	.w5(32'hbb269fdc),
	.w6(32'hba1e8c30),
	.w7(32'hb9d4d47a),
	.w8(32'hbb0afba6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1efe2),
	.w1(32'hbb43d100),
	.w2(32'hbb09283c),
	.w3(32'hbb272581),
	.w4(32'hbaf30d19),
	.w5(32'h3aec71e6),
	.w6(32'hbb575ae8),
	.w7(32'hbb3496ca),
	.w8(32'h3ba0cf03),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b726bce),
	.w1(32'h3ba97c3a),
	.w2(32'h3be082a6),
	.w3(32'h3a84b5a3),
	.w4(32'h3af0e948),
	.w5(32'hb8dc1121),
	.w6(32'h3b866a73),
	.w7(32'h3b98c99d),
	.w8(32'h3a070b1a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7fbf7),
	.w1(32'h3b30a99f),
	.w2(32'h3b2f2148),
	.w3(32'h391bb352),
	.w4(32'h390830f5),
	.w5(32'hbaabbae2),
	.w6(32'hba8993a8),
	.w7(32'hb9b4d810),
	.w8(32'hb9da207f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a7591),
	.w1(32'hba5fe2a1),
	.w2(32'hb9894084),
	.w3(32'hbacfd6bc),
	.w4(32'hba3aa3ea),
	.w5(32'hbb85fe28),
	.w6(32'hba7990b6),
	.w7(32'hba4d56b2),
	.w8(32'hbb82bffa),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb741480),
	.w1(32'hbbaa197a),
	.w2(32'hbba138dc),
	.w3(32'hbba8d09e),
	.w4(32'hbb970b0c),
	.w5(32'h3b46f7c3),
	.w6(32'hbba9578e),
	.w7(32'hbba4b6b0),
	.w8(32'h3b977c2e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87a105),
	.w1(32'h3ba5847d),
	.w2(32'h3b7f5778),
	.w3(32'h3b5bb91a),
	.w4(32'h3b1205fe),
	.w5(32'hbb16b826),
	.w6(32'h3b59cc42),
	.w7(32'h3b80c3e6),
	.w8(32'hbb108c78),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21ebf3),
	.w1(32'hbb541540),
	.w2(32'hbb21a85b),
	.w3(32'hbb3df220),
	.w4(32'hbb28627d),
	.w5(32'hb9e9a8d9),
	.w6(32'hbb3a8678),
	.w7(32'hbb2b1eac),
	.w8(32'hb80a34bb),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a251675),
	.w1(32'hba1d7929),
	.w2(32'hbad74407),
	.w3(32'hbaf09ba6),
	.w4(32'h37b17376),
	.w5(32'hbb01e647),
	.w6(32'hbac517da),
	.w7(32'hba4322c5),
	.w8(32'hba966cad),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae216d0),
	.w1(32'hba996ab1),
	.w2(32'hba4e8356),
	.w3(32'hbac88d44),
	.w4(32'hbabe2818),
	.w5(32'hb930e0a5),
	.w6(32'h3a33ed57),
	.w7(32'h39f26aef),
	.w8(32'hba9b127d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf15891),
	.w1(32'hbb422da4),
	.w2(32'hbad68b11),
	.w3(32'hba6f275e),
	.w4(32'h38405284),
	.w5(32'hbb167807),
	.w6(32'hbb12d563),
	.w7(32'hba64a8e6),
	.w8(32'hbae218cb),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf091d7),
	.w1(32'hba4ca9cd),
	.w2(32'h3956e1ca),
	.w3(32'hbaad4673),
	.w4(32'hbab60b25),
	.w5(32'hbb3fc538),
	.w6(32'hb9683058),
	.w7(32'h3a342a45),
	.w8(32'h39f5e1ca),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b244ecc),
	.w1(32'h3af054a6),
	.w2(32'hbab9dc07),
	.w3(32'hba184f0e),
	.w4(32'hb868f100),
	.w5(32'hbb03857b),
	.w6(32'h3a3f6118),
	.w7(32'h37f58ea0),
	.w8(32'hba7a3382),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9158c3),
	.w1(32'hbb2b7494),
	.w2(32'hbad513ac),
	.w3(32'hbb058869),
	.w4(32'hbb4f308a),
	.w5(32'h3b01c0bc),
	.w6(32'hbb0ea7b5),
	.w7(32'hbb192ddb),
	.w8(32'h3a6e512c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3eaf2),
	.w1(32'h39dab881),
	.w2(32'h3aa912ca),
	.w3(32'h3ab8c269),
	.w4(32'h3b2a39e7),
	.w5(32'h39642a92),
	.w6(32'h398792c7),
	.w7(32'h3aae89c0),
	.w8(32'h3a36100f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90c7d2),
	.w1(32'h391642bc),
	.w2(32'h39b033b8),
	.w3(32'h39f4deef),
	.w4(32'h3a53760a),
	.w5(32'h3a1c97f9),
	.w6(32'h3a8d22dc),
	.w7(32'hb7264319),
	.w8(32'hbad828a7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0295ca),
	.w1(32'hbabf7724),
	.w2(32'h3a98bc83),
	.w3(32'hbb45f3c4),
	.w4(32'hbb3a8350),
	.w5(32'hbb11d1e0),
	.w6(32'hba371b9a),
	.w7(32'hbadc7a75),
	.w8(32'hba2663a2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a222c77),
	.w1(32'hbab0a38d),
	.w2(32'hba1463b0),
	.w3(32'hbb11aad6),
	.w4(32'hbb05ce19),
	.w5(32'h3ba46786),
	.w6(32'hbb1ef483),
	.w7(32'hbabdeb09),
	.w8(32'h3b99b82f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9699fc),
	.w1(32'h3b873ab0),
	.w2(32'h3b8774c4),
	.w3(32'h3b5a054a),
	.w4(32'h3b4b044b),
	.w5(32'hbafb4360),
	.w6(32'h3b90d68f),
	.w7(32'h3b742596),
	.w8(32'hba92fb94),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a354c6),
	.w1(32'h3a7b8256),
	.w2(32'h3ac50c2e),
	.w3(32'hbaab8fac),
	.w4(32'hbb4e8593),
	.w5(32'h3a779da2),
	.w6(32'hbabadff6),
	.w7(32'h38e02d43),
	.w8(32'h3a7ffcc2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b8d6a),
	.w1(32'hba40159a),
	.w2(32'hb9799583),
	.w3(32'hba273a12),
	.w4(32'hba03a3d8),
	.w5(32'hba5f6c0f),
	.w6(32'hba51d0d4),
	.w7(32'hba9d6dfe),
	.w8(32'hba75c542),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba4ef3),
	.w1(32'hbb346382),
	.w2(32'hbad35c41),
	.w3(32'hbb0e1aa7),
	.w4(32'hb9a42f8b),
	.w5(32'hbac97d5c),
	.w6(32'hbaeae793),
	.w7(32'hba201795),
	.w8(32'hbae6e48f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e690d),
	.w1(32'hbad32e06),
	.w2(32'hbae504a2),
	.w3(32'hba666700),
	.w4(32'hba5765f1),
	.w5(32'h3966b6ee),
	.w6(32'hba60c0f0),
	.w7(32'hbabb98c3),
	.w8(32'hb985c10a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ba9e2),
	.w1(32'hba9d4f61),
	.w2(32'hbb108c08),
	.w3(32'hba9410b1),
	.w4(32'hba88dbe4),
	.w5(32'hbb888399),
	.w6(32'hbaf337b2),
	.w7(32'hbb072358),
	.w8(32'hbafc5282),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16189e),
	.w1(32'hb9e593ae),
	.w2(32'h39beb251),
	.w3(32'hbb4250f4),
	.w4(32'hbb310af9),
	.w5(32'hbae14268),
	.w6(32'hbaa650c7),
	.w7(32'hbb091a44),
	.w8(32'hbb659793),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860d7c),
	.w1(32'hbb8db6b4),
	.w2(32'hbba26c9a),
	.w3(32'hbb26e5a2),
	.w4(32'hbb13bb50),
	.w5(32'hbb2a9ff6),
	.w6(32'hbb76afb0),
	.w7(32'hbb63e9eb),
	.w8(32'hbb0ddf39),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ad290c),
	.w1(32'h3ad0bdd1),
	.w2(32'h3940cb48),
	.w3(32'hbab01b79),
	.w4(32'hbac680cf),
	.w5(32'h3a8573e8),
	.w6(32'hbaa72b2f),
	.w7(32'hbaaeae1c),
	.w8(32'h3a3bd954),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ef4af),
	.w1(32'h3a7790ee),
	.w2(32'h39f772ef),
	.w3(32'h3a8e64cc),
	.w4(32'h39bd014e),
	.w5(32'h3b06c928),
	.w6(32'h3a47c2f0),
	.w7(32'hb7b55801),
	.w8(32'h3b1e8a2c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6e40c),
	.w1(32'h3b08e197),
	.w2(32'h3b233762),
	.w3(32'h3add32b4),
	.w4(32'h3a5042ef),
	.w5(32'hb9cc33c0),
	.w6(32'h3b47c478),
	.w7(32'h3b10a386),
	.w8(32'hba443c65),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebbcd1),
	.w1(32'hba6d58bc),
	.w2(32'h3a5fbb97),
	.w3(32'hb9900de1),
	.w4(32'h3a1b11f7),
	.w5(32'hba9fc8e5),
	.w6(32'hb92c3826),
	.w7(32'h3906b5b7),
	.w8(32'h3a300afb),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule