module layer_8_featuremap_246(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb57c4),
	.w1(32'h3af5289c),
	.w2(32'hbc13b894),
	.w3(32'h3ca9e1a7),
	.w4(32'hb9d1d5d8),
	.w5(32'hbbe980c5),
	.w6(32'hbb2d6055),
	.w7(32'hbb2cd6af),
	.w8(32'hbb7fcb5e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac68759),
	.w1(32'h3c094bfe),
	.w2(32'hbb2a0231),
	.w3(32'hbbd08683),
	.w4(32'h3bc0df26),
	.w5(32'hbb9807f2),
	.w6(32'h3b53f053),
	.w7(32'hba854635),
	.w8(32'hbbb2ef96),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cd07b),
	.w1(32'h3ab241d4),
	.w2(32'h3a9d1181),
	.w3(32'hbc8c50f0),
	.w4(32'h3b354771),
	.w5(32'h3a8de9ec),
	.w6(32'hbbafee5f),
	.w7(32'h3988a8e9),
	.w8(32'h3b2c9732),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a557b1c),
	.w1(32'hbc0aa9eb),
	.w2(32'hbbd93077),
	.w3(32'hbb523550),
	.w4(32'hbbe06e2b),
	.w5(32'hbc006947),
	.w6(32'hbb42ae66),
	.w7(32'h3a38a758),
	.w8(32'hba24fda1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec8480),
	.w1(32'hbb38cce6),
	.w2(32'hba0070a8),
	.w3(32'hbaddd6e9),
	.w4(32'hba9fffcb),
	.w5(32'hbad9b0ea),
	.w6(32'hbb502c8d),
	.w7(32'h39f97558),
	.w8(32'hb9c06875),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65abe7),
	.w1(32'hba8fb183),
	.w2(32'hbb552b41),
	.w3(32'hbb5ac833),
	.w4(32'h3bca492f),
	.w5(32'hbbb35af7),
	.w6(32'hbbd30a82),
	.w7(32'h3b5007dc),
	.w8(32'h3b4dbd89),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba729f6),
	.w1(32'hbc2f6626),
	.w2(32'h3b5d0668),
	.w3(32'hba5c078c),
	.w4(32'hbc1353ad),
	.w5(32'h3b98c569),
	.w6(32'hbc3b7984),
	.w7(32'hbb597e8c),
	.w8(32'h3b8d35ad),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77d9ad),
	.w1(32'hbc1d42f9),
	.w2(32'hbc0309ff),
	.w3(32'h3b968906),
	.w4(32'hbc1e4f1b),
	.w5(32'hbbfb02d3),
	.w6(32'hbc4dbae5),
	.w7(32'hba87b17e),
	.w8(32'h39e568e1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1e2c6),
	.w1(32'hbc399eea),
	.w2(32'h3b898694),
	.w3(32'hbc590a67),
	.w4(32'hbc54e4de),
	.w5(32'h3b89a91e),
	.w6(32'hbcb79a76),
	.w7(32'hbc244923),
	.w8(32'hbad76c69),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fe801),
	.w1(32'hbc13e553),
	.w2(32'hbc62b1c7),
	.w3(32'h3c06f695),
	.w4(32'hbbe53140),
	.w5(32'hbc1ffad8),
	.w6(32'h3a37f4eb),
	.w7(32'hbc03f986),
	.w8(32'hbbf3d598),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca1250),
	.w1(32'hbac30d14),
	.w2(32'hbc057ae5),
	.w3(32'h3b8d075d),
	.w4(32'h3a250093),
	.w5(32'hbbcc95e2),
	.w6(32'h395dcc1b),
	.w7(32'hbb64dd7c),
	.w8(32'hb7705054),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a7c97),
	.w1(32'hba8e3a3c),
	.w2(32'hbc11ba3a),
	.w3(32'hb9e6479f),
	.w4(32'hbbb7bbe3),
	.w5(32'hbc0bccfa),
	.w6(32'h3b862236),
	.w7(32'h3b3bf7f9),
	.w8(32'hba75c87c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2557c),
	.w1(32'hbb656001),
	.w2(32'hbb2c17e3),
	.w3(32'hbb9a34a5),
	.w4(32'hbc3464f5),
	.w5(32'hbb2104e6),
	.w6(32'hbc0ef891),
	.w7(32'hbbebceaf),
	.w8(32'hbad99e57),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf472b),
	.w1(32'h398464e1),
	.w2(32'hba8435a8),
	.w3(32'h3aea95f4),
	.w4(32'hba9d9700),
	.w5(32'h395da509),
	.w6(32'h3a5c7b98),
	.w7(32'h38861326),
	.w8(32'h3b4690f4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49783b),
	.w1(32'h3bc6b206),
	.w2(32'hbc3456dd),
	.w3(32'hbb5f6bdd),
	.w4(32'h3b2a5161),
	.w5(32'hbc314f4e),
	.w6(32'h3bb77dcd),
	.w7(32'hbb8aa1ad),
	.w8(32'hbc5848da),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab7d97),
	.w1(32'h3b887e7e),
	.w2(32'h3bd9d3b2),
	.w3(32'hbca4fb66),
	.w4(32'h3b69f26e),
	.w5(32'h3b590894),
	.w6(32'hbaf6ba03),
	.w7(32'hbb4b187c),
	.w8(32'h3ba2414e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14602a),
	.w1(32'h3b8ce29a),
	.w2(32'h3b77f78c),
	.w3(32'h3be7b567),
	.w4(32'h3bebd8d7),
	.w5(32'h3b7f8531),
	.w6(32'h3ac32e1c),
	.w7(32'h3a7c3f00),
	.w8(32'h3ac7211b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a4683),
	.w1(32'hb9826018),
	.w2(32'hba8efd2f),
	.w3(32'hba3fd415),
	.w4(32'hbbed2d57),
	.w5(32'hbac83a99),
	.w6(32'hbafb5d20),
	.w7(32'h3b1fdff5),
	.w8(32'h3ae58a38),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccfabf1),
	.w1(32'hbc80d5e8),
	.w2(32'hbcf1454a),
	.w3(32'h3b53b09f),
	.w4(32'hbbdf0154),
	.w5(32'hbc9f9d5c),
	.w6(32'h3c6ce346),
	.w7(32'hbb60f3ca),
	.w8(32'hbc613531),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d9938),
	.w1(32'hbcd567cc),
	.w2(32'hbc82bebc),
	.w3(32'hba2fab90),
	.w4(32'hbc949181),
	.w5(32'hbc2709f5),
	.w6(32'hbc8548df),
	.w7(32'hbc12d3fc),
	.w8(32'hbbc5603d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b148f35),
	.w1(32'hb8949584),
	.w2(32'hb8ac5c93),
	.w3(32'h3c4a78c4),
	.w4(32'h3c0337d7),
	.w5(32'h3bacc44d),
	.w6(32'h3c11817b),
	.w7(32'h3c765fb5),
	.w8(32'h3b014de2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddb75a),
	.w1(32'hbb6766a2),
	.w2(32'hba283fd0),
	.w3(32'hbbc63a1f),
	.w4(32'hbc1b106b),
	.w5(32'h3b58e5aa),
	.w6(32'hbba755cc),
	.w7(32'hbbefeee6),
	.w8(32'h39d51cff),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5f8c1),
	.w1(32'hbbbc8b04),
	.w2(32'hbcfa6142),
	.w3(32'h3c613e4a),
	.w4(32'hbb9e64b7),
	.w5(32'hbc764be7),
	.w6(32'h3c7de16c),
	.w7(32'hbc56ba91),
	.w8(32'hbc8e15bd),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084428),
	.w1(32'hbb390571),
	.w2(32'h3b86a220),
	.w3(32'h3bc08a83),
	.w4(32'h3ba6bcbc),
	.w5(32'h3b562662),
	.w6(32'h3c186c16),
	.w7(32'h3c38828b),
	.w8(32'h3c1810e2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3a5f6),
	.w1(32'h38746914),
	.w2(32'h3adecd4b),
	.w3(32'h3c03c145),
	.w4(32'hbb30a88f),
	.w5(32'h3b17af2a),
	.w6(32'hbb2ed1f5),
	.w7(32'hba7f29eb),
	.w8(32'h394e0840),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b4398),
	.w1(32'h3b9a1266),
	.w2(32'hbc0e8c26),
	.w3(32'h3bb6b2f6),
	.w4(32'h3addb648),
	.w5(32'hbaa20ae2),
	.w6(32'h3b3682cc),
	.w7(32'h3af92ef8),
	.w8(32'hbb71e4b2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12d196),
	.w1(32'hbaf6daa8),
	.w2(32'h3a2606cd),
	.w3(32'hb90896a0),
	.w4(32'h3a47d161),
	.w5(32'h3b0b493b),
	.w6(32'hbb908e73),
	.w7(32'h3b3f4645),
	.w8(32'h3bc94555),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb580a),
	.w1(32'hba326dff),
	.w2(32'hbd0dcdea),
	.w3(32'hbca78037),
	.w4(32'hbc03ef5f),
	.w5(32'hbb2bd8b4),
	.w6(32'h3d890d52),
	.w7(32'h3cd3e185),
	.w8(32'hbd537652),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e9376),
	.w1(32'hbad49fbe),
	.w2(32'hbbb224af),
	.w3(32'h3bae3607),
	.w4(32'hbbbeec71),
	.w5(32'hbbb01b88),
	.w6(32'hbb9c85ac),
	.w7(32'h3a8a3872),
	.w8(32'hbb2df665),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d92d6),
	.w1(32'h3ad06c56),
	.w2(32'h384ef554),
	.w3(32'h3bf61180),
	.w4(32'hbb2ce16a),
	.w5(32'hbbc44c04),
	.w6(32'hbad14d1f),
	.w7(32'h3b349e2a),
	.w8(32'h3c42310a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6671b0),
	.w1(32'hbabb474e),
	.w2(32'hbabcd2db),
	.w3(32'h3c11f098),
	.w4(32'hbba6c906),
	.w5(32'h39ed854c),
	.w6(32'hbb3d817b),
	.w7(32'hb84a33b3),
	.w8(32'hb9c3dc4d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96f763),
	.w1(32'h3b2217f0),
	.w2(32'hbb7309b2),
	.w3(32'h3bc54751),
	.w4(32'h3a618462),
	.w5(32'hbbc23cd0),
	.w6(32'hb9966d8c),
	.w7(32'h3a7dee59),
	.w8(32'hb9a1198d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2173),
	.w1(32'h39e281fa),
	.w2(32'h3bccc042),
	.w3(32'hbbc5af11),
	.w4(32'hbac88c05),
	.w5(32'h3acfbe44),
	.w6(32'hbaa1e787),
	.w7(32'h3b8e6262),
	.w8(32'h3b370936),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8f160),
	.w1(32'h3b0d4c1f),
	.w2(32'h3ab07703),
	.w3(32'h3b5c2853),
	.w4(32'h3b852b1e),
	.w5(32'h3b49b40f),
	.w6(32'h3a60da95),
	.w7(32'hbace4913),
	.w8(32'h3b8c28fe),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aa219),
	.w1(32'hbbbd2f41),
	.w2(32'hb985a268),
	.w3(32'h3b072734),
	.w4(32'hba5bc456),
	.w5(32'h3bd0b510),
	.w6(32'hbbae35cb),
	.w7(32'h39f9743a),
	.w8(32'h3ac5aa6e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a3c25),
	.w1(32'h3bcc4fa1),
	.w2(32'hbba99ce4),
	.w3(32'h3ab0b50e),
	.w4(32'h3bb8f0b7),
	.w5(32'hbb0df019),
	.w6(32'h3b0f95d1),
	.w7(32'h3b1196ba),
	.w8(32'h3a90ad98),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aaeb11),
	.w1(32'h3a87bb82),
	.w2(32'h3b21c4f6),
	.w3(32'hbb4644dc),
	.w4(32'h3b0b64c2),
	.w5(32'h3b35ff67),
	.w6(32'h3b46bac5),
	.w7(32'h3b0ad2bb),
	.w8(32'h3b0e7c94),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99fb8d),
	.w1(32'h3c4bf2e3),
	.w2(32'hbc978cb0),
	.w3(32'hba8a6fba),
	.w4(32'h3b935b34),
	.w5(32'hbca6a600),
	.w6(32'h3c42d0d7),
	.w7(32'hbbb58b75),
	.w8(32'hbcae49d1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a6b27),
	.w1(32'hbb66da26),
	.w2(32'h3b734df5),
	.w3(32'hbcfd1f1e),
	.w4(32'hbb3fce3a),
	.w5(32'h3bd69e03),
	.w6(32'h3a22d852),
	.w7(32'h3acb7cf4),
	.w8(32'h3a1610ec),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390bda32),
	.w1(32'h3bcc5163),
	.w2(32'h3b0eabde),
	.w3(32'h3b8d83a7),
	.w4(32'h3af6ecac),
	.w5(32'h3a8288c7),
	.w6(32'h3be3933f),
	.w7(32'h3b07585d),
	.w8(32'h3b0ef1bd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84de15),
	.w1(32'hbc975140),
	.w2(32'hbcf6a717),
	.w3(32'hbc530408),
	.w4(32'hbcaa1f5f),
	.w5(32'hbcb636ab),
	.w6(32'hbbd510fd),
	.w7(32'hbc02c688),
	.w8(32'hbc4863fc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb2bab),
	.w1(32'hbc311094),
	.w2(32'hbb90adb6),
	.w3(32'hbb1f8d05),
	.w4(32'hbb337733),
	.w5(32'hbb815da1),
	.w6(32'hbbd720f1),
	.w7(32'hbb0431dc),
	.w8(32'h3b0245aa),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bc843),
	.w1(32'hbb651862),
	.w2(32'hbb858500),
	.w3(32'hbb45f83a),
	.w4(32'hbb836d0d),
	.w5(32'hbba68390),
	.w6(32'hbb8f6cfc),
	.w7(32'hbaef0df0),
	.w8(32'h3b289b4e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baec7aa),
	.w1(32'hbb8bb8a9),
	.w2(32'hbbe5fa7b),
	.w3(32'h3b291293),
	.w4(32'hbb4b4af9),
	.w5(32'hbb8480ea),
	.w6(32'hbb7d59ee),
	.w7(32'h3b077a9e),
	.w8(32'hbb53218f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c131a80),
	.w1(32'hbbaea0a8),
	.w2(32'hbc831dc7),
	.w3(32'h3bc8a0ea),
	.w4(32'h3a8f58de),
	.w5(32'hbc01bce3),
	.w6(32'h3b2a0a1f),
	.w7(32'hbb59113f),
	.w8(32'hbbe2df5a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81f505),
	.w1(32'hbbe13400),
	.w2(32'hbbba875b),
	.w3(32'hbbf5d6a7),
	.w4(32'hbbabfe28),
	.w5(32'hbb90fe22),
	.w6(32'hbb98e4a0),
	.w7(32'hbb76f53c),
	.w8(32'hbbff661d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfc202),
	.w1(32'hbb081316),
	.w2(32'hbb578a02),
	.w3(32'h3aaa2b66),
	.w4(32'hbb110d3d),
	.w5(32'hbb973dd1),
	.w6(32'hbadc3e0b),
	.w7(32'h3a4e3e3d),
	.w8(32'h3b76ce05),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4de022),
	.w1(32'hba7c9913),
	.w2(32'hbc2e77dd),
	.w3(32'h3b0c79a0),
	.w4(32'h3ac35982),
	.w5(32'hbb2e4dd6),
	.w6(32'h3ba81791),
	.w7(32'h3b4e511c),
	.w8(32'hbb9b7136),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc76b31),
	.w1(32'h3ab531c9),
	.w2(32'h3b94eb1c),
	.w3(32'h3b6ebbe0),
	.w4(32'hbbf159be),
	.w5(32'hbac6072e),
	.w6(32'hbab7c3c9),
	.w7(32'h3a44abe1),
	.w8(32'h3b6648ed),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc47a3),
	.w1(32'hbb80f1f4),
	.w2(32'hbbf95ecf),
	.w3(32'hba4aaed9),
	.w4(32'h3aea15eb),
	.w5(32'hbb0aebe6),
	.w6(32'hb98cdf97),
	.w7(32'h388b12f7),
	.w8(32'h3b2d053c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76818e),
	.w1(32'hbbae0bb8),
	.w2(32'hbc98a8b2),
	.w3(32'hbcb22f15),
	.w4(32'hbc5927cd),
	.w5(32'hbc856c2a),
	.w6(32'hbbdefe87),
	.w7(32'hbbf7f5a3),
	.w8(32'hbb452919),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8645c3),
	.w1(32'hbc896566),
	.w2(32'hbcf7c8b7),
	.w3(32'hbc687d1a),
	.w4(32'hbca54b15),
	.w5(32'hbcf705d7),
	.w6(32'hbba2c635),
	.w7(32'hbc607984),
	.w8(32'hbcab9ebf),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdff49),
	.w1(32'h3c8b3fa3),
	.w2(32'hbc9dbaa5),
	.w3(32'hbc3819cf),
	.w4(32'h3bbd8ada),
	.w5(32'hbcd7eabe),
	.w6(32'h3c768dbd),
	.w7(32'hbb666f4a),
	.w8(32'hbcbc1a6a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a6b6f),
	.w1(32'hbc13b422),
	.w2(32'hbc3519a5),
	.w3(32'hbd1c8ebe),
	.w4(32'hbc3720fb),
	.w5(32'hbc053c11),
	.w6(32'h3987830a),
	.w7(32'h3b5ba43c),
	.w8(32'hbb9372b2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b36ad),
	.w1(32'hbb70a018),
	.w2(32'h3b21e41d),
	.w3(32'hba45e1cf),
	.w4(32'h3a7c691d),
	.w5(32'h3b311405),
	.w6(32'hbbb295e9),
	.w7(32'hb9807766),
	.w8(32'h3a9b6af5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb01e06),
	.w1(32'hbb311fb4),
	.w2(32'hbc995237),
	.w3(32'h3b1c2ed0),
	.w4(32'hbb7bed15),
	.w5(32'hbba3d76f),
	.w6(32'h3bd1b658),
	.w7(32'hbac6a9b0),
	.w8(32'hbbd07290),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadab8c7),
	.w1(32'hb9149212),
	.w2(32'h3baa1817),
	.w3(32'h3b45aca8),
	.w4(32'h3bbb3280),
	.w5(32'h3bd6a82a),
	.w6(32'h3b5785d8),
	.w7(32'h3b6ea71a),
	.w8(32'hb9fb418b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76f9bd),
	.w1(32'hbbbac7e6),
	.w2(32'hbb3808d9),
	.w3(32'h3c53a34f),
	.w4(32'hbbbaeabd),
	.w5(32'hbb1caa60),
	.w6(32'hbbdd986c),
	.w7(32'hbb488253),
	.w8(32'h3bde4a86),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c04ba),
	.w1(32'h3bc4a8f4),
	.w2(32'hbc00762a),
	.w3(32'h3ca1a637),
	.w4(32'h3b98c698),
	.w5(32'hbc0018b4),
	.w6(32'h3c172323),
	.w7(32'h3a7797db),
	.w8(32'hbc0816ca),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23688c),
	.w1(32'h3b1ca6b2),
	.w2(32'hbba89750),
	.w3(32'hbbd6e401),
	.w4(32'hbb328722),
	.w5(32'hbb173fe6),
	.w6(32'h3a56c80d),
	.w7(32'hba5421ab),
	.w8(32'hbbb33996),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fbcc6),
	.w1(32'hbb8b9cce),
	.w2(32'hb9fd6e0a),
	.w3(32'hb9cbaad9),
	.w4(32'hbb79b466),
	.w5(32'h3b377df7),
	.w6(32'hbb7f97e1),
	.w7(32'hbb0ce297),
	.w8(32'h3be51e29),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b565e05),
	.w1(32'h39134f92),
	.w2(32'hb969135a),
	.w3(32'h3b92a6a6),
	.w4(32'hb9ff5e71),
	.w5(32'hbb54551d),
	.w6(32'h394f50e1),
	.w7(32'h3adbd850),
	.w8(32'h3ac39b33),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fa6a0),
	.w1(32'hbb392911),
	.w2(32'hbc2af573),
	.w3(32'hbc85ff9a),
	.w4(32'hbc55d552),
	.w5(32'hbc28eb3e),
	.w6(32'h3b2cb5de),
	.w7(32'h3adf8cbe),
	.w8(32'hba0134cc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc042d),
	.w1(32'h3bcacbdf),
	.w2(32'h3c07b9c5),
	.w3(32'h3c1a8a67),
	.w4(32'h3b6c764a),
	.w5(32'h3bba1a61),
	.w6(32'h3a114f38),
	.w7(32'h3b2033cd),
	.w8(32'h3ba865ce),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaac5d),
	.w1(32'h3c7ff6fa),
	.w2(32'hbbdc4789),
	.w3(32'h3b790924),
	.w4(32'h3c2a5442),
	.w5(32'hbc153830),
	.w6(32'h3c2fd8d1),
	.w7(32'h3a96abe5),
	.w8(32'hbc0c3ad8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab3cda),
	.w1(32'hbb2ff066),
	.w2(32'h3a8bd9c2),
	.w3(32'hbca6ffcd),
	.w4(32'hba40c90d),
	.w5(32'h3bac180d),
	.w6(32'h3a4a5256),
	.w7(32'h3b053739),
	.w8(32'h3bdd250b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b775d63),
	.w1(32'h3ace7e80),
	.w2(32'hb951fe0c),
	.w3(32'h3b5a5a3a),
	.w4(32'h3a02a956),
	.w5(32'hbbdea938),
	.w6(32'hbbaf1b47),
	.w7(32'hbb2dcaf6),
	.w8(32'hbb18918c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb602ac1),
	.w1(32'h3b53f5df),
	.w2(32'hbbbfbb22),
	.w3(32'hbaff5290),
	.w4(32'hbb24f13c),
	.w5(32'hbac3eb29),
	.w6(32'h3bf40517),
	.w7(32'h3c006c2f),
	.w8(32'h3bb61701),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b050cd3),
	.w1(32'h3b1b48c0),
	.w2(32'hbb39209a),
	.w3(32'hbb20164d),
	.w4(32'hbaf01289),
	.w5(32'hbad0fdaf),
	.w6(32'h3ad3254d),
	.w7(32'h3a87c47c),
	.w8(32'h3bc41d48),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d62c1),
	.w1(32'h3be7a58e),
	.w2(32'hbc5b8053),
	.w3(32'h3c138c2b),
	.w4(32'h3c0f64a5),
	.w5(32'hbbaba0c7),
	.w6(32'h3c031beb),
	.w7(32'h3bd3f2f3),
	.w8(32'hbc635861),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39fc13),
	.w1(32'hbbeba420),
	.w2(32'hbbd080f2),
	.w3(32'h39a6744c),
	.w4(32'hbbd71089),
	.w5(32'hbbfbeef1),
	.w6(32'hbc092dbd),
	.w7(32'hbbc77de5),
	.w8(32'hbc5ba183),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cf84d),
	.w1(32'hba807364),
	.w2(32'hbb1f1a95),
	.w3(32'hbca14da8),
	.w4(32'h3a3e0d82),
	.w5(32'hbc006587),
	.w6(32'h3baff888),
	.w7(32'hbaf9a2de),
	.w8(32'hbaeb7080),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae48f81),
	.w1(32'hbb0b9a0d),
	.w2(32'hbb448aa7),
	.w3(32'hbb61a1e7),
	.w4(32'h39ce2b41),
	.w5(32'hbb028864),
	.w6(32'hbbca37d6),
	.w7(32'hbba0f3c1),
	.w8(32'h3a07ae43),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6279d),
	.w1(32'hbc1755d1),
	.w2(32'hbc415140),
	.w3(32'hbc6fedb4),
	.w4(32'hbc5a5ac2),
	.w5(32'hbb5711a1),
	.w6(32'hbc0e22ad),
	.w7(32'hbba17bd8),
	.w8(32'hbba81166),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad877a3),
	.w1(32'hbc33fd96),
	.w2(32'hbc28a2a7),
	.w3(32'h3b2f7f7e),
	.w4(32'hbc131235),
	.w5(32'hbbefd112),
	.w6(32'hbc097dab),
	.w7(32'hbc08105d),
	.w8(32'hbc194e37),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a6a58),
	.w1(32'hbbe36e8a),
	.w2(32'hbbe699cb),
	.w3(32'hbbe5321f),
	.w4(32'hbb66d6c5),
	.w5(32'hbb35af91),
	.w6(32'h3ace0531),
	.w7(32'h3ac06f07),
	.w8(32'hbb7a8e64),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ae2eb),
	.w1(32'hbb9e38d2),
	.w2(32'hbb92cf1f),
	.w3(32'h3b9d8b50),
	.w4(32'hbbbf040c),
	.w5(32'h39309c7e),
	.w6(32'hbb93fb1d),
	.w7(32'hbb8d1d34),
	.w8(32'h3b7ed196),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c604146),
	.w1(32'hbbf68b2c),
	.w2(32'hbc42d934),
	.w3(32'h3be9e59d),
	.w4(32'hbbf0b5e4),
	.w5(32'hbba4a05f),
	.w6(32'h3ae634ec),
	.w7(32'hb9d3a264),
	.w8(32'h3b88d8ba),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f980d),
	.w1(32'hbc3a0f45),
	.w2(32'hbc676478),
	.w3(32'h3c58b9f9),
	.w4(32'hbc51fd3c),
	.w5(32'hbc0d2510),
	.w6(32'hba96e602),
	.w7(32'hbbb40285),
	.w8(32'hbbe73d16),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1094c1),
	.w1(32'h38819e8c),
	.w2(32'h3c1330e1),
	.w3(32'hbba92b97),
	.w4(32'h3b49282f),
	.w5(32'h3b8d1aa1),
	.w6(32'h39b28108),
	.w7(32'h3b4cd573),
	.w8(32'h3b593cd7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29a54f),
	.w1(32'h39cdcc93),
	.w2(32'h3a7c5bdb),
	.w3(32'h3b686a86),
	.w4(32'h39a633ba),
	.w5(32'h3b1ba245),
	.w6(32'hb99a20a1),
	.w7(32'hbb2fc864),
	.w8(32'hb7c9765d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc078734),
	.w1(32'hbba4b697),
	.w2(32'hbb3032b7),
	.w3(32'h3ac8905c),
	.w4(32'hb9f97d92),
	.w5(32'h3affa277),
	.w6(32'hb96e093d),
	.w7(32'hbaa0633f),
	.w8(32'hbb9cf91e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13fbb3),
	.w1(32'h3ae6a869),
	.w2(32'hbc1c29ef),
	.w3(32'hbb38ec05),
	.w4(32'h3a0c7da1),
	.w5(32'hbb300be2),
	.w6(32'h3c85ebb2),
	.w7(32'h3a558a14),
	.w8(32'hbb8b6723),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92cf23),
	.w1(32'hbcfbc8a4),
	.w2(32'hbcd7c5d1),
	.w3(32'hbd0b58ee),
	.w4(32'hbcebc37a),
	.w5(32'hbcc27453),
	.w6(32'hbc9e7da9),
	.w7(32'hba1aa14e),
	.w8(32'hbc67a4f8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5853ba),
	.w1(32'hbc1c7be9),
	.w2(32'hbccaa60d),
	.w3(32'hbbedeecf),
	.w4(32'hbc2be22a),
	.w5(32'hbc6e2229),
	.w6(32'hb9e27c8d),
	.w7(32'h3a8ac074),
	.w8(32'hba83c5f3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba271bf8),
	.w1(32'hbbaf1048),
	.w2(32'hbbed3a1b),
	.w3(32'hba9bd432),
	.w4(32'hbb3062f1),
	.w5(32'hbc3fb033),
	.w6(32'h3bab1f61),
	.w7(32'h3bd6e754),
	.w8(32'hbb209bc3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b180a90),
	.w1(32'hbb5c845c),
	.w2(32'h3a1e742f),
	.w3(32'h3abbe45e),
	.w4(32'hbaf70663),
	.w5(32'h3afb2654),
	.w6(32'hbb5556a4),
	.w7(32'hbad42a7f),
	.w8(32'h3b082d42),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92d370),
	.w1(32'hbb204126),
	.w2(32'hba5542b7),
	.w3(32'h3b884623),
	.w4(32'h3ab75ef6),
	.w5(32'h3a3a4ef9),
	.w6(32'hbb5be462),
	.w7(32'h3aec7bd3),
	.w8(32'h3aeeef3c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43f4f1),
	.w1(32'hba6933f4),
	.w2(32'h397b97ed),
	.w3(32'hbb383734),
	.w4(32'hbb8e4d5e),
	.w5(32'h3a9f8888),
	.w6(32'hbb22aa6b),
	.w7(32'hb9d02959),
	.w8(32'h3b045fa0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0ce0c),
	.w1(32'h39c60a37),
	.w2(32'h3b1d3d1f),
	.w3(32'h3c0b2383),
	.w4(32'h3abb88ad),
	.w5(32'h3a3bafdf),
	.w6(32'hbb0fa885),
	.w7(32'h3b0d1a0a),
	.w8(32'h3b0a5c53),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c8464),
	.w1(32'hbbb3e378),
	.w2(32'hbbb8013b),
	.w3(32'h39af0c98),
	.w4(32'hbb9847bc),
	.w5(32'hbbcd4e5e),
	.w6(32'h3aab73f8),
	.w7(32'hba36034c),
	.w8(32'hbb7d1142),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dca392),
	.w1(32'h3af1058f),
	.w2(32'h3ac1653c),
	.w3(32'hbb8415d1),
	.w4(32'h3a80868d),
	.w5(32'h3b03c2bc),
	.w6(32'h3b6d0093),
	.w7(32'h3a0336b5),
	.w8(32'h3a04a33f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3caa54),
	.w1(32'hbc02f5bd),
	.w2(32'h3ba62824),
	.w3(32'h3b4dde9c),
	.w4(32'hbb7d1328),
	.w5(32'h3c0cc080),
	.w6(32'hbc54b03f),
	.w7(32'hbb1f09b5),
	.w8(32'h3b80c9c8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59c2cc),
	.w1(32'hbb09c72e),
	.w2(32'hbb9c6b43),
	.w3(32'h3c643ff5),
	.w4(32'hbb4f4dd7),
	.w5(32'hbbbbb326),
	.w6(32'hb88ab287),
	.w7(32'h372b5fdf),
	.w8(32'hbb05ceab),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dbed0),
	.w1(32'hbb742c91),
	.w2(32'hbc0b732e),
	.w3(32'h39ad1aa6),
	.w4(32'hbb5a02b2),
	.w5(32'h3b7e6800),
	.w6(32'hba1531fe),
	.w7(32'hb8c9016b),
	.w8(32'h3b5097d7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fa50a),
	.w1(32'h3b8f1ac1),
	.w2(32'h3b35474c),
	.w3(32'h3b747984),
	.w4(32'h3bb0b504),
	.w5(32'h3b852009),
	.w6(32'h3bab78c7),
	.w7(32'h3baab9a0),
	.w8(32'h3b946770),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fb562),
	.w1(32'hbc0cdebd),
	.w2(32'hbc3470af),
	.w3(32'h3ba95b9e),
	.w4(32'hbc2c2992),
	.w5(32'hbbacf146),
	.w6(32'hbbcaa0d5),
	.w7(32'hbafc7ff5),
	.w8(32'hbbaad5c6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb54186),
	.w1(32'hba910ece),
	.w2(32'h3c0c35c6),
	.w3(32'h3bbb20ab),
	.w4(32'h3b6eb56b),
	.w5(32'h3bc24503),
	.w6(32'h3bb4f08a),
	.w7(32'h3ba6a689),
	.w8(32'h3b199fe3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dc73f),
	.w1(32'h3a5bf5b6),
	.w2(32'h3b958219),
	.w3(32'h3ac8a6d8),
	.w4(32'h3a2cf825),
	.w5(32'h3b84da55),
	.w6(32'hbb7d9dad),
	.w7(32'h3b7fd13d),
	.w8(32'hbb2ac28e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2297cb),
	.w1(32'hbb3ac6a9),
	.w2(32'hbb2c70ca),
	.w3(32'h3b8c7c52),
	.w4(32'hbba9909f),
	.w5(32'hbbbd6ac8),
	.w6(32'hba8f2262),
	.w7(32'hba561160),
	.w8(32'h38bf6bf0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed381a),
	.w1(32'hbc1660eb),
	.w2(32'h3a96b824),
	.w3(32'h3b6df7f7),
	.w4(32'hbc07afcd),
	.w5(32'hbb4667ee),
	.w6(32'h3bb7390b),
	.w7(32'h3af9efc6),
	.w8(32'h3aa1682f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb871770),
	.w1(32'hbc102ebb),
	.w2(32'h3b33993b),
	.w3(32'h3a5c711c),
	.w4(32'hbb930ac0),
	.w5(32'h3c0a025c),
	.w6(32'hbbf80996),
	.w7(32'hbb294f2c),
	.w8(32'hbb74a165),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dbee0),
	.w1(32'hbb05ac34),
	.w2(32'hbb150e2a),
	.w3(32'hb940994b),
	.w4(32'h3adcb0b8),
	.w5(32'hbb6dd2a8),
	.w6(32'hbbd089cf),
	.w7(32'hba516118),
	.w8(32'h3a36e836),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38c60c),
	.w1(32'hbb46b5e6),
	.w2(32'h3c151d54),
	.w3(32'hbad7b95a),
	.w4(32'hbb0ae5d8),
	.w5(32'h3c14c344),
	.w6(32'hbb8f02c0),
	.w7(32'hbbb7f229),
	.w8(32'h39941607),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2453b8),
	.w1(32'h3b320245),
	.w2(32'h3b35be48),
	.w3(32'h3b14e25d),
	.w4(32'h3b37b441),
	.w5(32'h394c9c2d),
	.w6(32'h3abaf9b1),
	.w7(32'h3b9e5635),
	.w8(32'h3bb4b444),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c306d3c),
	.w1(32'h3c537ae7),
	.w2(32'hbc1a3540),
	.w3(32'h3b91c397),
	.w4(32'h3bc18adb),
	.w5(32'hbc06fa42),
	.w6(32'h3c261840),
	.w7(32'h3b1270e2),
	.w8(32'hbc7cad72),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc408b74),
	.w1(32'hbb9a1262),
	.w2(32'hbb14981b),
	.w3(32'hbc496727),
	.w4(32'hbba01593),
	.w5(32'h3a335aee),
	.w6(32'hbb5ed474),
	.w7(32'hbb8dff42),
	.w8(32'hba8a2c91),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf0de0),
	.w1(32'h398ccb14),
	.w2(32'hb88021f2),
	.w3(32'h3c288a70),
	.w4(32'hba21b9aa),
	.w5(32'h3af8c505),
	.w6(32'hbb47637b),
	.w7(32'h3a38599c),
	.w8(32'h3a0c0ec9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fedab),
	.w1(32'h3ba3f48d),
	.w2(32'h3bc1605a),
	.w3(32'h39bfc04a),
	.w4(32'h3b4b81f5),
	.w5(32'h3bafb74f),
	.w6(32'h3b78881a),
	.w7(32'h3b9314a7),
	.w8(32'h3b7cd3d2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb088ab),
	.w1(32'h3c14951b),
	.w2(32'hbb70f725),
	.w3(32'h38bd7630),
	.w4(32'h3b9f037e),
	.w5(32'hbbddfb6a),
	.w6(32'h3c0c8509),
	.w7(32'hbabf9d4c),
	.w8(32'hbbcafa0e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6eedd9),
	.w1(32'h3a0fe9ce),
	.w2(32'hbb38b194),
	.w3(32'hbc6e4684),
	.w4(32'h3b9fb8af),
	.w5(32'h3aaddd6f),
	.w6(32'h3b5a628a),
	.w7(32'h3c184fbd),
	.w8(32'h3bafde99),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31dbd3),
	.w1(32'hbb593f82),
	.w2(32'h3b93cc33),
	.w3(32'hbb1a4897),
	.w4(32'h3491fe74),
	.w5(32'h3bc069d9),
	.w6(32'hbb8b7c5c),
	.w7(32'h3b85998a),
	.w8(32'h3be7280b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8998c4),
	.w1(32'h3bb33c86),
	.w2(32'h3bb447a0),
	.w3(32'h3ca1e97c),
	.w4(32'h3ba165ab),
	.w5(32'h3bf49f03),
	.w6(32'h3be5fffe),
	.w7(32'h3b068b85),
	.w8(32'h3ad63f83),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba868e05),
	.w1(32'hbb9406a8),
	.w2(32'hbbbdf50d),
	.w3(32'h3a2e4f3c),
	.w4(32'hbbd72df2),
	.w5(32'hbb5ca7fb),
	.w6(32'hba544e44),
	.w7(32'hbb42340f),
	.w8(32'hbb7fe1f0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd909b9),
	.w1(32'hbb335bf2),
	.w2(32'hbb7f0efb),
	.w3(32'h3b5109fd),
	.w4(32'hbb82f33e),
	.w5(32'hbb992b3e),
	.w6(32'hbad3ed68),
	.w7(32'hbb16d5d1),
	.w8(32'hbb38759e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58ec9c),
	.w1(32'h3c27a721),
	.w2(32'hbc283826),
	.w3(32'hbb74576e),
	.w4(32'h3be24493),
	.w5(32'hbc364ccc),
	.w6(32'h3c1b3f8e),
	.w7(32'hbb074c42),
	.w8(32'hbc37f61a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbcd5ff),
	.w1(32'hba033646),
	.w2(32'hbb7efc52),
	.w3(32'hbc9c9d4e),
	.w4(32'h3ab5e0af),
	.w5(32'hbba7a3fb),
	.w6(32'h3aded8ca),
	.w7(32'hbb0b2c7c),
	.w8(32'hba502eb1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e3ac5),
	.w1(32'h3aba7309),
	.w2(32'hbb30917d),
	.w3(32'hb7f7b524),
	.w4(32'hb9fbbd40),
	.w5(32'hba98e73a),
	.w6(32'hba4d2375),
	.w7(32'h3a7f37f0),
	.w8(32'hbaec066f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45be87),
	.w1(32'hbb9a7e50),
	.w2(32'hb9c92692),
	.w3(32'h39e724e1),
	.w4(32'h3b1c435f),
	.w5(32'h39ce10fd),
	.w6(32'hbaadd826),
	.w7(32'hba8fc514),
	.w8(32'h3a7dcb15),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba06b5c),
	.w1(32'hbbb0b0a3),
	.w2(32'hbb61f7dd),
	.w3(32'h3aada0fe),
	.w4(32'hbb42cbba),
	.w5(32'hba199b89),
	.w6(32'hbafb934d),
	.w7(32'hbad9c23a),
	.w8(32'hba857232),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9b87b),
	.w1(32'hbb6dea19),
	.w2(32'hbb77c6da),
	.w3(32'h3ba13b61),
	.w4(32'hbbbf9dea),
	.w5(32'hbaecb887),
	.w6(32'hbaec3ae5),
	.w7(32'h3b377412),
	.w8(32'hbaa8d7aa),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe6433),
	.w1(32'hbc0b72b2),
	.w2(32'hbbadba55),
	.w3(32'h39b138b3),
	.w4(32'h39a81b5e),
	.w5(32'hbb466b3e),
	.w6(32'hb9b135c5),
	.w7(32'h3a5119b3),
	.w8(32'h3a8d1b38),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba2780),
	.w1(32'hbbea6abe),
	.w2(32'h3b1a63e9),
	.w3(32'hbb7933a7),
	.w4(32'hbbaebd33),
	.w5(32'h3b275c54),
	.w6(32'hbc02ea71),
	.w7(32'hba89bd81),
	.w8(32'h3b534ee2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab0857),
	.w1(32'hbb6df9ac),
	.w2(32'hbabefa4d),
	.w3(32'h3bda2882),
	.w4(32'hba210924),
	.w5(32'h3aaa99ea),
	.w6(32'hbafe49de),
	.w7(32'h3b520126),
	.w8(32'h3ab4e4e8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bd356),
	.w1(32'hbbc6396f),
	.w2(32'hbbc44e4b),
	.w3(32'hbbd0e37b),
	.w4(32'hbbb8d785),
	.w5(32'hbbde5b7e),
	.w6(32'hbb321d34),
	.w7(32'hbb724d34),
	.w8(32'h3b0340fa),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c97d),
	.w1(32'h3b2b6a51),
	.w2(32'h3bc51c60),
	.w3(32'hbaab752d),
	.w4(32'h3bb0e9c9),
	.w5(32'hbb8f9da0),
	.w6(32'hba367287),
	.w7(32'h3b5c7c3c),
	.w8(32'h3b629277),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b547859),
	.w1(32'hbbd3941c),
	.w2(32'hbbd0f397),
	.w3(32'h3aca3291),
	.w4(32'hbb32dabc),
	.w5(32'hba0a88fe),
	.w6(32'h3a007aef),
	.w7(32'h3af78f03),
	.w8(32'h3a8d4430),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a167f4a),
	.w1(32'h3aa08f24),
	.w2(32'hb91117f2),
	.w3(32'h3bb20ce4),
	.w4(32'h3c010ecb),
	.w5(32'h39e47296),
	.w6(32'h3b9734ac),
	.w7(32'h3ba770cb),
	.w8(32'hbb721cf7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule