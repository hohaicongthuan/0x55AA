module layer_10_featuremap_360(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc6add),
	.w1(32'hba23cb82),
	.w2(32'hba8ef2b4),
	.w3(32'h3a608b91),
	.w4(32'hb9886509),
	.w5(32'h3a44d289),
	.w6(32'h3aa10a02),
	.w7(32'hbaa6c4ba),
	.w8(32'h3ae091da),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad7cb),
	.w1(32'h3ab0a3c6),
	.w2(32'h3a5c383f),
	.w3(32'h3b958dd7),
	.w4(32'h3b0ca6b2),
	.w5(32'h3b255e69),
	.w6(32'h3ae016c8),
	.w7(32'hba4d4fcb),
	.w8(32'h3b29f10c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c8015),
	.w1(32'hbb7fd3f3),
	.w2(32'hbb550abb),
	.w3(32'h3b2818fe),
	.w4(32'h3c0178f8),
	.w5(32'hba8c3cd6),
	.w6(32'h3bcf4cb3),
	.w7(32'h3a73f860),
	.w8(32'hb9a9e1e5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11be87),
	.w1(32'h3a073ea2),
	.w2(32'h39db5965),
	.w3(32'hba6d59fd),
	.w4(32'hba479b4e),
	.w5(32'hbb3ec920),
	.w6(32'h39f6e8c9),
	.w7(32'h3a4450b6),
	.w8(32'hbbacf86c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b9514),
	.w1(32'hbb89ac44),
	.w2(32'hbb168063),
	.w3(32'hbbc02b4f),
	.w4(32'hbbaa2038),
	.w5(32'h38630a31),
	.w6(32'hbbb7a72f),
	.w7(32'hbb44d391),
	.w8(32'h3a1c21f0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93375ea),
	.w1(32'hb9c37e2b),
	.w2(32'h3958f9da),
	.w3(32'h3a334920),
	.w4(32'h3a84d230),
	.w5(32'hb986785c),
	.w6(32'h3962726e),
	.w7(32'hb8b1f135),
	.w8(32'hba2476cd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b7e1f),
	.w1(32'hbae541e3),
	.w2(32'hbb07d7e4),
	.w3(32'h3a87a0f9),
	.w4(32'hbaac341d),
	.w5(32'h3a90bac3),
	.w6(32'h3930119f),
	.w7(32'hbaf22dd6),
	.w8(32'h3b322b77),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92a5cb),
	.w1(32'hbbdff98a),
	.w2(32'hbb958b54),
	.w3(32'hbb829e1c),
	.w4(32'hb9ec6078),
	.w5(32'hbb22780d),
	.w6(32'h3b0a3433),
	.w7(32'h3a8acea1),
	.w8(32'hbb674782),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f75d5),
	.w1(32'hbb1adbce),
	.w2(32'hbb1b0018),
	.w3(32'hbad06020),
	.w4(32'hb9f386a5),
	.w5(32'hba829502),
	.w6(32'hbafc9a78),
	.w7(32'hbaed6f3c),
	.w8(32'hb9a78975),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb014a74),
	.w1(32'hbac9e61a),
	.w2(32'hbb3821d8),
	.w3(32'hba6947b9),
	.w4(32'hbac71081),
	.w5(32'hbb4c342a),
	.w6(32'hbaac8b83),
	.w7(32'hb9899f32),
	.w8(32'hbafbf0c4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19ec74),
	.w1(32'hba26ec64),
	.w2(32'hba6ec9ed),
	.w3(32'hb9af8c79),
	.w4(32'h3a2fda1e),
	.w5(32'h3a129ea6),
	.w6(32'h3ad615e5),
	.w7(32'h3a80fb06),
	.w8(32'h3aba61d8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb2ec9),
	.w1(32'h3b07511b),
	.w2(32'hba11ca9f),
	.w3(32'h3ade8701),
	.w4(32'h3b1927bf),
	.w5(32'h3bcde777),
	.w6(32'h3b39e254),
	.w7(32'h399f3557),
	.w8(32'h3b9502bd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f2403),
	.w1(32'hba233d31),
	.w2(32'hbb09ff88),
	.w3(32'h3bec227a),
	.w4(32'h3ac0ce36),
	.w5(32'hbba12425),
	.w6(32'h3b7c4e18),
	.w7(32'hb957c76c),
	.w8(32'hbb572da5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06dad6),
	.w1(32'hbb5719c7),
	.w2(32'hba101fff),
	.w3(32'hbb3ca455),
	.w4(32'hba5956ff),
	.w5(32'hbb184c3d),
	.w6(32'hbb4cd095),
	.w7(32'hbac9defa),
	.w8(32'hbae8015b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fdf9d6),
	.w1(32'hb9b59a3f),
	.w2(32'hb9c856a6),
	.w3(32'hba592cc8),
	.w4(32'h3aff3d95),
	.w5(32'hba2ba046),
	.w6(32'hbb258f92),
	.w7(32'h398d0959),
	.w8(32'hbac0fc42),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f9e37),
	.w1(32'hbade3082),
	.w2(32'hba982828),
	.w3(32'hbb2a06d1),
	.w4(32'hbad39a60),
	.w5(32'h3aa32d1f),
	.w6(32'hbba8d387),
	.w7(32'hbb35b3d9),
	.w8(32'hb9b3627c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97a461),
	.w1(32'hbb6a266b),
	.w2(32'hbae3e016),
	.w3(32'h3a0fbe04),
	.w4(32'hb8cd9775),
	.w5(32'hb88c4899),
	.w6(32'hb9d8d78e),
	.w7(32'hba822bb5),
	.w8(32'h381e9b04),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09c429),
	.w1(32'hbc032545),
	.w2(32'hbc038bee),
	.w3(32'hbc02d33c),
	.w4(32'hbc0a9aa1),
	.w5(32'hbc0109c0),
	.w6(32'hbb4045b0),
	.w7(32'hbb972150),
	.w8(32'hbbf1f8eb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc9b56),
	.w1(32'hbc06d3bd),
	.w2(32'hbbfe5bf8),
	.w3(32'hbbb19c1b),
	.w4(32'hbbd3bf39),
	.w5(32'hbbadec22),
	.w6(32'hbc02c2e7),
	.w7(32'hbbf2012a),
	.w8(32'hbb76818c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb049735),
	.w1(32'hbadf20e9),
	.w2(32'h3b01f98b),
	.w3(32'hba855a50),
	.w4(32'hb9a9905a),
	.w5(32'h3a0bbb8c),
	.w6(32'hb9ea071b),
	.w7(32'h3a2c6202),
	.w8(32'hb9e7a0af),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4be88c),
	.w1(32'h3a06c57e),
	.w2(32'hba2a1038),
	.w3(32'h3ace1776),
	.w4(32'h3ab8edb4),
	.w5(32'hb982a17c),
	.w6(32'hbaa410e9),
	.w7(32'h39873be2),
	.w8(32'hb9ea2a5f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d3c84),
	.w1(32'hba59427a),
	.w2(32'hba9b2ee0),
	.w3(32'h39c7e3af),
	.w4(32'hba46ecd1),
	.w5(32'h3b04bf08),
	.w6(32'hba39a1f3),
	.w7(32'hbaaf7f32),
	.w8(32'h3acd95c6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc050b8b),
	.w1(32'hbb7b63e7),
	.w2(32'hbc0c6f0b),
	.w3(32'hbb9f3a22),
	.w4(32'hbb6a74b8),
	.w5(32'hbc32e841),
	.w6(32'hbb782cb2),
	.w7(32'hbbea155c),
	.w8(32'hbc0d5012),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8e996),
	.w1(32'hb877c68d),
	.w2(32'hbb16d9bf),
	.w3(32'hba2ba2b4),
	.w4(32'hbb78d9a9),
	.w5(32'hba229d90),
	.w6(32'hbb1069c6),
	.w7(32'hbb0e4bc9),
	.w8(32'h3b8306b5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc327ac),
	.w1(32'h3b5f490f),
	.w2(32'hba61eb83),
	.w3(32'h3b876531),
	.w4(32'h3bf5432e),
	.w5(32'hbaded893),
	.w6(32'hb9921f16),
	.w7(32'hba8cdd97),
	.w8(32'hbbcb41df),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6296a),
	.w1(32'hb9ec2ec1),
	.w2(32'h39c43569),
	.w3(32'hbae07bc0),
	.w4(32'hba9f7b69),
	.w5(32'h3b1e23e1),
	.w6(32'hbaefc980),
	.w7(32'h39acef57),
	.w8(32'h3ad912e7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a358e32),
	.w1(32'hb93bc117),
	.w2(32'hba1b0346),
	.w3(32'h3a208629),
	.w4(32'h39bd168b),
	.w5(32'hba5b861a),
	.w6(32'hb87fe620),
	.w7(32'hba852957),
	.w8(32'hba6e9f22),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b2be8),
	.w1(32'hb975ef37),
	.w2(32'hba9fe2b9),
	.w3(32'h3a40e008),
	.w4(32'h3a0a4e06),
	.w5(32'hbb4b1866),
	.w6(32'hba981c10),
	.w7(32'hbb36d840),
	.w8(32'hbb59f377),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92dda8d),
	.w1(32'h3ab12bf7),
	.w2(32'h3aac6e65),
	.w3(32'h3ab9b7e8),
	.w4(32'h3b72799e),
	.w5(32'h3b011519),
	.w6(32'hbac63047),
	.w7(32'h3a4ae588),
	.w8(32'h3b3c46ad),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f647f),
	.w1(32'h3b0dcce9),
	.w2(32'hbb1f63e3),
	.w3(32'hba118dbb),
	.w4(32'h39413154),
	.w5(32'hbb50c864),
	.w6(32'hb9b63c5f),
	.w7(32'hbad35ccb),
	.w8(32'hbb62c110),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0650d),
	.w1(32'h3b3ef4a3),
	.w2(32'h3b943407),
	.w3(32'hbb35442d),
	.w4(32'hbb7bf156),
	.w5(32'h3b13c98e),
	.w6(32'hbafdf1af),
	.w7(32'hb891ec9e),
	.w8(32'h3b1fe92e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16c94e),
	.w1(32'hbabf50c4),
	.w2(32'h3a0ae520),
	.w3(32'hb93d18ac),
	.w4(32'h3a26558c),
	.w5(32'h39a11d80),
	.w6(32'h3b3c6d78),
	.w7(32'h39ecfe1d),
	.w8(32'h39e09c0b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8be98),
	.w1(32'hb90d78f2),
	.w2(32'hbad666bd),
	.w3(32'hba153dca),
	.w4(32'hba804558),
	.w5(32'h3a893dd7),
	.w6(32'h3b08ca59),
	.w7(32'h3ac2aa21),
	.w8(32'h3a852dbb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2d39e),
	.w1(32'h3a682880),
	.w2(32'hb9c350a8),
	.w3(32'h3a948459),
	.w4(32'hb998de51),
	.w5(32'hb9bbfdf2),
	.w6(32'hbadd90ee),
	.w7(32'hba8dac73),
	.w8(32'h3ad7ceeb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e18d1),
	.w1(32'h3b176fe0),
	.w2(32'hb9a376fa),
	.w3(32'hba3ff60d),
	.w4(32'hbb391517),
	.w5(32'h3ad0505c),
	.w6(32'h388a9a81),
	.w7(32'h3a4b815a),
	.w8(32'h398a4694),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a882b53),
	.w1(32'hba33bfcf),
	.w2(32'hba0c89dc),
	.w3(32'h3b277712),
	.w4(32'h3b496c41),
	.w5(32'hbba12afb),
	.w6(32'hba6e439c),
	.w7(32'hba312333),
	.w8(32'hbb314ca9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b44ea),
	.w1(32'hbb4bdc84),
	.w2(32'hbb2d7c92),
	.w3(32'hbbb6f9e3),
	.w4(32'hbb8dbfbb),
	.w5(32'hb844f4a2),
	.w6(32'hbbe050d9),
	.w7(32'hbb8fdca8),
	.w8(32'hbb2b5c06),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a681f54),
	.w1(32'h3bc3f535),
	.w2(32'h3b8abd42),
	.w3(32'h3bc3ac5b),
	.w4(32'h3bf795c6),
	.w5(32'h3b3b04ed),
	.w6(32'hbb2a8e7c),
	.w7(32'hb981dcc9),
	.w8(32'hb94a0a98),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc4ce1),
	.w1(32'h3ba73bbb),
	.w2(32'h3b82c541),
	.w3(32'h3bedbd38),
	.w4(32'h3b9dd966),
	.w5(32'hbb70d19f),
	.w6(32'h3bbf2e03),
	.w7(32'h3ad435f3),
	.w8(32'hbbc4a4ac),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1593f8),
	.w1(32'hbaffbaf3),
	.w2(32'hbb9f74b5),
	.w3(32'hbb3b3f72),
	.w4(32'hbbcdda33),
	.w5(32'hba260d78),
	.w6(32'hbb4e1043),
	.w7(32'hbbc3a982),
	.w8(32'hb8cb0118),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26ac40),
	.w1(32'h3b6041e8),
	.w2(32'h39b0e6b7),
	.w3(32'hba3e1b66),
	.w4(32'hbaa34647),
	.w5(32'hba851960),
	.w6(32'h3a4a784d),
	.w7(32'h389a33cf),
	.w8(32'hbaa6e1b0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8d479),
	.w1(32'h38cc79a4),
	.w2(32'h39efda6e),
	.w3(32'h3a1ca1f5),
	.w4(32'hba54a0db),
	.w5(32'hbb7b5209),
	.w6(32'h3a55eb00),
	.w7(32'hba69b6c6),
	.w8(32'hba91f34f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b352f80),
	.w1(32'h3b1e2bf4),
	.w2(32'h3b5cd269),
	.w3(32'hbae1510d),
	.w4(32'h3ad20478),
	.w5(32'h3b9af161),
	.w6(32'hba93fc79),
	.w7(32'h3a9174c6),
	.w8(32'h3acd6ed4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb0138),
	.w1(32'hbb9ed2e0),
	.w2(32'hbb550dc8),
	.w3(32'h3b270ed6),
	.w4(32'h3b87938c),
	.w5(32'hbbb06135),
	.w6(32'hbb8a0547),
	.w7(32'hbafd0f33),
	.w8(32'hbb2b2809),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30aede),
	.w1(32'hba94d2da),
	.w2(32'hbb6a4386),
	.w3(32'hbabe1aa6),
	.w4(32'h39d177a4),
	.w5(32'hb987d074),
	.w6(32'hbb4b1d2e),
	.w7(32'hba1086f6),
	.w8(32'hbad9bdb4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab5ae6),
	.w1(32'h390abe36),
	.w2(32'hba42dadc),
	.w3(32'hb9704cb7),
	.w4(32'hbaee68f9),
	.w5(32'hbb08b63c),
	.w6(32'hbb28875e),
	.w7(32'hbaab9791),
	.w8(32'hbb034163),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc04073),
	.w1(32'hbbb598f6),
	.w2(32'hbc0743c7),
	.w3(32'hbb3715bb),
	.w4(32'hbae6b701),
	.w5(32'hbaf66c3e),
	.w6(32'hbbbec3f2),
	.w7(32'hbb9b8855),
	.w8(32'hbb74978b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeb450),
	.w1(32'hbc13ec09),
	.w2(32'hbc098f7f),
	.w3(32'hbbf85993),
	.w4(32'hbbd15202),
	.w5(32'hbb097eac),
	.w6(32'hbb2c36fa),
	.w7(32'hbb7e8aea),
	.w8(32'hbad9f250),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87f2ca),
	.w1(32'h3b8b8c77),
	.w2(32'h3b9c8b38),
	.w3(32'h3b8e1ad9),
	.w4(32'h3b230eb5),
	.w5(32'hba84e71a),
	.w6(32'h3b87bd78),
	.w7(32'h3b832728),
	.w8(32'hbaa0963b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11ce46),
	.w1(32'hbb440a41),
	.w2(32'hbb839cac),
	.w3(32'hbae8b5d1),
	.w4(32'hbb2ad131),
	.w5(32'hbbfb40a2),
	.w6(32'hbab258e6),
	.w7(32'hbb620b00),
	.w8(32'hbb787700),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba606477),
	.w1(32'hbb181dfd),
	.w2(32'hba83a880),
	.w3(32'hbb0bffaa),
	.w4(32'hbab3eea9),
	.w5(32'h39d57bdb),
	.w6(32'hbaad98c4),
	.w7(32'h39c7999f),
	.w8(32'hb9acf07e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e461a),
	.w1(32'hba0f1bf0),
	.w2(32'h3a0c2cca),
	.w3(32'hb94fefb8),
	.w4(32'hb9d5fb63),
	.w5(32'hbb7d0a42),
	.w6(32'h39f47857),
	.w7(32'h3a3cfce1),
	.w8(32'hbb785d62),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6179e),
	.w1(32'h3a9385d1),
	.w2(32'h3a8d86d0),
	.w3(32'hbb351a39),
	.w4(32'hbae14a76),
	.w5(32'hbaeaa278),
	.w6(32'h398efdc5),
	.w7(32'h3aa43ac5),
	.w8(32'h3992f00e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25a8fb),
	.w1(32'hbb07362b),
	.w2(32'hbb944e35),
	.w3(32'hbbd55063),
	.w4(32'hbb998113),
	.w5(32'hbb626f54),
	.w6(32'h399797e4),
	.w7(32'hbbc23338),
	.w8(32'hbb62ef7a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71990a),
	.w1(32'h39c526c0),
	.w2(32'h3ad05cfe),
	.w3(32'h38276fc4),
	.w4(32'h3918a3a5),
	.w5(32'hbaa6accd),
	.w6(32'h3a4f54c4),
	.w7(32'h3ad9a655),
	.w8(32'hb94f0da8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1800e7),
	.w1(32'h3af8083d),
	.w2(32'hb9ec72b0),
	.w3(32'hbb1da8a3),
	.w4(32'hbb214244),
	.w5(32'h3a01a454),
	.w6(32'hba737f35),
	.w7(32'hbaa8e3ed),
	.w8(32'h3a4e146f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d3ed4),
	.w1(32'h3b1307b2),
	.w2(32'hba0e4cd6),
	.w3(32'h39055ad8),
	.w4(32'hb9b1cc81),
	.w5(32'hba7ae9a6),
	.w6(32'hba989f92),
	.w7(32'hba87975f),
	.w8(32'h3ae59cdf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93f3c8),
	.w1(32'hba9841a5),
	.w2(32'h3af127b5),
	.w3(32'h39a2972d),
	.w4(32'h3b97804f),
	.w5(32'hbaae3322),
	.w6(32'h3b0ef47a),
	.w7(32'h3b1bf522),
	.w8(32'hbabd1067),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab33116),
	.w1(32'hba7bf41b),
	.w2(32'hba17bb58),
	.w3(32'hb9ff089e),
	.w4(32'hbaa130bc),
	.w5(32'h3b38f63b),
	.w6(32'hb6f8af65),
	.w7(32'hbaf4eec5),
	.w8(32'h3998112c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f1b2),
	.w1(32'hbba40cdb),
	.w2(32'hbac457ef),
	.w3(32'h3a8e4451),
	.w4(32'h3a649a1d),
	.w5(32'hbb09b753),
	.w6(32'h3a88b9fe),
	.w7(32'h3abbfa61),
	.w8(32'hbb124537),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e5daf),
	.w1(32'hbba48e4f),
	.w2(32'hbb888132),
	.w3(32'hbb9b774f),
	.w4(32'hbb85480d),
	.w5(32'hbb0c7d41),
	.w6(32'hbaaa0357),
	.w7(32'hb9060d35),
	.w8(32'hbae383ff),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc015a),
	.w1(32'hbb793723),
	.w2(32'hbaf3756a),
	.w3(32'hbb726149),
	.w4(32'hbb0a27c2),
	.w5(32'hbb85fa87),
	.w6(32'hbb225f01),
	.w7(32'hbaa23165),
	.w8(32'hbae0859c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5059ca),
	.w1(32'h38bf62df),
	.w2(32'h3a2aaa70),
	.w3(32'hbb368a06),
	.w4(32'hbba44462),
	.w5(32'hba8f6542),
	.w6(32'hbabf0182),
	.w7(32'h3a49eb64),
	.w8(32'h38a265b1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d315),
	.w1(32'h3b2fbf1d),
	.w2(32'hba83f7dc),
	.w3(32'hbabc5116),
	.w4(32'hba5414c4),
	.w5(32'h38cbf5b0),
	.w6(32'hbab523b2),
	.w7(32'hba97e9a0),
	.w8(32'hbabd8f74),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba131220),
	.w1(32'h3a37f612),
	.w2(32'hb960ad9b),
	.w3(32'h39159d6e),
	.w4(32'hbad769ca),
	.w5(32'hba82d7b6),
	.w6(32'hbab0e053),
	.w7(32'hba64b8f1),
	.w8(32'hbafd878f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac78034),
	.w1(32'h3b43f766),
	.w2(32'h3b532c80),
	.w3(32'hbb11cae5),
	.w4(32'hba80b147),
	.w5(32'hb8c7a85b),
	.w6(32'hba92bfc3),
	.w7(32'h3b44f1c0),
	.w8(32'h3aeba0a7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7e366),
	.w1(32'hbaaf0ef6),
	.w2(32'hba2f2dfe),
	.w3(32'hbb6b183b),
	.w4(32'hb93a22b1),
	.w5(32'h3a14df89),
	.w6(32'hba4fdc5b),
	.w7(32'hba42aa4e),
	.w8(32'hba59ce7e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf3fc3),
	.w1(32'h3af02736),
	.w2(32'h3b03f4cd),
	.w3(32'h3b587d0c),
	.w4(32'h3b726c9c),
	.w5(32'h3a7c3a50),
	.w6(32'h38dd1129),
	.w7(32'hb9af93e5),
	.w8(32'hbb090c57),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb848fe1),
	.w1(32'hbb8030f5),
	.w2(32'hbb8e2971),
	.w3(32'hb99f05ca),
	.w4(32'h3b599bf9),
	.w5(32'h3aaf6f7c),
	.w6(32'hb98d068a),
	.w7(32'hbb05eae9),
	.w8(32'hbad73b62),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80892f),
	.w1(32'h3a6c5ee5),
	.w2(32'h3a67e005),
	.w3(32'h3c3940c8),
	.w4(32'h3c0e14fd),
	.w5(32'hbb5e1491),
	.w6(32'hbb2be4c9),
	.w7(32'hb9545c48),
	.w8(32'hbb899059),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dec56),
	.w1(32'hba85bdc9),
	.w2(32'hbad81104),
	.w3(32'hbb5f53e7),
	.w4(32'hbac7c07e),
	.w5(32'h3b3fe163),
	.w6(32'hbb4c7ca9),
	.w7(32'hba8d9cb7),
	.w8(32'h3a083cfb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04bedd),
	.w1(32'h3b298e50),
	.w2(32'h39effcbc),
	.w3(32'hbb1f99f7),
	.w4(32'hba096d4e),
	.w5(32'hbaaa36b0),
	.w6(32'hba65726e),
	.w7(32'hb8d4150b),
	.w8(32'h39e3af61),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9be77),
	.w1(32'h3b388abe),
	.w2(32'h3a0cd2c0),
	.w3(32'h3aa102c6),
	.w4(32'h3a98f149),
	.w5(32'h3b098c08),
	.w6(32'h3a761c4a),
	.w7(32'hb953f6ac),
	.w8(32'h3ad84a4b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f0a76),
	.w1(32'h3b210dac),
	.w2(32'h3b8e37b1),
	.w3(32'h3b6285bd),
	.w4(32'h3b7a0ead),
	.w5(32'hbb1df937),
	.w6(32'h3a2bccc2),
	.w7(32'h3b0280ff),
	.w8(32'hb9cc4331),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee76b4),
	.w1(32'hba858c0c),
	.w2(32'hba352662),
	.w3(32'h3987679c),
	.w4(32'h3b1a5310),
	.w5(32'h3b5c2b31),
	.w6(32'h3a8b5313),
	.w7(32'h386f3da1),
	.w8(32'h3ae4e571),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2be56d),
	.w1(32'h3a782b59),
	.w2(32'h3a441633),
	.w3(32'h3a2b017b),
	.w4(32'h3a59d73a),
	.w5(32'hba838d7b),
	.w6(32'h3a5c4822),
	.w7(32'h3b25aa3d),
	.w8(32'hbb4f1d71),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b795f),
	.w1(32'hbb4cbe58),
	.w2(32'hbbc639e5),
	.w3(32'hbbb423d3),
	.w4(32'hbbb6b142),
	.w5(32'hbb9659f0),
	.w6(32'hbafc0ecb),
	.w7(32'hbb1cad43),
	.w8(32'hbb70779f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e656),
	.w1(32'hba113da0),
	.w2(32'hbad49304),
	.w3(32'h39d0f6a1),
	.w4(32'hb98c71e8),
	.w5(32'hba164503),
	.w6(32'hbaf0935f),
	.w7(32'hbae46b43),
	.w8(32'hb9bc1b3e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88bf8f),
	.w1(32'hbb300be3),
	.w2(32'hbb8193f6),
	.w3(32'hbaf6ed5a),
	.w4(32'hbb3c887a),
	.w5(32'hbb04e2f5),
	.w6(32'hb9e37185),
	.w7(32'hbaad0af6),
	.w8(32'hba28d108),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a9bed),
	.w1(32'hbb6cfca3),
	.w2(32'hbad8d9fe),
	.w3(32'hbadf36b5),
	.w4(32'hbb1474b4),
	.w5(32'h3b37a7fc),
	.w6(32'hbb05b59c),
	.w7(32'hbb77688d),
	.w8(32'h3ae3487f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97a177),
	.w1(32'h3b0b0894),
	.w2(32'h3aca9a7a),
	.w3(32'hba3ba9d4),
	.w4(32'h3b918d03),
	.w5(32'h3a705eef),
	.w6(32'hbae187d3),
	.w7(32'h3b76572b),
	.w8(32'hba239304),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98eb316),
	.w1(32'hba53f3de),
	.w2(32'hb97d8a89),
	.w3(32'hba314a68),
	.w4(32'hb8b4f3c7),
	.w5(32'hb9cbf5d0),
	.w6(32'hbb4450d0),
	.w7(32'hba52c0c3),
	.w8(32'hbae8faca),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb262a68),
	.w1(32'hba4097c1),
	.w2(32'hbb23c5fc),
	.w3(32'hb800e307),
	.w4(32'h3b0dad6d),
	.w5(32'h3bed83f0),
	.w6(32'h3adbc484),
	.w7(32'hbb04d0a3),
	.w8(32'h3b568e33),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40c783),
	.w1(32'h3b5742ae),
	.w2(32'h3b9b1c0f),
	.w3(32'h3b6608b4),
	.w4(32'h3b121a9b),
	.w5(32'h3b032dad),
	.w6(32'h3bb66f8f),
	.w7(32'h3b92afe3),
	.w8(32'h3a926d66),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe1272),
	.w1(32'hb9911863),
	.w2(32'hbb0a297c),
	.w3(32'h3b16e953),
	.w4(32'h3b2e23d2),
	.w5(32'hba2feec2),
	.w6(32'h3b0c2a29),
	.w7(32'hb9c13249),
	.w8(32'h3a854751),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71301f),
	.w1(32'hbb082a66),
	.w2(32'h3a6d633c),
	.w3(32'h3afe4d21),
	.w4(32'h3b08ce6b),
	.w5(32'hb9cfad13),
	.w6(32'h3b4cfeb6),
	.w7(32'h3b46073a),
	.w8(32'h3ad0d742),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1fa49),
	.w1(32'h38a6ac4c),
	.w2(32'hba0136c7),
	.w3(32'h3b849809),
	.w4(32'h3b9cdb08),
	.w5(32'h3a1f56a1),
	.w6(32'h3aea948b),
	.w7(32'hb9d7ab5a),
	.w8(32'hbae2c7a2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab5c7a),
	.w1(32'hbaa6c58b),
	.w2(32'h3aee6229),
	.w3(32'hbab44197),
	.w4(32'hbaa18f71),
	.w5(32'hba6c991f),
	.w6(32'hb964ac1b),
	.w7(32'h3b33bcfd),
	.w8(32'hba91460a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9caa90e),
	.w1(32'hbb0b0754),
	.w2(32'hbb04c03b),
	.w3(32'hba692e7e),
	.w4(32'hbb05f90d),
	.w5(32'hb99fb858),
	.w6(32'hbabc76df),
	.w7(32'hbb0b7bc5),
	.w8(32'h3a4087cd),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1abfc),
	.w1(32'hbb8c8d67),
	.w2(32'hbbb35481),
	.w3(32'hbc162e12),
	.w4(32'hbbb72dd5),
	.w5(32'hbb053cb0),
	.w6(32'hbb6ca5a1),
	.w7(32'hbba1c084),
	.w8(32'hbba8e44c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab10bdb),
	.w1(32'h3a2e8457),
	.w2(32'h3b4ad33f),
	.w3(32'h3b328998),
	.w4(32'hbad958b7),
	.w5(32'h3a130e15),
	.w6(32'h395cb241),
	.w7(32'hba6d7206),
	.w8(32'hbabd7471),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36c730),
	.w1(32'hbb27a248),
	.w2(32'h38b6d73d),
	.w3(32'hbaff96d9),
	.w4(32'hb98d50ee),
	.w5(32'h39685c8a),
	.w6(32'hbb650c30),
	.w7(32'hba057725),
	.w8(32'hbb103fc1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1ea94),
	.w1(32'hbace2d5b),
	.w2(32'hba7be46e),
	.w3(32'h3adab388),
	.w4(32'h39750385),
	.w5(32'h3b82a972),
	.w6(32'hb9a3013e),
	.w7(32'hba1e0cdc),
	.w8(32'h3b5aa1c9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e91ed),
	.w1(32'hbb2e3960),
	.w2(32'hba010d93),
	.w3(32'hba8dccf1),
	.w4(32'h3b85b8ca),
	.w5(32'h3a94a1bd),
	.w6(32'h3a80d301),
	.w7(32'h3a59e4d7),
	.w8(32'hbabe95ea),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef1cee),
	.w1(32'h3b20cbd3),
	.w2(32'h3a7228d0),
	.w3(32'h3b31c4de),
	.w4(32'h3b06b882),
	.w5(32'hba7b23ce),
	.w6(32'h3b00bdc7),
	.w7(32'hb9f449db),
	.w8(32'hbb634141),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9939c6d),
	.w1(32'hba374a12),
	.w2(32'hbac104d0),
	.w3(32'hb9b3c473),
	.w4(32'h3b1c08ba),
	.w5(32'hbb75a58c),
	.w6(32'hbabb390c),
	.w7(32'hbb2b0b82),
	.w8(32'hba258c29),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef651a),
	.w1(32'h3ba280f1),
	.w2(32'h3a094ad4),
	.w3(32'h39c7bb6d),
	.w4(32'hba973e08),
	.w5(32'h3a3127ae),
	.w6(32'h3a86ba5b),
	.w7(32'h3a3faf30),
	.w8(32'hbb391a64),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a483ab),
	.w1(32'hbad99c40),
	.w2(32'hbb4c8f7e),
	.w3(32'hbb7c4ef3),
	.w4(32'hbb6183d3),
	.w5(32'hbb553507),
	.w6(32'hbab9344b),
	.w7(32'hbb4da74d),
	.w8(32'hbb8e897a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8448dc),
	.w1(32'hbaeae989),
	.w2(32'hbaef01ec),
	.w3(32'h3ad8f258),
	.w4(32'h3abf3ee5),
	.w5(32'hbb7bdc59),
	.w6(32'hbaa9d4d2),
	.w7(32'hbb348c97),
	.w8(32'hbbfd9094),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f2ae7),
	.w1(32'hbbb9d445),
	.w2(32'hbb997065),
	.w3(32'hbbf7bc3f),
	.w4(32'hbb826b43),
	.w5(32'hbb39d665),
	.w6(32'hbb1d0900),
	.w7(32'hbb6ee5d4),
	.w8(32'hbb064565),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f45fc),
	.w1(32'h3c039d6c),
	.w2(32'h3b1fcbdb),
	.w3(32'h3ba0e879),
	.w4(32'h3c01917f),
	.w5(32'h39a05b04),
	.w6(32'hba98a4e8),
	.w7(32'h3a2b7213),
	.w8(32'hbb59a89b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4b900),
	.w1(32'h3abdd80f),
	.w2(32'hbae74a26),
	.w3(32'h3a6e04bd),
	.w4(32'hba47b1f7),
	.w5(32'hbaaf063a),
	.w6(32'hbb11c6b1),
	.w7(32'hbaa53488),
	.w8(32'hbac587ae),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade37d6),
	.w1(32'hbaefbf25),
	.w2(32'hbb4cfc84),
	.w3(32'hba07662a),
	.w4(32'hb8859d5a),
	.w5(32'hbbad55e9),
	.w6(32'h39c64c93),
	.w7(32'h3a4a912d),
	.w8(32'hbbc647e6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb176aa7),
	.w1(32'hba833214),
	.w2(32'hbac79180),
	.w3(32'hbacf1424),
	.w4(32'hb9d8227a),
	.w5(32'h3b2df874),
	.w6(32'hbb48597e),
	.w7(32'hb9eaf898),
	.w8(32'h3acb37b8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb836290),
	.w1(32'hbbf9a42c),
	.w2(32'hbc02c6fb),
	.w3(32'hbbf7ac06),
	.w4(32'hbbdadd32),
	.w5(32'hbbb74140),
	.w6(32'hba3ffd73),
	.w7(32'hb9ce04e6),
	.w8(32'hbbbfb558),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11ca56),
	.w1(32'hb9f414d7),
	.w2(32'hbb400fc2),
	.w3(32'h3b1f4dd2),
	.w4(32'h396bca04),
	.w5(32'hbb4924b9),
	.w6(32'h3af506c4),
	.w7(32'h393e2dc1),
	.w8(32'hbaf2c248),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a715980),
	.w1(32'hba1a7d71),
	.w2(32'hba81145b),
	.w3(32'hba3b2a5a),
	.w4(32'h3ab9ffe9),
	.w5(32'h391995e1),
	.w6(32'hba159ceb),
	.w7(32'hb9399366),
	.w8(32'h38853cd2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee296b),
	.w1(32'h3ab03616),
	.w2(32'h2f5b3000),
	.w3(32'hb9c6fdfb),
	.w4(32'h393157e4),
	.w5(32'hba31f852),
	.w6(32'h380e52db),
	.w7(32'hba3e5e62),
	.w8(32'hba7b2db0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2dfe1),
	.w1(32'h3ac4da5e),
	.w2(32'h39853efc),
	.w3(32'h3ad1e53b),
	.w4(32'h3a09f067),
	.w5(32'h3a2fbc1a),
	.w6(32'hba1c406e),
	.w7(32'h3a1e9e74),
	.w8(32'h39c90627),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a991270),
	.w1(32'h3ad487f3),
	.w2(32'hbaad7fc5),
	.w3(32'h3b29f3a2),
	.w4(32'h3ae528f6),
	.w5(32'h38de5a68),
	.w6(32'h3b303e65),
	.w7(32'h3b17c3e2),
	.w8(32'h39c3ab76),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15419f),
	.w1(32'h3b3a4255),
	.w2(32'hba83e80a),
	.w3(32'h3b05f241),
	.w4(32'h3b1bd70c),
	.w5(32'hbb450ada),
	.w6(32'h39deab3a),
	.w7(32'h3730562a),
	.w8(32'hbb12be94),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12d5af),
	.w1(32'h386d4b0c),
	.w2(32'hba4f8668),
	.w3(32'hbb12eb04),
	.w4(32'hbaca050d),
	.w5(32'hba2ec827),
	.w6(32'hbb11e639),
	.w7(32'hbb03feaa),
	.w8(32'hbaa926cc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8b534),
	.w1(32'h3a86cf5b),
	.w2(32'h3abe7baa),
	.w3(32'h3a4f9a7d),
	.w4(32'h3adaef35),
	.w5(32'h3a82f9d9),
	.w6(32'h3a7efc8c),
	.w7(32'h3ab69646),
	.w8(32'h3aee8349),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d0f57),
	.w1(32'hba353ed4),
	.w2(32'hba807c4c),
	.w3(32'hbb2a087b),
	.w4(32'hbaabb9f8),
	.w5(32'hbb1fc239),
	.w6(32'hbb096497),
	.w7(32'hbaa5656c),
	.w8(32'hbb145fce),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9ea1c),
	.w1(32'hba959215),
	.w2(32'hba15326c),
	.w3(32'hbaa69d98),
	.w4(32'h3a44e260),
	.w5(32'hba8dbd58),
	.w6(32'hba92485e),
	.w7(32'hb92dc563),
	.w8(32'hbabf370a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f2664),
	.w1(32'hba0eca14),
	.w2(32'hba1192c5),
	.w3(32'hbb14e205),
	.w4(32'hba944fe6),
	.w5(32'h3aa27ed1),
	.w6(32'hbac1ddb5),
	.w7(32'hba1d6e23),
	.w8(32'h3a92cc61),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abed401),
	.w1(32'h3a98cabf),
	.w2(32'h3a88b7f6),
	.w3(32'h3acaacb7),
	.w4(32'h3ae82b64),
	.w5(32'h3a92d920),
	.w6(32'h3a4c264e),
	.w7(32'h3aba6685),
	.w8(32'h39c7c119),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1416ce),
	.w1(32'hba5df92d),
	.w2(32'hba0c8cf3),
	.w3(32'hbaebd90a),
	.w4(32'hbb0b3783),
	.w5(32'h3aaab8c6),
	.w6(32'h3a86132e),
	.w7(32'hb9cf13e3),
	.w8(32'h3a9624b1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00debd),
	.w1(32'hb93d9879),
	.w2(32'h3ac30d46),
	.w3(32'h3a500dd4),
	.w4(32'h3af50c94),
	.w5(32'hba4f312f),
	.w6(32'h3a29b53e),
	.w7(32'h3b06664f),
	.w8(32'hbaf80540),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e70fa),
	.w1(32'h3a40eb97),
	.w2(32'hba61132f),
	.w3(32'h3a03953e),
	.w4(32'hbab55f38),
	.w5(32'hb79d789a),
	.w6(32'hbb1e4b13),
	.w7(32'hbb1a6f7a),
	.w8(32'hb89f372b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ddb44),
	.w1(32'hba6bd671),
	.w2(32'hbac7bc40),
	.w3(32'hbae47892),
	.w4(32'hba945fd0),
	.w5(32'h3a9e51aa),
	.w6(32'hbaf05673),
	.w7(32'h38ba6aae),
	.w8(32'h3a786056),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8392c9),
	.w1(32'hba9da6b5),
	.w2(32'hb9715202),
	.w3(32'h3a2dab81),
	.w4(32'h380d3379),
	.w5(32'hba079f70),
	.w6(32'h3a401978),
	.w7(32'h3ad143d1),
	.w8(32'hbade398b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04de04),
	.w1(32'h3babdd59),
	.w2(32'h3b2063e1),
	.w3(32'h3b0a20ff),
	.w4(32'h3af1cb75),
	.w5(32'hba92f376),
	.w6(32'hba68185e),
	.w7(32'hbb02c1ab),
	.w8(32'hbb676a1b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b586ae),
	.w1(32'h39dbbd2b),
	.w2(32'h39947251),
	.w3(32'h3aa1ff83),
	.w4(32'h399617bc),
	.w5(32'h3a5b6518),
	.w6(32'h3b07bfd6),
	.w7(32'h39f36aab),
	.w8(32'hb9ead4d3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ac26e),
	.w1(32'h3a88baa9),
	.w2(32'hba263396),
	.w3(32'h39838e22),
	.w4(32'h391690a7),
	.w5(32'hbb21ecee),
	.w6(32'h399c1db4),
	.w7(32'h392c2ad8),
	.w8(32'hbadecb15),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384edd6c),
	.w1(32'hbb175819),
	.w2(32'hbae63761),
	.w3(32'hbab69809),
	.w4(32'hba3c4993),
	.w5(32'h39881fba),
	.w6(32'hba67920a),
	.w7(32'hb9ff7d25),
	.w8(32'hb9a89820),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390341d4),
	.w1(32'h3a2b26f3),
	.w2(32'hb9ea090f),
	.w3(32'h3a4a5758),
	.w4(32'h373b068a),
	.w5(32'hbaabe127),
	.w6(32'h3a326cdd),
	.w7(32'hb9b7873a),
	.w8(32'hb9febc78),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a69a4),
	.w1(32'hbaa4003a),
	.w2(32'hbad78df7),
	.w3(32'hba8ca371),
	.w4(32'hba3c5862),
	.w5(32'hba8ac359),
	.w6(32'h3a3c30cf),
	.w7(32'hba9b7af0),
	.w8(32'hb9e56bfb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9930f6e),
	.w1(32'hbb0f45e5),
	.w2(32'hba9ffc37),
	.w3(32'hbaa7af9b),
	.w4(32'hbae0e201),
	.w5(32'h3aa0723a),
	.w6(32'hb9ebd1ca),
	.w7(32'hb9d616a2),
	.w8(32'h3a1007ec),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabc53c),
	.w1(32'hba36af3c),
	.w2(32'hba5d31a2),
	.w3(32'hba973e07),
	.w4(32'hbaa93964),
	.w5(32'hb8bb55bf),
	.w6(32'h397f550d),
	.w7(32'hbaa74b39),
	.w8(32'hb8f04d10),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277221),
	.w1(32'hbad6865e),
	.w2(32'hbadccfeb),
	.w3(32'hba939859),
	.w4(32'hb8512506),
	.w5(32'h3a09456f),
	.w6(32'hbae20c0b),
	.w7(32'hb9d63c4d),
	.w8(32'h39a76ca0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1d0fc),
	.w1(32'h3a3cbd36),
	.w2(32'h39f125e8),
	.w3(32'h3992a25e),
	.w4(32'h39d81ff5),
	.w5(32'hbabb5701),
	.w6(32'h39996f47),
	.w7(32'hb934bd1b),
	.w8(32'hbae77e8e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d03e2),
	.w1(32'hbb06d2e3),
	.w2(32'hbaf800ca),
	.w3(32'hbabd0539),
	.w4(32'hba971972),
	.w5(32'h3a7df14e),
	.w6(32'hbade3bea),
	.w7(32'hbab5b5ab),
	.w8(32'h3ac42fba),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ab862),
	.w1(32'h3ac4b5f5),
	.w2(32'h3a6dc931),
	.w3(32'h39099dfc),
	.w4(32'h3a961599),
	.w5(32'h3ad9ed8a),
	.w6(32'h3a022aa0),
	.w7(32'h3a32d0e3),
	.w8(32'hb9a92b73),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52e24e),
	.w1(32'hbb98db65),
	.w2(32'hbb9caa8e),
	.w3(32'hbb7dd689),
	.w4(32'hbb25e86f),
	.w5(32'hbb08dc9d),
	.w6(32'hbb3514e8),
	.w7(32'hbb644652),
	.w8(32'hbadc032d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981357e),
	.w1(32'hbab0b1d8),
	.w2(32'hba6a1dea),
	.w3(32'hb80785e6),
	.w4(32'hb98780c3),
	.w5(32'h3a6df6a7),
	.w6(32'hbacb0b87),
	.w7(32'hb9c0d399),
	.w8(32'h3a763d4f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee837a),
	.w1(32'h3aa51d83),
	.w2(32'hbaa292df),
	.w3(32'h39bb94a1),
	.w4(32'hb985d027),
	.w5(32'hbac96147),
	.w6(32'hba2cdc5d),
	.w7(32'hba46faec),
	.w8(32'hbac5654c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c930),
	.w1(32'hbb6cf7d8),
	.w2(32'hbb7af816),
	.w3(32'hbb28cc5c),
	.w4(32'hbaffdb56),
	.w5(32'hbad5741b),
	.w6(32'hb9b7428b),
	.w7(32'hbaa49b1c),
	.w8(32'hbab13a55),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a097e09),
	.w1(32'h3ab98f48),
	.w2(32'h3a76246e),
	.w3(32'h39c3f7e4),
	.w4(32'h3aaa3ab1),
	.w5(32'h3b0d3da1),
	.w6(32'hba29e278),
	.w7(32'hb9318aa9),
	.w8(32'h3aaa067f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af106f),
	.w1(32'h3aafa49a),
	.w2(32'hba2481dc),
	.w3(32'h3b054000),
	.w4(32'h3a3cf0e3),
	.w5(32'hbb241d0a),
	.w6(32'hb9acd482),
	.w7(32'hb94a4c28),
	.w8(32'hbb520a38),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4afed2),
	.w1(32'hbb3a65d3),
	.w2(32'hbb25a55f),
	.w3(32'hbad26e77),
	.w4(32'hbabf22b5),
	.w5(32'hbb2ae1cd),
	.w6(32'hbb0dd447),
	.w7(32'hbb2ddaee),
	.w8(32'hbb35ec45),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399db7a4),
	.w1(32'h3a41daca),
	.w2(32'hba330e9a),
	.w3(32'h3ab8c69b),
	.w4(32'h392c4a70),
	.w5(32'hb9b979f6),
	.w6(32'hbae1d64b),
	.w7(32'hbabba5c8),
	.w8(32'hba394b62),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92c4dd),
	.w1(32'h3acdb6df),
	.w2(32'h39edb491),
	.w3(32'h3ad329c4),
	.w4(32'h3af3d9dd),
	.w5(32'hba07de33),
	.w6(32'h3ac372a2),
	.w7(32'h3ad587e8),
	.w8(32'hba2cd453),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53d79d),
	.w1(32'hba648414),
	.w2(32'hba8c76fd),
	.w3(32'hbabd2f35),
	.w4(32'hbb02f6c0),
	.w5(32'h3a814ee4),
	.w6(32'hb9289400),
	.w7(32'hbb1731a3),
	.w8(32'h3a7dd24e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06bb2b),
	.w1(32'h3a9e0743),
	.w2(32'h39d67696),
	.w3(32'h3a17b4b8),
	.w4(32'h3a898f64),
	.w5(32'hba0c734a),
	.w6(32'h3a99f889),
	.w7(32'h3a21fe13),
	.w8(32'hba71f6b5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e4d89),
	.w1(32'hba2f8c91),
	.w2(32'hb9c056f3),
	.w3(32'h3798d1ce),
	.w4(32'hb801d658),
	.w5(32'hbaa4d327),
	.w6(32'hb9854649),
	.w7(32'hba093247),
	.w8(32'hbad97563),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b075974),
	.w1(32'h3a36f7dd),
	.w2(32'hb9e1d5a8),
	.w3(32'h3a5ea814),
	.w4(32'h39513769),
	.w5(32'hbad9263a),
	.w6(32'hbaaa7f98),
	.w7(32'hbaad49b9),
	.w8(32'hbafb816d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba369589),
	.w1(32'hbb7b18a3),
	.w2(32'hbb2c7acf),
	.w3(32'hbaf6e378),
	.w4(32'hba88daf1),
	.w5(32'hba9b8eeb),
	.w6(32'hb9efea68),
	.w7(32'hba6b1d3e),
	.w8(32'hba7a9665),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f4172),
	.w1(32'hba80d91d),
	.w2(32'hbab87214),
	.w3(32'hba733724),
	.w4(32'hbb0f71e2),
	.w5(32'h3ad2f04b),
	.w6(32'h39d0e74a),
	.w7(32'hbb1c9640),
	.w8(32'h3aa06f05),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a42c53),
	.w1(32'hba14f9c5),
	.w2(32'hb9546448),
	.w3(32'h3ab94c85),
	.w4(32'h3a78a337),
	.w5(32'h377c7eed),
	.w6(32'hb9e4ff84),
	.w7(32'h3a86944e),
	.w8(32'h372f1591),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1297a6),
	.w1(32'h3a7e5382),
	.w2(32'hb8d7a357),
	.w3(32'h3b539cf0),
	.w4(32'h3964e664),
	.w5(32'hbb00e89d),
	.w6(32'h3adf1290),
	.w7(32'hb9626db8),
	.w8(32'hbac7af46),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33cc4f),
	.w1(32'hbb95b347),
	.w2(32'hbba62857),
	.w3(32'hbb55fe3f),
	.w4(32'hbb86abb2),
	.w5(32'hbb4e8f66),
	.w6(32'hbb4e993f),
	.w7(32'hbb7044dd),
	.w8(32'hbb1c5681),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5570d),
	.w1(32'h3b061f28),
	.w2(32'hbb254389),
	.w3(32'h3b16a218),
	.w4(32'h3ab628fd),
	.w5(32'hba091c83),
	.w6(32'h39ddd134),
	.w7(32'hba5d5a44),
	.w8(32'hba7f5c14),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4219f6),
	.w1(32'h3b40c160),
	.w2(32'h3abb992b),
	.w3(32'h3b51f487),
	.w4(32'h3b064cb3),
	.w5(32'h3a7b39c0),
	.w6(32'h3b0f1728),
	.w7(32'hb9d43736),
	.w8(32'hb92ea321),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08e6cc),
	.w1(32'h3aa32439),
	.w2(32'h3af908e7),
	.w3(32'h3b35a4a9),
	.w4(32'h3b446876),
	.w5(32'h3ae3cd39),
	.w6(32'h3b2c5c9c),
	.w7(32'h3b2d73dd),
	.w8(32'h3aeb200c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad24a29),
	.w1(32'hba64d90c),
	.w2(32'hbb277ff2),
	.w3(32'hbabafb5f),
	.w4(32'hba7ae1b0),
	.w5(32'hbb0a8212),
	.w6(32'hba6ecc7f),
	.w7(32'hb9f70cd5),
	.w8(32'hbb63f961),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba704682),
	.w1(32'hb9cbd032),
	.w2(32'h38f434a7),
	.w3(32'h3b02f437),
	.w4(32'h3a902630),
	.w5(32'h3ab40842),
	.w6(32'h391b6765),
	.w7(32'hbaad8348),
	.w8(32'hbaf81bd9),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97276f),
	.w1(32'h3af5110e),
	.w2(32'h3a331e61),
	.w3(32'h3ae0b6fa),
	.w4(32'h3aaff88f),
	.w5(32'hba8ab851),
	.w6(32'h3a96db3b),
	.w7(32'hb8d689e8),
	.w8(32'h3a56999e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392362be),
	.w1(32'hbae4b61e),
	.w2(32'hb9abef50),
	.w3(32'hbb79afce),
	.w4(32'hbb3d5d16),
	.w5(32'h394af9b1),
	.w6(32'hbabd9571),
	.w7(32'hb92570d6),
	.w8(32'h3858d734),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba638f37),
	.w1(32'h3a023f19),
	.w2(32'hbaa95cc3),
	.w3(32'h3ac23cd6),
	.w4(32'h3ac20962),
	.w5(32'hbadda5b1),
	.w6(32'h3a83f86b),
	.w7(32'h3993b927),
	.w8(32'h3a5ca3d7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa763f8),
	.w1(32'hb9a634e0),
	.w2(32'h3a8d518a),
	.w3(32'hba9bd4b0),
	.w4(32'hba16c5b0),
	.w5(32'hbaa32b8c),
	.w6(32'h39a6e4e9),
	.w7(32'hba256f68),
	.w8(32'hbb258a38),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371c0be4),
	.w1(32'hb9924ae7),
	.w2(32'hb9bd310d),
	.w3(32'hba33819a),
	.w4(32'hb9b4bb6f),
	.w5(32'h3b19ed4f),
	.w6(32'h39215247),
	.w7(32'hb9e72cf6),
	.w8(32'h3ae4db67),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb4dfb),
	.w1(32'h3b35da0e),
	.w2(32'h3ac55787),
	.w3(32'h3b247e72),
	.w4(32'h3a57396a),
	.w5(32'hba9ba127),
	.w6(32'h3b3e3803),
	.w7(32'h3ad33540),
	.w8(32'hbaa660fd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60233a),
	.w1(32'hbac850b0),
	.w2(32'hba9add3b),
	.w3(32'hbace1611),
	.w4(32'hbad6129a),
	.w5(32'h3801745a),
	.w6(32'hba89feb9),
	.w7(32'hbab40462),
	.w8(32'h3a5c696b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac467e),
	.w1(32'h3a810331),
	.w2(32'h3ad305dc),
	.w3(32'h3b80b427),
	.w4(32'hb95d5746),
	.w5(32'h3b02db42),
	.w6(32'h3b95393d),
	.w7(32'h3abd5b8f),
	.w8(32'h3ae54fdb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a3071),
	.w1(32'h3a851789),
	.w2(32'h3a5fa726),
	.w3(32'h3abb44ea),
	.w4(32'h3a974c37),
	.w5(32'hb9a686d2),
	.w6(32'h3ab373c4),
	.w7(32'h3aa30ceb),
	.w8(32'hb99cb357),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393157f6),
	.w1(32'h39cc9e1b),
	.w2(32'h39f46954),
	.w3(32'h3a2c4161),
	.w4(32'h39e7259a),
	.w5(32'hba4cc106),
	.w6(32'h3ab24201),
	.w7(32'h3aa6ab95),
	.w8(32'hba626558),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ec938),
	.w1(32'h3ac7ac79),
	.w2(32'h3a80bc3b),
	.w3(32'h3acab0e2),
	.w4(32'h3a916812),
	.w5(32'h3b0b2d5a),
	.w6(32'hb917baf7),
	.w7(32'h3b14060f),
	.w8(32'h3ab7d53a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7c857),
	.w1(32'hba94b818),
	.w2(32'hbb5600f1),
	.w3(32'hbb467b59),
	.w4(32'hbb6ec678),
	.w5(32'hba954bd9),
	.w6(32'hbbaee156),
	.w7(32'hbb8fa839),
	.w8(32'hbb46d3c5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25117e),
	.w1(32'h3afa5aa3),
	.w2(32'h3ac60c50),
	.w3(32'h3b31452e),
	.w4(32'h3adc7ac0),
	.w5(32'h3af8746f),
	.w6(32'h3b20c10e),
	.w7(32'h3ac5388f),
	.w8(32'h3aff336b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12e00e),
	.w1(32'h39932661),
	.w2(32'hba833f08),
	.w3(32'h3ad19542),
	.w4(32'h3a2f5ca5),
	.w5(32'hbab2fac4),
	.w6(32'h3abf4dd0),
	.w7(32'h3a8dd8de),
	.w8(32'hbaf36fce),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9736573),
	.w1(32'h39e73c5b),
	.w2(32'hba3244bb),
	.w3(32'hbb19d099),
	.w4(32'h38f8a47f),
	.w5(32'hba5a67a5),
	.w6(32'hba81580a),
	.w7(32'hba3fb5b1),
	.w8(32'h399e7db7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb115c5d),
	.w1(32'hba4518a1),
	.w2(32'hba477ce4),
	.w3(32'hba6a76eb),
	.w4(32'hb9f2b354),
	.w5(32'hbaf24e8a),
	.w6(32'h39fc9a46),
	.w7(32'h399f5797),
	.w8(32'hba6dd01e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f2b30),
	.w1(32'hbb0ffa0c),
	.w2(32'hbb445f5c),
	.w3(32'hbb3c1a6b),
	.w4(32'hbabc339e),
	.w5(32'hbb0f8c29),
	.w6(32'hbb2b0efb),
	.w7(32'hbb071abf),
	.w8(32'hbb3ce570),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb751019),
	.w1(32'hbaa8dc7e),
	.w2(32'hbb1fa859),
	.w3(32'hbb2a7ff2),
	.w4(32'hba198c6b),
	.w5(32'h3a277739),
	.w6(32'hbb0a749e),
	.w7(32'hbacca03e),
	.w8(32'hb72ae53b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6701c),
	.w1(32'h3a9ed567),
	.w2(32'h3abecde8),
	.w3(32'h3b30bffe),
	.w4(32'h3b293617),
	.w5(32'h3a9b31ec),
	.w6(32'h3aeea88d),
	.w7(32'h3b4ed6e1),
	.w8(32'h3ab46ae2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79f0dd),
	.w1(32'hb9840eb7),
	.w2(32'hb9749167),
	.w3(32'hba578d07),
	.w4(32'hb9e761c9),
	.w5(32'h3b05c261),
	.w6(32'hba67f86c),
	.w7(32'h39ad2a16),
	.w8(32'h3aa41065),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc153f),
	.w1(32'h3a8a650b),
	.w2(32'h3ac4888e),
	.w3(32'h3b376993),
	.w4(32'h3b060602),
	.w5(32'hba197728),
	.w6(32'h3ab54baa),
	.w7(32'h3b01143e),
	.w8(32'hb78e37cf),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9265f8),
	.w1(32'h3a735518),
	.w2(32'hb9598361),
	.w3(32'hba53a95b),
	.w4(32'hb8eeb986),
	.w5(32'h39bd02d6),
	.w6(32'h36335c79),
	.w7(32'hb91b25a6),
	.w8(32'h3984ccb9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba873310),
	.w1(32'hbaa3fcc3),
	.w2(32'hb7846e3d),
	.w3(32'hbaf24437),
	.w4(32'hba9116af),
	.w5(32'h3aa26f44),
	.w6(32'hba7448ef),
	.w7(32'hba16c52d),
	.w8(32'h39b05e05),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee5b7a),
	.w1(32'hba1db6c7),
	.w2(32'hba9ed10a),
	.w3(32'hba6920c3),
	.w4(32'hba8bdefc),
	.w5(32'hba80f0a7),
	.w6(32'hbb175c40),
	.w7(32'hbb14e5f8),
	.w8(32'hba015096),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45843b),
	.w1(32'h3a9ed76a),
	.w2(32'h3a880178),
	.w3(32'h3b2f3954),
	.w4(32'hba711202),
	.w5(32'hbadf501a),
	.w6(32'h3b4f0dd4),
	.w7(32'h393f3a79),
	.w8(32'hbae1d54e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8eb5be),
	.w1(32'hbb2333cc),
	.w2(32'hbafac451),
	.w3(32'hbae1d3a5),
	.w4(32'hba3daea7),
	.w5(32'h3a76621a),
	.w6(32'hba6db5ee),
	.w7(32'hba3ce96e),
	.w8(32'hb80e9284),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cdd16),
	.w1(32'h3ab5dfc6),
	.w2(32'hb9ca174a),
	.w3(32'h3a04763b),
	.w4(32'hb9c68cd3),
	.w5(32'h3a6672f3),
	.w6(32'h3a11ac3f),
	.w7(32'hbaaf0b07),
	.w8(32'hb9beada2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c36768),
	.w1(32'h390396c2),
	.w2(32'hbac86525),
	.w3(32'h3b09e96b),
	.w4(32'hb8b74ae1),
	.w5(32'hb96a36a1),
	.w6(32'h3b007de3),
	.w7(32'hbb026546),
	.w8(32'hbb2edb02),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36583328),
	.w1(32'hba163c2d),
	.w2(32'h38b4ce70),
	.w3(32'hbaf18a92),
	.w4(32'hb91bd811),
	.w5(32'h3ad71bd5),
	.w6(32'hba190c12),
	.w7(32'hb9d7d2c4),
	.w8(32'h39b150af),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e374e),
	.w1(32'h39f3c878),
	.w2(32'h3a2f20ff),
	.w3(32'h3b094bdd),
	.w4(32'h3ae49b5a),
	.w5(32'hba742385),
	.w6(32'h3aef961b),
	.w7(32'h3ab2340c),
	.w8(32'hba166678),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2105a),
	.w1(32'hbc01bdda),
	.w2(32'hbbcad05a),
	.w3(32'hbb1f6138),
	.w4(32'hbab999d8),
	.w5(32'hbb4d9b5a),
	.w6(32'hbb0619f6),
	.w7(32'h391e6f5e),
	.w8(32'hba177912),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efdd3a),
	.w1(32'h3b293d4f),
	.w2(32'h396e5372),
	.w3(32'h3b6cce92),
	.w4(32'h3b8ca935),
	.w5(32'hbad58810),
	.w6(32'h3901193a),
	.w7(32'h3b24cbd5),
	.w8(32'hbb878e18),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c6a05d),
	.w1(32'hb98424e4),
	.w2(32'hba59af24),
	.w3(32'hba13036d),
	.w4(32'hb968a921),
	.w5(32'hb97cc029),
	.w6(32'hb975fa07),
	.w7(32'hba513580),
	.w8(32'h3949a335),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa89905),
	.w1(32'hba74c862),
	.w2(32'hbab9a925),
	.w3(32'hb960f5c2),
	.w4(32'hba9ca576),
	.w5(32'h3ad8f797),
	.w6(32'h3a183955),
	.w7(32'hb9dd8302),
	.w8(32'h39cd2fc7),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80ed12f),
	.w1(32'h3aaf7030),
	.w2(32'h3a0adfa2),
	.w3(32'h3aa48e88),
	.w4(32'hba20002b),
	.w5(32'h3b10acce),
	.w6(32'h3b42e107),
	.w7(32'h399971be),
	.w8(32'h3aaae35c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e30378),
	.w1(32'h3a0bc2de),
	.w2(32'h39dbac2c),
	.w3(32'h3a53e5fe),
	.w4(32'hb93a6ec2),
	.w5(32'h3a954359),
	.w6(32'h3aee3cc8),
	.w7(32'h3970c648),
	.w8(32'h395c4511),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a055bef),
	.w1(32'h393100bc),
	.w2(32'hbabb8e08),
	.w3(32'h3a94cd0a),
	.w4(32'h39b61193),
	.w5(32'hba81b9d7),
	.w6(32'h39644325),
	.w7(32'hb9e2bcc2),
	.w8(32'h37b52557),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2ca1d),
	.w1(32'hba8bfcf6),
	.w2(32'hbad26295),
	.w3(32'h3a18063e),
	.w4(32'hb9e65533),
	.w5(32'hba4168d4),
	.w6(32'h39838e9b),
	.w7(32'hba121e22),
	.w8(32'hbaa5e86c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88cb21),
	.w1(32'h3a74b21a),
	.w2(32'h3a8e2b79),
	.w3(32'h3a61b003),
	.w4(32'h3a60fb97),
	.w5(32'h3a3c8710),
	.w6(32'h3a1d9034),
	.w7(32'h3a94b8d1),
	.w8(32'h3aaedb8f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a827d7f),
	.w1(32'hbaea0b08),
	.w2(32'hba3927c1),
	.w3(32'hbaa825ab),
	.w4(32'hba99bc50),
	.w5(32'hba182207),
	.w6(32'hba0fb828),
	.w7(32'hbad0f5c3),
	.w8(32'hba4981c6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395fdae0),
	.w1(32'h3a489bfb),
	.w2(32'hbaec947b),
	.w3(32'h394c1535),
	.w4(32'h3a807363),
	.w5(32'hbab206cd),
	.w6(32'h39306683),
	.w7(32'hb97123dd),
	.w8(32'hb8bf1650),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0353f6),
	.w1(32'hb99c3cb7),
	.w2(32'h395f0004),
	.w3(32'h392a5fa0),
	.w4(32'hba13f9dd),
	.w5(32'hbac3cb56),
	.w6(32'h39c57625),
	.w7(32'h3a826e5a),
	.w8(32'hba95ff05),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ded6c),
	.w1(32'hb9b4fc12),
	.w2(32'hba833957),
	.w3(32'hba4fa5c3),
	.w4(32'hbaba1183),
	.w5(32'hba3ae161),
	.w6(32'hb8a9ba99),
	.w7(32'hbaf5d130),
	.w8(32'hba3c4ab5),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb0e88),
	.w1(32'hbaf89359),
	.w2(32'hba3d64b3),
	.w3(32'hba5a32bd),
	.w4(32'hb9ae03f2),
	.w5(32'h393da7ae),
	.w6(32'hb9ad86e5),
	.w7(32'h3ab1a992),
	.w8(32'hba9398b2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38326c06),
	.w1(32'hba78b60e),
	.w2(32'hbaa761a7),
	.w3(32'hba1df4ae),
	.w4(32'hbb1ef3b5),
	.w5(32'h394b99d3),
	.w6(32'h3a124c14),
	.w7(32'hbad84a42),
	.w8(32'h3a023363),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb6048),
	.w1(32'h3a4d4818),
	.w2(32'hb8f0bbc6),
	.w3(32'h3a34c8b8),
	.w4(32'h3a98a55b),
	.w5(32'hbb30ce35),
	.w6(32'h3ae4cea9),
	.w7(32'h3aaeeba4),
	.w8(32'hbb54f6e4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45fded),
	.w1(32'hb9a274df),
	.w2(32'hba8bb64a),
	.w3(32'h3aaa4c22),
	.w4(32'h37c2ff74),
	.w5(32'h3af344c3),
	.w6(32'hbb185ac8),
	.w7(32'hbb506b70),
	.w8(32'h3a59febf),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09c8d8),
	.w1(32'h3b01c2ca),
	.w2(32'hb946991b),
	.w3(32'h3b102976),
	.w4(32'h3a78c2bf),
	.w5(32'hbac7c379),
	.w6(32'h3a75b7c3),
	.w7(32'h395b83da),
	.w8(32'hbb055862),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3815fac1),
	.w1(32'hb9f2f4f5),
	.w2(32'h3a403994),
	.w3(32'hba31d1b4),
	.w4(32'h3a6fcd7b),
	.w5(32'hba30e1b4),
	.w6(32'hb9d637c8),
	.w7(32'h39f282c1),
	.w8(32'hba987af8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94dfdb6),
	.w1(32'h398e86ea),
	.w2(32'hbabbe9f4),
	.w3(32'h39e279f0),
	.w4(32'h39803f99),
	.w5(32'hb9065362),
	.w6(32'hbb198307),
	.w7(32'hba3cf962),
	.w8(32'h396cec88),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e5f9b),
	.w1(32'hb973573d),
	.w2(32'hba481e68),
	.w3(32'hbaa3480b),
	.w4(32'hba78d9a0),
	.w5(32'hbac76f8a),
	.w6(32'h39bd9ade),
	.w7(32'hb8a858a4),
	.w8(32'hbafdbe26),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8c545),
	.w1(32'hbba28601),
	.w2(32'hbb8efd53),
	.w3(32'hbb35416e),
	.w4(32'hbb47b0ef),
	.w5(32'hbb179a90),
	.w6(32'hbb584038),
	.w7(32'hbb392402),
	.w8(32'hbafb1fa0),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ebe160),
	.w1(32'hba9e1478),
	.w2(32'hba9e018a),
	.w3(32'hba9e2f89),
	.w4(32'hba7bf535),
	.w5(32'hba6d59cf),
	.w6(32'hbab21fef),
	.w7(32'hbaaef85a),
	.w8(32'h399c6dc7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d977f8),
	.w1(32'hb9a49ab0),
	.w2(32'hb91edd1c),
	.w3(32'hbab07ff9),
	.w4(32'hbab84218),
	.w5(32'h3a835cc3),
	.w6(32'hba081a48),
	.w7(32'hbabf9e90),
	.w8(32'h3a62738b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af51424),
	.w1(32'h3ade6e6b),
	.w2(32'h3a4fbbcc),
	.w3(32'h3b54f6d5),
	.w4(32'h3acebf7a),
	.w5(32'h392c97fc),
	.w6(32'h3ac9dd5d),
	.w7(32'h39ff3d4e),
	.w8(32'hb9a25cec),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad32145),
	.w1(32'hbb4aa5d3),
	.w2(32'hbb7e76b3),
	.w3(32'hbaadcbd5),
	.w4(32'hbaf612a9),
	.w5(32'hbae17a65),
	.w6(32'hbb7509c7),
	.w7(32'hbb61fae3),
	.w8(32'hbb831659),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978a5c3),
	.w1(32'h3a72dd1b),
	.w2(32'hba61a0a2),
	.w3(32'h3a26da9b),
	.w4(32'h3a0f8003),
	.w5(32'hb9cb7b0f),
	.w6(32'hba61c6d8),
	.w7(32'hb9b64724),
	.w8(32'hba04782c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a870e11),
	.w1(32'h3a8cc21f),
	.w2(32'h38c050da),
	.w3(32'h3a775ed8),
	.w4(32'h3b11c77d),
	.w5(32'hb70a9de4),
	.w6(32'h3a11e95f),
	.w7(32'hb99a2c0e),
	.w8(32'hba0d6211),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa967c1),
	.w1(32'hb9e324b1),
	.w2(32'hb98b94fe),
	.w3(32'hb9cd2694),
	.w4(32'h397e72b8),
	.w5(32'h3aa52f3a),
	.w6(32'h39d93ce8),
	.w7(32'h3a270450),
	.w8(32'h3a9e5418),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a05a9),
	.w1(32'h3a033213),
	.w2(32'h388a0d00),
	.w3(32'hb9f4828c),
	.w4(32'h381baf8f),
	.w5(32'hb969fa8e),
	.w6(32'h39a1f02d),
	.w7(32'hba09f6da),
	.w8(32'hbaa6f9d0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea7f4e),
	.w1(32'h3ab5a501),
	.w2(32'hbb073859),
	.w3(32'hba60390f),
	.w4(32'hbaeff001),
	.w5(32'hbae004bb),
	.w6(32'h37b11714),
	.w7(32'hbaaa5a63),
	.w8(32'hb615b48c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c1d42),
	.w1(32'hbbbeecdd),
	.w2(32'hbb4c96a3),
	.w3(32'hbb5fe189),
	.w4(32'hbb4fa9a0),
	.w5(32'hba7fc8ad),
	.w6(32'h3a2c4754),
	.w7(32'hb9dcf3f2),
	.w8(32'h3a02434b),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed9c48),
	.w1(32'hbaf6c8fb),
	.w2(32'hbac047b4),
	.w3(32'hba9355d7),
	.w4(32'hbb282059),
	.w5(32'hb9a82195),
	.w6(32'hbafc1d16),
	.w7(32'hbade1bcf),
	.w8(32'h3a024dcc),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7dd915),
	.w1(32'h3b16b4a2),
	.w2(32'h39972c21),
	.w3(32'h3ab2e3eb),
	.w4(32'h3b15ab25),
	.w5(32'h3aab4d16),
	.w6(32'h3a8b7954),
	.w7(32'h39102bf6),
	.w8(32'hb5079394),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b98dc),
	.w1(32'h3aa8ff22),
	.w2(32'h38ee73e6),
	.w3(32'h3aa0a66c),
	.w4(32'h3aad04e1),
	.w5(32'hba1bc2ad),
	.w6(32'hb9637467),
	.w7(32'h39c5a0bb),
	.w8(32'hbab8908d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1667fe),
	.w1(32'hba45b7d9),
	.w2(32'hba347b49),
	.w3(32'hba32ad6f),
	.w4(32'hbae2694d),
	.w5(32'h3af20fed),
	.w6(32'hb932ba6e),
	.w7(32'hbaac121b),
	.w8(32'h3b018c66),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b5d78),
	.w1(32'h39346913),
	.w2(32'h39a978f4),
	.w3(32'h389eed45),
	.w4(32'h3ac7c434),
	.w5(32'hba61ea55),
	.w6(32'h3a319399),
	.w7(32'h3a5716a4),
	.w8(32'hbad2b5c6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb9cc2),
	.w1(32'hba8f3394),
	.w2(32'hb6271ffa),
	.w3(32'hba25e66f),
	.w4(32'hba923737),
	.w5(32'h3a1f221b),
	.w6(32'hbab32a9a),
	.w7(32'hba80684b),
	.w8(32'h3b08cd7d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3f8bd),
	.w1(32'h3a191110),
	.w2(32'h399f5ec8),
	.w3(32'h3a0a8554),
	.w4(32'hba749ac5),
	.w5(32'h3abfc431),
	.w6(32'h3af0b738),
	.w7(32'hb9e0d884),
	.w8(32'hb74551b7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b350620),
	.w1(32'hbb7e66ac),
	.w2(32'h3b0a9d07),
	.w3(32'h3a2a03fc),
	.w4(32'h3ba995f8),
	.w5(32'hbbda7f93),
	.w6(32'hbc2439fd),
	.w7(32'hbacbda3a),
	.w8(32'hbbe3d619),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d6139),
	.w1(32'hbc64f024),
	.w2(32'hbc6517f4),
	.w3(32'hbc2d71d9),
	.w4(32'hbc3ca187),
	.w5(32'hbaca6e40),
	.w6(32'hbc15031d),
	.w7(32'hbc86e418),
	.w8(32'h38aa354e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be80e4b),
	.w1(32'h39f2faf8),
	.w2(32'hbb6558be),
	.w3(32'hb856a6ce),
	.w4(32'hbae92e6d),
	.w5(32'h3ad31a4a),
	.w6(32'hbb98b1bd),
	.w7(32'hbb20bd5d),
	.w8(32'hb9d522c3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a933b94),
	.w1(32'h3b0b35c3),
	.w2(32'hb9e09e0d),
	.w3(32'h3aed9e65),
	.w4(32'h3b1a93b0),
	.w5(32'hba8e5c99),
	.w6(32'hba33877a),
	.w7(32'h3b669eba),
	.w8(32'h3ad1cf10),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4a9f),
	.w1(32'hbb918a5d),
	.w2(32'hbc0075c8),
	.w3(32'hbae52332),
	.w4(32'hbbb05943),
	.w5(32'h3c542863),
	.w6(32'hbb7201f4),
	.w7(32'hbb9e2e88),
	.w8(32'h3c887db1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7311c3),
	.w1(32'h3c621d62),
	.w2(32'h3c0f6feb),
	.w3(32'h3c91288a),
	.w4(32'h3c45fc24),
	.w5(32'h3b44ddd2),
	.w6(32'hbc0d287d),
	.w7(32'h3c786057),
	.w8(32'hbb996e0e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba08519),
	.w1(32'h3baedd2e),
	.w2(32'h3b8dd9b2),
	.w3(32'h3c6ad693),
	.w4(32'h3ab0204e),
	.w5(32'hbb969d33),
	.w6(32'h3cdfdbb3),
	.w7(32'h3c2fb9bb),
	.w8(32'hbac28c6a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc43395),
	.w1(32'hbaad6693),
	.w2(32'hba161408),
	.w3(32'hbbf84fc9),
	.w4(32'hbbced9c7),
	.w5(32'hbc8023cd),
	.w6(32'h3c437d92),
	.w7(32'h3b395acb),
	.w8(32'hbc3d5f1a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2241a7),
	.w1(32'h3b90dc11),
	.w2(32'hbb565d1a),
	.w3(32'hbc5e5ffd),
	.w4(32'hbae9816d),
	.w5(32'h390a70ff),
	.w6(32'hbbd47b37),
	.w7(32'h3b954db9),
	.w8(32'hbbbc3ee1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77d0f58),
	.w1(32'hbaa14899),
	.w2(32'hbacc35e8),
	.w3(32'hbc2f8b5d),
	.w4(32'hbba408c7),
	.w5(32'hbc132c9c),
	.w6(32'h3bb29a3c),
	.w7(32'hbb594b9e),
	.w8(32'hbc4cc1de),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeba7cd),
	.w1(32'hbcaaf804),
	.w2(32'hbc0905f1),
	.w3(32'hbc185227),
	.w4(32'h3ae5a6c6),
	.w5(32'h3ab5363f),
	.w6(32'hbca5ef85),
	.w7(32'hbc10e759),
	.w8(32'hbaa52376),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a893360),
	.w1(32'hbbb6d5f1),
	.w2(32'hbb3afc66),
	.w3(32'hbbaf8247),
	.w4(32'hbb5c681d),
	.w5(32'hbb9fb591),
	.w6(32'hbb1ad28d),
	.w7(32'hbbada5ca),
	.w8(32'hbc46fc66),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fc0d7),
	.w1(32'hbc7e7ad4),
	.w2(32'hbc5d1e32),
	.w3(32'hbc6a0938),
	.w4(32'hbbd0b160),
	.w5(32'hbb95b352),
	.w6(32'hbcaa7d6a),
	.w7(32'hbc9b4a7d),
	.w8(32'h3a7d90b5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e22dc1),
	.w1(32'hbbb21a40),
	.w2(32'hbaa8a7cf),
	.w3(32'hbbb347a4),
	.w4(32'hbb799c0f),
	.w5(32'hbc55ec5f),
	.w6(32'hbaa53cc3),
	.w7(32'hb92a7794),
	.w8(32'hbc2cf089),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9851d8),
	.w1(32'hbc2131de),
	.w2(32'hbc0dfe80),
	.w3(32'hbc5e9b0b),
	.w4(32'hbc6c88f5),
	.w5(32'hbb928ece),
	.w6(32'h3c0c9f2c),
	.w7(32'hbbd8147f),
	.w8(32'hba9fdb58),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9743896),
	.w1(32'hba69cab2),
	.w2(32'hbb33a961),
	.w3(32'hb9ac227b),
	.w4(32'hbad81b57),
	.w5(32'h3bd2667e),
	.w6(32'hbbb08526),
	.w7(32'h3994189d),
	.w8(32'h3d146f6a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c491696),
	.w1(32'h3d13bf15),
	.w2(32'h3c256e9c),
	.w3(32'h3b9e5e96),
	.w4(32'h3baf3aea),
	.w5(32'hbb8d3809),
	.w6(32'h3c533b42),
	.w7(32'hb9be1deb),
	.w8(32'h3a089a2e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ef0a1),
	.w1(32'hbb2ac0d4),
	.w2(32'hbaecb203),
	.w3(32'hbb8c7ee1),
	.w4(32'hbb37acf7),
	.w5(32'hbbdffc1c),
	.w6(32'h3bb2caee),
	.w7(32'h38ddda3b),
	.w8(32'hbb79776f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd5968),
	.w1(32'hbbaf6ddc),
	.w2(32'hbb2f727a),
	.w3(32'hbc227a9a),
	.w4(32'hbb901f1a),
	.w5(32'h3b79ccff),
	.w6(32'hbc035b6e),
	.w7(32'h39a3d946),
	.w8(32'hbc2bb073),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bece626),
	.w1(32'hbc0618e6),
	.w2(32'h3ba79bdf),
	.w3(32'h3cd81746),
	.w4(32'h3c2279dc),
	.w5(32'h3b5dd594),
	.w6(32'h3c855558),
	.w7(32'h3c98ae19),
	.w8(32'h3b89646e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a9897),
	.w1(32'h3bb5a82f),
	.w2(32'h3c1f89b3),
	.w3(32'h3bbf2aed),
	.w4(32'h3c2ef033),
	.w5(32'h3caef0fb),
	.w6(32'hbb757dd1),
	.w7(32'h3be902c1),
	.w8(32'h3cf432bb),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce8f1ed),
	.w1(32'h3c8f0d06),
	.w2(32'h3ca31ffb),
	.w3(32'h3ce47945),
	.w4(32'h3d132559),
	.w5(32'hbb082aff),
	.w6(32'hbc20df8d),
	.w7(32'h3cfb4473),
	.w8(32'hb995d953),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea3e72),
	.w1(32'h3b7a293d),
	.w2(32'hb99a967b),
	.w3(32'h3bfa7418),
	.w4(32'h3b6d996b),
	.w5(32'h3a86b6f0),
	.w6(32'h3c088392),
	.w7(32'h3c081b2e),
	.w8(32'hbbc47643),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b954d56),
	.w1(32'hbbbb23df),
	.w2(32'hbaf14a89),
	.w3(32'hba06d693),
	.w4(32'h3b65ecee),
	.w5(32'hbc351366),
	.w6(32'h3b595e75),
	.w7(32'h3b034c20),
	.w8(32'hb86954a2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c71a),
	.w1(32'h3c0cc7e6),
	.w2(32'hbb2269b8),
	.w3(32'hbb94c404),
	.w4(32'hbb64653f),
	.w5(32'h3bbb61a6),
	.w6(32'h3bf52dba),
	.w7(32'hbba683f4),
	.w8(32'hbae6b7b1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f1ac),
	.w1(32'hbad7f0a3),
	.w2(32'hbbb7ab05),
	.w3(32'hbc027083),
	.w4(32'hbb7efb58),
	.w5(32'hbb801172),
	.w6(32'h3c7290fe),
	.w7(32'hbc0dc503),
	.w8(32'h3acf240a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cefb5),
	.w1(32'h3b878d0d),
	.w2(32'hba843d23),
	.w3(32'hb9c754d7),
	.w4(32'h3b6abd35),
	.w5(32'h3b2fb245),
	.w6(32'hb966414f),
	.w7(32'hbbb18809),
	.w8(32'hbbb577e9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0225b),
	.w1(32'hbb8c9937),
	.w2(32'h3b27170d),
	.w3(32'hbb50b590),
	.w4(32'hbadf459e),
	.w5(32'h3a95a3dd),
	.w6(32'hbbff34be),
	.w7(32'h3bdfcf3e),
	.w8(32'hbb5a6da2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6a7f4),
	.w1(32'h3b3a466d),
	.w2(32'h3b996c79),
	.w3(32'hbbccc4c2),
	.w4(32'h3aa516b5),
	.w5(32'hbbf5e9b1),
	.w6(32'h3c57037c),
	.w7(32'hba1375f1),
	.w8(32'h3a9299f9),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2658c),
	.w1(32'hbb89783a),
	.w2(32'hbbb90008),
	.w3(32'h38ebbda2),
	.w4(32'hbb5d909e),
	.w5(32'hbbc4331a),
	.w6(32'hbb81e853),
	.w7(32'h3b497d5c),
	.w8(32'hbc320644),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule