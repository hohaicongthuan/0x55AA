module layer_10_featuremap_14(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba8cff),
	.w1(32'h3c880353),
	.w2(32'h3bd79fcc),
	.w3(32'hbb88e01c),
	.w4(32'h3bf7f121),
	.w5(32'h3bdb7c5c),
	.w6(32'h3ac705ce),
	.w7(32'h3b33b090),
	.w8(32'h3c918789),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51feb2),
	.w1(32'h3c013fcf),
	.w2(32'h3c09f909),
	.w3(32'h3ced7abd),
	.w4(32'h3c880c61),
	.w5(32'h3b3b3141),
	.w6(32'h3c86b99e),
	.w7(32'h3bbad282),
	.w8(32'hbb9ca4e4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7181ff),
	.w1(32'h3a316bb9),
	.w2(32'h3c692b60),
	.w3(32'h3c147ce2),
	.w4(32'h3c12ee0b),
	.w5(32'h3c8eaafd),
	.w6(32'hb93d1345),
	.w7(32'hbc42ce61),
	.w8(32'h3c83e46a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80a859),
	.w1(32'hbc93b624),
	.w2(32'hbc137301),
	.w3(32'hbb4bf233),
	.w4(32'hbcab4005),
	.w5(32'hb99ac358),
	.w6(32'h3bb33543),
	.w7(32'hbc8c74b5),
	.w8(32'hbc0bfa16),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d70ca),
	.w1(32'h3c54979b),
	.w2(32'h3a801786),
	.w3(32'h3b84656c),
	.w4(32'h3c86ef15),
	.w5(32'h3ae00910),
	.w6(32'h3b56dbd0),
	.w7(32'h3c34e8e9),
	.w8(32'hbb35f05e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b3af3),
	.w1(32'hbb844903),
	.w2(32'h39b13bda),
	.w3(32'hbc170e07),
	.w4(32'hbc04346b),
	.w5(32'hba497212),
	.w6(32'hbb28fccc),
	.w7(32'hbb79e9d6),
	.w8(32'h3a0c93c1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b29762),
	.w1(32'hbaa20068),
	.w2(32'h3b852475),
	.w3(32'h3aa4ba18),
	.w4(32'h3b0cea00),
	.w5(32'hb9c3416f),
	.w6(32'hbb145b2a),
	.w7(32'h3b005cd9),
	.w8(32'hbc11fc44),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beaf220),
	.w1(32'h3c1924a3),
	.w2(32'h3c013226),
	.w3(32'h3b4a9842),
	.w4(32'h3aa4fae2),
	.w5(32'h3affa661),
	.w6(32'hbb641083),
	.w7(32'hbab8584a),
	.w8(32'h377cfee2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f152c),
	.w1(32'h3b94cc24),
	.w2(32'h3bc641b6),
	.w3(32'h3b58045c),
	.w4(32'h3c089078),
	.w5(32'h3c104b59),
	.w6(32'hbb7c6b79),
	.w7(32'h3b608f5c),
	.w8(32'h3c49e861),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e750b),
	.w1(32'hbb08c73a),
	.w2(32'h3b88cb36),
	.w3(32'h3ad6988e),
	.w4(32'hbacc6b1b),
	.w5(32'h3b98e52b),
	.w6(32'h3c07cbf0),
	.w7(32'hbb344e23),
	.w8(32'h3ba15fef),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46db20),
	.w1(32'h3afd1b8e),
	.w2(32'h3bdb431b),
	.w3(32'h3acdaed1),
	.w4(32'h3a563ba0),
	.w5(32'h3c7bd90f),
	.w6(32'h3ae83ee4),
	.w7(32'h3b0f3e84),
	.w8(32'h3ca644a5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80cee3),
	.w1(32'hbbf4e6c7),
	.w2(32'h3ad96168),
	.w3(32'h3b86b38c),
	.w4(32'hbcc34970),
	.w5(32'h3b8bc4df),
	.w6(32'h3c14bd86),
	.w7(32'hbcd5365e),
	.w8(32'h3a62420c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81a35e),
	.w1(32'h3ba0e372),
	.w2(32'h3bbd25e6),
	.w3(32'hba1bc838),
	.w4(32'h3b30dfc8),
	.w5(32'h3c31c003),
	.w6(32'hbaf17251),
	.w7(32'hb9779d07),
	.w8(32'h3b0b6c85),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b783a32),
	.w1(32'h3c208554),
	.w2(32'hbb9f222d),
	.w3(32'h3c281c3f),
	.w4(32'h3bdf1dd6),
	.w5(32'hbbe46b7c),
	.w6(32'hbb083e27),
	.w7(32'h3bb162ed),
	.w8(32'hbc04056e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88414c),
	.w1(32'h3bd239c3),
	.w2(32'hbb56f0c3),
	.w3(32'hba759425),
	.w4(32'h3c1702ec),
	.w5(32'hba94b15e),
	.w6(32'h3b1564ca),
	.w7(32'h3c1ce7f3),
	.w8(32'h3a38f885),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98211c),
	.w1(32'hb925320e),
	.w2(32'h3b7fe074),
	.w3(32'hba4c1fff),
	.w4(32'hbb148315),
	.w5(32'h3b8b6327),
	.w6(32'h3b552825),
	.w7(32'h3abb92f4),
	.w8(32'h3ba12376),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9617965),
	.w1(32'h3ab67b60),
	.w2(32'h3a28348d),
	.w3(32'h3a97c710),
	.w4(32'h3a8f22cf),
	.w5(32'hbb19b71f),
	.w6(32'h3a2125eb),
	.w7(32'h3b1358aa),
	.w8(32'h3b0987f9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac20a85),
	.w1(32'h3bd8a124),
	.w2(32'h3c69d4fa),
	.w3(32'h3a560d73),
	.w4(32'h3ad49fb7),
	.w5(32'h3c154ab9),
	.w6(32'hbb47efb1),
	.w7(32'hbb36e3f5),
	.w8(32'h3c2d880a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9890f),
	.w1(32'h3c13ad1d),
	.w2(32'h3c8682e6),
	.w3(32'h3c0a7a1c),
	.w4(32'h3b56ef94),
	.w5(32'h3b6576c6),
	.w6(32'h3bbfd17c),
	.w7(32'hba36916e),
	.w8(32'h3b16f035),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57911f),
	.w1(32'hba5273fa),
	.w2(32'h3aa8f335),
	.w3(32'h3c01be44),
	.w4(32'hb98b7056),
	.w5(32'hbabf86d2),
	.w6(32'hbc1502af),
	.w7(32'hbbd821c9),
	.w8(32'h3ae9d590),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd106e),
	.w1(32'h3b460ecd),
	.w2(32'hbaf02667),
	.w3(32'h3b867973),
	.w4(32'h3b295b34),
	.w5(32'hbbab84fd),
	.w6(32'h3b92f57e),
	.w7(32'h3b35c148),
	.w8(32'h3b2e920f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7ba92),
	.w1(32'hbc9c1dc7),
	.w2(32'h3b826919),
	.w3(32'h3a6fe721),
	.w4(32'hbc239e60),
	.w5(32'h384a74e8),
	.w6(32'hbbb68629),
	.w7(32'hbbdc1ea0),
	.w8(32'hbb5cf85c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc00911),
	.w1(32'h3b8bf1ee),
	.w2(32'h3bbbd90f),
	.w3(32'h3bb16b58),
	.w4(32'hbb4af355),
	.w5(32'h3bd923ac),
	.w6(32'hbb89202a),
	.w7(32'hbbc793c2),
	.w8(32'h3c02d5e3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952b1a2),
	.w1(32'hba7da901),
	.w2(32'h3af80d6a),
	.w3(32'hbad6b723),
	.w4(32'hbb35d42d),
	.w5(32'hbaad21b0),
	.w6(32'hbb437d3c),
	.w7(32'hbb1a4d16),
	.w8(32'hb9bf2e35),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c4cf4),
	.w1(32'h3c3b1bb2),
	.w2(32'h3bd1ca0a),
	.w3(32'h3a8a640e),
	.w4(32'h3ba4fdd5),
	.w5(32'h3bdd227f),
	.w6(32'h3bd99cd6),
	.w7(32'h3b6002d7),
	.w8(32'h3c059668),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04a365),
	.w1(32'hbc313198),
	.w2(32'hbc219553),
	.w3(32'h3c42827f),
	.w4(32'hb9bb6506),
	.w5(32'hbc3565be),
	.w6(32'hb888c8d5),
	.w7(32'hbbf9e080),
	.w8(32'hbc8eaa5f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41089e),
	.w1(32'h3cc670e4),
	.w2(32'h39dbc969),
	.w3(32'hbba24df5),
	.w4(32'h3ceab7bc),
	.w5(32'h3ab0771b),
	.w6(32'hbc2438bd),
	.w7(32'h3cbad848),
	.w8(32'h383017aa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba72057),
	.w1(32'hbb5f16ab),
	.w2(32'hbb9464d0),
	.w3(32'hbb104915),
	.w4(32'h36f20e05),
	.w5(32'hbbcb4c64),
	.w6(32'hba8ffa77),
	.w7(32'hba9988f0),
	.w8(32'hbba224ac),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72a7f1),
	.w1(32'h3b2e18b7),
	.w2(32'h3a5a7263),
	.w3(32'hba1c657f),
	.w4(32'h3b174599),
	.w5(32'h3c47ae8b),
	.w6(32'h3a8b57e1),
	.w7(32'h3b8eb779),
	.w8(32'hbbc24943),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b87b0),
	.w1(32'hbc4679c6),
	.w2(32'hbbe8d115),
	.w3(32'h3ba87a02),
	.w4(32'hbca37fcf),
	.w5(32'hbbcbc331),
	.w6(32'h3c2e916e),
	.w7(32'h3bba7325),
	.w8(32'hbbc25d66),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d9425),
	.w1(32'hba06a7ed),
	.w2(32'h3b42d752),
	.w3(32'hba69523b),
	.w4(32'hbb25d82f),
	.w5(32'h3ba66a5a),
	.w6(32'hba74a8fd),
	.w7(32'hbb88a92f),
	.w8(32'hbbf76f70),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f1420),
	.w1(32'hbc2e35e0),
	.w2(32'hbacc4c37),
	.w3(32'h3c0c94c3),
	.w4(32'hbc13fcfd),
	.w5(32'h3bba4862),
	.w6(32'h3c7314a2),
	.w7(32'h3bbc4b21),
	.w8(32'hba8b2400),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6731c4),
	.w1(32'h3c73b926),
	.w2(32'h3b87738a),
	.w3(32'h3bcdabad),
	.w4(32'hbb3ddb1b),
	.w5(32'h3a612002),
	.w6(32'h3ba6f2de),
	.w7(32'hb8766967),
	.w8(32'hbb11968b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f35e01),
	.w1(32'h3a2da1ff),
	.w2(32'hbb130eb4),
	.w3(32'hba5af3d3),
	.w4(32'h3b0b81ea),
	.w5(32'hbb98138d),
	.w6(32'hba39d2e4),
	.w7(32'h3a91c3ab),
	.w8(32'h3c6557f5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ea9a4),
	.w1(32'h3c4e6adb),
	.w2(32'h3b35b6f8),
	.w3(32'hbcacf186),
	.w4(32'hbc5604fb),
	.w5(32'h385edd7e),
	.w6(32'h3c1265fe),
	.w7(32'hbc485ad5),
	.w8(32'hb99dcac2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd983ab),
	.w1(32'h3b3d7002),
	.w2(32'hbba9de20),
	.w3(32'h3aaf0c46),
	.w4(32'h3b3c4991),
	.w5(32'h3ce995d6),
	.w6(32'hb8baebab),
	.w7(32'hba4a6031),
	.w8(32'h3d2e9342),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cbe4a),
	.w1(32'h3c15b06b),
	.w2(32'h3be5c03a),
	.w3(32'hbd0fc8cc),
	.w4(32'hbd14da11),
	.w5(32'h3b53ff9a),
	.w6(32'h3d27e90b),
	.w7(32'hbcb25526),
	.w8(32'h3b2f6a64),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc293f3),
	.w1(32'hbc14d246),
	.w2(32'hbc6c630f),
	.w3(32'hbbceaa0b),
	.w4(32'hbb3f4a23),
	.w5(32'hbca9b6f9),
	.w6(32'hbabfe7e6),
	.w7(32'hbb0462c4),
	.w8(32'hbca85ed9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4321ad),
	.w1(32'hbb82a0ae),
	.w2(32'hbc36d92e),
	.w3(32'h3c36a9ce),
	.w4(32'h3c846a4f),
	.w5(32'hbbecd278),
	.w6(32'hbc01efa6),
	.w7(32'h3bffa6a0),
	.w8(32'hbc12bf34),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10a998),
	.w1(32'hbc0daa74),
	.w2(32'hbbf0253b),
	.w3(32'h3b844915),
	.w4(32'hbc122f9a),
	.w5(32'hbbaeef7c),
	.w6(32'h3c47793f),
	.w7(32'h3c707a5c),
	.w8(32'h3990cae8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9b331),
	.w1(32'hbbc14dbd),
	.w2(32'hba9ae6c7),
	.w3(32'hbb37e6f3),
	.w4(32'hbb9a1811),
	.w5(32'h3b86e885),
	.w6(32'hbb000aea),
	.w7(32'hba1d492a),
	.w8(32'hbb490dc0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03a174),
	.w1(32'h3b4e3824),
	.w2(32'hbba6c39b),
	.w3(32'hbadbc6da),
	.w4(32'h3b965b55),
	.w5(32'hbbf727b0),
	.w6(32'hbc0080ba),
	.w7(32'hbbc7ffac),
	.w8(32'hbc6c56ae),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66f608),
	.w1(32'h3a8a466b),
	.w2(32'h3ba47ec7),
	.w3(32'h3b12aa3f),
	.w4(32'h3bee62ed),
	.w5(32'h3ad2637b),
	.w6(32'hbb9308dd),
	.w7(32'h3ba58175),
	.w8(32'h3ac9cbf9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54650b),
	.w1(32'hb97390d8),
	.w2(32'hbacc6642),
	.w3(32'h3a945375),
	.w4(32'hbb0bf09d),
	.w5(32'hbc6439ff),
	.w6(32'hb914085a),
	.w7(32'hba7461b9),
	.w8(32'hbc6be9bd),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c707f26),
	.w1(32'hbbcac45a),
	.w2(32'hbccdabfc),
	.w3(32'h3c85070b),
	.w4(32'h3c519630),
	.w5(32'h3c6f3ebe),
	.w6(32'hbc43e2a6),
	.w7(32'h3bff07e8),
	.w8(32'h3c999e28),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd12f520),
	.w1(32'hbb3b5f7c),
	.w2(32'h3bb0cfbc),
	.w3(32'hbcd1b551),
	.w4(32'hbc37d121),
	.w5(32'h395da7b2),
	.w6(32'hbbae36a3),
	.w7(32'h3c047ebb),
	.w8(32'h3c29ec4a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7770ae),
	.w1(32'hbc8de59e),
	.w2(32'h3ab0c773),
	.w3(32'h3b44fbba),
	.w4(32'h3b8bf734),
	.w5(32'h3a9ce2cb),
	.w6(32'hbc155674),
	.w7(32'hbbb9f871),
	.w8(32'h3b9c2f09),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11d804),
	.w1(32'h3c248142),
	.w2(32'h3c3fc5c2),
	.w3(32'hbbea1233),
	.w4(32'hbb86d14a),
	.w5(32'h3c1c55b1),
	.w6(32'h3bc8e4fc),
	.w7(32'hbbb76233),
	.w8(32'h3c18f249),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90d3ab),
	.w1(32'h3b756d9b),
	.w2(32'hbbc3892d),
	.w3(32'h3b51ad50),
	.w4(32'h3b4082a6),
	.w5(32'hbb63ba43),
	.w6(32'hba018d1a),
	.w7(32'h3a9631d1),
	.w8(32'h3b2ba2a7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dfe59),
	.w1(32'h3937b336),
	.w2(32'hbbbd06a5),
	.w3(32'h3b9419c0),
	.w4(32'h3b8f111b),
	.w5(32'hbb026b73),
	.w6(32'hbb929221),
	.w7(32'h3b386da8),
	.w8(32'h3cb8c709),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb579a50),
	.w1(32'h3ca03b07),
	.w2(32'hbb768b22),
	.w3(32'hbcffcea3),
	.w4(32'hbbe0a80b),
	.w5(32'h3b278ba2),
	.w6(32'hb71f1677),
	.w7(32'hbc80b788),
	.w8(32'h3c874cc5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84912e),
	.w1(32'h3c932f6e),
	.w2(32'hbc0dcbf8),
	.w3(32'hbb056968),
	.w4(32'h3ab592bb),
	.w5(32'hbbfd4b27),
	.w6(32'h3c0f872c),
	.w7(32'h3c41aa6d),
	.w8(32'h3c96431f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0f65e),
	.w1(32'h3cd0ca97),
	.w2(32'h3ac8988f),
	.w3(32'hbd08ee08),
	.w4(32'hbbf6db59),
	.w5(32'h3afdd112),
	.w6(32'hbadea404),
	.w7(32'hbc2e2694),
	.w8(32'h3ae1f905),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb898531),
	.w1(32'h3b1205a7),
	.w2(32'h3c67fe09),
	.w3(32'h3c2eb17c),
	.w4(32'h3b275e56),
	.w5(32'h3c86f35c),
	.w6(32'hbac9282c),
	.w7(32'hbb5481f3),
	.w8(32'h3c066cb5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76b192),
	.w1(32'hbb8f4317),
	.w2(32'h38f0501c),
	.w3(32'hbbf195bb),
	.w4(32'hbc828e7b),
	.w5(32'h3c090d14),
	.w6(32'h3c3e7198),
	.w7(32'h3b2cec90),
	.w8(32'h3bb2cf37),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb11365),
	.w1(32'h3bf873c5),
	.w2(32'hbabbf10c),
	.w3(32'h3bc02fb6),
	.w4(32'hbc394068),
	.w5(32'h3a76d4eb),
	.w6(32'h3c5531d8),
	.w7(32'hbc11b535),
	.w8(32'hbb08c3f1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd311d),
	.w1(32'hbbef33bf),
	.w2(32'h38c60a55),
	.w3(32'h3c9cb01c),
	.w4(32'h3a58d213),
	.w5(32'hbbe91b7e),
	.w6(32'h3c0b2318),
	.w7(32'h3c057429),
	.w8(32'hbb8e9a50),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff8d83),
	.w1(32'h3b0ee6a5),
	.w2(32'h38acf91a),
	.w3(32'h3b1d93d3),
	.w4(32'h3b810323),
	.w5(32'hbb707fb4),
	.w6(32'hbad54c14),
	.w7(32'hbb5e7990),
	.w8(32'hbb54683c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba500c4),
	.w1(32'h3b82d8a2),
	.w2(32'h3ac7a7e9),
	.w3(32'hbb4b6370),
	.w4(32'h3b5ea9d2),
	.w5(32'h3b0fc131),
	.w6(32'hbb0ba54e),
	.w7(32'h3b40c0bd),
	.w8(32'h39a79a3d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf0bbf),
	.w1(32'hba87afbf),
	.w2(32'hbc168feb),
	.w3(32'h3a126940),
	.w4(32'h3b11e8ec),
	.w5(32'hbb6f546a),
	.w6(32'hbb5038b6),
	.w7(32'hbbb9e95a),
	.w8(32'hbbc89937),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe50101),
	.w1(32'h3b2148c3),
	.w2(32'hbb6701fe),
	.w3(32'hbb8d7721),
	.w4(32'hbbdb2a58),
	.w5(32'hbb47b981),
	.w6(32'h3ad694f5),
	.w7(32'h3b8cbd9e),
	.w8(32'h3c572192),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fa48c),
	.w1(32'hbb92c811),
	.w2(32'h3bd9327b),
	.w3(32'h3b3c25fe),
	.w4(32'h3b64e223),
	.w5(32'h3b6a1092),
	.w6(32'hbc14d6ff),
	.w7(32'h3ba66923),
	.w8(32'h3b087849),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17cb90),
	.w1(32'hbafabf42),
	.w2(32'hb9532080),
	.w3(32'h3b673210),
	.w4(32'h3bcdc302),
	.w5(32'hbadf8e0e),
	.w6(32'h3a86f5be),
	.w7(32'h3c8b4349),
	.w8(32'h3b3b1f5a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb646fc2),
	.w1(32'hbb43eb2c),
	.w2(32'hba6091c9),
	.w3(32'h3ada88b5),
	.w4(32'hba0a47e2),
	.w5(32'h3c7acb7e),
	.w6(32'hbadab433),
	.w7(32'hbbad5f86),
	.w8(32'h3b9f614d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5b911),
	.w1(32'hbc349db9),
	.w2(32'h3b372519),
	.w3(32'h3bb7e2f0),
	.w4(32'hbcb4a568),
	.w5(32'h3a8153e3),
	.w6(32'h3c9622b4),
	.w7(32'hbc18b34f),
	.w8(32'h3aa97948),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba524909),
	.w1(32'hbb95f20c),
	.w2(32'h3bfebc18),
	.w3(32'hbb79421c),
	.w4(32'hbbb5eeb7),
	.w5(32'h3b49dc28),
	.w6(32'hba318556),
	.w7(32'hbb6119a5),
	.w8(32'h3a9e6030),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b203632),
	.w1(32'h3b466295),
	.w2(32'hbbc2c04f),
	.w3(32'h3aa137e1),
	.w4(32'h3a9d3f30),
	.w5(32'hbc495c35),
	.w6(32'hbb2216cb),
	.w7(32'hbbd56d4f),
	.w8(32'h3954b13c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfde0d9),
	.w1(32'h3cbf9f3a),
	.w2(32'h3b0bf52f),
	.w3(32'hbcc47e96),
	.w4(32'h3bb153fc),
	.w5(32'h3a702e0d),
	.w6(32'hbc7858b1),
	.w7(32'hbc5df9b3),
	.w8(32'h3c502ed9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6088f),
	.w1(32'h3a8cb885),
	.w2(32'h3b5d8fea),
	.w3(32'hbc991f3e),
	.w4(32'hbc80c989),
	.w5(32'h3aa7700c),
	.w6(32'h3b714ca3),
	.w7(32'hbb5dee2a),
	.w8(32'h39bb48a5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf42969),
	.w1(32'hbc0b20d8),
	.w2(32'hb9d12438),
	.w3(32'hbba4179d),
	.w4(32'hbc13f9f7),
	.w5(32'hbb9d48c7),
	.w6(32'hbb1cc977),
	.w7(32'hbb9995a2),
	.w8(32'h3a3a2bb2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be192e4),
	.w1(32'h3b8875c2),
	.w2(32'h3c29f0ad),
	.w3(32'h3b71f76e),
	.w4(32'h3b3f40ab),
	.w5(32'hba74bdcc),
	.w6(32'hba9a5af5),
	.w7(32'h3a31471b),
	.w8(32'h3a81661b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ce61f),
	.w1(32'h3b9ca707),
	.w2(32'h3af72c6f),
	.w3(32'h3b889ba6),
	.w4(32'h3add4fc4),
	.w5(32'h3a9321d5),
	.w6(32'hbadb2c05),
	.w7(32'hbb734db8),
	.w8(32'h3bde5ae5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7bff8),
	.w1(32'hbb033a4f),
	.w2(32'h3ba1f6e4),
	.w3(32'h39688d84),
	.w4(32'h3c1e59f2),
	.w5(32'h3c56cd4c),
	.w6(32'hbb99e8e2),
	.w7(32'hbc1559de),
	.w8(32'hbc2244ff),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad2ab2),
	.w1(32'hbc9d9643),
	.w2(32'hbb1c5e71),
	.w3(32'h3c19ea39),
	.w4(32'hbcf54010),
	.w5(32'h3ab37890),
	.w6(32'h3c4fafe9),
	.w7(32'h3ba686d2),
	.w8(32'h3a38eaae),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae575ab),
	.w1(32'hbb05de76),
	.w2(32'h3b993abe),
	.w3(32'h3a87aa05),
	.w4(32'hbb3d5076),
	.w5(32'h3b349929),
	.w6(32'hb9224689),
	.w7(32'hbb4c27de),
	.w8(32'hba966f8c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b017146),
	.w1(32'h3b8f9712),
	.w2(32'h3c689a81),
	.w3(32'h3bb51224),
	.w4(32'h3bfe3652),
	.w5(32'h3cbbc49c),
	.w6(32'hb9b7751e),
	.w7(32'h3b8ca96f),
	.w8(32'h3c8215ab),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ca8d0),
	.w1(32'hbc39b142),
	.w2(32'h3c3c9cb1),
	.w3(32'h3bafc774),
	.w4(32'hbcade7b6),
	.w5(32'h3cb60bdc),
	.w6(32'h3cb7cdae),
	.w7(32'h3ab80853),
	.w8(32'h3c85f03c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58c963),
	.w1(32'hbc708d92),
	.w2(32'hbbc44f2b),
	.w3(32'h3c2cc450),
	.w4(32'hbca30b52),
	.w5(32'hbb028396),
	.w6(32'h3cb93e2d),
	.w7(32'h3c348a16),
	.w8(32'h3bbd224a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b510f7a),
	.w1(32'h3bb3ca10),
	.w2(32'h3b812289),
	.w3(32'h39fa09c9),
	.w4(32'h3c10da44),
	.w5(32'hba17c933),
	.w6(32'hbb550605),
	.w7(32'h3a736998),
	.w8(32'h3a6d28a6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b6ca0),
	.w1(32'hb955ad16),
	.w2(32'hbae066ad),
	.w3(32'hbad1bfe2),
	.w4(32'hba87ad7a),
	.w5(32'h3a840f10),
	.w6(32'hbad4eb72),
	.w7(32'hbb3cbf36),
	.w8(32'h3b2c0596),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35b316),
	.w1(32'h3c02f583),
	.w2(32'h3bb813b2),
	.w3(32'hbb603ab8),
	.w4(32'h3b443f57),
	.w5(32'h3b102fe6),
	.w6(32'h3b89d5d5),
	.w7(32'hbabbdc78),
	.w8(32'h37f406e3),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1e39c),
	.w1(32'h3b9afa6f),
	.w2(32'hbbb7bedb),
	.w3(32'h3bb4d477),
	.w4(32'h3afa5422),
	.w5(32'h3bed6b13),
	.w6(32'h3b34a1c7),
	.w7(32'h391bc238),
	.w8(32'h3cbb5bf4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60e1f3),
	.w1(32'h3c55d76b),
	.w2(32'hbbd8a9f7),
	.w3(32'hbcdce707),
	.w4(32'hbba04476),
	.w5(32'h3aa711e4),
	.w6(32'h3c5553ed),
	.w7(32'hbc102829),
	.w8(32'h3c2d7900),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3f6f8),
	.w1(32'hbb85afb9),
	.w2(32'hbbcad40b),
	.w3(32'hbbaad9f9),
	.w4(32'hbb5b9587),
	.w5(32'h3b4cce12),
	.w6(32'h3b1f4723),
	.w7(32'hbbe2352a),
	.w8(32'h3bb2c2e0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45ec01),
	.w1(32'hbc7702c3),
	.w2(32'hbb92a1d2),
	.w3(32'h3b70f044),
	.w4(32'h3b150d5c),
	.w5(32'hbcae9dcb),
	.w6(32'hbba2cbd0),
	.w7(32'h3c019134),
	.w8(32'h3a8c64bb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd59aa),
	.w1(32'h3c82e5ca),
	.w2(32'h3b1391d3),
	.w3(32'hbbc0286f),
	.w4(32'h3c30611d),
	.w5(32'hba90a862),
	.w6(32'hbca743db),
	.w7(32'h3a233df9),
	.w8(32'h3b038276),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0609fe),
	.w1(32'hbac77f5b),
	.w2(32'h3b019e8b),
	.w3(32'hbb803cb0),
	.w4(32'hbb5b0b07),
	.w5(32'h39257430),
	.w6(32'hba218a67),
	.w7(32'hbb92545b),
	.w8(32'h3b34c0fb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5421c),
	.w1(32'hbb2b8ab4),
	.w2(32'hbb00e8e8),
	.w3(32'hba2040c8),
	.w4(32'hbbb5e665),
	.w5(32'hbb05428e),
	.w6(32'hba4cba08),
	.w7(32'hbba27c14),
	.w8(32'h3c8c719a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c2f22),
	.w1(32'h3cd55157),
	.w2(32'h3c0398e1),
	.w3(32'hbcff9408),
	.w4(32'hba2ebda7),
	.w5(32'hbb67f516),
	.w6(32'hbb631e89),
	.w7(32'hbbd0aa52),
	.w8(32'hbb3bb3db),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fccce),
	.w1(32'h3c516c79),
	.w2(32'h3b9fb171),
	.w3(32'h3bef1b77),
	.w4(32'h3b0ed172),
	.w5(32'hbbf676ff),
	.w6(32'h3b9dc86f),
	.w7(32'hbc20f641),
	.w8(32'hbb33e7f9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59129f),
	.w1(32'h3af88477),
	.w2(32'hbb788a4a),
	.w3(32'hbba77ea2),
	.w4(32'hbb4c5896),
	.w5(32'hbb99fca6),
	.w6(32'hba1f220e),
	.w7(32'h3b156943),
	.w8(32'hbb2207a7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab55db1),
	.w1(32'h3a791c2d),
	.w2(32'h3a627d78),
	.w3(32'hb91c21a0),
	.w4(32'h3bc218ff),
	.w5(32'h3aa83068),
	.w6(32'hbbf2778c),
	.w7(32'hba173ae0),
	.w8(32'h3aac8326),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94fd38),
	.w1(32'hbc1ed04c),
	.w2(32'hbbb79d8c),
	.w3(32'hbbc0c247),
	.w4(32'hbbf5474f),
	.w5(32'hbb9fe73b),
	.w6(32'hba49c344),
	.w7(32'hba5d7963),
	.w8(32'h3abeaf08),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6faa),
	.w1(32'hba6b534f),
	.w2(32'h3b335663),
	.w3(32'hbb98310d),
	.w4(32'hbbb185d2),
	.w5(32'h3ad23d78),
	.w6(32'hbac630d7),
	.w7(32'hbb705595),
	.w8(32'h3c32afbe),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55e323),
	.w1(32'h3ad8a33a),
	.w2(32'hb915b647),
	.w3(32'hbcd8403d),
	.w4(32'hbc2e613c),
	.w5(32'hbb8414d5),
	.w6(32'hbb8b9bfe),
	.w7(32'hbb4701f6),
	.w8(32'hbc59f55d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900efe),
	.w1(32'hbc91f0a2),
	.w2(32'hbc4a2a93),
	.w3(32'h3b7ed706),
	.w4(32'h3b98a3ff),
	.w5(32'h3b69e899),
	.w6(32'hbcaeaac5),
	.w7(32'hbba3d049),
	.w8(32'hba02f236),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b0cc9),
	.w1(32'h3c0a8dc8),
	.w2(32'hbb472829),
	.w3(32'hbc5999eb),
	.w4(32'hbbad1c7f),
	.w5(32'hbc465d7a),
	.w6(32'h392bbbd1),
	.w7(32'hbc1a4d5a),
	.w8(32'h3bf0d7e7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f7983),
	.w1(32'h3b857adf),
	.w2(32'h3c1db809),
	.w3(32'hbc2b257e),
	.w4(32'h3bf41be4),
	.w5(32'h3c13373f),
	.w6(32'hbbee6e97),
	.w7(32'h3c3499c1),
	.w8(32'h3c78768d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83c5ff),
	.w1(32'hbae69fae),
	.w2(32'h38b7bef6),
	.w3(32'hbabea365),
	.w4(32'hbca8a6ff),
	.w5(32'h3b6049b5),
	.w6(32'h3c859dbc),
	.w7(32'hbb02ddcb),
	.w8(32'h3bfcf3bd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baefbc6),
	.w1(32'hba17078f),
	.w2(32'h3caaafd2),
	.w3(32'h3c086ef4),
	.w4(32'hb9d41c87),
	.w5(32'h3ad7dbe2),
	.w6(32'h3c6db698),
	.w7(32'hbb639e39),
	.w8(32'hbc8b52a0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beae247),
	.w1(32'hbca1e197),
	.w2(32'hbbe61a51),
	.w3(32'h3c6946c6),
	.w4(32'hbc76a208),
	.w5(32'h3c178ea4),
	.w6(32'h39e2fd65),
	.w7(32'hbb8742e2),
	.w8(32'hbca091ee),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30a335),
	.w1(32'hbc4b22d8),
	.w2(32'hbb61460b),
	.w3(32'h3c8aa97c),
	.w4(32'hbc9dd26a),
	.w5(32'hbb183dbc),
	.w6(32'h3c43fcc6),
	.w7(32'hbb3535f7),
	.w8(32'hba9f17e4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fdb19),
	.w1(32'h3ba40eea),
	.w2(32'h3c1210e5),
	.w3(32'h3c233817),
	.w4(32'h3b527af5),
	.w5(32'h3a753629),
	.w6(32'h3b838cd7),
	.w7(32'hb9f2bee6),
	.w8(32'h3bebe68b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b712e62),
	.w1(32'h3c00d382),
	.w2(32'hbc084e83),
	.w3(32'h3b11220b),
	.w4(32'hb9a9db0f),
	.w5(32'hbca2614a),
	.w6(32'h3b9d50f5),
	.w7(32'hbb827a96),
	.w8(32'hbabfc692),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46db47),
	.w1(32'h3bcbe4fb),
	.w2(32'hba404b60),
	.w3(32'hbc0e5ef0),
	.w4(32'h3c518843),
	.w5(32'hbab6fcb5),
	.w6(32'hbc3c2753),
	.w7(32'hbc09db61),
	.w8(32'h3bea9d8c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe1738),
	.w1(32'hba88317b),
	.w2(32'hb9dbfb96),
	.w3(32'hba5250fd),
	.w4(32'hbb328a68),
	.w5(32'hbb3a1179),
	.w6(32'h3bc77028),
	.w7(32'hbbc1ed72),
	.w8(32'hb81fb292),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1ecd4),
	.w1(32'h3bb67995),
	.w2(32'h3acc0b25),
	.w3(32'h3a6aad2c),
	.w4(32'h3b5fd75a),
	.w5(32'hba48f05b),
	.w6(32'hb9fe372e),
	.w7(32'hbb8f6ed6),
	.w8(32'h3bd96e0d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaeb92),
	.w1(32'hbbffc4c3),
	.w2(32'h3ba8f10f),
	.w3(32'h3bf2d95a),
	.w4(32'h3ae4cdb1),
	.w5(32'hbbaea47d),
	.w6(32'h3b20e30b),
	.w7(32'hbb88ffbf),
	.w8(32'hbba67960),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82fbe67),
	.w1(32'hbca87d99),
	.w2(32'h3c159fd5),
	.w3(32'h3c398470),
	.w4(32'h3bd18e23),
	.w5(32'h3b7f6b4f),
	.w6(32'h3bf64241),
	.w7(32'h3c2ad67f),
	.w8(32'hbc230e18),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25e7bc),
	.w1(32'hbc627ba8),
	.w2(32'hbbde3c2d),
	.w3(32'h3c641ae6),
	.w4(32'hbbdadd38),
	.w5(32'hbc9ca7f2),
	.w6(32'h3aadb669),
	.w7(32'h3b87dcaa),
	.w8(32'h3aa7552a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4268a4),
	.w1(32'hba05f031),
	.w2(32'hbc2ac78b),
	.w3(32'h3b28db00),
	.w4(32'h3c3490c0),
	.w5(32'hbc2f40b4),
	.w6(32'hbc26f7b0),
	.w7(32'h3bc51c85),
	.w8(32'h3b1495cc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06fbff),
	.w1(32'h3c4905a3),
	.w2(32'h3ab2aba0),
	.w3(32'hbc37e33f),
	.w4(32'h3b9f786b),
	.w5(32'h3bf02076),
	.w6(32'hbc23298e),
	.w7(32'hbb7b80f3),
	.w8(32'h3c6610fc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee4a28),
	.w1(32'h3c7d3345),
	.w2(32'h3ad9aebe),
	.w3(32'hbc8f115c),
	.w4(32'hbba04a84),
	.w5(32'hbc2b1b02),
	.w6(32'h3a23f20e),
	.w7(32'hbc1229a1),
	.w8(32'hbc417f6c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb699d0c),
	.w1(32'h3b953d4c),
	.w2(32'h3c1e7e61),
	.w3(32'h3b6aaa63),
	.w4(32'hba9b7caf),
	.w5(32'h3bc1e9db),
	.w6(32'hba849221),
	.w7(32'h3926da17),
	.w8(32'h3bb48ae2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936a2c),
	.w1(32'h3ac2b2b9),
	.w2(32'hba60584f),
	.w3(32'h3c1e0777),
	.w4(32'hbc69ff33),
	.w5(32'hba0d7b22),
	.w6(32'h3c8f5ecf),
	.w7(32'h3b4aa897),
	.w8(32'hb9ffe9f9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3698b),
	.w1(32'hbafbc239),
	.w2(32'hb9d2ae5d),
	.w3(32'hbbbbc73a),
	.w4(32'hbbc00d1a),
	.w5(32'hba90cedf),
	.w6(32'hbbd869c9),
	.w7(32'hbbb7f43d),
	.w8(32'h3bccfc22),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb574662),
	.w1(32'h3a0fa01b),
	.w2(32'hbaefb5b0),
	.w3(32'hbc179892),
	.w4(32'hbba1f7f2),
	.w5(32'hba8203d8),
	.w6(32'h3a0feeb3),
	.w7(32'hbb39f28b),
	.w8(32'hb9d69553),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10444c),
	.w1(32'h39b68330),
	.w2(32'h3bcb1d61),
	.w3(32'hb9ee1db1),
	.w4(32'h39c89130),
	.w5(32'h3c700531),
	.w6(32'h3a4ac29b),
	.w7(32'h381bbf02),
	.w8(32'hb9fe991a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb24d1a),
	.w1(32'hbc87706b),
	.w2(32'h3bff88ee),
	.w3(32'h3c14da48),
	.w4(32'hbcbd5701),
	.w5(32'h3c2406f6),
	.w6(32'h3cabd88c),
	.w7(32'hba03942d),
	.w8(32'hbc4527fd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27e2ee),
	.w1(32'hbc2f1903),
	.w2(32'hbb13c758),
	.w3(32'h3cad3b71),
	.w4(32'hbc06f7b6),
	.w5(32'hbbb8368b),
	.w6(32'h3c0e0064),
	.w7(32'hba9b93f2),
	.w8(32'h3a8669de),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ac8ab),
	.w1(32'h3bafe382),
	.w2(32'h3924ff3d),
	.w3(32'hbaa983c6),
	.w4(32'h3c4db5ba),
	.w5(32'hba9ea542),
	.w6(32'hbc1cdddd),
	.w7(32'h3bfa1434),
	.w8(32'hbab9c975),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9273b),
	.w1(32'hbaa50520),
	.w2(32'h3991103d),
	.w3(32'h3aadb0ac),
	.w4(32'hba87b0a2),
	.w5(32'h3a429639),
	.w6(32'hbb4bdf61),
	.w7(32'hbbb920b0),
	.w8(32'hba08fea8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba042dd1),
	.w1(32'hbaa2fe66),
	.w2(32'hbc04626b),
	.w3(32'hbb9adb54),
	.w4(32'hbba42769),
	.w5(32'h3a64c18b),
	.w6(32'hbb637916),
	.w7(32'hbb459720),
	.w8(32'h3bd50311),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d7ca4),
	.w1(32'h3c219226),
	.w2(32'h3bb2958d),
	.w3(32'hbc4cc39f),
	.w4(32'hbc12898c),
	.w5(32'h3b50aea7),
	.w6(32'h3c11175d),
	.w7(32'hbc66af0c),
	.w8(32'hba839ce5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc03b90),
	.w1(32'h3bc5b79c),
	.w2(32'hbc43c3f3),
	.w3(32'h3b8c7ce9),
	.w4(32'h3b33856a),
	.w5(32'hbb4651fe),
	.w6(32'h3b4a92f1),
	.w7(32'h3b16125a),
	.w8(32'h3c8e6a71),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8476e7),
	.w1(32'h3c7ac3e0),
	.w2(32'hbb3ba40b),
	.w3(32'hbcbb655a),
	.w4(32'h3b40b93a),
	.w5(32'hbc4e7b37),
	.w6(32'h3b8599dd),
	.w7(32'hbb88ebe8),
	.w8(32'h3bc3c9fc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9290ba),
	.w1(32'h3c9f9d09),
	.w2(32'hbc117ba5),
	.w3(32'hbc57707a),
	.w4(32'h3c3e9942),
	.w5(32'hbbe5317f),
	.w6(32'hbc9ece45),
	.w7(32'hbc49626f),
	.w8(32'h3afcd170),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccf202b),
	.w1(32'h3c31dd31),
	.w2(32'h3bb9393e),
	.w3(32'h3b126a6d),
	.w4(32'h3c89c1d5),
	.w5(32'h3bf51a15),
	.w6(32'hbc88f15c),
	.w7(32'hbc7fa069),
	.w8(32'hbbf76784),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2923a6),
	.w1(32'hbbd2a084),
	.w2(32'hbba08ace),
	.w3(32'h3be0ab73),
	.w4(32'hba271266),
	.w5(32'hbc4a10de),
	.w6(32'hbb151ae0),
	.w7(32'h3aa97aa4),
	.w8(32'h3c45971d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06a91d),
	.w1(32'h3c44129f),
	.w2(32'h3c8e9318),
	.w3(32'hbbfd3640),
	.w4(32'h3c923918),
	.w5(32'h3c28d3c1),
	.w6(32'hbc83fd61),
	.w7(32'hbaeea2b5),
	.w8(32'hbc2ebeed),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86751be),
	.w1(32'hbbd0e149),
	.w2(32'h3baad8f1),
	.w3(32'h3bd0c5ed),
	.w4(32'hbc1c660f),
	.w5(32'hbc7b1a19),
	.w6(32'h3c239e30),
	.w7(32'hbb6483ed),
	.w8(32'hbc683d06),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4315d),
	.w1(32'h3c15061e),
	.w2(32'h3c02d01e),
	.w3(32'h3ad05b33),
	.w4(32'h3c3383ae),
	.w5(32'h3d0a818a),
	.w6(32'hbc3c9767),
	.w7(32'h3c5bdc7b),
	.w8(32'h3bec0a79),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd59613),
	.w1(32'hbc5fab06),
	.w2(32'h3cc8039e),
	.w3(32'h3c6edf22),
	.w4(32'hbbd9c1c2),
	.w5(32'hbc2df7dd),
	.w6(32'h3c4c492f),
	.w7(32'hbb755a7b),
	.w8(32'hbbfd920f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03dc0a),
	.w1(32'h3c241282),
	.w2(32'hb8adf80f),
	.w3(32'h3cf6b54b),
	.w4(32'h3cddb159),
	.w5(32'h3af23534),
	.w6(32'hbc1abc1a),
	.w7(32'h3a8d5484),
	.w8(32'hb9be4da4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac53b2a),
	.w1(32'hba7e86c5),
	.w2(32'h3bf4eaf9),
	.w3(32'h3b0a9531),
	.w4(32'hbb94f8c0),
	.w5(32'h3bf506fe),
	.w6(32'hbb266c78),
	.w7(32'hbc0ee5c5),
	.w8(32'h3b4061d2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc681f8e),
	.w1(32'hbc1c2227),
	.w2(32'h3c2d7d59),
	.w3(32'hbc08a055),
	.w4(32'hbc133f47),
	.w5(32'hbaa8aef5),
	.w6(32'hbad10223),
	.w7(32'hbc1b1741),
	.w8(32'h3a87dae3),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b952f8f),
	.w1(32'h3b887f65),
	.w2(32'hba001d85),
	.w3(32'h3b66d39a),
	.w4(32'hb9ab01d9),
	.w5(32'hbb9a85ca),
	.w6(32'hbc03dcde),
	.w7(32'hbbb004a8),
	.w8(32'hbba08f0a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb95ce),
	.w1(32'hbad950c6),
	.w2(32'h3b84afe1),
	.w3(32'hbb17d290),
	.w4(32'hbb9cefcf),
	.w5(32'h3bbbf948),
	.w6(32'hbb67ca2a),
	.w7(32'hbbaecce1),
	.w8(32'h3ba1016e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94542fc),
	.w1(32'hbb3aaa28),
	.w2(32'hba6ec81d),
	.w3(32'hbaa023ff),
	.w4(32'hbb0ceb07),
	.w5(32'hbaf8bf90),
	.w6(32'h3ae55cb3),
	.w7(32'h392f3c7b),
	.w8(32'hbc826b83),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ad0e0),
	.w1(32'h3c0b7050),
	.w2(32'hbab5f06d),
	.w3(32'h3c2a0b3f),
	.w4(32'h3c23d7b3),
	.w5(32'h3a34a84a),
	.w6(32'hbc400296),
	.w7(32'h3bde4ee2),
	.w8(32'h3adc633a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3fe0e),
	.w1(32'h39ce0ce6),
	.w2(32'h3bde7f3e),
	.w3(32'hbb23d45c),
	.w4(32'hbb37e8fc),
	.w5(32'h3bbf49da),
	.w6(32'h3af34e23),
	.w7(32'hbadc4fe3),
	.w8(32'h3c1cd2d3),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23ff5b),
	.w1(32'hbaac4b13),
	.w2(32'h3c481c76),
	.w3(32'hbb0aef43),
	.w4(32'h3b3363c2),
	.w5(32'h3b9a3a4d),
	.w6(32'h3c065351),
	.w7(32'h3c15a877),
	.w8(32'hbc770894),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b4651),
	.w1(32'hbd119e21),
	.w2(32'h3b4cd3f5),
	.w3(32'h3d22b1a6),
	.w4(32'h3c221556),
	.w5(32'h3b08a0e9),
	.w6(32'h3a54598a),
	.w7(32'h3c2d57d6),
	.w8(32'h3b2b61e0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85f1fd),
	.w1(32'hbb1670bb),
	.w2(32'h3ac06eff),
	.w3(32'hb99f9a64),
	.w4(32'hb8193d70),
	.w5(32'h3a4f513c),
	.w6(32'hbaeb6c10),
	.w7(32'hb9f0a6e6),
	.w8(32'h3aeeb5bb),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe9504),
	.w1(32'h3ac3d698),
	.w2(32'hbb808c28),
	.w3(32'h3992de81),
	.w4(32'h3b059795),
	.w5(32'hbbd4872e),
	.w6(32'h3a44ed22),
	.w7(32'h3a9885ec),
	.w8(32'hbc027399),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6eac22),
	.w1(32'hbbed501e),
	.w2(32'h3baffdda),
	.w3(32'hbb5b0eae),
	.w4(32'hbb9bcf95),
	.w5(32'h3a89fa74),
	.w6(32'hbbc3b150),
	.w7(32'hbbb637cf),
	.w8(32'h3ba1ce47),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5c76b),
	.w1(32'h3b9710a3),
	.w2(32'hbc3e6268),
	.w3(32'h3b660390),
	.w4(32'h3bee891b),
	.w5(32'hbc6270a3),
	.w6(32'h3bd9b8a0),
	.w7(32'h3c26d0db),
	.w8(32'hbb21208d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b2a41),
	.w1(32'hbb63628a),
	.w2(32'h3bbac03c),
	.w3(32'hb5e10352),
	.w4(32'h3b4e816e),
	.w5(32'hb844b319),
	.w6(32'hbbdd3dd6),
	.w7(32'h3c2c3dfb),
	.w8(32'h3b156a06),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba831023),
	.w1(32'h3b5ec305),
	.w2(32'hbb89ffce),
	.w3(32'h3a0eb016),
	.w4(32'h3a6b73a1),
	.w5(32'hbb01104d),
	.w6(32'h3c001f2c),
	.w7(32'h3b66a300),
	.w8(32'hb92fc353),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b6b6),
	.w1(32'hbc2aaa78),
	.w2(32'hb607cfdc),
	.w3(32'hbbb3b952),
	.w4(32'h390c9feb),
	.w5(32'h3b2abb58),
	.w6(32'h3b46e22c),
	.w7(32'h3bd1c23e),
	.w8(32'h3abfa36e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea969f),
	.w1(32'hbbb932f3),
	.w2(32'h3b7c7e22),
	.w3(32'h3b0eb7c8),
	.w4(32'hbc72bb19),
	.w5(32'hba643a3c),
	.w6(32'h3a22a940),
	.w7(32'hba881be7),
	.w8(32'hbb071845),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c095a61),
	.w1(32'h3b6d720c),
	.w2(32'h3bef6ca4),
	.w3(32'h3ba417f9),
	.w4(32'h3a1a04bc),
	.w5(32'h3c044542),
	.w6(32'hba55ec74),
	.w7(32'hba72a616),
	.w8(32'h3c369de5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5aaf30),
	.w1(32'h3b80031c),
	.w2(32'hba831245),
	.w3(32'hbbbfebfa),
	.w4(32'hbab22f04),
	.w5(32'hbcd418c4),
	.w6(32'h3bacd730),
	.w7(32'h3b89d761),
	.w8(32'hbbc4fd3c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb7bc13),
	.w1(32'h3be31c66),
	.w2(32'h3b10255e),
	.w3(32'hbc21c76d),
	.w4(32'h3c97fcfb),
	.w5(32'h3ca38bf2),
	.w6(32'hbc6a4893),
	.w7(32'hbae5e821),
	.w8(32'h3c9e032a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6399d3),
	.w1(32'hbc53b609),
	.w2(32'h3af024b7),
	.w3(32'hbb24ba77),
	.w4(32'hbca51090),
	.w5(32'hbb3149eb),
	.w6(32'h3cb4cd8a),
	.w7(32'h3b8cf03b),
	.w8(32'h3ac5dc7b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da8107),
	.w1(32'h3960a5f2),
	.w2(32'hbbad50c0),
	.w3(32'hbc064009),
	.w4(32'hbb6e22fa),
	.w5(32'hbc1a081d),
	.w6(32'hbb380a1f),
	.w7(32'hb7d3ff89),
	.w8(32'hbc1b9e8d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd9f48),
	.w1(32'h3c21b0f6),
	.w2(32'hbb8e1dfd),
	.w3(32'h38abe2b1),
	.w4(32'h3c4c241a),
	.w5(32'hbc127018),
	.w6(32'h3aa58f63),
	.w7(32'h3c1b00cb),
	.w8(32'hbb5bcad7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd019a8),
	.w1(32'h3aaedb94),
	.w2(32'hba6b0dde),
	.w3(32'h39d5f110),
	.w4(32'hbc067acc),
	.w5(32'h3ab2408c),
	.w6(32'hbaa4fa9c),
	.w7(32'h3b00e320),
	.w8(32'h3b9946af),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a004e),
	.w1(32'hbb2708dc),
	.w2(32'h3a340ec0),
	.w3(32'hbb0a41f7),
	.w4(32'hbb01c73d),
	.w5(32'h3c4b2426),
	.w6(32'h3b360d03),
	.w7(32'h3a0b5dec),
	.w8(32'h3c8c04de),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c114b2f),
	.w1(32'h3b9394f8),
	.w2(32'hbb8583c1),
	.w3(32'h3cb7574c),
	.w4(32'h3c1390b1),
	.w5(32'hbbc6f559),
	.w6(32'h3c594358),
	.w7(32'hbae260be),
	.w8(32'h3bc4e02e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0190ca),
	.w1(32'hb9832347),
	.w2(32'h3a7c5029),
	.w3(32'h3bcdc025),
	.w4(32'hbaa5b87b),
	.w5(32'h3b1d1722),
	.w6(32'hba3088d8),
	.w7(32'hbc0d9720),
	.w8(32'h3ac00d60),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba230f3),
	.w1(32'hbbd7a4a1),
	.w2(32'h3c8affdc),
	.w3(32'h3a0905b4),
	.w4(32'h3b631b54),
	.w5(32'h3a15fa14),
	.w6(32'h39993015),
	.w7(32'h3baa7c9e),
	.w8(32'h3bb6ea6f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b116f86),
	.w1(32'h397eb395),
	.w2(32'hbb85f150),
	.w3(32'hbc75e767),
	.w4(32'hbc187a36),
	.w5(32'hbb96c1b2),
	.w6(32'hbc2a1d26),
	.w7(32'hbb508b47),
	.w8(32'hbb930faa),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396512c2),
	.w1(32'h38e32c85),
	.w2(32'hbae53ba1),
	.w3(32'h39d1e0a1),
	.w4(32'h3a9077b7),
	.w5(32'h3b9c1c9c),
	.w6(32'hbb4fbee6),
	.w7(32'hb9ae7486),
	.w8(32'hbab38445),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9c24a),
	.w1(32'hbc13a504),
	.w2(32'h3a7e1674),
	.w3(32'hbb6112b1),
	.w4(32'hbc611002),
	.w5(32'hb9ea44d5),
	.w6(32'hbc0bf828),
	.w7(32'hbbeb49e2),
	.w8(32'hbbb12ea3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3dbb43),
	.w1(32'h3b04ff51),
	.w2(32'h3b5e0f06),
	.w3(32'h3b9df4f6),
	.w4(32'h3c220c89),
	.w5(32'h3c3e0226),
	.w6(32'hba225a6c),
	.w7(32'h3c271d77),
	.w8(32'h3aee5c3c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c826154),
	.w1(32'h3c5c0dd8),
	.w2(32'hbaecec55),
	.w3(32'h3c861591),
	.w4(32'h3ab50b19),
	.w5(32'hb847475b),
	.w6(32'hbba684c1),
	.w7(32'hbbca6e38),
	.w8(32'h3c30be50),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb234b9),
	.w1(32'hbbc0d203),
	.w2(32'hbb3d7458),
	.w3(32'hbcc7cce1),
	.w4(32'hbc84f364),
	.w5(32'hbb830093),
	.w6(32'hbc16a45f),
	.w7(32'hbc319da9),
	.w8(32'hbbd152c1),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeb553),
	.w1(32'hbbf87136),
	.w2(32'h3b40bedc),
	.w3(32'hbbf1d752),
	.w4(32'hbc4c5086),
	.w5(32'h3c07bd92),
	.w6(32'hbb069b63),
	.w7(32'hbc2491a4),
	.w8(32'h3ca0e4c0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb017c98),
	.w1(32'h3ae80831),
	.w2(32'hbb803d9a),
	.w3(32'h3c94a2b6),
	.w4(32'h3c6089fe),
	.w5(32'hbbf526dc),
	.w6(32'h3ca191e2),
	.w7(32'h3c1ec053),
	.w8(32'hbc1fad28),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48c721),
	.w1(32'hbc655598),
	.w2(32'hb742609d),
	.w3(32'hbcb27f3a),
	.w4(32'hbcb07916),
	.w5(32'hbb8deb44),
	.w6(32'hbc90fc23),
	.w7(32'hbcb6127a),
	.w8(32'hbc0b2c79),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ea97f),
	.w1(32'h3ba14aad),
	.w2(32'hbb08adab),
	.w3(32'hba947db5),
	.w4(32'hbab2998d),
	.w5(32'hbbc3155c),
	.w6(32'hbc3bef6e),
	.w7(32'hbbe146f1),
	.w8(32'hbc1165b2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaf205),
	.w1(32'h3b9f4afa),
	.w2(32'hbb8bbe78),
	.w3(32'h3b5c0e5e),
	.w4(32'h3c0d6469),
	.w5(32'h3b026372),
	.w6(32'h3a07c8b8),
	.w7(32'h3b6489cc),
	.w8(32'h3b0a6348),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa1462),
	.w1(32'hbb84e58f),
	.w2(32'hbbe73cfb),
	.w3(32'hbc254762),
	.w4(32'h3c4485d7),
	.w5(32'hbc1048bd),
	.w6(32'h3ae6a6ac),
	.w7(32'h3acaf49d),
	.w8(32'hbbc22a21),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb654079),
	.w1(32'hbbab3d58),
	.w2(32'hb9d6c9c4),
	.w3(32'h3ba154f5),
	.w4(32'hbc149cef),
	.w5(32'h3b640d18),
	.w6(32'hbb2c0f29),
	.w7(32'hbc044c6c),
	.w8(32'h3c90e42c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d0b76),
	.w1(32'hbaef742c),
	.w2(32'h3b0ca72a),
	.w3(32'h3b6ee02c),
	.w4(32'hbbb2a4a5),
	.w5(32'h3ac6cc28),
	.w6(32'h3ca06e5a),
	.w7(32'h3c298a13),
	.w8(32'hbb3d14fc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd73fc0),
	.w1(32'h3c1dae51),
	.w2(32'h3c23b738),
	.w3(32'h3b9de610),
	.w4(32'h3bf33f76),
	.w5(32'h3b2578d3),
	.w6(32'hbb213f45),
	.w7(32'hb811c621),
	.w8(32'h383051e1),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c1250),
	.w1(32'h3b21bf67),
	.w2(32'hbaf022a0),
	.w3(32'h3b6e7ca3),
	.w4(32'hb9dc0514),
	.w5(32'hba82a93e),
	.w6(32'hbae3c71e),
	.w7(32'hb926391a),
	.w8(32'h3b5838ef),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c1082),
	.w1(32'hbc0b8a30),
	.w2(32'h3ba35648),
	.w3(32'hbb3d9cde),
	.w4(32'h3b0f8605),
	.w5(32'hbbede34f),
	.w6(32'hbb21aee4),
	.w7(32'h3c1bed53),
	.w8(32'hbb989c4b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bc0d0),
	.w1(32'hbba6bedd),
	.w2(32'h3c209151),
	.w3(32'hbc14d2a7),
	.w4(32'h3a1d83e0),
	.w5(32'hb959e085),
	.w6(32'h3b90cd00),
	.w7(32'h3c43d36f),
	.w8(32'hbaa6d088),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf059d),
	.w1(32'hbc49bf07),
	.w2(32'h3bb232d5),
	.w3(32'hbbfa304e),
	.w4(32'h399d3b76),
	.w5(32'h3b6be8c8),
	.w6(32'hbbefcbf8),
	.w7(32'h3c051cde),
	.w8(32'h3bb71c5b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab46d23),
	.w1(32'h390ea099),
	.w2(32'hba035527),
	.w3(32'hbbbe302f),
	.w4(32'hbbb50168),
	.w5(32'h3ba7c83a),
	.w6(32'hbb113d9e),
	.w7(32'hbb154454),
	.w8(32'hbb1655a4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d3cbe),
	.w1(32'hbc022be8),
	.w2(32'h3c02e62d),
	.w3(32'hbbc813af),
	.w4(32'hbc29d222),
	.w5(32'h3ba7e676),
	.w6(32'hbb0c6077),
	.w7(32'hbbbc2bc9),
	.w8(32'h3b9693ae),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0da3dc),
	.w1(32'h3b624bb0),
	.w2(32'hbc10be43),
	.w3(32'h3b8da6f0),
	.w4(32'hbbe10d57),
	.w5(32'hbc47edfa),
	.w6(32'h3b71fc2b),
	.w7(32'hbbcb10a5),
	.w8(32'hbb9f833f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddd1b5),
	.w1(32'h3b16ba73),
	.w2(32'h3b5bc69b),
	.w3(32'hbb200f93),
	.w4(32'hbb504638),
	.w5(32'hb8485948),
	.w6(32'hbbfc4588),
	.w7(32'hbbbb4d2b),
	.w8(32'h3b848a26),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27b432),
	.w1(32'h3b4742d4),
	.w2(32'hba5336bb),
	.w3(32'hba9f0596),
	.w4(32'hbb644aa8),
	.w5(32'h3a8cc976),
	.w6(32'h3b9a67de),
	.w7(32'hbbac150e),
	.w8(32'h3b62cf62),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e320b),
	.w1(32'h3c680bb2),
	.w2(32'h3b1d957c),
	.w3(32'hbaeeb9dd),
	.w4(32'h3ca6880a),
	.w5(32'h3b5cf270),
	.w6(32'h3a89a9c9),
	.w7(32'h3ce88e1c),
	.w8(32'hbb7676e5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2426d3),
	.w1(32'h3c0decba),
	.w2(32'h3c324e7f),
	.w3(32'h3c4978d3),
	.w4(32'h3b3b72c7),
	.w5(32'h3c236908),
	.w6(32'h3a271d28),
	.w7(32'hba5117d4),
	.w8(32'h3c69c200),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a315b),
	.w1(32'hbc0b3ca7),
	.w2(32'hbcb165f3),
	.w3(32'hbc2054cf),
	.w4(32'hba899bd9),
	.w5(32'hbc84feae),
	.w6(32'h3b7ed013),
	.w7(32'hbb50a2ae),
	.w8(32'hbc6eb6fa),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc097d34),
	.w1(32'hbbd291a2),
	.w2(32'hbb9acb64),
	.w3(32'hbc7d0a33),
	.w4(32'hbbf93004),
	.w5(32'hbc0216b8),
	.w6(32'hbc5be416),
	.w7(32'hbbff5490),
	.w8(32'hbad45264),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ae178),
	.w1(32'hbbf2b502),
	.w2(32'h3b45aedb),
	.w3(32'hbcb81ce4),
	.w4(32'hbc8aa285),
	.w5(32'h3b7c0bc7),
	.w6(32'hbc58db83),
	.w7(32'hbc244c53),
	.w8(32'hb9a3af93),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ee6a5),
	.w1(32'h3b456f62),
	.w2(32'h3b8b6bd7),
	.w3(32'h3c2d5bb2),
	.w4(32'h3c7d934d),
	.w5(32'h3c68b349),
	.w6(32'h3b43f819),
	.w7(32'h3bd190fe),
	.w8(32'h3baf3f3b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d68d3),
	.w1(32'h3bff0d41),
	.w2(32'h3b1a38b9),
	.w3(32'h3ce0e95a),
	.w4(32'h3cb840f2),
	.w5(32'hbb910e43),
	.w6(32'h3cbb1c27),
	.w7(32'h3bd9e3cf),
	.w8(32'hbc06b37c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e2b8d),
	.w1(32'h3c207f56),
	.w2(32'h3b892080),
	.w3(32'hbbab7de8),
	.w4(32'h3b851245),
	.w5(32'h3a157923),
	.w6(32'hbc1b914a),
	.w7(32'hbb8e7528),
	.w8(32'hbc03a2cb),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05239e),
	.w1(32'h3bf5420b),
	.w2(32'h3c4a7f50),
	.w3(32'h3b607478),
	.w4(32'h3bb9d819),
	.w5(32'h3cc2a032),
	.w6(32'hbbd70ac9),
	.w7(32'h3a3ded5d),
	.w8(32'h3cbd7932),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca317dc),
	.w1(32'h3cbed66f),
	.w2(32'h3bb6d512),
	.w3(32'h3d29a0e8),
	.w4(32'h3cd24360),
	.w5(32'h3ae67e13),
	.w6(32'h3ce43aa5),
	.w7(32'h3cb6bec1),
	.w8(32'hbbc312e7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88be932),
	.w1(32'hbb32173a),
	.w2(32'h3b4d20ea),
	.w3(32'hbc6b451d),
	.w4(32'hbc2c298c),
	.w5(32'h394120f6),
	.w6(32'h3a1f6192),
	.w7(32'h3be8d442),
	.w8(32'h3b364424),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ed577),
	.w1(32'h3bd21853),
	.w2(32'h3be7e868),
	.w3(32'h3b50314f),
	.w4(32'h3b033b67),
	.w5(32'h3bf305b6),
	.w6(32'h3bd812fd),
	.w7(32'h3b71ef14),
	.w8(32'h3b89f522),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82bf2e),
	.w1(32'hbb805da6),
	.w2(32'h3b226d87),
	.w3(32'h3c6d5e01),
	.w4(32'hbb776a4f),
	.w5(32'hbb8e5239),
	.w6(32'h3c25b0b9),
	.w7(32'hba7c2bfa),
	.w8(32'hbbc202f4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915d799),
	.w1(32'h3b130959),
	.w2(32'hba51344a),
	.w3(32'hbc968f06),
	.w4(32'hbb997360),
	.w5(32'h3aab0e11),
	.w6(32'hbc6030ed),
	.w7(32'hbc030bc5),
	.w8(32'hbb0e667c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca7ca9),
	.w1(32'h3b80ef4b),
	.w2(32'hbc03a106),
	.w3(32'h3bdc3651),
	.w4(32'hbb8317ee),
	.w5(32'hbc8f744e),
	.w6(32'hbbfd3d51),
	.w7(32'hbc122383),
	.w8(32'hbc569c09),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19384c),
	.w1(32'hbca7c100),
	.w2(32'h3a072dd2),
	.w3(32'hbcb0be28),
	.w4(32'hbcd61b3b),
	.w5(32'hbad40914),
	.w6(32'hbc507c3b),
	.w7(32'hbc380ce1),
	.w8(32'hbae72b9b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29acf8),
	.w1(32'h3b4f3916),
	.w2(32'hbc03e6ec),
	.w3(32'hbafc9332),
	.w4(32'h3a9d35f3),
	.w5(32'hbbaa93d6),
	.w6(32'hbb15c869),
	.w7(32'h398b7f4c),
	.w8(32'h3bca157b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f6fdb),
	.w1(32'hbc8798a5),
	.w2(32'h3b3e3612),
	.w3(32'hbc8b9cc7),
	.w4(32'hbc935ecd),
	.w5(32'hbb2d96a5),
	.w6(32'hbbaaa924),
	.w7(32'hbbe9753b),
	.w8(32'h3b5f7418),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4efbcf),
	.w1(32'hbbd6a3b1),
	.w2(32'h3ab761de),
	.w3(32'h3b0fe782),
	.w4(32'hbc3c1788),
	.w5(32'h3c362141),
	.w6(32'hba0724a3),
	.w7(32'h3bd2fad6),
	.w8(32'h3c28f73d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87ddec),
	.w1(32'hbb98a5a6),
	.w2(32'hbc3f83b5),
	.w3(32'h3c961f7d),
	.w4(32'h3bd6d76d),
	.w5(32'h3b239b0f),
	.w6(32'h3c5c802a),
	.w7(32'h3b9d652f),
	.w8(32'hbaa09531),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe3b7e),
	.w1(32'hbc5c1b03),
	.w2(32'hba7818ca),
	.w3(32'hba566152),
	.w4(32'hbc350228),
	.w5(32'hbc2f87ef),
	.w6(32'h3b8286e5),
	.w7(32'hbc5e1b2f),
	.w8(32'hbaa13921),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1485c9),
	.w1(32'h3b0266e7),
	.w2(32'h3befa298),
	.w3(32'hbc3f0bae),
	.w4(32'hbc20f3df),
	.w5(32'h3c093356),
	.w6(32'h3b8d6a8b),
	.w7(32'hbacf1d98),
	.w8(32'h3c1468f4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38f438),
	.w1(32'hbbf5a9f9),
	.w2(32'h3bddce87),
	.w3(32'h3c2f9950),
	.w4(32'h3a55395e),
	.w5(32'h3b092d09),
	.w6(32'h3c6cfcbb),
	.w7(32'h3bc52afb),
	.w8(32'h3b276eb2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b794ca5),
	.w1(32'h3b5cefd4),
	.w2(32'h3a9ef442),
	.w3(32'hbb739526),
	.w4(32'hba19ad73),
	.w5(32'h3b330cac),
	.w6(32'hbb852994),
	.w7(32'hb9316db0),
	.w8(32'hbb9b43cb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb041b5),
	.w1(32'hbc08afc3),
	.w2(32'hbb9fa45d),
	.w3(32'hbc299741),
	.w4(32'hba8b1280),
	.w5(32'hbc3584a9),
	.w6(32'hbc8605ca),
	.w7(32'hbafe1e66),
	.w8(32'hbc804858),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc78a50),
	.w1(32'h3a7f74ab),
	.w2(32'hbc2fcdf1),
	.w3(32'hbc1fed32),
	.w4(32'hbbb54d65),
	.w5(32'hbcc39ae3),
	.w6(32'hbc0c9daf),
	.w7(32'hbbc81b08),
	.w8(32'hbc3fdc39),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93f7c1),
	.w1(32'hbcb57dac),
	.w2(32'h3bc6deb5),
	.w3(32'hbcdc4882),
	.w4(32'hbce997bb),
	.w5(32'hbb99b410),
	.w6(32'hbcbaf7bb),
	.w7(32'hbcd46148),
	.w8(32'hbb8693dd),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba453c35),
	.w1(32'h3b2e1869),
	.w2(32'h3b025096),
	.w3(32'hbbc59081),
	.w4(32'h3bf73d94),
	.w5(32'hba01b96b),
	.w6(32'h3b3c2e88),
	.w7(32'h3c3e0d7e),
	.w8(32'h38822770),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba173aa),
	.w1(32'h3bcd6fb4),
	.w2(32'h3b6280b6),
	.w3(32'hbc831e18),
	.w4(32'hba4c8da2),
	.w5(32'h3b86decf),
	.w6(32'hbcb2cfa1),
	.w7(32'hbbce8686),
	.w8(32'h3b1f7483),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea75a2),
	.w1(32'h39c256d4),
	.w2(32'hbb7b113e),
	.w3(32'hbb8be9e8),
	.w4(32'hbb537f5a),
	.w5(32'hbba20d04),
	.w6(32'hbaa94be2),
	.w7(32'hbad88bcd),
	.w8(32'hbc31454b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48c51a),
	.w1(32'hbbe7ccad),
	.w2(32'h3bd06f39),
	.w3(32'hbc9c0703),
	.w4(32'hbc333181),
	.w5(32'h3c076400),
	.w6(32'hbbfbe317),
	.w7(32'h3b92c3f2),
	.w8(32'h3bb7cf5a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2b62a),
	.w1(32'hbb151b0d),
	.w2(32'h3bdf0ba3),
	.w3(32'h3b918ed2),
	.w4(32'hbc22d5ec),
	.w5(32'hbb014eba),
	.w6(32'h3a492915),
	.w7(32'hbc6e1ba8),
	.w8(32'hbc129605),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4a258),
	.w1(32'h3c262583),
	.w2(32'h3c5aa7e3),
	.w3(32'hbb31b0eb),
	.w4(32'h3b9bb7ff),
	.w5(32'h3c684c63),
	.w6(32'hbc9af89c),
	.w7(32'hbbff94e3),
	.w8(32'h3bdba87d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9432cc),
	.w1(32'h3c894788),
	.w2(32'h3b96d475),
	.w3(32'h3c877ea3),
	.w4(32'h3ca2be10),
	.w5(32'h3ac2b813),
	.w6(32'h3c2207e2),
	.w7(32'h3be1523b),
	.w8(32'h3aa1ce47),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d5d25),
	.w1(32'hbb4a6a14),
	.w2(32'h3a69f0e1),
	.w3(32'hbb88171f),
	.w4(32'hbb963614),
	.w5(32'h3a6212a2),
	.w6(32'h3a5f7094),
	.w7(32'hbac05e09),
	.w8(32'h3b10c779),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cd2ee),
	.w1(32'hb9d4355a),
	.w2(32'h3baab596),
	.w3(32'hbb696e7b),
	.w4(32'hbbacc270),
	.w5(32'hbbd19c64),
	.w6(32'h3ae2e048),
	.w7(32'hbaeee04f),
	.w8(32'hbbbcfa95),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d62cc5),
	.w1(32'hbbc2c841),
	.w2(32'hba8c1f0a),
	.w3(32'hbc072d3a),
	.w4(32'hbb780202),
	.w5(32'hbbf0d2dc),
	.w6(32'hbb879d33),
	.w7(32'h3c4d5d0d),
	.w8(32'hbc26f205),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9995a3d),
	.w1(32'h3a8aa789),
	.w2(32'hbb22a56f),
	.w3(32'hbbfb6d32),
	.w4(32'hbb316ec8),
	.w5(32'hbbb31b1a),
	.w6(32'hbc33a87e),
	.w7(32'hba49cafa),
	.w8(32'hbabcfec6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41d5c6),
	.w1(32'hbb853ccc),
	.w2(32'hbbe74c82),
	.w3(32'hbc29e244),
	.w4(32'hbbf4a049),
	.w5(32'hbc5c66e0),
	.w6(32'hbbc4ffea),
	.w7(32'hba5ef448),
	.w8(32'hbb2d5f43),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90d66b),
	.w1(32'hbc3a6c7d),
	.w2(32'h3b47cb13),
	.w3(32'hbcb9b7f8),
	.w4(32'hbcab9ba4),
	.w5(32'hbb816c78),
	.w6(32'hbc708162),
	.w7(32'hbc3b4681),
	.w8(32'hba8395ae),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade7279),
	.w1(32'hbc1ff192),
	.w2(32'h3b912bcb),
	.w3(32'hbc1bbddd),
	.w4(32'hbbc1499b),
	.w5(32'h3acec7cd),
	.w6(32'hbabc8981),
	.w7(32'h3b065810),
	.w8(32'hbba8ac68),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7f56),
	.w1(32'hbc388f98),
	.w2(32'h3c352cfb),
	.w3(32'h3c195145),
	.w4(32'hbc211d97),
	.w5(32'h3c549379),
	.w6(32'h3b7b00ec),
	.w7(32'hbaa6807d),
	.w8(32'h3c7ae291),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6164a4),
	.w1(32'h3c5319ab),
	.w2(32'h3bc39325),
	.w3(32'h3cabd8f1),
	.w4(32'h3c463496),
	.w5(32'h3ce256b4),
	.w6(32'h3c8c3d80),
	.w7(32'h3b477e51),
	.w8(32'h3c92d65b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdd5cbe),
	.w1(32'h3cdce398),
	.w2(32'h3b112593),
	.w3(32'h3d0c4f1b),
	.w4(32'h3caa0251),
	.w5(32'hb96b779e),
	.w6(32'h3cc8fc58),
	.w7(32'h3be6cf54),
	.w8(32'h3abda564),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf09725),
	.w1(32'h3b4be3b5),
	.w2(32'h3ca429b6),
	.w3(32'hbb16f5d1),
	.w4(32'hbaad3946),
	.w5(32'h3c09409b),
	.w6(32'hbc61d96f),
	.w7(32'hbc13ef1e),
	.w8(32'h3c179db5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc1a04),
	.w1(32'h3bcb25aa),
	.w2(32'h3c1a5a3b),
	.w3(32'h3bf07a06),
	.w4(32'h3b320d56),
	.w5(32'h3c9c481b),
	.w6(32'h38a4b077),
	.w7(32'h3991f15b),
	.w8(32'h3c093fdf),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2de60c),
	.w1(32'h3b517f4b),
	.w2(32'h3b800dd9),
	.w3(32'h3c984b06),
	.w4(32'h3c64d679),
	.w5(32'hbb61ac64),
	.w6(32'h3c382e03),
	.w7(32'h3c09a76e),
	.w8(32'hbb3556e7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25a64b),
	.w1(32'h39d125fd),
	.w2(32'hba5b5204),
	.w3(32'hbb9bff0a),
	.w4(32'h3aab3af4),
	.w5(32'hbb87dc35),
	.w6(32'hbb14a69b),
	.w7(32'h3b03ba1e),
	.w8(32'hbb9256c5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e07864),
	.w1(32'hb9daa47c),
	.w2(32'hbada278a),
	.w3(32'hbb524126),
	.w4(32'h3b41f74d),
	.w5(32'h3bf1b3e8),
	.w6(32'hbb52ea73),
	.w7(32'hbb146a00),
	.w8(32'h3c43a345),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7b206),
	.w1(32'hbc300ce4),
	.w2(32'hbc4f6344),
	.w3(32'h3c74d11d),
	.w4(32'hbba10040),
	.w5(32'hbc895793),
	.w6(32'h3c83df28),
	.w7(32'hbae240ae),
	.w8(32'hbc85f7fd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7aa47),
	.w1(32'hbcd542f2),
	.w2(32'hbbe70caf),
	.w3(32'hbd00450b),
	.w4(32'hbceffd94),
	.w5(32'h3bd56625),
	.w6(32'hbcaef4c0),
	.w7(32'hbcd6e3e2),
	.w8(32'h3c056c13),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac8570),
	.w1(32'h3be24617),
	.w2(32'hba0ab4c6),
	.w3(32'h3c4ad912),
	.w4(32'h3c0af9ab),
	.w5(32'hbc1fd65f),
	.w6(32'h3c3f296e),
	.w7(32'h3aa75da7),
	.w8(32'hbb134100),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc589334),
	.w1(32'hbb828d82),
	.w2(32'h39d1e82b),
	.w3(32'hbc6bce27),
	.w4(32'hbc67bea1),
	.w5(32'hba2a53df),
	.w6(32'hba003c47),
	.w7(32'hbb5ba156),
	.w8(32'hbb8dd6f6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d5bbb),
	.w1(32'h3c82bd2f),
	.w2(32'h3c1c3093),
	.w3(32'h3c435e8a),
	.w4(32'h3c09ea53),
	.w5(32'h3beda8dd),
	.w6(32'h3b668212),
	.w7(32'h3be0eeb3),
	.w8(32'h3b0eecb6),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7329d),
	.w1(32'hbb54b33b),
	.w2(32'hbc60b334),
	.w3(32'h3be19986),
	.w4(32'h3b5c46a0),
	.w5(32'hbb93ccf6),
	.w6(32'h3c00eb2c),
	.w7(32'h3bb6ffb7),
	.w8(32'h3bfaf5ba),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbec17),
	.w1(32'hbca49dd8),
	.w2(32'h3bbfa3a5),
	.w3(32'hbc4fb68a),
	.w4(32'hbcf6fa68),
	.w5(32'h3b216e56),
	.w6(32'hbb5ce06f),
	.w7(32'hbc70aedb),
	.w8(32'hba4880ad),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92c933),
	.w1(32'hb9cb33f0),
	.w2(32'h3bd7bd35),
	.w3(32'h3a73f5c8),
	.w4(32'hbb9a4111),
	.w5(32'h3c224838),
	.w6(32'h3c427422),
	.w7(32'h3c2d0ad7),
	.w8(32'h3b5f50e9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8732f),
	.w1(32'hbae14491),
	.w2(32'h3b85363c),
	.w3(32'h3c54daea),
	.w4(32'h3aa38dd1),
	.w5(32'h3acbc1d6),
	.w6(32'h3c2dc437),
	.w7(32'h3bdfa0eb),
	.w8(32'h3c06f69c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38f345),
	.w1(32'h3b9c7a8e),
	.w2(32'h3b992a8e),
	.w3(32'hbbcd8a36),
	.w4(32'h3bda7c1e),
	.w5(32'h3b97f5c8),
	.w6(32'hbafcc2c6),
	.w7(32'hbb428cc3),
	.w8(32'h3b7044cb),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9ef5b),
	.w1(32'h3b2d5f54),
	.w2(32'h3c526d0c),
	.w3(32'h3c0a5354),
	.w4(32'h3b7788b4),
	.w5(32'h3ca18986),
	.w6(32'h3bc2c6db),
	.w7(32'h3b5e3568),
	.w8(32'h3c2922c3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1288e0),
	.w1(32'h3c1d6f9a),
	.w2(32'h3c423961),
	.w3(32'h3cae9105),
	.w4(32'h3c4ec7a5),
	.w5(32'h3cb3695e),
	.w6(32'h3c05f3d4),
	.w7(32'h3b60611c),
	.w8(32'h3cb9de91),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93a95f),
	.w1(32'h3caeb698),
	.w2(32'hbba337e3),
	.w3(32'h3cd4bb5e),
	.w4(32'h3ca7d874),
	.w5(32'hbc50901e),
	.w6(32'h3cc3eba8),
	.w7(32'h3c10bab4),
	.w8(32'hba16a93f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f61b0),
	.w1(32'hbc137237),
	.w2(32'h3a866290),
	.w3(32'hbce97e9c),
	.w4(32'hbc642837),
	.w5(32'h3ac39757),
	.w6(32'hbc84b43b),
	.w7(32'hbc209adf),
	.w8(32'h3b679713),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac438f9),
	.w1(32'hbb4c0b30),
	.w2(32'hbb88c0aa),
	.w3(32'hbaaca725),
	.w4(32'hba1d7ef1),
	.w5(32'hbad1299f),
	.w6(32'h3ad28e12),
	.w7(32'h3ad2c20f),
	.w8(32'h3b4592b0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc34f2),
	.w1(32'hbc1126d9),
	.w2(32'h3be03f0f),
	.w3(32'hbbe35f22),
	.w4(32'hbbfb2ef8),
	.w5(32'h3ad8d164),
	.w6(32'hb936fc70),
	.w7(32'hbb31d603),
	.w8(32'hbc481009),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50f307),
	.w1(32'h3c167dac),
	.w2(32'h3a31c465),
	.w3(32'hbc996a39),
	.w4(32'h3bd61ccd),
	.w5(32'h39cb4958),
	.w6(32'hbcaa7889),
	.w7(32'hbbdda78d),
	.w8(32'h3b87c07b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95e741),
	.w1(32'h3bde2086),
	.w2(32'h3b8341cd),
	.w3(32'h3b849f78),
	.w4(32'h3a89fcc6),
	.w5(32'hbb9a5cad),
	.w6(32'h3b6f3094),
	.w7(32'hbaf01674),
	.w8(32'h39a2b943),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf576fb),
	.w1(32'hbae3a2eb),
	.w2(32'h3b898847),
	.w3(32'hb8a046a6),
	.w4(32'h3c524838),
	.w5(32'h3ca6675b),
	.w6(32'h3bd02f37),
	.w7(32'h3c1eed63),
	.w8(32'h3c771c95),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c600fd2),
	.w1(32'h3cad5e83),
	.w2(32'h3c01b254),
	.w3(32'h3cfa6e4d),
	.w4(32'h3cfe12de),
	.w5(32'h3ca20e43),
	.w6(32'h3cb905c1),
	.w7(32'h3cab0bdf),
	.w8(32'h3c8dd114),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf3e0d5),
	.w1(32'h3cb9bc00),
	.w2(32'hbc0211af),
	.w3(32'h3d29089c),
	.w4(32'h3d0345f9),
	.w5(32'hbc199dea),
	.w6(32'h3ccf3296),
	.w7(32'h3c6282ca),
	.w8(32'hbc244964),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule