module layer_8_featuremap_51(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b6dc0),
	.w1(32'hbb9d4afd),
	.w2(32'hbc165cdc),
	.w3(32'h3a09c88c),
	.w4(32'hbbb6a2e3),
	.w5(32'hbc35871c),
	.w6(32'hbadda1a2),
	.w7(32'hbc31e2a9),
	.w8(32'hbb532094),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1bb6f),
	.w1(32'hbacb55b6),
	.w2(32'hbbb33c5d),
	.w3(32'h3bb7fb85),
	.w4(32'hba9e2bdb),
	.w5(32'hbb950c73),
	.w6(32'hbb1dd22d),
	.w7(32'hbbecee80),
	.w8(32'h3b516815),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13bcae),
	.w1(32'h3b061dbf),
	.w2(32'hbbb4f26b),
	.w3(32'h3c08febc),
	.w4(32'h3ac71711),
	.w5(32'hbb899d25),
	.w6(32'hbafa153e),
	.w7(32'hbc27d42a),
	.w8(32'hbc08e072),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba4606),
	.w1(32'h3b378869),
	.w2(32'hbb7b4071),
	.w3(32'h3b3aefa4),
	.w4(32'h3b778ac6),
	.w5(32'hbaa825d5),
	.w6(32'hba613356),
	.w7(32'hbaa42207),
	.w8(32'h3bed3834),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3f176),
	.w1(32'hbb6aae90),
	.w2(32'hbc2e58f9),
	.w3(32'h3b7cdf26),
	.w4(32'hbb1e3bb4),
	.w5(32'hbc18dbe1),
	.w6(32'hbb848b30),
	.w7(32'hbc3f45f5),
	.w8(32'h3d1f01d0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d87639e),
	.w1(32'h3b894625),
	.w2(32'hbd162ea4),
	.w3(32'h3d485bcd),
	.w4(32'hb9e255d8),
	.w5(32'hbcd8b2b8),
	.w6(32'hbc76dd35),
	.w7(32'hbd252e1d),
	.w8(32'h3c39358f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfed9fd),
	.w1(32'hba190fc1),
	.w2(32'hbbed4768),
	.w3(32'h3bd3e93b),
	.w4(32'h399890b5),
	.w5(32'hbbb9db93),
	.w6(32'hba7f3ed8),
	.w7(32'hbbb8d53e),
	.w8(32'h3bbb37c2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb4ed8),
	.w1(32'h3aafa842),
	.w2(32'hbbf9ec7b),
	.w3(32'h3b55c84d),
	.w4(32'hb9b89c40),
	.w5(32'hbb9db3e1),
	.w6(32'hbb5242e8),
	.w7(32'hbc5edf3a),
	.w8(32'h3bf4e25a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c798f31),
	.w1(32'h3c11c54e),
	.w2(32'hbaeb745d),
	.w3(32'h3c81be1a),
	.w4(32'h3bfef373),
	.w5(32'hba734555),
	.w6(32'h38e0b622),
	.w7(32'hbc1a2752),
	.w8(32'hbc85f49c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f99d1),
	.w1(32'hbc3bfde0),
	.w2(32'hbc2f01a4),
	.w3(32'h3a07ca41),
	.w4(32'hbbf7d5fd),
	.w5(32'hbc6c4a34),
	.w6(32'hbc446158),
	.w7(32'hbc6d8467),
	.w8(32'h3b8acccf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49c346),
	.w1(32'hbbaa6097),
	.w2(32'hbc920d6c),
	.w3(32'h3b41aa07),
	.w4(32'hbb0f5caf),
	.w5(32'hbc56c336),
	.w6(32'hbab749c0),
	.w7(32'hbc90fbd0),
	.w8(32'hbb008c47),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c29ae),
	.w1(32'h3aca35e8),
	.w2(32'hbbafc28b),
	.w3(32'h3c0549b9),
	.w4(32'hba31cee7),
	.w5(32'hbb9e3e81),
	.w6(32'h3af8f203),
	.w7(32'hbbf6cef2),
	.w8(32'hb93112a5),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffa46a),
	.w1(32'h3985158a),
	.w2(32'hbb992e95),
	.w3(32'h3bc0fecb),
	.w4(32'hbb203234),
	.w5(32'hbbe69617),
	.w6(32'hbb8fbe14),
	.w7(32'hbc430c24),
	.w8(32'h3d3c3b6f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8d2951),
	.w1(32'hba4c12cd),
	.w2(32'hbd2f7939),
	.w3(32'h3d66fbab),
	.w4(32'hba065f99),
	.w5(32'hbd0c8e86),
	.w6(32'hbc6aa498),
	.w7(32'hbd3413c1),
	.w8(32'h3ca1b010),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d022aa2),
	.w1(32'hbb2def26),
	.w2(32'hbccef1af),
	.w3(32'h3cdd5871),
	.w4(32'hb9c9dd56),
	.w5(32'hbc96dfba),
	.w6(32'hbc0854fd),
	.w7(32'hbccbf7a6),
	.w8(32'h39cf7501),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad823b9),
	.w1(32'hbb5631dc),
	.w2(32'hbb9b9e86),
	.w3(32'h395d27cf),
	.w4(32'hbb403f17),
	.w5(32'hbb5cb87f),
	.w6(32'hbb6ac43f),
	.w7(32'hbb986294),
	.w8(32'h3b6920a0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51eead),
	.w1(32'h3b89d47e),
	.w2(32'hbbcb3da6),
	.w3(32'h3ad84864),
	.w4(32'h3a915f74),
	.w5(32'hbc0c84f8),
	.w6(32'h3b86970a),
	.w7(32'h36994860),
	.w8(32'h3b1381bf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab6c45),
	.w1(32'hb9899c89),
	.w2(32'hbbc97faa),
	.w3(32'h3bb122a5),
	.w4(32'hbb3f974b),
	.w5(32'hbbdf7fca),
	.w6(32'hbb5e53b9),
	.w7(32'hbc2c1e5b),
	.w8(32'hbaae79b3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba27d16),
	.w1(32'hbbe26c5f),
	.w2(32'hbbee413b),
	.w3(32'hbae594a9),
	.w4(32'hbbb78fc6),
	.w5(32'hbbd505dd),
	.w6(32'h3c5b1949),
	.w7(32'hbca097fa),
	.w8(32'hbc8f9b9f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52652b),
	.w1(32'hbae172dd),
	.w2(32'hbca79a96),
	.w3(32'hbc9b02a6),
	.w4(32'hbbd47589),
	.w5(32'hbc886e18),
	.w6(32'hbbd46c82),
	.w7(32'hbcc512f6),
	.w8(32'hbbd01139),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc404cae),
	.w1(32'h3b85defe),
	.w2(32'h3c88ad9d),
	.w3(32'hbc336f53),
	.w4(32'h3b167e49),
	.w5(32'h3c62af48),
	.w6(32'h3c3342cd),
	.w7(32'h3cabd398),
	.w8(32'h3c5afc2e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8dab6),
	.w1(32'hbb8fea68),
	.w2(32'hbc4ce2ab),
	.w3(32'h3bd17734),
	.w4(32'hbb7d6cbe),
	.w5(32'hbc47a52c),
	.w6(32'hbb8e72fc),
	.w7(32'hbc6a1fd3),
	.w8(32'hbcdc17b4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd44d638),
	.w1(32'hbb745e25),
	.w2(32'h3d72486a),
	.w3(32'hbd2b0eb5),
	.w4(32'hbc6d8502),
	.w5(32'h3d131f42),
	.w6(32'h3bda04c0),
	.w7(32'h3d162713),
	.w8(32'hbc5f3fc2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a7c78),
	.w1(32'hbadf4e1d),
	.w2(32'hbb6214ab),
	.w3(32'hba9e8bfe),
	.w4(32'hbb9d511b),
	.w5(32'hbb1983c0),
	.w6(32'hbbccf7f5),
	.w7(32'hbbcd0e13),
	.w8(32'hb78a8734),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19d0a1),
	.w1(32'hbb02eac6),
	.w2(32'hbb3270a3),
	.w3(32'hbbfa047b),
	.w4(32'hbbcf35c7),
	.w5(32'hbbba2160),
	.w6(32'h3ac92709),
	.w7(32'hba1d1bf1),
	.w8(32'hbcc9073d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd17f2c3),
	.w1(32'hbacac38c),
	.w2(32'h3d52007d),
	.w3(32'hbd0d01be),
	.w4(32'hbc2f9839),
	.w5(32'h3d13b083),
	.w6(32'h3bb4c365),
	.w7(32'h3d182b61),
	.w8(32'hbceac5d1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec25dd),
	.w1(32'h39491b23),
	.w2(32'h3d27bcfa),
	.w3(32'hbce79937),
	.w4(32'hbc0f2063),
	.w5(32'h3ce09d9f),
	.w6(32'h3ab42493),
	.w7(32'h3d0e3645),
	.w8(32'hbc382024),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1464fe),
	.w1(32'hbbdb82e0),
	.w2(32'h3d83a74f),
	.w3(32'hbd0325eb),
	.w4(32'h3918b54e),
	.w5(32'h3d637c0e),
	.w6(32'h3d783c95),
	.w7(32'h3d6f0dc7),
	.w8(32'hbd3450a4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca372d6),
	.w1(32'hbc68cc7a),
	.w2(32'hbc5314f4),
	.w3(32'hbcb25325),
	.w4(32'hbca13617),
	.w5(32'hbc9bc66d),
	.w6(32'hbc720b0f),
	.w7(32'hbcb8215b),
	.w8(32'h3a74b292),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b6a1a),
	.w1(32'h39873913),
	.w2(32'hbbaa49ba),
	.w3(32'h3b91a542),
	.w4(32'h3a95f0cb),
	.w5(32'hbb3a28fc),
	.w6(32'hba55d209),
	.w7(32'hbbaf8b9c),
	.w8(32'h3c0f1dec),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad385e1),
	.w1(32'h3a6ddb9e),
	.w2(32'hbc28fa92),
	.w3(32'hbc2cf9f3),
	.w4(32'h3c32e501),
	.w5(32'h3c025e45),
	.w6(32'h3b12b5d9),
	.w7(32'hbc01cc6e),
	.w8(32'hbca10abf),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce4396f),
	.w1(32'hbb3fb4ef),
	.w2(32'h3c72dcea),
	.w3(32'hbcc2869d),
	.w4(32'hbbca5920),
	.w5(32'h3c33245e),
	.w6(32'h3b825320),
	.w7(32'h3c889e1e),
	.w8(32'h3a36b526),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b4c87),
	.w1(32'h3b31329b),
	.w2(32'hbae2a52a),
	.w3(32'hbb934dcf),
	.w4(32'hbaf26cfc),
	.w5(32'h3bafa775),
	.w6(32'hbb04334a),
	.w7(32'h3ba13c0f),
	.w8(32'h3b087f20),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070272),
	.w1(32'hb8481ba4),
	.w2(32'h3b70de5e),
	.w3(32'hbb1a7f2b),
	.w4(32'h3acf20d2),
	.w5(32'h3b86739b),
	.w6(32'hbb8761d5),
	.w7(32'hbbb55844),
	.w8(32'h3d23a6a2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d85832c),
	.w1(32'h3b83e4ee),
	.w2(32'hbd01b294),
	.w3(32'h3d553253),
	.w4(32'h3a3b4661),
	.w5(32'hbcdb6bef),
	.w6(32'hbc2366e5),
	.w7(32'hbd036a9a),
	.w8(32'h3c3f8856),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae952e4),
	.w1(32'hbbadcc63),
	.w2(32'hbbc48979),
	.w3(32'h3b5e7170),
	.w4(32'hba571b15),
	.w5(32'hbb568186),
	.w6(32'h3b119ca7),
	.w7(32'hbbba980f),
	.w8(32'hbc0dcdaa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ccae2),
	.w1(32'hbb8d5b3e),
	.w2(32'h3b1177f0),
	.w3(32'hbc072f47),
	.w4(32'hbbc0f240),
	.w5(32'hbb6625ae),
	.w6(32'hbae7b6f3),
	.w7(32'h3b275480),
	.w8(32'h3bca0618),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b810aff),
	.w1(32'hbad1d78c),
	.w2(32'hbc1ae688),
	.w3(32'h3b806edf),
	.w4(32'hb9a41e0a),
	.w5(32'hbbe959d7),
	.w6(32'hbb4ed804),
	.w7(32'hbc147062),
	.w8(32'h3ce353d6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d513e2d),
	.w1(32'hbbf8b1b9),
	.w2(32'hbd2aeb86),
	.w3(32'h3d2b7be3),
	.w4(32'hbb5ffd95),
	.w5(32'hbcfa5079),
	.w6(32'hbc825a0a),
	.w7(32'hbd2740be),
	.w8(32'hbc4a136d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c9e19),
	.w1(32'hbbbcee64),
	.w2(32'h3c41e723),
	.w3(32'hbc8fe9a5),
	.w4(32'hbc0b63f2),
	.w5(32'h3bdaeb88),
	.w6(32'hba99089e),
	.w7(32'h3c5bcbec),
	.w8(32'hbc2e7a16),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59e70a),
	.w1(32'h3ad443fb),
	.w2(32'h3cd4d4c7),
	.w3(32'hbc7bbb77),
	.w4(32'hbc3b1fad),
	.w5(32'h3bb153fe),
	.w6(32'h3bc65e0c),
	.w7(32'h3bfb6a8e),
	.w8(32'hbc68a9cf),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba250592),
	.w1(32'hb97b3989),
	.w2(32'h3b115220),
	.w3(32'hb94781c5),
	.w4(32'hb925e196),
	.w5(32'h3ad50a1c),
	.w6(32'h3aa39dc9),
	.w7(32'hb9d15ea7),
	.w8(32'h39cf0412),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d578c8),
	.w1(32'h379def5e),
	.w2(32'h3afd7b3d),
	.w3(32'hb9a805d8),
	.w4(32'hb96b1790),
	.w5(32'h3a79c29e),
	.w6(32'hba3b0e7b),
	.w7(32'h3ad28e3b),
	.w8(32'h39d7c709),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad4a3e),
	.w1(32'hbac515ab),
	.w2(32'hb92b8834),
	.w3(32'hbb1eba2e),
	.w4(32'hbb0cf6da),
	.w5(32'hbaaa8b9c),
	.w6(32'h3a365531),
	.w7(32'hbb5cdfbc),
	.w8(32'hbbcc1c20),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8be41),
	.w1(32'hba833891),
	.w2(32'h3b729868),
	.w3(32'hbb81ad16),
	.w4(32'hbacd70e3),
	.w5(32'h3b58d5e2),
	.w6(32'h3b2525fa),
	.w7(32'hbbed1d30),
	.w8(32'hbc0186e7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aacd9d),
	.w1(32'h3b04cd0c),
	.w2(32'h3b809724),
	.w3(32'h3aadff74),
	.w4(32'h3abd78cd),
	.w5(32'h3b28ab6a),
	.w6(32'h3b40b764),
	.w7(32'hb9328e10),
	.w8(32'h39eba948),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b547a),
	.w1(32'h39d25167),
	.w2(32'hba329fa7),
	.w3(32'hb9e6b9da),
	.w4(32'hbab9b082),
	.w5(32'hbaf777da),
	.w6(32'hba3a7ad8),
	.w7(32'hba255954),
	.w8(32'h3a924602),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39794a),
	.w1(32'hb94df86a),
	.w2(32'h3b86f2d3),
	.w3(32'hbad29c26),
	.w4(32'h3b1b2308),
	.w5(32'h3bc77584),
	.w6(32'h3bbc1b1b),
	.w7(32'h38a45762),
	.w8(32'hbb2a043c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c5749),
	.w1(32'hbb415c16),
	.w2(32'hbaebc0d5),
	.w3(32'h3a22d682),
	.w4(32'hbb3d89b5),
	.w5(32'hbb18ccdc),
	.w6(32'hbafe4860),
	.w7(32'hbb471ec2),
	.w8(32'hbb6674b3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9939c5a),
	.w1(32'h39c625f6),
	.w2(32'h3806cba4),
	.w3(32'h398e05db),
	.w4(32'hb9a7e72c),
	.w5(32'hb83ff57a),
	.w6(32'h3b28b27a),
	.w7(32'hbb898e5b),
	.w8(32'hbb9541ce),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e775),
	.w1(32'h3ae7cfef),
	.w2(32'h3ba71d55),
	.w3(32'hbb573849),
	.w4(32'hbaa27e65),
	.w5(32'hba646d7a),
	.w6(32'hbb451dab),
	.w7(32'h3aab36ee),
	.w8(32'h3a78db68),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a8197),
	.w1(32'hbbcec5fa),
	.w2(32'h3b180f7a),
	.w3(32'hbc5060b7),
	.w4(32'hbbc53942),
	.w5(32'h3b2bab4a),
	.w6(32'hbaa6d615),
	.w7(32'hbc85c7cb),
	.w8(32'hbc518207),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad28e3),
	.w1(32'hb9fca7f9),
	.w2(32'h3a4d4bf5),
	.w3(32'hbabadd5b),
	.w4(32'h39eb26be),
	.w5(32'h3ac15d8d),
	.w6(32'h3b3b3a77),
	.w7(32'h3a0207ba),
	.w8(32'hbb79933b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c4d8c),
	.w1(32'hbaffe7f9),
	.w2(32'hba98f4bb),
	.w3(32'hba8f8ee8),
	.w4(32'hbb8731f4),
	.w5(32'hbc12d747),
	.w6(32'hbaf2c03a),
	.w7(32'hbb4047b6),
	.w8(32'hbb3fbeb9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aade32),
	.w1(32'h3a91f0a9),
	.w2(32'h388695d4),
	.w3(32'hb981c5ad),
	.w4(32'h3994cc7c),
	.w5(32'hb9dde65d),
	.w6(32'h3aae7d3c),
	.w7(32'h3a70bf36),
	.w8(32'hbade929d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6ec93),
	.w1(32'h393bf9a2),
	.w2(32'h3c33e857),
	.w3(32'hbaecc107),
	.w4(32'hb9bfc4f0),
	.w5(32'h3c005499),
	.w6(32'h3bb373d6),
	.w7(32'h3a8a7f28),
	.w8(32'hbbee98e7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ffe38f),
	.w1(32'h3b6804f9),
	.w2(32'h3b8e11bc),
	.w3(32'h3a8b7ac4),
	.w4(32'h3aeaf68f),
	.w5(32'h3ab4c0c6),
	.w6(32'h39ff51fb),
	.w7(32'h3b443d05),
	.w8(32'h3ba5f44d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8dc34),
	.w1(32'h3a87b4aa),
	.w2(32'h3b191102),
	.w3(32'hba4eb6ae),
	.w4(32'hba44a796),
	.w5(32'h3b042be7),
	.w6(32'h3a5511c9),
	.w7(32'hbc179b45),
	.w8(32'hbae89bdc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4e3ae),
	.w1(32'hbb96ba66),
	.w2(32'hba223282),
	.w3(32'hba7d3bca),
	.w4(32'hbb52cf5c),
	.w5(32'hba194843),
	.w6(32'hb8ea558e),
	.w7(32'hba923540),
	.w8(32'hbbe9ddbf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedffc7),
	.w1(32'hbb5dde77),
	.w2(32'hbabf131b),
	.w3(32'hbaa4d3aa),
	.w4(32'hbb84d6b5),
	.w5(32'hbb42e974),
	.w6(32'hbb79bcd8),
	.w7(32'hb9e32996),
	.w8(32'h3a726927),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074132),
	.w1(32'hbade091a),
	.w2(32'hba0c6506),
	.w3(32'hbab182be),
	.w4(32'hba367752),
	.w5(32'hbab3cf7c),
	.w6(32'hba90e276),
	.w7(32'hba094bac),
	.w8(32'h3a7f6145),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b279f),
	.w1(32'h3a9b1fb9),
	.w2(32'h3a091c1c),
	.w3(32'h395f62c1),
	.w4(32'h39a437d6),
	.w5(32'hb779ee3e),
	.w6(32'h3a5b52dc),
	.w7(32'hb83e8d4f),
	.w8(32'hba5ec82c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33bde3),
	.w1(32'h3b2a5eb4),
	.w2(32'h3bc2988c),
	.w3(32'hba79e37f),
	.w4(32'hbbaf126a),
	.w5(32'hbb5ac8ab),
	.w6(32'h3b104bcc),
	.w7(32'hbb68ecf3),
	.w8(32'hbb1087fc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc12990),
	.w1(32'h3b4ff6e3),
	.w2(32'h3af238bc),
	.w3(32'h3b4e8555),
	.w4(32'h3a9e16c9),
	.w5(32'h3b14db7e),
	.w6(32'h3b05f467),
	.w7(32'hba693caf),
	.w8(32'hbaa8af24),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27cd16),
	.w1(32'h3ae54b11),
	.w2(32'h3958e7f6),
	.w3(32'hb9e43c35),
	.w4(32'h39b3f235),
	.w5(32'hb9ebab15),
	.w6(32'h3a626e28),
	.w7(32'h3977f16c),
	.w8(32'hba64f81d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49b798),
	.w1(32'hba76a2b2),
	.w2(32'h3b3bcf9f),
	.w3(32'hbb263a0d),
	.w4(32'hbaece4ad),
	.w5(32'h3a9ef895),
	.w6(32'hba0a4210),
	.w7(32'hbb8fe019),
	.w8(32'hbb6aafcd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9492d93),
	.w1(32'hbaac0bce),
	.w2(32'h3a60cd32),
	.w3(32'hbaa6f207),
	.w4(32'hbaf68751),
	.w5(32'h383804d4),
	.w6(32'hbb2dda2a),
	.w7(32'hbb73caf1),
	.w8(32'hba215128),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b96d4),
	.w1(32'h3b8e6cac),
	.w2(32'h3c0654f7),
	.w3(32'h3ba95883),
	.w4(32'h3b22769a),
	.w5(32'h3b69ac07),
	.w6(32'h3bcecd88),
	.w7(32'h3b742117),
	.w8(32'h3af435ef),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba434b2b),
	.w1(32'hba1e777a),
	.w2(32'hba33ab1a),
	.w3(32'hba1840c1),
	.w4(32'hba16c928),
	.w5(32'hba1f95f1),
	.w6(32'hba059f7b),
	.w7(32'hba2cd6ef),
	.w8(32'h3ba925f5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003c49),
	.w1(32'hbbedf67a),
	.w2(32'h3aa1858d),
	.w3(32'h3ab96b25),
	.w4(32'h3baec5f0),
	.w5(32'h3c0b64de),
	.w6(32'h3c67170c),
	.w7(32'h3b91da3c),
	.w8(32'hbc8b2197),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba916f25),
	.w1(32'hba82f13c),
	.w2(32'hba50d7d8),
	.w3(32'hba974f78),
	.w4(32'hba80be50),
	.w5(32'hba4ac84e),
	.w6(32'hba826a73),
	.w7(32'hba6606bf),
	.w8(32'hba8b64d1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb297855),
	.w1(32'hbb2212d0),
	.w2(32'hb9e32a6c),
	.w3(32'hbb23087a),
	.w4(32'hbb1f83b3),
	.w5(32'hbada5b34),
	.w6(32'hba794315),
	.w7(32'hbb7f4bfe),
	.w8(32'hbb93ae6e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17cae7),
	.w1(32'hbb1804cc),
	.w2(32'hbaeaed24),
	.w3(32'hbb062018),
	.w4(32'hbb0736da),
	.w5(32'hbad9b6cc),
	.w6(32'hbaf9751a),
	.w7(32'hbad353b5),
	.w8(32'h3a865081),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfc47e),
	.w1(32'h3ba5a875),
	.w2(32'h3c00d4bc),
	.w3(32'h3b9fdc23),
	.w4(32'hb9ee552d),
	.w5(32'h3b1e544b),
	.w6(32'h3b985fe2),
	.w7(32'h3b70cb84),
	.w8(32'hba403aa2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba974dac),
	.w1(32'hbab59447),
	.w2(32'hba473803),
	.w3(32'hbaa33cd6),
	.w4(32'hbaa4a817),
	.w5(32'hba4ac2de),
	.w6(32'hbaa10705),
	.w7(32'hba31902b),
	.w8(32'hba454dc9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb950cb4),
	.w1(32'hbb7652ef),
	.w2(32'hba59dfbe),
	.w3(32'hbb5f68b0),
	.w4(32'hbb5063ab),
	.w5(32'hba9dee77),
	.w6(32'hba2bca6a),
	.w7(32'hbb2868a8),
	.w8(32'hbb123508),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba955ce3),
	.w1(32'hba9d2fa2),
	.w2(32'hba72efa9),
	.w3(32'hba9bee63),
	.w4(32'hbaa1b987),
	.w5(32'hba6a41b5),
	.w6(32'hba982996),
	.w7(32'hba6f0bab),
	.w8(32'h3bd58f13),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03c38f),
	.w1(32'hbb5d613d),
	.w2(32'h3b8be263),
	.w3(32'h39ff8f22),
	.w4(32'hba6e9ca3),
	.w5(32'h3b559a8e),
	.w6(32'h3c0b14ce),
	.w7(32'h3b176141),
	.w8(32'hbbf0e843),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb65778),
	.w1(32'h3bcd02cd),
	.w2(32'h3c31cf1e),
	.w3(32'h3b8316a5),
	.w4(32'h3bc867ab),
	.w5(32'h3c2c0511),
	.w6(32'h3bec5721),
	.w7(32'h3bec134b),
	.w8(32'h3b8995c5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e61c52),
	.w1(32'h3931e2a6),
	.w2(32'h3911624f),
	.w3(32'h398000cf),
	.w4(32'hb87e7475),
	.w5(32'h38840ac8),
	.w6(32'h3a1090a5),
	.w7(32'hb86d1c48),
	.w8(32'h3a973539),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fa97d),
	.w1(32'h39a02647),
	.w2(32'h3a9be72d),
	.w3(32'h3ae447c6),
	.w4(32'h38ac6303),
	.w5(32'h385fc1cb),
	.w6(32'h3a729dca),
	.w7(32'h3a539d1a),
	.w8(32'hb9c17be1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caa0b3),
	.w1(32'hbb2629d0),
	.w2(32'hbbad0cc2),
	.w3(32'hbb5405a4),
	.w4(32'hbb5dfb1a),
	.w5(32'hbb14e090),
	.w6(32'hbb8fe817),
	.w7(32'hbb87d3cf),
	.w8(32'hbb2fada5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b43c24),
	.w1(32'h3ae8ba75),
	.w2(32'h3b946838),
	.w3(32'h385f9c41),
	.w4(32'hb88cc5eb),
	.w5(32'h3af3e54c),
	.w6(32'h3bb7a8f9),
	.w7(32'hbaf25fc4),
	.w8(32'hbb39d61c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca581f8),
	.w1(32'h3caf5372),
	.w2(32'h3c539f7f),
	.w3(32'h3c7ff650),
	.w4(32'h3c239fc5),
	.w5(32'hbb6dfa84),
	.w6(32'h3bed4c40),
	.w7(32'h3a307704),
	.w8(32'h3af4b36e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9ac9b),
	.w1(32'hb99d1316),
	.w2(32'h3bc63d73),
	.w3(32'hbb561a74),
	.w4(32'hbaaab77e),
	.w5(32'h3ab2febb),
	.w6(32'h3bb4fc26),
	.w7(32'hbc3124f8),
	.w8(32'hbc6d3acf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c0fa7),
	.w1(32'hbb741263),
	.w2(32'hbbba9402),
	.w3(32'hbb1949b4),
	.w4(32'hbb288e84),
	.w5(32'hbb547ae7),
	.w6(32'hbb4cdabc),
	.w7(32'hbba44cf2),
	.w8(32'hba9324df),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a33228),
	.w1(32'hbb1aee48),
	.w2(32'hbb0815ca),
	.w3(32'h3a5b232b),
	.w4(32'hbaa200b0),
	.w5(32'hba8744df),
	.w6(32'hbaaa69c1),
	.w7(32'hba071112),
	.w8(32'hba41ef14),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3edcf6),
	.w1(32'hb8f3ddd1),
	.w2(32'hb99aad3d),
	.w3(32'hba1c6b68),
	.w4(32'hb908c29a),
	.w5(32'hb9ccaf33),
	.w6(32'hb91ba586),
	.w7(32'hb9b30278),
	.w8(32'hbaa17df0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f6e54),
	.w1(32'hb983651a),
	.w2(32'hb8e39adf),
	.w3(32'hb93aeea4),
	.w4(32'h36b4cae1),
	.w5(32'hb93b50e2),
	.w6(32'hba92cab3),
	.w7(32'hba26f119),
	.w8(32'h3af8f94a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33a3aa),
	.w1(32'hbb9c7aff),
	.w2(32'hbb99e519),
	.w3(32'hb99a7942),
	.w4(32'hbb0f87be),
	.w5(32'hbb263b1e),
	.w6(32'hbaca4373),
	.w7(32'hbaddb4b3),
	.w8(32'h38fe7a25),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b663823),
	.w1(32'h3a7032e3),
	.w2(32'hba3401c7),
	.w3(32'h3a4c9ffb),
	.w4(32'hbb2c9b8c),
	.w5(32'hbaace111),
	.w6(32'hba0f0081),
	.w7(32'h3a4f91e2),
	.w8(32'hbb1698dd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb540aae),
	.w1(32'hbb137764),
	.w2(32'hbb126b7e),
	.w3(32'hbb3f628a),
	.w4(32'hbb1227a3),
	.w5(32'hbb26e545),
	.w6(32'hbb4047a9),
	.w7(32'hbb2e6ad4),
	.w8(32'hbad27d9c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93f4a5),
	.w1(32'h3b8a0b58),
	.w2(32'h3b097383),
	.w3(32'h3af2e5d1),
	.w4(32'h3b891d38),
	.w5(32'h3b914483),
	.w6(32'h3b5abc52),
	.w7(32'h3b8bcc5f),
	.w8(32'h3b35f60b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8448a6),
	.w1(32'h39eb4f94),
	.w2(32'h3a269b8b),
	.w3(32'h3a98f341),
	.w4(32'hba568eaf),
	.w5(32'hba947c80),
	.w6(32'h3b0b1278),
	.w7(32'hbaa930d2),
	.w8(32'hbb544063),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d8b5d),
	.w1(32'h3ba9b884),
	.w2(32'h3bbcd7f7),
	.w3(32'h3a0bb538),
	.w4(32'h39d1d8b2),
	.w5(32'h3b0d0bf9),
	.w6(32'hba543461),
	.w7(32'hb993c415),
	.w8(32'hb9bd9353),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb532234),
	.w1(32'hbacafcd3),
	.w2(32'h3aea18f6),
	.w3(32'hb616e360),
	.w4(32'h3a065e6e),
	.w5(32'h398e9a30),
	.w6(32'h3ad4f44b),
	.w7(32'hba88ee93),
	.w8(32'h3b13dbb7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a67e3),
	.w1(32'h3b632b06),
	.w2(32'h3bfa27ff),
	.w3(32'hbac6c99f),
	.w4(32'h3b1d2522),
	.w5(32'h3b93354a),
	.w6(32'h3b74cc21),
	.w7(32'hba9ede58),
	.w8(32'h3b1fda9a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91353e0),
	.w1(32'hb96ca1e5),
	.w2(32'hba222cfc),
	.w3(32'hba2a478d),
	.w4(32'hbaaa3855),
	.w5(32'hbab0bf8d),
	.w6(32'hb9976dc5),
	.w7(32'hba6795c0),
	.w8(32'h3bbabde6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5122e4),
	.w1(32'h3a8cb306),
	.w2(32'h3b4614e5),
	.w3(32'h3b919910),
	.w4(32'h3b094079),
	.w5(32'h3b856f5e),
	.w6(32'h3b643e2d),
	.w7(32'h3bafcb76),
	.w8(32'hba968fc5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab858ac),
	.w1(32'hba3b472a),
	.w2(32'hba4bcd4f),
	.w3(32'hbaa2984d),
	.w4(32'hba4eb162),
	.w5(32'hba6f259f),
	.w6(32'hba248c4c),
	.w7(32'hba367edd),
	.w8(32'hba05f3a5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e255a1),
	.w1(32'h39ed4339),
	.w2(32'h397de105),
	.w3(32'h39a738e1),
	.w4(32'h39ac5fba),
	.w5(32'hb9835c84),
	.w6(32'hba1322e6),
	.w7(32'hb95f46db),
	.w8(32'hb9b8fab5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fd442),
	.w1(32'hb9e8f6fb),
	.w2(32'h3832d692),
	.w3(32'hba541220),
	.w4(32'hba535999),
	.w5(32'hba21fd7d),
	.w6(32'hbac4b7e0),
	.w7(32'hbadd2cb7),
	.w8(32'h3ac785d8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c61d2),
	.w1(32'h3b15de62),
	.w2(32'h3b7466bd),
	.w3(32'h3b30e6e7),
	.w4(32'h3b2488bc),
	.w5(32'h3b859bd7),
	.w6(32'h3b5ce50f),
	.w7(32'h3b85b9fa),
	.w8(32'hbb25c9fb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae40e86),
	.w1(32'hbb44f361),
	.w2(32'hbb1a2ad2),
	.w3(32'hbaeaa104),
	.w4(32'hbaf16260),
	.w5(32'hbb22c87b),
	.w6(32'hbb8ddaaa),
	.w7(32'hb890d367),
	.w8(32'h3b3be1b6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc018d),
	.w1(32'hba9912d5),
	.w2(32'hbaceb567),
	.w3(32'h3a2f45d9),
	.w4(32'hbab88f64),
	.w5(32'hba85cd0c),
	.w6(32'hba521ad3),
	.w7(32'hba363d9b),
	.w8(32'h3a4283d3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cb67b),
	.w1(32'hbb881790),
	.w2(32'hbb1abc3e),
	.w3(32'hbb9639ba),
	.w4(32'hbb19b23f),
	.w5(32'h38502037),
	.w6(32'h3afbb1e8),
	.w7(32'hbbbbc9d8),
	.w8(32'hbc3ee12b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc51e),
	.w1(32'hbb4b6486),
	.w2(32'hba88c3b6),
	.w3(32'hba4e73f8),
	.w4(32'hbadec0a3),
	.w5(32'hb9c3e893),
	.w6(32'h38a666a1),
	.w7(32'hba9981ab),
	.w8(32'hba38e375),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28fb0d),
	.w1(32'hba5f21f1),
	.w2(32'hb92c6cae),
	.w3(32'hba58ce4a),
	.w4(32'hbac7b7a6),
	.w5(32'hbab1929c),
	.w6(32'hbaa2f188),
	.w7(32'hbaa7f887),
	.w8(32'hb9be596b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c3330),
	.w1(32'hba143be4),
	.w2(32'hbabecd95),
	.w3(32'h3998a0cf),
	.w4(32'hba4c3833),
	.w5(32'hbaf6ab3e),
	.w6(32'hba9b4793),
	.w7(32'hba1256fc),
	.w8(32'hba829947),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa6553),
	.w1(32'h39b85c27),
	.w2(32'h3af8b5ea),
	.w3(32'hba10d794),
	.w4(32'h3a8674fe),
	.w5(32'h3b51e643),
	.w6(32'hba89fe4d),
	.w7(32'hbb043fa0),
	.w8(32'hbb29d3dc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24a2b2),
	.w1(32'h3b30937e),
	.w2(32'h3bb62abe),
	.w3(32'h3a9973d7),
	.w4(32'h3a2d2af7),
	.w5(32'h3b066dc2),
	.w6(32'h3b0ecf0a),
	.w7(32'h3ac091db),
	.w8(32'h3b64f4de),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cb6ad),
	.w1(32'h3ae7cf2c),
	.w2(32'h3b7b8743),
	.w3(32'h3b297f49),
	.w4(32'hb9fb289e),
	.w5(32'h3adf2093),
	.w6(32'h3b204530),
	.w7(32'hbb10fde5),
	.w8(32'hb9a86378),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4aedd9),
	.w1(32'h3a0dd5b8),
	.w2(32'hb8e1be69),
	.w3(32'h3b1e848e),
	.w4(32'h39f76dbe),
	.w5(32'h3a7c4c2a),
	.w6(32'hb9f87609),
	.w7(32'hb9752c28),
	.w8(32'h3a6a038e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a880ff),
	.w1(32'hb9354fc5),
	.w2(32'hb8e9d978),
	.w3(32'hb966a1d1),
	.w4(32'hb938dbfa),
	.w5(32'hb94469e5),
	.w6(32'hb799f3f6),
	.w7(32'h3832def3),
	.w8(32'hb99a17ff),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39085a18),
	.w1(32'h3a2f6c7c),
	.w2(32'h3a378a7b),
	.w3(32'h3962b75b),
	.w4(32'h3ac38723),
	.w5(32'h3a3fcf1a),
	.w6(32'h39f6f00f),
	.w7(32'h3a212ce8),
	.w8(32'h3a9c88fb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d6672),
	.w1(32'h3aade66e),
	.w2(32'h3ace2dcd),
	.w3(32'h3aa1861f),
	.w4(32'h3acd4345),
	.w5(32'h3a93722d),
	.w6(32'h3a8732cf),
	.w7(32'h3a8affaf),
	.w8(32'h39df6efd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac3120),
	.w1(32'hb98c6514),
	.w2(32'h39840a9e),
	.w3(32'hba074101),
	.w4(32'hbaa3eae6),
	.w5(32'hba41b3fa),
	.w6(32'h3a703726),
	.w7(32'hbadec6ef),
	.w8(32'hba5a1c99),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba043ae4),
	.w1(32'hb8e75a5a),
	.w2(32'h3b558162),
	.w3(32'hbab21ac8),
	.w4(32'hbaa8a6cd),
	.w5(32'h3af8d2da),
	.w6(32'h3b368d9a),
	.w7(32'hba0b2b3e),
	.w8(32'hbb716cfc),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75f6d57),
	.w1(32'h397e4ae7),
	.w2(32'h391ad38a),
	.w3(32'hba078137),
	.w4(32'h3a38be84),
	.w5(32'h3a2a83c5),
	.w6(32'hb96160ad),
	.w7(32'hb9f71b56),
	.w8(32'hb9cfef4a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba624796),
	.w1(32'hba220637),
	.w2(32'hb9b3698d),
	.w3(32'hba35d13c),
	.w4(32'hba592080),
	.w5(32'hb9a0eb3e),
	.w6(32'hba090457),
	.w7(32'hb9a3d9e0),
	.w8(32'h3847a54f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b954d4c),
	.w1(32'h3b8f3f58),
	.w2(32'h3b830411),
	.w3(32'h3ad3d6c9),
	.w4(32'hbb24a6e3),
	.w5(32'hbae6028a),
	.w6(32'hbae14e9a),
	.w7(32'h3b333271),
	.w8(32'h3b9bbb3b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30b59d),
	.w1(32'hbb3a1162),
	.w2(32'hba93f24f),
	.w3(32'h3afd79eb),
	.w4(32'hbaf8c9b5),
	.w5(32'hbb15741c),
	.w6(32'h3b9f070d),
	.w7(32'hbaec4e43),
	.w8(32'hbb69dc68),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0662ea),
	.w1(32'hb9c2ae1f),
	.w2(32'h39d0d7d7),
	.w3(32'h39255559),
	.w4(32'hb96ea6ca),
	.w5(32'hb7a4eee5),
	.w6(32'h3908618a),
	.w7(32'h39b985cd),
	.w8(32'hba634a07),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac98b52),
	.w1(32'hbb0b90fc),
	.w2(32'hbb3dec24),
	.w3(32'hbabd92d7),
	.w4(32'hbac4501f),
	.w5(32'hbb2a260a),
	.w6(32'hbb070910),
	.w7(32'hbb031e26),
	.w8(32'hbb14b2d9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ce288),
	.w1(32'hbb3a69e4),
	.w2(32'hbad933fa),
	.w3(32'hbb72c63e),
	.w4(32'hbb1846aa),
	.w5(32'hbb0b9507),
	.w6(32'hbb14c1ab),
	.w7(32'hbb10f771),
	.w8(32'hbad98504),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab17658),
	.w1(32'h39faa6fc),
	.w2(32'h3a956afa),
	.w3(32'h3a8a75db),
	.w4(32'h3acaf6db),
	.w5(32'h3a896799),
	.w6(32'h3ac57c04),
	.w7(32'h3aa3c373),
	.w8(32'hb83d0f84),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e5c9a),
	.w1(32'h38fd17de),
	.w2(32'h3afd33a5),
	.w3(32'h3a92472e),
	.w4(32'hbaaa50d5),
	.w5(32'h38f7aaed),
	.w6(32'h3b38cbdc),
	.w7(32'h3a8e8795),
	.w8(32'h3a707853),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed9bf6),
	.w1(32'hbb01aeff),
	.w2(32'h3ac5eb9d),
	.w3(32'hbaec674d),
	.w4(32'h38da7830),
	.w5(32'h3afea0e1),
	.w6(32'h3b43c047),
	.w7(32'h3af7bdd5),
	.w8(32'h3a4c9737),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule