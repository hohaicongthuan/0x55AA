module layer_6_featuremap_22(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3c0f4),
	.w1(32'hbbad2ee7),
	.w2(32'hbb209f40),
	.w3(32'hbb956a4a),
	.w4(32'hbc0618e2),
	.w5(32'hbbdaa59c),
	.w6(32'hbb6615a1),
	.w7(32'hbc39c615),
	.w8(32'hbbcfc3df),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c7f48),
	.w1(32'hba112462),
	.w2(32'hb8b727b8),
	.w3(32'h36b865a7),
	.w4(32'hb96c8349),
	.w5(32'h3a46727e),
	.w6(32'hb9b79d74),
	.w7(32'h39b6be64),
	.w8(32'h390da9dc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badddd6),
	.w1(32'h3cb8d970),
	.w2(32'h3cb34180),
	.w3(32'h3c3f8743),
	.w4(32'hbb6c1906),
	.w5(32'h3be266c8),
	.w6(32'h3cc78062),
	.w7(32'h3c26e76c),
	.w8(32'h3886d498),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47d605),
	.w1(32'hbc2f884a),
	.w2(32'hbc74d3bb),
	.w3(32'hb70d2890),
	.w4(32'h3be0a984),
	.w5(32'hbb907ab2),
	.w6(32'hbb9eb086),
	.w7(32'hbb630810),
	.w8(32'hbc306b79),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c246c40),
	.w1(32'h3c0a0b0d),
	.w2(32'h3b627271),
	.w3(32'h3c90db0a),
	.w4(32'h3c3f050c),
	.w5(32'h3bca29b5),
	.w6(32'h3c462b72),
	.w7(32'h3bba4d3a),
	.w8(32'h3a67f5c2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1baec4),
	.w1(32'h3b8e48ed),
	.w2(32'h3ba49f8f),
	.w3(32'h393bd5b9),
	.w4(32'hb9d94098),
	.w5(32'h3b0d855f),
	.w6(32'h3b527b0f),
	.w7(32'h39f3fb3e),
	.w8(32'hb868aac9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e65a4),
	.w1(32'h3b9556ac),
	.w2(32'h3c0929d2),
	.w3(32'h3b077f47),
	.w4(32'h3b803b3a),
	.w5(32'h3bdbbcae),
	.w6(32'h3ad88dfb),
	.w7(32'h3b8fefc2),
	.w8(32'h3bf07999),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7eaeaa),
	.w1(32'h3b0b4a4e),
	.w2(32'h3a98cb94),
	.w3(32'h3b306113),
	.w4(32'h3b0e9eff),
	.w5(32'h3b3797ce),
	.w6(32'h3b354aa3),
	.w7(32'h3b1a8865),
	.w8(32'h3a347ffb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3635df),
	.w1(32'h3b579217),
	.w2(32'hb986863e),
	.w3(32'h3a0d8b27),
	.w4(32'hbb67166d),
	.w5(32'hba4ceeba),
	.w6(32'h3be05426),
	.w7(32'hba6a9221),
	.w8(32'hbb893193),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf28f31),
	.w1(32'h3bf912ec),
	.w2(32'h3c476593),
	.w3(32'h3b1a1654),
	.w4(32'h3be83bb1),
	.w5(32'h3c625909),
	.w6(32'h3b8e2fef),
	.w7(32'h3ba1ac16),
	.w8(32'h3c4b8641),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c812836),
	.w1(32'h3c00c31c),
	.w2(32'h3c0b6849),
	.w3(32'h3cbc167e),
	.w4(32'h3c266a13),
	.w5(32'h3c8995a8),
	.w6(32'h3cc016c3),
	.w7(32'h3c3fff68),
	.w8(32'h3c2b45fb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba9395),
	.w1(32'hbb022cf0),
	.w2(32'hbaf9aa24),
	.w3(32'hbaa11543),
	.w4(32'h3a0ccabc),
	.w5(32'h3a749c8a),
	.w6(32'h3a376e79),
	.w7(32'h392c3450),
	.w8(32'h38fe57ac),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae50858),
	.w1(32'h3a8e1d2f),
	.w2(32'hba54039c),
	.w3(32'h3b044d50),
	.w4(32'h3b26175a),
	.w5(32'h3b55d18b),
	.w6(32'h3b41a294),
	.w7(32'h3b22970b),
	.w8(32'hba7259c2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47bde3),
	.w1(32'h3ca463e7),
	.w2(32'h3cd8e21b),
	.w3(32'h3d2f17f6),
	.w4(32'h3d213c1f),
	.w5(32'h3d0df081),
	.w6(32'h3d1c77d2),
	.w7(32'h3d23dc80),
	.w8(32'h3d00095d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e2195),
	.w1(32'h3aaf3ba5),
	.w2(32'h3a72caab),
	.w3(32'hb907f211),
	.w4(32'h3ab9a3e5),
	.w5(32'h3a293b44),
	.w6(32'hbaae601c),
	.w7(32'h3ac5480a),
	.w8(32'h3bc6b4bf),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb397b),
	.w1(32'h3bae3289),
	.w2(32'h3b9b13a6),
	.w3(32'h3bd60deb),
	.w4(32'h3b741fa3),
	.w5(32'h3c0559a9),
	.w6(32'h3c2141c2),
	.w7(32'h3bd84eab),
	.w8(32'h3b34591f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d840a23),
	.w1(32'h3d3ff7df),
	.w2(32'h3d0b70fa),
	.w3(32'h3d4f1379),
	.w4(32'h3d158b98),
	.w5(32'h3d160a3e),
	.w6(32'h3cdacd18),
	.w7(32'h3bfbf71c),
	.w8(32'h3c9a36df),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905a86a),
	.w1(32'hba124ac3),
	.w2(32'hb7b8684f),
	.w3(32'hb93cc6b7),
	.w4(32'hb8c67956),
	.w5(32'h3ae95599),
	.w6(32'h3966d483),
	.w7(32'hb8d4deaa),
	.w8(32'hb946d26b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d86f58),
	.w1(32'h3c174fc7),
	.w2(32'h3c015535),
	.w3(32'h3bd95419),
	.w4(32'h3c3f12bc),
	.w5(32'h3c042893),
	.w6(32'h3bb9e67f),
	.w7(32'h3bfa4dae),
	.w8(32'h3bcba72e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9214dc),
	.w1(32'h3c8a254f),
	.w2(32'h3c92437f),
	.w3(32'h3c21812e),
	.w4(32'h3bf8d0fb),
	.w5(32'h3c1d0d5a),
	.w6(32'h3bf8f3f6),
	.w7(32'h3ba6e3f3),
	.w8(32'h3c2673dc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50dfe0),
	.w1(32'hbb916b6d),
	.w2(32'hbb759462),
	.w3(32'hb9f43c4b),
	.w4(32'h378c0671),
	.w5(32'hbace5c0b),
	.w6(32'hbad6f914),
	.w7(32'hbb414555),
	.w8(32'hbad62967),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4700fd),
	.w1(32'h3ce1538e),
	.w2(32'h3cc410c0),
	.w3(32'h3cc8ce35),
	.w4(32'h3cadc748),
	.w5(32'h3cb3172f),
	.w6(32'h3d15159e),
	.w7(32'h3cf93f9a),
	.w8(32'h3ca24969),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc564ccf),
	.w1(32'hbc972dad),
	.w2(32'hbc8f81c7),
	.w3(32'hbc6b12ab),
	.w4(32'hbcb6a164),
	.w5(32'hbca142a6),
	.w6(32'hbc59c2a1),
	.w7(32'hbc82ef22),
	.w8(32'hbc853d2f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68e8e3),
	.w1(32'h3c874f37),
	.w2(32'h3d0f0b96),
	.w3(32'h3d5831f1),
	.w4(32'h3ce07d39),
	.w5(32'h3c990116),
	.w6(32'h3d63bd3e),
	.w7(32'h3d26736c),
	.w8(32'h3c9ae913),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d5895),
	.w1(32'h3bc8a31f),
	.w2(32'hba27ce79),
	.w3(32'hbb92ac23),
	.w4(32'h3bdfc683),
	.w5(32'hb9ad2581),
	.w6(32'h3c190677),
	.w7(32'hbbeb6626),
	.w8(32'hbd2d200e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ff831),
	.w1(32'h3ccb81cb),
	.w2(32'h3ce15b7d),
	.w3(32'h3c8d02e4),
	.w4(32'h3d0f35ae),
	.w5(32'h3cb9d769),
	.w6(32'h3cd6c24b),
	.w7(32'h3d0792b7),
	.w8(32'h3ce562b9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90e3bf),
	.w1(32'h3c1f576b),
	.w2(32'h3ce67064),
	.w3(32'h3cd9f6f2),
	.w4(32'h3ca7677c),
	.w5(32'h3c9ab4dd),
	.w6(32'h3cde5cb3),
	.w7(32'h3cc2915c),
	.w8(32'h3c95489b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0b36),
	.w1(32'h3c4594a7),
	.w2(32'h3bf3ed35),
	.w3(32'hbb804cca),
	.w4(32'h3ac5326d),
	.w5(32'h3c1122cb),
	.w6(32'h3bd7fb28),
	.w7(32'h3bc846e2),
	.w8(32'h3bf2431f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab96f1f),
	.w1(32'h3a7ca8f3),
	.w2(32'hbaae1ff9),
	.w3(32'h3bace4cf),
	.w4(32'h3ac58ec6),
	.w5(32'h3ac5a120),
	.w6(32'h3bdfcc00),
	.w7(32'h3b9db777),
	.w8(32'h3b963a9b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8b60a7),
	.w1(32'hbc9c9bea),
	.w2(32'hbcc3f7a5),
	.w3(32'h3d53fb36),
	.w4(32'h3c77d7d7),
	.w5(32'h3a0dc3e8),
	.w6(32'h3d955278),
	.w7(32'h3d85406b),
	.w8(32'h3d7287cb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8494cf),
	.w1(32'hb9b95df2),
	.w2(32'hb9409068),
	.w3(32'h394c7bac),
	.w4(32'hb94955e3),
	.w5(32'hb95398e7),
	.w6(32'h3880da7b),
	.w7(32'hb88d5501),
	.w8(32'hb9225ef4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90d41a),
	.w1(32'h3c87379c),
	.w2(32'h3c906bde),
	.w3(32'h3c9902a0),
	.w4(32'h3c81016b),
	.w5(32'h3c8f00ac),
	.w6(32'h3c5ab9b6),
	.w7(32'h3c5d0303),
	.w8(32'h3c8deb0e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19510e),
	.w1(32'h3b09a6b9),
	.w2(32'h3afeb5d0),
	.w3(32'h3af46b09),
	.w4(32'h3af2c422),
	.w5(32'h3adcb7ed),
	.w6(32'h3b187a7c),
	.w7(32'h3b1659de),
	.w8(32'h3b0bd1a9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f5d1b4),
	.w1(32'hba2fd891),
	.w2(32'hb9939c74),
	.w3(32'hb930dd12),
	.w4(32'hba1249cb),
	.w5(32'hba005e05),
	.w6(32'h392e0ef2),
	.w7(32'hb98559b3),
	.w8(32'hba33a9c5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97fa29),
	.w1(32'h3a747cf0),
	.w2(32'h3a6cc59a),
	.w3(32'h3a7df08e),
	.w4(32'h3a1522bc),
	.w5(32'h39ef091a),
	.w6(32'h3a254ddc),
	.w7(32'h3aa45cf3),
	.w8(32'h3a036666),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc70066),
	.w1(32'h3cddc5d6),
	.w2(32'h3c921e20),
	.w3(32'h3ca7ea6d),
	.w4(32'h3d00bbab),
	.w5(32'h3cb94c69),
	.w6(32'h3d3916ab),
	.w7(32'h3d45b524),
	.w8(32'h3d197e32),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09a389),
	.w1(32'h3b2b14c7),
	.w2(32'h3b47eee6),
	.w3(32'h3aa79c2a),
	.w4(32'h3ad84f1e),
	.w5(32'h3b392462),
	.w6(32'h3a2259ce),
	.w7(32'h3abf2346),
	.w8(32'h3b30c950),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c1b37),
	.w1(32'h3c6e7e1c),
	.w2(32'h3c13d6a8),
	.w3(32'h3c5746e9),
	.w4(32'h3cccb8c4),
	.w5(32'h3c27c771),
	.w6(32'h3c89b9df),
	.w7(32'h3c88547a),
	.w8(32'h3c120584),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d7fb9),
	.w1(32'h3b1e8fd9),
	.w2(32'h3b245c1c),
	.w3(32'h3adf39ad),
	.w4(32'h3a9df7b3),
	.w5(32'h3b122dc7),
	.w6(32'h3aa59e69),
	.w7(32'h3a3cbc28),
	.w8(32'h3a8ee53c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1fda32),
	.w1(32'h3d6f3201),
	.w2(32'h3d0690d0),
	.w3(32'h3d5f67df),
	.w4(32'h3d757b0c),
	.w5(32'h3d4c2668),
	.w6(32'h3d57cda3),
	.w7(32'h3d3227f9),
	.w8(32'h3c9bdca5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c727fc5),
	.w1(32'h3cba91d6),
	.w2(32'h3d00276c),
	.w3(32'h3bcee735),
	.w4(32'h3c7e8dbb),
	.w5(32'h3d0725ad),
	.w6(32'h3b4089ac),
	.w7(32'h3b9c0c29),
	.w8(32'h3cc94344),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad8e20),
	.w1(32'h3bbd1108),
	.w2(32'h3c0f1a76),
	.w3(32'h3bf07799),
	.w4(32'h3c643d69),
	.w5(32'h3c956529),
	.w6(32'h3ca58ca8),
	.w7(32'h3cacc978),
	.w8(32'h3cb566cd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b768fe),
	.w1(32'h35dda159),
	.w2(32'hb8407677),
	.w3(32'h36f288c9),
	.w4(32'hb7f17458),
	.w5(32'hb708ae65),
	.w6(32'hb7ae9d22),
	.w7(32'hb85d74e3),
	.w8(32'hb81d121f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d892e8a),
	.w1(32'h3d5603e0),
	.w2(32'h3c84e388),
	.w3(32'h3d5cb3c3),
	.w4(32'h3dc01020),
	.w5(32'h3d25385a),
	.w6(32'h3da3b1d8),
	.w7(32'h3df7b5aa),
	.w8(32'h3d96ce84),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fe0f3),
	.w1(32'h3d119c03),
	.w2(32'h3cd85cfa),
	.w3(32'h3cdf0da6),
	.w4(32'h3c97d434),
	.w5(32'h3c82054c),
	.w6(32'h3ca27932),
	.w7(32'h3c24e422),
	.w8(32'h3b85673d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397edbef),
	.w1(32'h39858067),
	.w2(32'h39a2362e),
	.w3(32'h3948ceb9),
	.w4(32'h39abad7e),
	.w5(32'h3a00a4ab),
	.w6(32'h38f69c43),
	.w7(32'h398e0f05),
	.w8(32'h3a0969ca),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a291e8),
	.w1(32'h38d030d9),
	.w2(32'hb7da5ea0),
	.w3(32'h38e10c34),
	.w4(32'h38cc7d72),
	.w5(32'hb8dca231),
	.w6(32'h39006fa5),
	.w7(32'h3897dbf0),
	.w8(32'hb93dc4a7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ae44f),
	.w1(32'hbb83ef37),
	.w2(32'hbc97ae84),
	.w3(32'h3c575c3f),
	.w4(32'h3ca384be),
	.w5(32'hbc84fc1e),
	.w6(32'h3bef1be6),
	.w7(32'h3c5713aa),
	.w8(32'hbcac6c49),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76f9b9),
	.w1(32'h3c5a6eea),
	.w2(32'h3c6b425f),
	.w3(32'h3c8ec4df),
	.w4(32'h3c7b15ff),
	.w5(32'h3c91fe45),
	.w6(32'h3c650e52),
	.w7(32'h3c4b90b6),
	.w8(32'h3c6fab09),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6958be),
	.w1(32'hbb7676c9),
	.w2(32'h3b6deff3),
	.w3(32'hbbbbe361),
	.w4(32'h3c47ab7b),
	.w5(32'h3c55a350),
	.w6(32'hbc453efb),
	.w7(32'hbbc3b721),
	.w8(32'hbbb90f8b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392df9b1),
	.w1(32'hb8e0e87a),
	.w2(32'h3b9f3cc4),
	.w3(32'h3b2aa367),
	.w4(32'h3bbc444f),
	.w5(32'h3bc3567b),
	.w6(32'hbac82637),
	.w7(32'hbabedab0),
	.w8(32'hbb6fa050),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13c06e),
	.w1(32'h3c8b2ddf),
	.w2(32'h3cab53ae),
	.w3(32'hbbcc0ba7),
	.w4(32'h3c6ca1a9),
	.w5(32'h3cdf5b08),
	.w6(32'hbbf1467a),
	.w7(32'h3b97fb98),
	.w8(32'h3cbb0d9a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca02b44),
	.w1(32'h3d1194aa),
	.w2(32'h3c45f304),
	.w3(32'h3ce0baee),
	.w4(32'h3c75f7a0),
	.w5(32'hbb0a8bfb),
	.w6(32'h3cff73a6),
	.w7(32'h3c6f5280),
	.w8(32'hbc9d44c1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be585ed),
	.w1(32'h3c0e043b),
	.w2(32'h3c3211da),
	.w3(32'h3c28c334),
	.w4(32'h3c392fad),
	.w5(32'h3c85a9eb),
	.w6(32'h38606546),
	.w7(32'hbc49b722),
	.w8(32'hbb4209de),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2100bb),
	.w1(32'h3bfbe969),
	.w2(32'h3bf4cef3),
	.w3(32'h3aa6814c),
	.w4(32'h3be9c2d6),
	.w5(32'h3c00e01c),
	.w6(32'h3aa82175),
	.w7(32'h3b96256c),
	.w8(32'h3be1f2f9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd856d),
	.w1(32'hbcb4f431),
	.w2(32'hbd05a601),
	.w3(32'hbcb03056),
	.w4(32'hbbf9445a),
	.w5(32'hbcbbb6c7),
	.w6(32'hbc3eb537),
	.w7(32'hbbe2058f),
	.w8(32'hbc8e16e9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b916c),
	.w1(32'h3c9c953a),
	.w2(32'h3cda082b),
	.w3(32'h3c688f53),
	.w4(32'h3c6b09dd),
	.w5(32'h3ccc501b),
	.w6(32'h3c5e97d4),
	.w7(32'h3c59fac5),
	.w8(32'h3cbbc51c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4a8446),
	.w1(32'h3d4f1ec1),
	.w2(32'h3d38b0c0),
	.w3(32'h3d4d13a8),
	.w4(32'h3d5f7957),
	.w5(32'h3d3c1f97),
	.w6(32'h3d39f9de),
	.w7(32'h3d4b0af0),
	.w8(32'h3d3c5263),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c3df2),
	.w1(32'h3ce1194e),
	.w2(32'h3cc9c8ae),
	.w3(32'h3c9bf030),
	.w4(32'h3cf0450c),
	.w5(32'h3cb51970),
	.w6(32'h3cb6a30b),
	.w7(32'h3ce54dde),
	.w8(32'h3cdcfb4a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce6ad59),
	.w1(32'h3d1a29f5),
	.w2(32'h3cfc3e4a),
	.w3(32'h3cbb1915),
	.w4(32'h3cd46ab7),
	.w5(32'h3d0b7a7e),
	.w6(32'h3c3c708a),
	.w7(32'hbb47be72),
	.w8(32'h3bb1833e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc81360),
	.w1(32'h39839550),
	.w2(32'hbcedf81e),
	.w3(32'hbb86aecd),
	.w4(32'hbaab594b),
	.w5(32'hbca66ab7),
	.w6(32'hbb0f45c5),
	.w7(32'hbc6f96cb),
	.w8(32'hbc394887),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c583f9d),
	.w1(32'h3cf2cfb7),
	.w2(32'h3ca20019),
	.w3(32'h3c8d05f7),
	.w4(32'h3d07b1b0),
	.w5(32'h3cb33f77),
	.w6(32'h3cc0cadc),
	.w7(32'h3d021d84),
	.w8(32'h3c934373),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdc9e911),
	.w1(32'hbdcd776e),
	.w2(32'h3c919e52),
	.w3(32'hbd7fb958),
	.w4(32'h3ca8ec66),
	.w5(32'h3d3600da),
	.w6(32'h3c0d54c8),
	.w7(32'h3d45873c),
	.w8(32'h3cac2927),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6d68b1),
	.w1(32'h3caab2ca),
	.w2(32'h3cbcfa67),
	.w3(32'hbd13d858),
	.w4(32'h3b90a470),
	.w5(32'hbc1ac3bc),
	.w6(32'hbd3b443f),
	.w7(32'h3d937207),
	.w8(32'hbba47b91),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule