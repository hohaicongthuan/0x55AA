module layer_10_featuremap_320(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9b24d),
	.w1(32'hb9cc8e2c),
	.w2(32'hb94c1197),
	.w3(32'hb9a49b33),
	.w4(32'hb95e8347),
	.w5(32'h38fd1600),
	.w6(32'hba3e5056),
	.w7(32'hb9fe34eb),
	.w8(32'h399af0db),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e6411),
	.w1(32'h3b0a29cd),
	.w2(32'h3b67a7bd),
	.w3(32'h3a4b3849),
	.w4(32'h3b08b05d),
	.w5(32'h3a7ae7bc),
	.w6(32'hb89a4bed),
	.w7(32'hba255260),
	.w8(32'hba180d69),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bb94b),
	.w1(32'h3a245d80),
	.w2(32'h3959d320),
	.w3(32'h39b3bfb2),
	.w4(32'h392b60a7),
	.w5(32'hb6967b6a),
	.w6(32'h393e6a3e),
	.w7(32'h39a7821e),
	.w8(32'hb889b128),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3c29a),
	.w1(32'h3a4cf978),
	.w2(32'hba0c656b),
	.w3(32'h3994c68d),
	.w4(32'h39cd0e24),
	.w5(32'hba465f66),
	.w6(32'h39a9d8f3),
	.w7(32'h3a00816d),
	.w8(32'hb9a3bb86),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39122e2e),
	.w1(32'hb937f3df),
	.w2(32'h396288ba),
	.w3(32'hb9f351f9),
	.w4(32'h39468c67),
	.w5(32'h39314d93),
	.w6(32'h391aa3c2),
	.w7(32'h3a1d6f60),
	.w8(32'h398433f3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e06e27),
	.w1(32'h399cd1a9),
	.w2(32'h39a371fe),
	.w3(32'hb8d7f560),
	.w4(32'hb8faab21),
	.w5(32'h3a8dd02d),
	.w6(32'h383f8e69),
	.w7(32'hb8b00453),
	.w8(32'h3a881077),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3587e),
	.w1(32'h3ae0246e),
	.w2(32'hbb01d316),
	.w3(32'h3b9e4b60),
	.w4(32'h3b2b0fdd),
	.w5(32'hbb1f8db3),
	.w6(32'h3b95d4a2),
	.w7(32'h39a9d45a),
	.w8(32'hbb9296c4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb823dfd),
	.w1(32'hbab0dddd),
	.w2(32'hbbc91279),
	.w3(32'hbb8eb162),
	.w4(32'hbb80f0b2),
	.w5(32'hbb60d57b),
	.w6(32'hbacf1f92),
	.w7(32'hbaa03bb7),
	.w8(32'hbb34a085),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d8229),
	.w1(32'hba59f1c9),
	.w2(32'hbab46821),
	.w3(32'hb9a31ade),
	.w4(32'hba3a5b0e),
	.w5(32'hba511444),
	.w6(32'h3a39fc86),
	.w7(32'hb9e3855d),
	.w8(32'hba9234d4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa72b9),
	.w1(32'hbb0d6761),
	.w2(32'hbb3b8db1),
	.w3(32'h39d13692),
	.w4(32'hbb0b2a95),
	.w5(32'hbb6d5153),
	.w6(32'h3b0abde7),
	.w7(32'hba0481ea),
	.w8(32'hbb952b30),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a288cce),
	.w1(32'h3a0fa715),
	.w2(32'hb9714e89),
	.w3(32'hb8d77043),
	.w4(32'hb9d0998d),
	.w5(32'hba3dd40f),
	.w6(32'h3a027a90),
	.w7(32'hb9d1770c),
	.w8(32'hba7c0927),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2a45f),
	.w1(32'h3b927893),
	.w2(32'hbb5f535e),
	.w3(32'h3b93289d),
	.w4(32'h3b487e87),
	.w5(32'hbb0da7ef),
	.w6(32'h3b8d7a0e),
	.w7(32'h3b5e2bf0),
	.w8(32'hb9745202),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b157e54),
	.w1(32'hba2b84e1),
	.w2(32'hbb3899e8),
	.w3(32'h3a88d1db),
	.w4(32'hbaccae7f),
	.w5(32'hbb87425d),
	.w6(32'h3b856d0d),
	.w7(32'h3a137b17),
	.w8(32'hbb60ec61),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a201111),
	.w1(32'h3a4fe80b),
	.w2(32'h39f61898),
	.w3(32'h3947e9a0),
	.w4(32'h39dd33bd),
	.w5(32'h3a88d478),
	.w6(32'hba523257),
	.w7(32'hb9db3a01),
	.w8(32'hb8c344c7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92722f),
	.w1(32'h3a06a6a1),
	.w2(32'h3a61e283),
	.w3(32'h3b048de6),
	.w4(32'h3b3072fe),
	.w5(32'h3ac63277),
	.w6(32'h3b149565),
	.w7(32'h3a8c70c6),
	.w8(32'h391b4a10),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad10c86),
	.w1(32'hbafec27c),
	.w2(32'h39361eab),
	.w3(32'h39b9497c),
	.w4(32'hba8295f4),
	.w5(32'hbb35fd52),
	.w6(32'hbb25b046),
	.w7(32'hbb847e25),
	.w8(32'hbb85fb03),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fa4ca),
	.w1(32'h3a89389d),
	.w2(32'h3a45ab9d),
	.w3(32'hb996248a),
	.w4(32'hba10bc4b),
	.w5(32'hba4592bf),
	.w6(32'hba1d46d7),
	.w7(32'hbad08728),
	.w8(32'hba4d389c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d853d0),
	.w1(32'hbbfd81e9),
	.w2(32'hbc2d5ffc),
	.w3(32'hbb935203),
	.w4(32'hbc12f1e3),
	.w5(32'hbbdb0850),
	.w6(32'hbb05af63),
	.w7(32'hbc2fdb52),
	.w8(32'hbbc0509f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bdce4),
	.w1(32'hbafb3fbb),
	.w2(32'hbb81efa1),
	.w3(32'hba8bd950),
	.w4(32'hbb80b453),
	.w5(32'hbb336ee1),
	.w6(32'h3a9a3527),
	.w7(32'hbb5e504e),
	.w8(32'hbb1878b2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9811819),
	.w1(32'h39986a45),
	.w2(32'h39e20152),
	.w3(32'h3a0849af),
	.w4(32'h3957cd51),
	.w5(32'h39b9c187),
	.w6(32'h391fb097),
	.w7(32'h399debfe),
	.w8(32'hb8e31aff),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398557bb),
	.w1(32'h3a03cb74),
	.w2(32'h39b721e8),
	.w3(32'h39bed52f),
	.w4(32'h3899f846),
	.w5(32'h3a9027f9),
	.w6(32'hb8b9547d),
	.w7(32'hb8769d81),
	.w8(32'h3a854787),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00cf1e),
	.w1(32'h3b196e96),
	.w2(32'h3b0f3c70),
	.w3(32'h3b2f73d2),
	.w4(32'h3b5fa49e),
	.w5(32'h3adb53a2),
	.w6(32'h3a8e27e6),
	.w7(32'h3adf4884),
	.w8(32'h3a75cca1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d2a7b),
	.w1(32'hbbb92227),
	.w2(32'hbc602ca2),
	.w3(32'hbb05c392),
	.w4(32'hbb3e7623),
	.w5(32'hbc010b1c),
	.w6(32'hbbe12afb),
	.w7(32'hbbb5c6d9),
	.w8(32'hbbfc4238),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acebf04),
	.w1(32'hbac23d9c),
	.w2(32'hb9177159),
	.w3(32'h3b0d8a5b),
	.w4(32'h3a2ba522),
	.w5(32'h39aac93a),
	.w6(32'h3b4c23cd),
	.w7(32'h3a519896),
	.w8(32'hba94f4fa),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02df37),
	.w1(32'h3a395c53),
	.w2(32'h3b5efd18),
	.w3(32'h3a7c1a27),
	.w4(32'h3bbb69f1),
	.w5(32'h3ba8532c),
	.w6(32'hba758316),
	.w7(32'h370f3dba),
	.w8(32'hbabf4433),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4dc26b),
	.w1(32'h39f46cfc),
	.w2(32'h38737c9b),
	.w3(32'hb8679970),
	.w4(32'h394f71e7),
	.w5(32'h39bd4439),
	.w6(32'hb9779c73),
	.w7(32'h395aeb21),
	.w8(32'h38ca8a5b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b1322),
	.w1(32'hb9c758cc),
	.w2(32'h39cb4fbb),
	.w3(32'hb9129433),
	.w4(32'h39aa76e0),
	.w5(32'hba4e7752),
	.w6(32'hba0c6379),
	.w7(32'h381b88df),
	.w8(32'hba85f106),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a6669),
	.w1(32'hbb19a86f),
	.w2(32'h39f7775f),
	.w3(32'h3b3382d7),
	.w4(32'h3ac12c57),
	.w5(32'h3908508a),
	.w6(32'h3a5598fc),
	.w7(32'hbb151c7a),
	.w8(32'hbb1c092e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d8623),
	.w1(32'hb90e2faa),
	.w2(32'h3a94247d),
	.w3(32'h3a3547f1),
	.w4(32'h3aab3098),
	.w5(32'h3ad42764),
	.w6(32'hb9c5671b),
	.w7(32'h3a714ac0),
	.w8(32'h3a81c8de),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2011c5),
	.w1(32'h3a1b98b9),
	.w2(32'h3b45d8c7),
	.w3(32'h3b305ec8),
	.w4(32'h3b70a260),
	.w5(32'h3b3d8d5e),
	.w6(32'h3b0bf9e5),
	.w7(32'h3aa69c10),
	.w8(32'hba5c7160),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64eac9),
	.w1(32'hba0bff2f),
	.w2(32'hb96dc1f4),
	.w3(32'h39567834),
	.w4(32'h3911d15d),
	.w5(32'h3a01dc41),
	.w6(32'h3a624e52),
	.w7(32'h3975eb19),
	.w8(32'h3a806adc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a170c80),
	.w1(32'h3a46d6cd),
	.w2(32'h39b5e5e4),
	.w3(32'h3a3ca7c9),
	.w4(32'h39d336a0),
	.w5(32'h39e2c52c),
	.w6(32'h3a696ff8),
	.w7(32'h3a029fa5),
	.w8(32'h3a819679),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0596c8),
	.w1(32'hba5a307d),
	.w2(32'hbb267518),
	.w3(32'h3b082be0),
	.w4(32'h3907cb68),
	.w5(32'hbaed4f24),
	.w6(32'h3b2261e3),
	.w7(32'h39d1e28f),
	.w8(32'hbaf1a0cb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d9b6a),
	.w1(32'hb96490e0),
	.w2(32'h3a1cc662),
	.w3(32'hba4db37f),
	.w4(32'h3a24169d),
	.w5(32'h3a7af289),
	.w6(32'hba584ab2),
	.w7(32'hb7f4a076),
	.w8(32'hb9660f6c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a719eac),
	.w1(32'hb7419be1),
	.w2(32'h3a15d99c),
	.w3(32'h39eab737),
	.w4(32'h399083e1),
	.w5(32'hb967b95d),
	.w6(32'h3a404c01),
	.w7(32'hb95c3528),
	.w8(32'hb9cb3c97),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3766da),
	.w1(32'h3b05214d),
	.w2(32'hb9e623e7),
	.w3(32'h3a84bdd0),
	.w4(32'h3a673e17),
	.w5(32'hbaae3619),
	.w6(32'h3b289d8a),
	.w7(32'h3b0d22b4),
	.w8(32'hba5e5967),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac18a0b),
	.w1(32'h3c54ccc0),
	.w2(32'hbc4debc1),
	.w3(32'h3b1de13e),
	.w4(32'h3bd0e60a),
	.w5(32'hbbb56ec3),
	.w6(32'hba8f1d13),
	.w7(32'h3bd87367),
	.w8(32'hbbaf37aa),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc05878),
	.w1(32'h3bb4a3ff),
	.w2(32'h3c1a2f20),
	.w3(32'h3a1c39ff),
	.w4(32'h3c2e9b40),
	.w5(32'h3c1bc6fd),
	.w6(32'hbb791e9a),
	.w7(32'h39eaad08),
	.w8(32'h3a2859d6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d15a),
	.w1(32'h3ab7800e),
	.w2(32'h3b991620),
	.w3(32'h3b6a0c16),
	.w4(32'h3ba718e2),
	.w5(32'h3bc02ddb),
	.w6(32'h3b86ef2b),
	.w7(32'hb8da948d),
	.w8(32'h3aa5d424),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38adb76e),
	.w1(32'h3a91de2d),
	.w2(32'h3a9921ca),
	.w3(32'h3a9ec9d4),
	.w4(32'h3ad77ebf),
	.w5(32'h3a91b958),
	.w6(32'h3a3cd141),
	.w7(32'h3a44a9c5),
	.w8(32'hb6a5bbf5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385f726b),
	.w1(32'h38d25548),
	.w2(32'h399e1b57),
	.w3(32'h384e4ebc),
	.w4(32'h38da5724),
	.w5(32'hb9a2670f),
	.w6(32'hb9bf1d69),
	.w7(32'h39903c7a),
	.w8(32'hba0d74da),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb0319),
	.w1(32'hba49acde),
	.w2(32'hb9c5a8f9),
	.w3(32'hba66efde),
	.w4(32'hb9d6e5a6),
	.w5(32'h392659ad),
	.w6(32'hba88fa49),
	.w7(32'hba479b1e),
	.w8(32'hb9335149),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c3e03),
	.w1(32'hba486bb1),
	.w2(32'h398d06c0),
	.w3(32'hba484793),
	.w4(32'h3910b11c),
	.w5(32'h3a06e95d),
	.w6(32'hbaca6547),
	.w7(32'hb9b90a2a),
	.w8(32'hb823fd2c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99afe0f),
	.w1(32'hbb904477),
	.w2(32'hbad4c2bf),
	.w3(32'hbb587cc7),
	.w4(32'hbb72a2f9),
	.w5(32'hbba1481e),
	.w6(32'h3937eede),
	.w7(32'hbb260a9f),
	.w8(32'hbb51959c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cff8e),
	.w1(32'hbb6cdc33),
	.w2(32'hbb2fda65),
	.w3(32'hba438355),
	.w4(32'hb96a735a),
	.w5(32'hb92847f3),
	.w6(32'h390a491e),
	.w7(32'hba4787ac),
	.w8(32'hbade617d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2553b),
	.w1(32'hbb448d51),
	.w2(32'hb9d6fe8a),
	.w3(32'h3adde310),
	.w4(32'h3a808733),
	.w5(32'hbb0a1d09),
	.w6(32'h3b29e0a9),
	.w7(32'h3a3b8837),
	.w8(32'hbb87daf9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb109e6d),
	.w1(32'hbb612730),
	.w2(32'hbadf5081),
	.w3(32'hba9e8ed2),
	.w4(32'hbad53d53),
	.w5(32'h3ab32d7e),
	.w6(32'hbb8ec428),
	.w7(32'hbb55faca),
	.w8(32'hba821b41),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd5f77),
	.w1(32'hbad90a1d),
	.w2(32'hbc25c6ae),
	.w3(32'hb99ef60d),
	.w4(32'hbbaedf9c),
	.w5(32'hbc02330c),
	.w6(32'h38142ecc),
	.w7(32'hbba573b8),
	.w8(32'hbba7d8ed),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0c626),
	.w1(32'hba0ea27f),
	.w2(32'hb9c2623a),
	.w3(32'hba3890b2),
	.w4(32'hb9cb5758),
	.w5(32'h3aab11d7),
	.w6(32'hba1e5a61),
	.w7(32'h37eb4ab4),
	.w8(32'h3a87add1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93da0c0),
	.w1(32'hb94b505e),
	.w2(32'h39a05758),
	.w3(32'h36e9b74d),
	.w4(32'h393bd39e),
	.w5(32'hb9d1f14d),
	.w6(32'h39bbc45d),
	.w7(32'h3a09ea26),
	.w8(32'hb9982e17),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abe428),
	.w1(32'h39536f63),
	.w2(32'h3a37e771),
	.w3(32'h3972eaf2),
	.w4(32'h3aa9fd40),
	.w5(32'hb94cb5da),
	.w6(32'h3932d220),
	.w7(32'h3a9eb879),
	.w8(32'h388f81a4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a19f9),
	.w1(32'hbb091559),
	.w2(32'hba94e358),
	.w3(32'hbaa3397a),
	.w4(32'hba5473c7),
	.w5(32'hbac2384f),
	.w6(32'hb978fad2),
	.w7(32'hba57716b),
	.w8(32'hbb3475bd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6c9c7),
	.w1(32'hb9dae368),
	.w2(32'hbaa52d6c),
	.w3(32'hba941b5a),
	.w4(32'hba418686),
	.w5(32'hbaaa840c),
	.w6(32'hb93a67a5),
	.w7(32'h3a270bed),
	.w8(32'hbaa266c3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac30470),
	.w1(32'hbbbe9350),
	.w2(32'hbbe3071d),
	.w3(32'hbb8f6d03),
	.w4(32'hbbc2a584),
	.w5(32'hbb5a812b),
	.w6(32'hba99e03c),
	.w7(32'hbb5afb57),
	.w8(32'hbb5f8ac0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37660a),
	.w1(32'hba2d1fa5),
	.w2(32'hba8dc39b),
	.w3(32'hba17628b),
	.w4(32'hba4db4c5),
	.w5(32'hba60286c),
	.w6(32'h3865b22e),
	.w7(32'hb7dabae1),
	.w8(32'h391a2386),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f40ba),
	.w1(32'h39a0688e),
	.w2(32'h3a26e943),
	.w3(32'hb85270c5),
	.w4(32'h38b2c1e3),
	.w5(32'h392f6629),
	.w6(32'hb9415fc2),
	.w7(32'hb88c3b47),
	.w8(32'h38ef232f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7043ea6),
	.w1(32'h3908ec9a),
	.w2(32'h391b56f9),
	.w3(32'h390c0b62),
	.w4(32'hb8e37211),
	.w5(32'h37db7265),
	.w6(32'hb906ffae),
	.w7(32'hb924a500),
	.w8(32'hb9e9d7f8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc1a7b),
	.w1(32'hb98bbaa5),
	.w2(32'h39a89ea8),
	.w3(32'h3a429fdf),
	.w4(32'hb826d851),
	.w5(32'h3a701778),
	.w6(32'h39936368),
	.w7(32'h393dddf4),
	.w8(32'h39eba06d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa43830),
	.w1(32'h3a9cf330),
	.w2(32'h3a841a76),
	.w3(32'h3aabf0be),
	.w4(32'h3ad5a77c),
	.w5(32'h3aab41f8),
	.w6(32'h39e2c6b0),
	.w7(32'h3a736343),
	.w8(32'h3aeeb4e0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb3e75),
	.w1(32'h3aa4b872),
	.w2(32'h3acce880),
	.w3(32'h3a717290),
	.w4(32'h3a0edd62),
	.w5(32'h39932255),
	.w6(32'h3b5d2dde),
	.w7(32'h3ab6cf7d),
	.w8(32'h39ced5d9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78ef1f),
	.w1(32'hbac69daf),
	.w2(32'hbb2324ae),
	.w3(32'hb954eb82),
	.w4(32'hbad77eae),
	.w5(32'hbb01f664),
	.w6(32'h3a4cf6f9),
	.w7(32'hbacfdd33),
	.w8(32'hbab733fa),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd7106),
	.w1(32'hbb2e5dae),
	.w2(32'hb9bfbe19),
	.w3(32'hbb863023),
	.w4(32'hbb2845d2),
	.w5(32'hbadbc020),
	.w6(32'hbb35f168),
	.w7(32'hbb429919),
	.w8(32'hb9bf5742),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b1e61),
	.w1(32'h37eec3ef),
	.w2(32'h39ef1f4b),
	.w3(32'h3730fe78),
	.w4(32'h3a1b1eaf),
	.w5(32'h38835796),
	.w6(32'h39644893),
	.w7(32'h3a2e7382),
	.w8(32'h3854457b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38410938),
	.w1(32'h398354e2),
	.w2(32'h3a61e65f),
	.w3(32'h399fc71e),
	.w4(32'h39e8de72),
	.w5(32'h39a91261),
	.w6(32'hb93194a6),
	.w7(32'h39ff86f8),
	.w8(32'h392513df),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a929f2),
	.w1(32'h396d668c),
	.w2(32'h3a14437c),
	.w3(32'h3a0277ba),
	.w4(32'h39f2469d),
	.w5(32'hb9f01101),
	.w6(32'h38fbf95b),
	.w7(32'h397ddbe3),
	.w8(32'h38a1eb13),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fc0a0),
	.w1(32'hb9801868),
	.w2(32'h388905d5),
	.w3(32'hba6627e5),
	.w4(32'hba3a4416),
	.w5(32'h399210fb),
	.w6(32'h39e9c00d),
	.w7(32'h39894d18),
	.w8(32'h38a3aaf3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baacefd),
	.w1(32'hb8dfb420),
	.w2(32'hba4cc0cf),
	.w3(32'h3b362b61),
	.w4(32'hba4b8d2f),
	.w5(32'h3a1014af),
	.w6(32'h398a40df),
	.w7(32'hbb57941f),
	.w8(32'hbb4da441),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b150974),
	.w1(32'hbb157465),
	.w2(32'hbb3c52e9),
	.w3(32'h3b59a6a8),
	.w4(32'h3ac749ab),
	.w5(32'hbb552ef5),
	.w6(32'h3ad463c4),
	.w7(32'h3aade9d0),
	.w8(32'hbb22e251),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9dfcf),
	.w1(32'hbba0b35d),
	.w2(32'hbbaec110),
	.w3(32'hbabf6cd6),
	.w4(32'hbb13f39a),
	.w5(32'hbb4bd5c6),
	.w6(32'hbb224971),
	.w7(32'hbb7984e8),
	.w8(32'hbb8717c7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb553b7a),
	.w1(32'h3aade440),
	.w2(32'h3b9a4357),
	.w3(32'h3afdaf94),
	.w4(32'h3bdbb679),
	.w5(32'h3b9e264f),
	.w6(32'h3a1a3704),
	.w7(32'hb97699d1),
	.w8(32'hbb4a25eb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942efba),
	.w1(32'hba08ef39),
	.w2(32'hb9b1aa33),
	.w3(32'h381deaf6),
	.w4(32'hb8f889a5),
	.w5(32'h37dd429f),
	.w6(32'hb9afd8d8),
	.w7(32'hb98428a4),
	.w8(32'hb7ead3d6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7ac3d),
	.w1(32'h3a139ec0),
	.w2(32'h3a1fffb1),
	.w3(32'h397d7553),
	.w4(32'h3a0dcd09),
	.w5(32'h3900cc04),
	.w6(32'h3a097ab3),
	.w7(32'h398b1854),
	.w8(32'h39f91a28),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a629783),
	.w1(32'h3a9609ed),
	.w2(32'h3a89f714),
	.w3(32'h38b7aaa2),
	.w4(32'h39317ee9),
	.w5(32'h39a0012e),
	.w6(32'h3a969ef3),
	.w7(32'h3a1cc982),
	.w8(32'h385c2236),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ea951),
	.w1(32'hba1ff596),
	.w2(32'hba870661),
	.w3(32'h3a1ab06f),
	.w4(32'hba145605),
	.w5(32'hbabcd33e),
	.w6(32'h3899e7e7),
	.w7(32'hba83bc39),
	.w8(32'hbad2f397),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395215fc),
	.w1(32'h3a04f000),
	.w2(32'h3a008028),
	.w3(32'h376b5cf9),
	.w4(32'h38cdcb0c),
	.w5(32'hb993d99b),
	.w6(32'hb7786c41),
	.w7(32'h38e1006d),
	.w8(32'h37f5b5f3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28c3b9),
	.w1(32'hbb2a67c5),
	.w2(32'hbbabe7f7),
	.w3(32'hb9d0aa60),
	.w4(32'hbb8b25eb),
	.w5(32'hbb584bce),
	.w6(32'hba7e0972),
	.w7(32'hbb0d180f),
	.w8(32'hbb7dd527),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac429e0),
	.w1(32'hba984599),
	.w2(32'hbbe39d43),
	.w3(32'h3a11f82f),
	.w4(32'hbb8f7c13),
	.w5(32'hbbd3ab80),
	.w6(32'hbab80fb6),
	.w7(32'hbb8b3987),
	.w8(32'hbbd01e04),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff7197),
	.w1(32'h3a7e5955),
	.w2(32'h3a91fdc9),
	.w3(32'h384ef528),
	.w4(32'h3add74d7),
	.w5(32'hb9caf048),
	.w6(32'h3a5ee2bf),
	.w7(32'h3a4acfd7),
	.w8(32'hbad99421),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e47b8),
	.w1(32'hbade3434),
	.w2(32'hbb39ab4d),
	.w3(32'hb913a32a),
	.w4(32'hbaafbaec),
	.w5(32'hba9dead4),
	.w6(32'h3acb06f1),
	.w7(32'hbab3b6aa),
	.w8(32'hbb0b81fa),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c0211),
	.w1(32'h39a94979),
	.w2(32'hba1ac616),
	.w3(32'h3aad26d9),
	.w4(32'h3a005905),
	.w5(32'hba94847f),
	.w6(32'h3b223277),
	.w7(32'hbaaca902),
	.w8(32'hbb596a20),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41afaf),
	.w1(32'hbb8ec551),
	.w2(32'hbb43c986),
	.w3(32'hbac7fb37),
	.w4(32'hba278804),
	.w5(32'hbae8132e),
	.w6(32'hbb0dd6da),
	.w7(32'hbaea1575),
	.w8(32'hbaf75162),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada6d4e),
	.w1(32'hbab81f11),
	.w2(32'hbb99320f),
	.w3(32'hb8194f96),
	.w4(32'hbb1908e1),
	.w5(32'hbb35d761),
	.w6(32'hb8fce424),
	.w7(32'hbb25ada6),
	.w8(32'hbb091541),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01f0f7),
	.w1(32'h3a1825db),
	.w2(32'h3a47823a),
	.w3(32'h3a154416),
	.w4(32'h3a3d905d),
	.w5(32'hba20d795),
	.w6(32'h3a4309f9),
	.w7(32'h3a538331),
	.w8(32'hb80316a4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395049e1),
	.w1(32'h39ae981e),
	.w2(32'h3782d28c),
	.w3(32'hba64b615),
	.w4(32'hba18ce6a),
	.w5(32'h395aa940),
	.w6(32'h395b7d44),
	.w7(32'hb927fbed),
	.w8(32'h39f5b545),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4135f9),
	.w1(32'h3a54407c),
	.w2(32'h3ab21e8c),
	.w3(32'h3a308b93),
	.w4(32'h3a5fa1c7),
	.w5(32'h3a20f407),
	.w6(32'h3a7037cc),
	.w7(32'h3a977879),
	.w8(32'h3a620af8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3892dee3),
	.w1(32'hb98aad0f),
	.w2(32'h398ec5a4),
	.w3(32'hb9455fc1),
	.w4(32'hb9d724bd),
	.w5(32'h39e7b2bd),
	.w6(32'h3a7dac8f),
	.w7(32'h3732bcb3),
	.w8(32'hb9501ffb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d30dd),
	.w1(32'h3a7dae37),
	.w2(32'h3ac2f4a2),
	.w3(32'h382799bd),
	.w4(32'h3b223082),
	.w5(32'h3ae1a9f1),
	.w6(32'hbb2d2ae5),
	.w7(32'hbaabe5b1),
	.w8(32'hbafcd56a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcc54b),
	.w1(32'hb8b196b8),
	.w2(32'h3932bf8c),
	.w3(32'hb9df8895),
	.w4(32'h38d9c226),
	.w5(32'h3a789c4e),
	.w6(32'h39813365),
	.w7(32'h3a304aae),
	.w8(32'h3a6b97ed),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85c48c),
	.w1(32'hba598cfa),
	.w2(32'hba3f43f2),
	.w3(32'h39479f4a),
	.w4(32'h3a6b032b),
	.w5(32'hba825631),
	.w6(32'h39a895f5),
	.w7(32'h3a4a961b),
	.w8(32'hbb0f24be),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b6fa6),
	.w1(32'hbbb4e9cf),
	.w2(32'hbbd730f4),
	.w3(32'hbba3df00),
	.w4(32'hbbfaaa66),
	.w5(32'hbb9ab402),
	.w6(32'hbbdec482),
	.w7(32'hbc000f1b),
	.w8(32'hbbbc3170),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba843673),
	.w1(32'h3ac395b9),
	.w2(32'h3a85340c),
	.w3(32'h3a278f33),
	.w4(32'h3b147ad3),
	.w5(32'h3b045c02),
	.w6(32'hb907ff64),
	.w7(32'h392d72be),
	.w8(32'h38af0f4a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b272897),
	.w1(32'h3a3f18a3),
	.w2(32'hbbf4e367),
	.w3(32'h3bb8b9fd),
	.w4(32'h3a94d47a),
	.w5(32'hbba67536),
	.w6(32'h3b423fa7),
	.w7(32'hba828911),
	.w8(32'hbbc7ac83),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49afda),
	.w1(32'h3a1599a0),
	.w2(32'h3ab15c95),
	.w3(32'h3ad238d6),
	.w4(32'h3acb125d),
	.w5(32'h3abe7b37),
	.w6(32'h39208458),
	.w7(32'h39bcf75d),
	.w8(32'h3a522032),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb563a4f),
	.w1(32'hbbcbff4a),
	.w2(32'hbb7a9da6),
	.w3(32'hb34c4800),
	.w4(32'hbb383df4),
	.w5(32'hbab7489e),
	.w6(32'hba011b40),
	.w7(32'hbb8bdc8e),
	.w8(32'hbbad37ae),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb189cc0),
	.w1(32'h399327cd),
	.w2(32'h3ab83ce4),
	.w3(32'h3ae3acf3),
	.w4(32'h3ae26510),
	.w5(32'h3913affe),
	.w6(32'h3a590056),
	.w7(32'h39b490b1),
	.w8(32'hb9837304),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9beeb3),
	.w1(32'h3acd62c7),
	.w2(32'h3b3a7424),
	.w3(32'h3ad15435),
	.w4(32'h3b5ef9d4),
	.w5(32'h3b5d7f50),
	.w6(32'h3ac56f2d),
	.w7(32'h3a9ab883),
	.w8(32'h3aa8133e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a087a46),
	.w1(32'h39e78dd0),
	.w2(32'hbacf6c4e),
	.w3(32'h3a822863),
	.w4(32'hbaa25e9c),
	.w5(32'hba8eb336),
	.w6(32'h3b076e66),
	.w7(32'hb91be6a7),
	.w8(32'h3a005398),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88d453),
	.w1(32'hbb97d07b),
	.w2(32'hbbc5e790),
	.w3(32'hba074f61),
	.w4(32'hbb51d9aa),
	.w5(32'hbb6a080e),
	.w6(32'h39a9ec3e),
	.w7(32'hbb35689f),
	.w8(32'hbb748037),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f924a),
	.w1(32'hba9c8b8f),
	.w2(32'hbb220153),
	.w3(32'hbb2446d7),
	.w4(32'h3999aa25),
	.w5(32'hbaba3df8),
	.w6(32'hbb8373a0),
	.w7(32'hbb3ee8eb),
	.w8(32'hbbde6a8a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fa3f4),
	.w1(32'hbb2370af),
	.w2(32'hbc384bef),
	.w3(32'hbbad0df6),
	.w4(32'h3aba814a),
	.w5(32'h3aa0d922),
	.w6(32'hbc3d44f4),
	.w7(32'hba8c479e),
	.w8(32'h3b13887c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b070bcf),
	.w1(32'h3c5d19b0),
	.w2(32'h3bb8c434),
	.w3(32'h3bed10e9),
	.w4(32'h3c34f7ab),
	.w5(32'h3be53e65),
	.w6(32'h3b94672e),
	.w7(32'h3c22391a),
	.w8(32'hbb86a83c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8841e4),
	.w1(32'hbbbed7cf),
	.w2(32'hbb80ce09),
	.w3(32'hbae2c0c5),
	.w4(32'h3b531474),
	.w5(32'h3abb5208),
	.w6(32'hbb4007d2),
	.w7(32'hbafe94d1),
	.w8(32'hba6b0a8b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ade18),
	.w1(32'h38b292e1),
	.w2(32'hbc447df6),
	.w3(32'h3b214659),
	.w4(32'hba250117),
	.w5(32'h3bae383d),
	.w6(32'h3a938e3f),
	.w7(32'hbaa62892),
	.w8(32'h3b213cb3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6abc61),
	.w1(32'h3aaaa25c),
	.w2(32'h3c0771d1),
	.w3(32'h3ac2f986),
	.w4(32'h3c1c643a),
	.w5(32'hbb056b0e),
	.w6(32'hbc0f0277),
	.w7(32'h3bf9af0f),
	.w8(32'hbbad05a3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3977c),
	.w1(32'h38eb5ed8),
	.w2(32'hbc9f0164),
	.w3(32'hbc69a357),
	.w4(32'hbc4a2b28),
	.w5(32'hbc8a6fa7),
	.w6(32'hbcb82bce),
	.w7(32'hbc6eec26),
	.w8(32'hbc61f6c7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb998c6e),
	.w1(32'hbb48373b),
	.w2(32'hbc244f5b),
	.w3(32'hbba7ce43),
	.w4(32'hbb275495),
	.w5(32'hbbd10b50),
	.w6(32'h3b9462a6),
	.w7(32'hba568281),
	.w8(32'hbc0325ca),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bf5f2),
	.w1(32'h390b9d97),
	.w2(32'hbb50252b),
	.w3(32'hbbea5e15),
	.w4(32'hbb9ddbe8),
	.w5(32'h3ab37bba),
	.w6(32'h3a6f52f7),
	.w7(32'hbbdda225),
	.w8(32'h3b24875e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23a7a1),
	.w1(32'hbb3d8958),
	.w2(32'hba1c9b80),
	.w3(32'hbab59a70),
	.w4(32'h3a004899),
	.w5(32'h3b5fde7f),
	.w6(32'hbb8d5633),
	.w7(32'hbae3c300),
	.w8(32'h39465902),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b524f24),
	.w1(32'hbb3cb12d),
	.w2(32'h3aa24cc4),
	.w3(32'hbb790dd1),
	.w4(32'h3a537da5),
	.w5(32'hbb80c80d),
	.w6(32'hbbf450e7),
	.w7(32'hbaa8fb4b),
	.w8(32'hbb1dc232),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6cf46),
	.w1(32'hbb71d44e),
	.w2(32'hbbd498dd),
	.w3(32'hbb2c4c56),
	.w4(32'hbbb7236e),
	.w5(32'hbab52ac7),
	.w6(32'h3b17b265),
	.w7(32'hbb57e239),
	.w8(32'hbb10c608),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd782e),
	.w1(32'hbc180a24),
	.w2(32'hbb9427d6),
	.w3(32'hbb95eb23),
	.w4(32'hbb25aaba),
	.w5(32'hbbb90781),
	.w6(32'hbaec9614),
	.w7(32'hbb8ed8c4),
	.w8(32'hba9bf44b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b97116),
	.w1(32'h3ad0faae),
	.w2(32'h3b128666),
	.w3(32'hbb99978b),
	.w4(32'h3b3bad93),
	.w5(32'hbaca7c25),
	.w6(32'hb85c7d38),
	.w7(32'h3a335a7c),
	.w8(32'hbba4616c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba467ff),
	.w1(32'h3b3ab28f),
	.w2(32'hbb82beab),
	.w3(32'hba9b2a24),
	.w4(32'hbb883c3b),
	.w5(32'hba973df1),
	.w6(32'h3b6d3669),
	.w7(32'hbb23cddd),
	.w8(32'h3baa6923),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f97574),
	.w1(32'h3abede7c),
	.w2(32'hbb63b300),
	.w3(32'hba8b1ce1),
	.w4(32'h392ee4dc),
	.w5(32'hbbf436b7),
	.w6(32'h3aa190f3),
	.w7(32'h3b105318),
	.w8(32'hbc03fee8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac65517),
	.w1(32'hbbd318f7),
	.w2(32'h3abb0bac),
	.w3(32'hbbd678ad),
	.w4(32'h3ae2109a),
	.w5(32'hbbad2e0d),
	.w6(32'h3ad7a76e),
	.w7(32'hbb9d4033),
	.w8(32'hbb529a40),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e53aa),
	.w1(32'hbb038881),
	.w2(32'h3a3b8de7),
	.w3(32'hbbb22cdc),
	.w4(32'h3b032765),
	.w5(32'hb896bb64),
	.w6(32'h39fca104),
	.w7(32'h3aff5c64),
	.w8(32'h3a8edcf9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2e48c),
	.w1(32'h3bdc4270),
	.w2(32'h3b51be40),
	.w3(32'h3b187840),
	.w4(32'h3ae81eb0),
	.w5(32'h3a95ec66),
	.w6(32'h3b6c089d),
	.w7(32'h3b83636e),
	.w8(32'hbb21b224),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e4862),
	.w1(32'hbbbb43d9),
	.w2(32'hbb5da23d),
	.w3(32'hbaf31b3e),
	.w4(32'h391a72d9),
	.w5(32'hba8e25ee),
	.w6(32'hbb2ea6ce),
	.w7(32'hbb66afda),
	.w8(32'hbb7d85d9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c29314),
	.w1(32'hbb9456ab),
	.w2(32'hbac33ff0),
	.w3(32'hbbc24ae2),
	.w4(32'hbaa8cb97),
	.w5(32'hb926f747),
	.w6(32'hbc292559),
	.w7(32'hbb6f5e81),
	.w8(32'hba6599b8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b876ddd),
	.w1(32'hb9da4cd6),
	.w2(32'h3b554bf2),
	.w3(32'hbbbcc82b),
	.w4(32'hba1be52e),
	.w5(32'hbbb30c1a),
	.w6(32'hbb04a3a6),
	.w7(32'h3b1f097e),
	.w8(32'h3a64f774),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcb699),
	.w1(32'h3b83baa0),
	.w2(32'hba796ef6),
	.w3(32'hbb86fa9b),
	.w4(32'h39a8ddea),
	.w5(32'hbb867a3b),
	.w6(32'h3c116bc1),
	.w7(32'h3b948b8e),
	.w8(32'hbb6aad38),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcb2ce),
	.w1(32'h3ad43a5b),
	.w2(32'hbb779f5b),
	.w3(32'h3a3744c8),
	.w4(32'hb9da4c61),
	.w5(32'hbb65fcb5),
	.w6(32'h38b5fce8),
	.w7(32'hbaf041ab),
	.w8(32'hbb8e3d9f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95574),
	.w1(32'hbba78501),
	.w2(32'hbb274af3),
	.w3(32'hbbcd32b7),
	.w4(32'h3981d8e9),
	.w5(32'h3b4a9850),
	.w6(32'h3b21930b),
	.w7(32'hbba41874),
	.w8(32'hbb9c20a1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca0e38),
	.w1(32'hbb08e779),
	.w2(32'hba728b9f),
	.w3(32'hbb269948),
	.w4(32'hbb85af49),
	.w5(32'hbb1538d2),
	.w6(32'hbade16bb),
	.w7(32'hbb8a4730),
	.w8(32'hbb8c5ab5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77b9ac),
	.w1(32'hbb64eb0a),
	.w2(32'hbb606c03),
	.w3(32'hbb555f11),
	.w4(32'hb9a6e432),
	.w5(32'h3afe94c9),
	.w6(32'hbb194a45),
	.w7(32'hbb4d1baa),
	.w8(32'h3ab777b1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb42335),
	.w1(32'hbb5e4265),
	.w2(32'hb872f303),
	.w3(32'hb87607cf),
	.w4(32'hba480a86),
	.w5(32'h3aca17e0),
	.w6(32'h3b8b5ed0),
	.w7(32'h3b7cbf80),
	.w8(32'h3b96bf93),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4ab4f),
	.w1(32'hba74ed20),
	.w2(32'hbb0969a6),
	.w3(32'hbb1bdec6),
	.w4(32'hba99b962),
	.w5(32'h397ba84e),
	.w6(32'hba8cb6f0),
	.w7(32'h3a046a72),
	.w8(32'h3a5e3a0f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b371a96),
	.w1(32'h3ae47aa9),
	.w2(32'h396a719a),
	.w3(32'h3b8f850c),
	.w4(32'h3aad3968),
	.w5(32'hbc6fbbff),
	.w6(32'h3c0e4d3f),
	.w7(32'h3b1cfcc2),
	.w8(32'hbc2bf8e3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11c238),
	.w1(32'hbc34707c),
	.w2(32'hbc92ee64),
	.w3(32'hbc2c8603),
	.w4(32'hbc4534b8),
	.w5(32'hbaed9030),
	.w6(32'hb9deda06),
	.w7(32'hbc287be9),
	.w8(32'hbb31fa5e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb100ec6),
	.w1(32'hbb339f21),
	.w2(32'hbaf387ab),
	.w3(32'hbb39d1d8),
	.w4(32'hbb56e83f),
	.w5(32'hbbf608af),
	.w6(32'h3a66379a),
	.w7(32'hbb181642),
	.w8(32'hbb90f2e2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66dc4f),
	.w1(32'hbb5347b1),
	.w2(32'hbbbe1cc9),
	.w3(32'hbbf49abc),
	.w4(32'hba6caeb9),
	.w5(32'hbafc0a85),
	.w6(32'h3a679922),
	.w7(32'h3a8d8a01),
	.w8(32'hbb185b48),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a926357),
	.w1(32'h3b210665),
	.w2(32'h3b314702),
	.w3(32'hba54be5e),
	.w4(32'h3afdb52c),
	.w5(32'h3b8e9a11),
	.w6(32'hbbb41943),
	.w7(32'hbaaa5539),
	.w8(32'hbbb1cb9d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae3d65),
	.w1(32'hbb8232ee),
	.w2(32'h39ccfa2e),
	.w3(32'hbaa54225),
	.w4(32'h3b937595),
	.w5(32'hb9909d0a),
	.w6(32'hbc317ca3),
	.w7(32'hbbb31b16),
	.w8(32'hba3f579b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb95ad8),
	.w1(32'h398c724f),
	.w2(32'hbab6533a),
	.w3(32'hb983a15a),
	.w4(32'hba0a7c63),
	.w5(32'hbac66931),
	.w6(32'hba980c67),
	.w7(32'hbb3635c6),
	.w8(32'hba88de23),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b652235),
	.w1(32'h395e7c4f),
	.w2(32'hbc21209d),
	.w3(32'h39df052c),
	.w4(32'hbb4f1e29),
	.w5(32'hbc24344e),
	.w6(32'h3b52e4b0),
	.w7(32'hbba43359),
	.w8(32'hbc23c1c2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23d9d5),
	.w1(32'h3b030807),
	.w2(32'hbb7d070e),
	.w3(32'h399be773),
	.w4(32'h3b703ddb),
	.w5(32'h3a41a855),
	.w6(32'h3aa3417c),
	.w7(32'h392ae44c),
	.w8(32'hba0454a2),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83a64e),
	.w1(32'h3a75cf7b),
	.w2(32'hbb9374b1),
	.w3(32'h3ac9c44d),
	.w4(32'hba8e3281),
	.w5(32'hba81b427),
	.w6(32'h3b3ec16f),
	.w7(32'hba6c4cc1),
	.w8(32'hbb09ce4d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62efbb),
	.w1(32'h39246202),
	.w2(32'hbc03eb25),
	.w3(32'h3b1f464d),
	.w4(32'hbb5a8e2e),
	.w5(32'hbb91e456),
	.w6(32'h3aa4c606),
	.w7(32'hbb0c629c),
	.w8(32'hbbba92d0),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb769f7b),
	.w1(32'h3b83a50c),
	.w2(32'h39b6aa29),
	.w3(32'h3a33af20),
	.w4(32'h3b487324),
	.w5(32'h3ac81364),
	.w6(32'hbb67530f),
	.w7(32'h3a98e0dc),
	.w8(32'hbadb8c05),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada9f61),
	.w1(32'hbb9b3579),
	.w2(32'hbc646b36),
	.w3(32'hbb716f9c),
	.w4(32'hbb000ecb),
	.w5(32'hbb84ca1a),
	.w6(32'h3b8a2858),
	.w7(32'hbab20068),
	.w8(32'hbc0fbd02),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba024c9),
	.w1(32'hbbea2b4b),
	.w2(32'hbc12ca1a),
	.w3(32'hbb15f429),
	.w4(32'hb9d84a68),
	.w5(32'h3af994ac),
	.w6(32'hbaac3362),
	.w7(32'hbbef5ea5),
	.w8(32'hba06f4f8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a8f9d),
	.w1(32'hba2a4a72),
	.w2(32'h3b6a1cbd),
	.w3(32'h3b182595),
	.w4(32'h3bbaad66),
	.w5(32'h3ab629bb),
	.w6(32'h3af95b9b),
	.w7(32'h3900c5d8),
	.w8(32'hbabefc7a),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b5722),
	.w1(32'hbaa812f8),
	.w2(32'hbac5c13f),
	.w3(32'hb92c4ead),
	.w4(32'h3a765465),
	.w5(32'h3ac6d8b1),
	.w6(32'h3a4d0914),
	.w7(32'hba7edadb),
	.w8(32'hbb11e1dc),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9400f),
	.w1(32'h396daea8),
	.w2(32'hbaf4c2ed),
	.w3(32'hbaa918fc),
	.w4(32'hbb801fb7),
	.w5(32'h3b168a97),
	.w6(32'hba470ef1),
	.w7(32'hbbb92aab),
	.w8(32'h3b11e4eb),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399078ac),
	.w1(32'hbab0c27a),
	.w2(32'hbb601798),
	.w3(32'h38995ff2),
	.w4(32'hba9febe4),
	.w5(32'hbabfca2b),
	.w6(32'h3a96ec75),
	.w7(32'hbaedccb6),
	.w8(32'hbb136605),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c67ef9),
	.w1(32'hba927e9d),
	.w2(32'h38fba498),
	.w3(32'hbb1e78c2),
	.w4(32'h3afc2437),
	.w5(32'h3adf1bc8),
	.w6(32'h3a460576),
	.w7(32'hb9eca59c),
	.w8(32'hbadef8ff),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b91fd),
	.w1(32'hbb415ee7),
	.w2(32'h398e5db1),
	.w3(32'h3938c9ba),
	.w4(32'h3ba611aa),
	.w5(32'hb9248dc8),
	.w6(32'hbb8fcce8),
	.w7(32'hbb2b0f48),
	.w8(32'hbb98d17d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ff35),
	.w1(32'hba660ecb),
	.w2(32'h3b84de4a),
	.w3(32'hba218b11),
	.w4(32'hba2e00fa),
	.w5(32'hbb8d4261),
	.w6(32'h3bb1f202),
	.w7(32'h3acceb23),
	.w8(32'hbb94ad83),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88f7d8),
	.w1(32'h3a9a0be5),
	.w2(32'hbac2dafa),
	.w3(32'h3a8ffd4f),
	.w4(32'hbbb88125),
	.w5(32'hb9bd8ec4),
	.w6(32'h39839ca3),
	.w7(32'hbbbe4c5b),
	.w8(32'h3abac4a3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b9d98),
	.w1(32'h3b59ec21),
	.w2(32'h3b66636d),
	.w3(32'h3ae5376c),
	.w4(32'h39d123cf),
	.w5(32'hbbbdaf02),
	.w6(32'h3a8cb741),
	.w7(32'h3bab18d2),
	.w8(32'hbb8a84e4),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23d1b9),
	.w1(32'hbade5af8),
	.w2(32'hbb92db0b),
	.w3(32'h3899f6f2),
	.w4(32'hbb15410b),
	.w5(32'hbba55f79),
	.w6(32'h3b457b54),
	.w7(32'h383cf825),
	.w8(32'hbc1a02dc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4b664),
	.w1(32'h3ab9c2a4),
	.w2(32'hbc663ce3),
	.w3(32'h3b1cf10b),
	.w4(32'hbbd94bca),
	.w5(32'hbc03ff06),
	.w6(32'hba0d4a38),
	.w7(32'hbc4273e2),
	.w8(32'hbbafb70f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb649134),
	.w1(32'hbb56cc2f),
	.w2(32'hbb386972),
	.w3(32'hbb09d5c0),
	.w4(32'hbac2208f),
	.w5(32'h3a1aee14),
	.w6(32'h3c0166d3),
	.w7(32'hbb83c248),
	.w8(32'h3a70e1fb),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc30a6),
	.w1(32'h3b9bb1c8),
	.w2(32'h3b1ddfd2),
	.w3(32'h3b880b70),
	.w4(32'h3a5412fd),
	.w5(32'h3bdb72d3),
	.w6(32'h3b578c88),
	.w7(32'h3b5c36e3),
	.w8(32'h3be8730c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf30f7b),
	.w1(32'h3c0b5674),
	.w2(32'h3bf7b421),
	.w3(32'h3bb4395c),
	.w4(32'h3bb33958),
	.w5(32'hbb8e3c07),
	.w6(32'h3b5ddccc),
	.w7(32'h3bf39d5c),
	.w8(32'hbb436149),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b6e34),
	.w1(32'hbbc8ee4d),
	.w2(32'hbc17130a),
	.w3(32'hbbb72d4e),
	.w4(32'hbc1bee4a),
	.w5(32'h3b18c2a2),
	.w6(32'hb99cb7f3),
	.w7(32'hbbf5a57b),
	.w8(32'hba27ea79),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc110224),
	.w1(32'h3aebed53),
	.w2(32'h3b32cd2e),
	.w3(32'hb9794ec2),
	.w4(32'h3ab1fc99),
	.w5(32'hbb873ef2),
	.w6(32'hb9e63f39),
	.w7(32'hba3416d0),
	.w8(32'hbc1f3db4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8acf85),
	.w1(32'h3b37b4b5),
	.w2(32'h3af964a0),
	.w3(32'h38c22770),
	.w4(32'h3afc0a8d),
	.w5(32'hbaaac9e3),
	.w6(32'hba7eb832),
	.w7(32'hbb7117f2),
	.w8(32'hbb3a17b7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd99fb5),
	.w1(32'hbc4ffd27),
	.w2(32'hbc03cfb9),
	.w3(32'hbb84beea),
	.w4(32'hbbc7cfcd),
	.w5(32'hbb7a0f12),
	.w6(32'hbba428f4),
	.w7(32'hbbf93113),
	.w8(32'hbb99e010),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed1487),
	.w1(32'hbb963715),
	.w2(32'hbc0221f7),
	.w3(32'hbc4aa505),
	.w4(32'hba8d6448),
	.w5(32'hbbbdd9c0),
	.w6(32'hbb2df549),
	.w7(32'hbbebf9f7),
	.w8(32'hbbf9f04a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1875d),
	.w1(32'h39c507d7),
	.w2(32'hbb664744),
	.w3(32'hb988f34a),
	.w4(32'hbb262507),
	.w5(32'h3a96f06a),
	.w6(32'h3c1a0b3e),
	.w7(32'hbbb2b1c9),
	.w8(32'hbba2a37b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c72d6),
	.w1(32'hb99e09e8),
	.w2(32'hbb0fccf8),
	.w3(32'h3a7f8545),
	.w4(32'hbb38be3a),
	.w5(32'hb94ecbf2),
	.w6(32'h3b5742ba),
	.w7(32'hbbc0381f),
	.w8(32'hbb39bc53),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfad34c),
	.w1(32'hbb2948d1),
	.w2(32'h3b28955f),
	.w3(32'hb9900c86),
	.w4(32'hbc017e78),
	.w5(32'hbc0495cc),
	.w6(32'h3bd753b1),
	.w7(32'h3ac85c11),
	.w8(32'hbbb672d4),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76889c),
	.w1(32'hbb80a9fe),
	.w2(32'hbbbd0d2c),
	.w3(32'hbb4a2c92),
	.w4(32'hbb14ed41),
	.w5(32'hbb9f8fe5),
	.w6(32'h3a78deb6),
	.w7(32'hbbcb892d),
	.w8(32'hbb91e4e1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b623f0e),
	.w1(32'hbb44239c),
	.w2(32'h3aec5954),
	.w3(32'hb862d547),
	.w4(32'hbc360bf6),
	.w5(32'h3b2d8edd),
	.w6(32'h3be7997e),
	.w7(32'hba5fe528),
	.w8(32'h3b4c56f4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8747d6),
	.w1(32'h3bb9e494),
	.w2(32'hbaf3e9a0),
	.w3(32'h3bc36882),
	.w4(32'h37e6b2be),
	.w5(32'hb9c83689),
	.w6(32'h3aaeaded),
	.w7(32'hbaa8a27b),
	.w8(32'hbb46203a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c5d4b),
	.w1(32'hbb666f32),
	.w2(32'hbb36f89d),
	.w3(32'hbb2e5ef9),
	.w4(32'hbbdfb389),
	.w5(32'h3b905dd6),
	.w6(32'h3a020321),
	.w7(32'hbb391889),
	.w8(32'h3c1d4fd2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c875c1c),
	.w1(32'h3c0b9056),
	.w2(32'h3c0e6a1b),
	.w3(32'h3bb73e4b),
	.w4(32'h3c14a740),
	.w5(32'h3a79cf93),
	.w6(32'hbc14c86d),
	.w7(32'h3c163a46),
	.w8(32'h3a6cdef6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefb760),
	.w1(32'hbb072685),
	.w2(32'hbc3e5a4f),
	.w3(32'hbb566525),
	.w4(32'hbbcc1219),
	.w5(32'hb90a92b4),
	.w6(32'h3b252c96),
	.w7(32'hbb80bb50),
	.w8(32'h3b75a0f7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb7491),
	.w1(32'h3c0f2751),
	.w2(32'h3ba04dd5),
	.w3(32'h3bcff927),
	.w4(32'h3b842866),
	.w5(32'hbb9f4c5f),
	.w6(32'h3b77362b),
	.w7(32'h3bd7fbb4),
	.w8(32'hbb9460fe),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdedf01),
	.w1(32'hbacb8edc),
	.w2(32'hb9b82702),
	.w3(32'hbba138da),
	.w4(32'hbb8ae990),
	.w5(32'h3ad1b2c3),
	.w6(32'h390c2aa3),
	.w7(32'hbb872e69),
	.w8(32'hbb6fc882),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba509d7),
	.w1(32'hbc33bf9d),
	.w2(32'hbad1709b),
	.w3(32'hbbe09c15),
	.w4(32'h3a5ed76a),
	.w5(32'h3a8e5ba5),
	.w6(32'hbc2ce599),
	.w7(32'hbbf9b9fd),
	.w8(32'h3aafe5d6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dbf2c),
	.w1(32'h3ba1a829),
	.w2(32'h3b66f2c2),
	.w3(32'h3abb0c35),
	.w4(32'hbb0a9e23),
	.w5(32'hbb97fc9a),
	.w6(32'h3b37d118),
	.w7(32'hba80be99),
	.w8(32'h39645865),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b6915),
	.w1(32'hbbdfd897),
	.w2(32'hbbfe27c0),
	.w3(32'hbb9efc33),
	.w4(32'hbb9c8c0f),
	.w5(32'h3b815126),
	.w6(32'hbbc1c579),
	.w7(32'hb75004ee),
	.w8(32'h3b41c24f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2e8fd),
	.w1(32'hbb0ee353),
	.w2(32'hbb59f28c),
	.w3(32'hb75f35c0),
	.w4(32'hbb4eafee),
	.w5(32'hbaa8cbca),
	.w6(32'hbb99fd0c),
	.w7(32'h3990afcc),
	.w8(32'h37d83c3c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cc72a),
	.w1(32'h3bdbe177),
	.w2(32'h3b909879),
	.w3(32'h3b837b1a),
	.w4(32'h3ad4f8e8),
	.w5(32'hbbea6ca4),
	.w6(32'h3b95d0e8),
	.w7(32'h3b8f4bbc),
	.w8(32'hbb155bfa),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7e15a),
	.w1(32'hbbc077f0),
	.w2(32'hbbc075f5),
	.w3(32'hbb6371ce),
	.w4(32'hbb938604),
	.w5(32'hba6bb6b2),
	.w6(32'h3bbf7318),
	.w7(32'hbbb04738),
	.w8(32'h3a56cc63),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b621c2f),
	.w1(32'h3bea867a),
	.w2(32'h3b8d69a2),
	.w3(32'h3acff690),
	.w4(32'hba6380e9),
	.w5(32'h3b93c444),
	.w6(32'h3b3f4284),
	.w7(32'h3b80301b),
	.w8(32'h3b02199e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba36920),
	.w1(32'hbba46b9e),
	.w2(32'hbb208713),
	.w3(32'hbc0826fb),
	.w4(32'h39c9f470),
	.w5(32'h3a9443d2),
	.w6(32'hbbed2ac1),
	.w7(32'hbb0e8feb),
	.w8(32'hbaf0fc5d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb832a5b),
	.w1(32'hbc0622fc),
	.w2(32'h373dd820),
	.w3(32'hbbab70f6),
	.w4(32'h3b5a6712),
	.w5(32'hbbc4caa3),
	.w6(32'hbb6029f2),
	.w7(32'hbae0d4c9),
	.w8(32'hbbdf8f9b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad7732),
	.w1(32'h393d547e),
	.w2(32'hba9a7186),
	.w3(32'hbb959ba3),
	.w4(32'h3b5cccc5),
	.w5(32'hba14ab5c),
	.w6(32'hbba487c2),
	.w7(32'h3adddad3),
	.w8(32'hba7c4c06),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b412753),
	.w1(32'h3afd1799),
	.w2(32'hbc0c5947),
	.w3(32'h3aa9691d),
	.w4(32'hbc1eb82d),
	.w5(32'hb9dacaac),
	.w6(32'h3b5b645e),
	.w7(32'hbbb12a91),
	.w8(32'hbabf8c57),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd15cc),
	.w1(32'hbac6c85e),
	.w2(32'h3b25eec6),
	.w3(32'h39d61520),
	.w4(32'h3a97a479),
	.w5(32'h3ac4772a),
	.w6(32'h3aff6899),
	.w7(32'h3a9e6ff4),
	.w8(32'hb9baaa1f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d60d2),
	.w1(32'hbb01aabb),
	.w2(32'hbb3cf27a),
	.w3(32'hbba1ad27),
	.w4(32'hbbb68038),
	.w5(32'h3b13b204),
	.w6(32'hba8d4b6d),
	.w7(32'hbbf40ca3),
	.w8(32'h3af0974c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4da3d1),
	.w1(32'hba397792),
	.w2(32'hbba5991f),
	.w3(32'hb835b8e4),
	.w4(32'hbb75b483),
	.w5(32'hbb7485f6),
	.w6(32'h3b9d9cd5),
	.w7(32'hbbbd6a23),
	.w8(32'hbc28ad4e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3bd6c),
	.w1(32'h3bbf3b0d),
	.w2(32'hbba96851),
	.w3(32'hba7cb6cc),
	.w4(32'hbb0740e9),
	.w5(32'hb83ab069),
	.w6(32'hbadfa8c0),
	.w7(32'hbaa2bd75),
	.w8(32'h3adf35d0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b238c7d),
	.w1(32'h3bf08ae7),
	.w2(32'h3aec89a2),
	.w3(32'h3b60e527),
	.w4(32'h3a3cd798),
	.w5(32'h3b6b2459),
	.w6(32'h3bdcfff0),
	.w7(32'h3b5d9c71),
	.w8(32'h3bcdd176),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d7390),
	.w1(32'hbbd9c422),
	.w2(32'hb8cc3b4b),
	.w3(32'h39efe1fe),
	.w4(32'h3a81de36),
	.w5(32'hbc140eeb),
	.w6(32'hbbd148d2),
	.w7(32'h3c363bb4),
	.w8(32'hbbab0e2e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc036e8e),
	.w1(32'hbb9e1b0b),
	.w2(32'h3acf3c01),
	.w3(32'hbb4c60ae),
	.w4(32'hba508b1f),
	.w5(32'hba82c856),
	.w6(32'hbb5c74bc),
	.w7(32'hbb5040fd),
	.w8(32'hbaa2689c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9ca61),
	.w1(32'hbb8692cd),
	.w2(32'hbbf224f9),
	.w3(32'hbb7656b7),
	.w4(32'hbba5172b),
	.w5(32'hbb455581),
	.w6(32'hb86ee4ba),
	.w7(32'hbb031fa2),
	.w8(32'hbc066619),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91edee),
	.w1(32'hbb9d1018),
	.w2(32'h3ae131ca),
	.w3(32'hbb458206),
	.w4(32'hbb5cc689),
	.w5(32'h3b7de082),
	.w6(32'hbb066798),
	.w7(32'hbb083572),
	.w8(32'h3b5496a3),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c5e45),
	.w1(32'h3b00fa37),
	.w2(32'h3a8e6e02),
	.w3(32'h39760f33),
	.w4(32'hbbbe354d),
	.w5(32'h3aa1d590),
	.w6(32'h3beec9df),
	.w7(32'hbaf4ea34),
	.w8(32'h3a6aea99),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f2b9e),
	.w1(32'hba9e6d62),
	.w2(32'hbaeb3f5a),
	.w3(32'h3989638e),
	.w4(32'hbb5b63d7),
	.w5(32'hb9ac5bc2),
	.w6(32'h3b451d89),
	.w7(32'hbb701796),
	.w8(32'hbb8b3441),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954ab2d),
	.w1(32'hbb49db5c),
	.w2(32'hbbac7646),
	.w3(32'hba47c067),
	.w4(32'h3b29da3e),
	.w5(32'hbbe2eb28),
	.w6(32'hbab2073b),
	.w7(32'hb92059df),
	.w8(32'hbbbb6061),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b5fb1),
	.w1(32'hbb246b50),
	.w2(32'hbbe6a481),
	.w3(32'hbb736b83),
	.w4(32'hbb8deecb),
	.w5(32'h3bd8f3e4),
	.w6(32'h3ac3972c),
	.w7(32'hbb5f56d1),
	.w8(32'h3bc591d1),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cc361),
	.w1(32'h3c671c87),
	.w2(32'h3c72a2e8),
	.w3(32'h3c30c924),
	.w4(32'h3c0d760b),
	.w5(32'hbb29db0c),
	.w6(32'h3c26f13d),
	.w7(32'h3c1661d1),
	.w8(32'hbb7ae4a5),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f96ce),
	.w1(32'hbb4ab9b5),
	.w2(32'hba466080),
	.w3(32'h3a18fe10),
	.w4(32'h3b429c59),
	.w5(32'hbc1876c8),
	.w6(32'h3b447351),
	.w7(32'hbaa4729e),
	.w8(32'hbc0f358f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1efff),
	.w1(32'hbc1accd3),
	.w2(32'hbc4a9702),
	.w3(32'hbc15c2c6),
	.w4(32'hbb989be9),
	.w5(32'hbbb0fb9c),
	.w6(32'hbb10a74d),
	.w7(32'hbbf5ea2a),
	.w8(32'hbb947282),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39974142),
	.w1(32'h3b23b41f),
	.w2(32'h388b7cfb),
	.w3(32'h394eff63),
	.w4(32'hb8235c55),
	.w5(32'hbb7ccb3e),
	.w6(32'h389449ab),
	.w7(32'h3aee647a),
	.w8(32'hbb5504c4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a468d80),
	.w1(32'hba9148c5),
	.w2(32'hbaf48458),
	.w3(32'h3b9522f8),
	.w4(32'h3aaf6b2b),
	.w5(32'hbaca3d9d),
	.w6(32'hbabfdb67),
	.w7(32'hba02f18f),
	.w8(32'hbb301113),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16defd),
	.w1(32'hbbc1d51b),
	.w2(32'hbbe173d6),
	.w3(32'hbb92a5d5),
	.w4(32'hbb65943b),
	.w5(32'h3a862009),
	.w6(32'hbb75dc98),
	.w7(32'hbb8b5c1d),
	.w8(32'hba079c14),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9853baa),
	.w1(32'h3adc6fa8),
	.w2(32'h3aed6898),
	.w3(32'h3b610e3b),
	.w4(32'hbb5299c9),
	.w5(32'hbb0ec5ef),
	.w6(32'h3bd1b84e),
	.w7(32'h3a8eb9ab),
	.w8(32'hbb3e4670),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba86caa),
	.w1(32'hbb40259c),
	.w2(32'hbc11d8b1),
	.w3(32'hbb7e8683),
	.w4(32'hbbb3af87),
	.w5(32'h3b1f52ea),
	.w6(32'h3a4485dc),
	.w7(32'hbbc44ae3),
	.w8(32'hba65a245),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87cc20),
	.w1(32'hbb942ed2),
	.w2(32'hb9dd9ff5),
	.w3(32'h393a1ce1),
	.w4(32'h3ba9baa5),
	.w5(32'h3b1482d1),
	.w6(32'hbaa55ce3),
	.w7(32'hbbabff10),
	.w8(32'hbb0f7db9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c51a23),
	.w1(32'hbaba02d9),
	.w2(32'hbbe07f2f),
	.w3(32'hba512961),
	.w4(32'h3b10030a),
	.w5(32'h3ac1d3c1),
	.w6(32'h3b03f029),
	.w7(32'h3a7cd824),
	.w8(32'hbb1e5b71),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b610ca0),
	.w1(32'hbb4851ab),
	.w2(32'hbaa07b10),
	.w3(32'hbb8595f7),
	.w4(32'h3ac0ab62),
	.w5(32'h3c20866b),
	.w6(32'hbbe5e399),
	.w7(32'hbbe3840b),
	.w8(32'h3bf13331),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18cc0d),
	.w1(32'h39f1df17),
	.w2(32'h3bab7f7b),
	.w3(32'h3bb53b23),
	.w4(32'h3c7b00e2),
	.w5(32'hbb7a0ae9),
	.w6(32'hbb1cad1c),
	.w7(32'h3be1f6f7),
	.w8(32'hbb94c9d8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca9f40),
	.w1(32'hbbb86b04),
	.w2(32'hbbfd50c2),
	.w3(32'hbb5a0b4d),
	.w4(32'hbbfede10),
	.w5(32'hbab3ff8e),
	.w6(32'h3969300d),
	.w7(32'hbba4f238),
	.w8(32'h3ac2027b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e0631),
	.w1(32'h3bf367ba),
	.w2(32'h3bbae998),
	.w3(32'h3b18d8d8),
	.w4(32'h3b0ec31b),
	.w5(32'hbbc04c0e),
	.w6(32'h3b11bead),
	.w7(32'h3b9189fd),
	.w8(32'hbb1d0306),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb065e0d),
	.w1(32'hbbbe2329),
	.w2(32'hbb6ea0a1),
	.w3(32'hbb7d8bc8),
	.w4(32'hbb12516d),
	.w5(32'hbb8628e3),
	.w6(32'h3b14764b),
	.w7(32'hbb08428f),
	.w8(32'hba8939c9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cbb1b),
	.w1(32'h3ab9322b),
	.w2(32'hbba4e6e0),
	.w3(32'hb996abba),
	.w4(32'h3b02b0bc),
	.w5(32'h3c139ea6),
	.w6(32'h3b1de87f),
	.w7(32'h3abb4ba3),
	.w8(32'h3bdb2534),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c161e1c),
	.w1(32'h3c0b90ee),
	.w2(32'h3c5f0a03),
	.w3(32'h3bfe717a),
	.w4(32'h3c16df32),
	.w5(32'hbc22ac5d),
	.w6(32'hb9c4489a),
	.w7(32'h3c43c020),
	.w8(32'hbb8e327a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2457f4),
	.w1(32'hbb9fd694),
	.w2(32'hbc336232),
	.w3(32'hbb8cad10),
	.w4(32'hbb8fa704),
	.w5(32'hbbf279bf),
	.w6(32'h338b5ca0),
	.w7(32'h3a6ac9f8),
	.w8(32'hbb9840d8),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9a902),
	.w1(32'hbc1582e4),
	.w2(32'hbba9e414),
	.w3(32'hbbe4088d),
	.w4(32'h393dfbaf),
	.w5(32'h3b1850c1),
	.w6(32'hbb7420a2),
	.w7(32'hbb9fcf96),
	.w8(32'hbaa7065a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb202fc),
	.w1(32'hba9ac2c1),
	.w2(32'hbc1fbad4),
	.w3(32'h39f7b84d),
	.w4(32'h38e03c90),
	.w5(32'h3b5f31e6),
	.w6(32'h3b5add3b),
	.w7(32'hbbba2a56),
	.w8(32'hbbba2748),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60f113),
	.w1(32'hbbcb893f),
	.w2(32'hbb89062d),
	.w3(32'h3a90c1c5),
	.w4(32'hbab57ce6),
	.w5(32'hb8dbc589),
	.w6(32'hbad51e15),
	.w7(32'hbb200d77),
	.w8(32'hba48694a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49f4a7),
	.w1(32'hb9b4507f),
	.w2(32'hbb728dd3),
	.w3(32'hba2a3f47),
	.w4(32'hbb270a36),
	.w5(32'hbbbd46d2),
	.w6(32'hb9913cbe),
	.w7(32'hbabfbe92),
	.w8(32'hbbb2006a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba639969),
	.w1(32'h3c484521),
	.w2(32'hbc4b8a2d),
	.w3(32'h3be892b3),
	.w4(32'h3c14122b),
	.w5(32'hbc30e8b0),
	.w6(32'h3c06a3af),
	.w7(32'h3aa6cbd5),
	.w8(32'hbb839598),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf46562),
	.w1(32'hbb1a779d),
	.w2(32'hbc26b9d9),
	.w3(32'hbb426f6b),
	.w4(32'hbc1d1e0f),
	.w5(32'hbc13ef57),
	.w6(32'h3a572083),
	.w7(32'hbc313c0e),
	.w8(32'hbc4c8359),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b7e27),
	.w1(32'h3be4d4be),
	.w2(32'hbb3e3bec),
	.w3(32'h3bc34cc0),
	.w4(32'h3aa88dac),
	.w5(32'hbbc0eb23),
	.w6(32'h3b10e2c1),
	.w7(32'hbacab42f),
	.w8(32'hbc26be9c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4f677),
	.w1(32'hbad21cb8),
	.w2(32'h3a8173dd),
	.w3(32'hbb1b0b5c),
	.w4(32'h3b20152b),
	.w5(32'h3b2b7343),
	.w6(32'h3ae78698),
	.w7(32'hbbb13e63),
	.w8(32'hbabba551),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc501d8),
	.w1(32'hbae65fac),
	.w2(32'hbb0b9b95),
	.w3(32'hbb3dee33),
	.w4(32'hb8b8e9f1),
	.w5(32'hbb0a9d6c),
	.w6(32'hbb352ccc),
	.w7(32'hbba90d15),
	.w8(32'hbbb6163b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b6d3d),
	.w1(32'h3b4153d9),
	.w2(32'hbbaf3a5c),
	.w3(32'h3b3c2cc0),
	.w4(32'hbb346a35),
	.w5(32'hbbfe271f),
	.w6(32'h3acb70d6),
	.w7(32'hbb90376f),
	.w8(32'hbbd161b9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52c89),
	.w1(32'hba8293ff),
	.w2(32'hbb047475),
	.w3(32'hbc65af09),
	.w4(32'hbb78e689),
	.w5(32'h3c8ba5ab),
	.w6(32'hbb85baf6),
	.w7(32'hbb84a996),
	.w8(32'h3c86f892),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c904b08),
	.w1(32'h3bb74aee),
	.w2(32'h3c413729),
	.w3(32'h3c05b74f),
	.w4(32'h3c6f6c9f),
	.w5(32'h3ab60fb5),
	.w6(32'hbb7df43a),
	.w7(32'h3c4ea571),
	.w8(32'hbb13eea8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4250a2),
	.w1(32'h3b081582),
	.w2(32'hbb01bbda),
	.w3(32'h3b617e9f),
	.w4(32'h3b613c52),
	.w5(32'hb97d6de8),
	.w6(32'h3c228f34),
	.w7(32'hba36c3ba),
	.w8(32'hba848669),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398533fd),
	.w1(32'hba19fb53),
	.w2(32'hbb1e1184),
	.w3(32'h3943972a),
	.w4(32'hb8d7c892),
	.w5(32'hb9cbae85),
	.w6(32'hba82f660),
	.w7(32'hb97e3558),
	.w8(32'hbae4a5e7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d1f95),
	.w1(32'hbab3b7e2),
	.w2(32'hbaafe3a3),
	.w3(32'h3ab61863),
	.w4(32'hbb197db8),
	.w5(32'hbb39ec3e),
	.w6(32'h3885e4a0),
	.w7(32'h3a7cd246),
	.w8(32'hbb882f3e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90e077),
	.w1(32'hbaa3d75a),
	.w2(32'hba936bc8),
	.w3(32'hba081feb),
	.w4(32'hba68283a),
	.w5(32'hbab151be),
	.w6(32'h3aa211bf),
	.w7(32'h3ae6a720),
	.w8(32'hbb48912e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe8d1e),
	.w1(32'hba99efc1),
	.w2(32'hbab5dc03),
	.w3(32'hba394aa4),
	.w4(32'hb8fcf8f1),
	.w5(32'h39e94978),
	.w6(32'hbad33593),
	.w7(32'hbb100bfe),
	.w8(32'h3a18b77b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe8257),
	.w1(32'h3b2e4036),
	.w2(32'hbbc039c7),
	.w3(32'h3a0988a8),
	.w4(32'h39770869),
	.w5(32'hbbee5500),
	.w6(32'hbb0222e8),
	.w7(32'hb9ed79b0),
	.w8(32'hbbc74521),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5fd58),
	.w1(32'hbb9b2cd2),
	.w2(32'hbb7ff23e),
	.w3(32'hbb68fc10),
	.w4(32'hbb98ebd8),
	.w5(32'h3996aed9),
	.w6(32'hbb782c04),
	.w7(32'hbb483540),
	.w8(32'h3aee2950),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a938b31),
	.w1(32'hb89b142f),
	.w2(32'h3ac7546a),
	.w3(32'hb7ed5fb6),
	.w4(32'hbacd8052),
	.w5(32'hb9e2cee9),
	.w6(32'h3bbe845f),
	.w7(32'h3b11de91),
	.w8(32'hbab76894),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d7d784),
	.w1(32'hbb0a84a2),
	.w2(32'hbb52c474),
	.w3(32'h3ac6269b),
	.w4(32'hbb3640d5),
	.w5(32'h37afa529),
	.w6(32'h3aba06a7),
	.w7(32'hbb17ce26),
	.w8(32'hbacf9af7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae51bf4),
	.w1(32'h3a61ac73),
	.w2(32'h3a8aa427),
	.w3(32'hb9fd9ef9),
	.w4(32'hba96490c),
	.w5(32'h3a9a5711),
	.w6(32'h3a8905e4),
	.w7(32'hba0cf164),
	.w8(32'h3a684e87),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f3ee9d),
	.w1(32'hba339839),
	.w2(32'hbaf24c14),
	.w3(32'hb9cab284),
	.w4(32'h394cf46a),
	.w5(32'h39b03c75),
	.w6(32'h3a24f2e3),
	.w7(32'h39be4082),
	.w8(32'h3a890a64),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9146f73),
	.w1(32'hb616c10e),
	.w2(32'hb9b44371),
	.w3(32'h38f6394f),
	.w4(32'h3a7e0999),
	.w5(32'hba4e21d9),
	.w6(32'hbadd4c3b),
	.w7(32'hb83ecaec),
	.w8(32'hba43fac7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4da6d3),
	.w1(32'hb9c7e350),
	.w2(32'hbad7d8da),
	.w3(32'hbaf5e8ee),
	.w4(32'hbb1e3c1a),
	.w5(32'h3b231c5c),
	.w6(32'hba0c61fc),
	.w7(32'hbacbd4d1),
	.w8(32'h3a56b8d9),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac903ff),
	.w1(32'h3b3378d1),
	.w2(32'h3b116e52),
	.w3(32'h3aae056b),
	.w4(32'h3b6d5b6b),
	.w5(32'hba6d8ca2),
	.w6(32'h3a59e784),
	.w7(32'h3ad9038a),
	.w8(32'hbb106a12),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1d0c6),
	.w1(32'hbb228fea),
	.w2(32'hbb441267),
	.w3(32'hbaca8913),
	.w4(32'hbadda73e),
	.w5(32'hbb1ba9df),
	.w6(32'hbabdfbad),
	.w7(32'hbb1b3e21),
	.w8(32'hbba33ce0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57fe5a),
	.w1(32'hbb3e597e),
	.w2(32'hbb5b69c3),
	.w3(32'hba1b4384),
	.w4(32'hbb079313),
	.w5(32'hb9b5506a),
	.w6(32'h3a88f87b),
	.w7(32'hbaeb2006),
	.w8(32'hb9d74eff),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6bf16),
	.w1(32'hbb4b6c86),
	.w2(32'hbb5cde1e),
	.w3(32'h3a906fba),
	.w4(32'hbad3cce4),
	.w5(32'hba05d236),
	.w6(32'h3ac876a6),
	.w7(32'hbb0f4623),
	.w8(32'hbb50a7f6),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6695ca),
	.w1(32'h3a94b115),
	.w2(32'h39c97937),
	.w3(32'h3b174a31),
	.w4(32'h3a17fe3b),
	.w5(32'hba9ee0d9),
	.w6(32'h3ab0abbc),
	.w7(32'h3a7fdf4d),
	.w8(32'hba84b5f1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa55640),
	.w1(32'h39ebcfde),
	.w2(32'hba308243),
	.w3(32'hba719e84),
	.w4(32'hb92ecb3b),
	.w5(32'hba9ec1a3),
	.w6(32'hba966a16),
	.w7(32'hb90f28bf),
	.w8(32'hbaedecc4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0beb),
	.w1(32'hba601079),
	.w2(32'h390d1200),
	.w3(32'hb9297be4),
	.w4(32'h39b37412),
	.w5(32'hbb117c80),
	.w6(32'hbae6d86a),
	.w7(32'h37bbe333),
	.w8(32'h3942bb34),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6941d),
	.w1(32'h3a039d1e),
	.w2(32'hb95e19e0),
	.w3(32'hbb04597d),
	.w4(32'hb9e09ef1),
	.w5(32'h397a3de1),
	.w6(32'h3b047ca3),
	.w7(32'hbb082800),
	.w8(32'hba94b25f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba844581),
	.w1(32'hbb4238b6),
	.w2(32'hbb2988c7),
	.w3(32'h3926c2d4),
	.w4(32'hbb08a6f7),
	.w5(32'hbb99e7c1),
	.w6(32'hbb3c4dc5),
	.w7(32'hbae59859),
	.w8(32'hbb8dff7e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a8024),
	.w1(32'hbb948491),
	.w2(32'hbb83b019),
	.w3(32'hbb2be5e9),
	.w4(32'hbb289463),
	.w5(32'hbb103076),
	.w6(32'hbb641f0c),
	.w7(32'hbb214dee),
	.w8(32'hbae76552),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0241dc),
	.w1(32'h3a50bac5),
	.w2(32'h3856ea03),
	.w3(32'hbacedd00),
	.w4(32'hbab1f312),
	.w5(32'h3b16012c),
	.w6(32'hbb101473),
	.w7(32'hba8557dd),
	.w8(32'h3993f7f9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0e9f2),
	.w1(32'h3abc85ef),
	.w2(32'h3b16d999),
	.w3(32'h3a1df6b1),
	.w4(32'h3b583885),
	.w5(32'hba923af4),
	.w6(32'h3ab12d1b),
	.w7(32'h3b2f9f13),
	.w8(32'hbb33e64d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdf11e),
	.w1(32'h3b0805dd),
	.w2(32'h3a19954d),
	.w3(32'h3996d26b),
	.w4(32'hbace1e84),
	.w5(32'h3b0c8ae2),
	.w6(32'hba0a5c95),
	.w7(32'hbb83caef),
	.w8(32'h3aa1deb2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6fbd),
	.w1(32'h3a1f4cad),
	.w2(32'h3aebac05),
	.w3(32'h3b314197),
	.w4(32'h3b2d7421),
	.w5(32'hb68e4a68),
	.w6(32'h3bb27303),
	.w7(32'h3b4b1c30),
	.w8(32'hbb4e4dc2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72c0da8),
	.w1(32'h3a209565),
	.w2(32'hba94f40a),
	.w3(32'h399c6ece),
	.w4(32'hb911fdde),
	.w5(32'hbb291d38),
	.w6(32'hb9cacce5),
	.w7(32'hbb4909c3),
	.w8(32'hba8fb7c4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b7f3f),
	.w1(32'hbb71a956),
	.w2(32'hbb0b3a3a),
	.w3(32'hbac474d6),
	.w4(32'hbb036b89),
	.w5(32'h3a802517),
	.w6(32'hbb983a47),
	.w7(32'hbbc4ab31),
	.w8(32'hbb179a4c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84543bb),
	.w1(32'hba96366f),
	.w2(32'hb9a169a9),
	.w3(32'h39617910),
	.w4(32'h3918e8e9),
	.w5(32'hbaf673d1),
	.w6(32'h39bd6026),
	.w7(32'hba0d30f7),
	.w8(32'hbaf78c6d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb795acd),
	.w1(32'hbb88f91f),
	.w2(32'hba93739e),
	.w3(32'hbb8882c5),
	.w4(32'hba6a2ce6),
	.w5(32'h3a9c9822),
	.w6(32'hbb30ac45),
	.w7(32'hbaad2c50),
	.w8(32'hbae23eab),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule