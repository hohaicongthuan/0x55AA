module layer_8_featuremap_162(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b3ebd),
	.w1(32'h3c2037d4),
	.w2(32'h3b1e11ea),
	.w3(32'hbc0e1d56),
	.w4(32'hbb5d4a54),
	.w5(32'hbbc3a8f1),
	.w6(32'h3bd16587),
	.w7(32'h3b942c35),
	.w8(32'h3baa61c3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83bbd2),
	.w1(32'h3a8c2f7e),
	.w2(32'h3c065fd0),
	.w3(32'h3b98afad),
	.w4(32'h3adfa12e),
	.w5(32'h3bc5d428),
	.w6(32'h3b1c895f),
	.w7(32'h3b94d926),
	.w8(32'h3bae0a38),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23db30),
	.w1(32'hb9d59a3f),
	.w2(32'h3c00746c),
	.w3(32'h3c12a492),
	.w4(32'hb9b9e032),
	.w5(32'h3b321f1e),
	.w6(32'h3b4b62ae),
	.w7(32'h3bdc87e1),
	.w8(32'h3bbb1d8f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50cfea),
	.w1(32'hbb379862),
	.w2(32'h3abc8dfe),
	.w3(32'h3c2428e5),
	.w4(32'hbba13ff5),
	.w5(32'h3bd5ff88),
	.w6(32'hbb00bd46),
	.w7(32'h3a021ac1),
	.w8(32'h3c056b4b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c113530),
	.w1(32'hbbe4e395),
	.w2(32'hbbe4b79e),
	.w3(32'h3c30ca96),
	.w4(32'hbbf68b89),
	.w5(32'hbb83594a),
	.w6(32'hbb9dea7e),
	.w7(32'hbb9e6ddd),
	.w8(32'h3a1ba727),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf2fab),
	.w1(32'hbb665b18),
	.w2(32'h3bf8fd13),
	.w3(32'h3a8141e2),
	.w4(32'hbc010447),
	.w5(32'h3c1dd9ab),
	.w6(32'hbc07c138),
	.w7(32'h3b92c540),
	.w8(32'h3c66ee15),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83b9d6),
	.w1(32'hb9e9cc3a),
	.w2(32'hbba1798e),
	.w3(32'h3be38286),
	.w4(32'hbb27a48e),
	.w5(32'hbb33ae0f),
	.w6(32'hb9b260f6),
	.w7(32'hbb20c41f),
	.w8(32'hbae7660f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81fbbd),
	.w1(32'h3bcee95b),
	.w2(32'h3b34b8a1),
	.w3(32'h3abb48e1),
	.w4(32'hba57076d),
	.w5(32'hbbdaf789),
	.w6(32'h3bd4796d),
	.w7(32'hba8d0364),
	.w8(32'hbbe1b4ce),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc91c8a),
	.w1(32'h3b105281),
	.w2(32'hbbe832c7),
	.w3(32'hbbd3fcee),
	.w4(32'h3b5f722e),
	.w5(32'hbb6812dc),
	.w6(32'h3bf2164c),
	.w7(32'hbb4f57c1),
	.w8(32'h3b4bc9f9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc9233),
	.w1(32'hbb3032c0),
	.w2(32'h3aaab02f),
	.w3(32'h3b97f5b5),
	.w4(32'hbc27b87f),
	.w5(32'hbb1c7509),
	.w6(32'hbb1ab73a),
	.w7(32'hbaee6471),
	.w8(32'hb9388740),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c320b05),
	.w1(32'h3b561b4d),
	.w2(32'hbb81cb32),
	.w3(32'h3c026e3c),
	.w4(32'h3b717aac),
	.w5(32'hbc0d4d6b),
	.w6(32'hbb5a34e3),
	.w7(32'hba24ea6d),
	.w8(32'h3bba04d3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf81d6),
	.w1(32'hbb7ed611),
	.w2(32'hba5947cc),
	.w3(32'hbba6b77d),
	.w4(32'hbc06b2d0),
	.w5(32'hbbe4b426),
	.w6(32'hbacdb9f6),
	.w7(32'hbb113331),
	.w8(32'h399e5f2c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fae2d),
	.w1(32'hbc0f2a78),
	.w2(32'hbb5f4f6d),
	.w3(32'h3b046311),
	.w4(32'hbbbac194),
	.w5(32'hba9f65d8),
	.w6(32'hbbb5649f),
	.w7(32'hbaf260b7),
	.w8(32'h3be44768),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3efdd),
	.w1(32'h3bb584ca),
	.w2(32'h3b9450f1),
	.w3(32'h3c525e78),
	.w4(32'hb8efa2e8),
	.w5(32'h3b2dfa18),
	.w6(32'h3b53324e),
	.w7(32'h3be2dd53),
	.w8(32'h3b9fadfb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01958f),
	.w1(32'h3bbb2790),
	.w2(32'hbb7cea11),
	.w3(32'h3c0fe32f),
	.w4(32'h3b534960),
	.w5(32'hbb34a4f3),
	.w6(32'h3b971009),
	.w7(32'hbb4386ff),
	.w8(32'hbbd0ef09),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fda43),
	.w1(32'h3adb8b04),
	.w2(32'h3c1af025),
	.w3(32'hbb542b4a),
	.w4(32'h3b7486d8),
	.w5(32'h3b3829f1),
	.w6(32'hb9b17fb5),
	.w7(32'h3c08cc0d),
	.w8(32'h3cc78963),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc03a52),
	.w1(32'h3c3978a4),
	.w2(32'h3bab57a2),
	.w3(32'h3c910335),
	.w4(32'h3b9bb350),
	.w5(32'h3c7250ed),
	.w6(32'h3b23e6a9),
	.w7(32'h3ae7f3ed),
	.w8(32'h3be21504),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c468b91),
	.w1(32'h3b2152b7),
	.w2(32'h3b98cec3),
	.w3(32'h3c4eb546),
	.w4(32'hb94867f8),
	.w5(32'h3bdfb58e),
	.w6(32'hbadd2fef),
	.w7(32'hbbc58946),
	.w8(32'h3c3f5f4a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c892e25),
	.w1(32'hba853cc3),
	.w2(32'h3c0812d7),
	.w3(32'h3c2b9ff9),
	.w4(32'hbc337457),
	.w5(32'hbaa2b617),
	.w6(32'hbc99600e),
	.w7(32'hbc51e00e),
	.w8(32'h3b438cf6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca82e29),
	.w1(32'h3b636c2d),
	.w2(32'h3b00d5aa),
	.w3(32'h3c760ed1),
	.w4(32'hbb391ebc),
	.w5(32'hbb9b1a81),
	.w6(32'h3c077670),
	.w7(32'hba784790),
	.w8(32'hba904256),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e3a8b),
	.w1(32'h3c660b15),
	.w2(32'h3bcdbd96),
	.w3(32'hbaec6926),
	.w4(32'h3ba9254d),
	.w5(32'h3c09aca2),
	.w6(32'h3a3e5a61),
	.w7(32'hbc0ff1fc),
	.w8(32'hbb5e7e90),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95d5d8),
	.w1(32'h3b7b36d5),
	.w2(32'h3aaf3ca7),
	.w3(32'h3baf6631),
	.w4(32'h3b945518),
	.w5(32'h3b81faf6),
	.w6(32'hba64e1cd),
	.w7(32'h3a1e1ee2),
	.w8(32'h3ab629e3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd8cab),
	.w1(32'h3b99d92e),
	.w2(32'hbaf19d7c),
	.w3(32'h3bba1683),
	.w4(32'hbc2070be),
	.w5(32'hbb7feae6),
	.w6(32'hbbbac924),
	.w7(32'hbc3fd832),
	.w8(32'hbbb0e486),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13932e),
	.w1(32'h3ba12390),
	.w2(32'hbbcb0e4d),
	.w3(32'h3c5da093),
	.w4(32'h3c1ef058),
	.w5(32'hba44590c),
	.w6(32'h3b1d1bbe),
	.w7(32'hbb1e7640),
	.w8(32'h3a260a3f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb228dd2),
	.w1(32'hbbc2972d),
	.w2(32'h3b9d9a8e),
	.w3(32'h3aded379),
	.w4(32'hbb47e1f4),
	.w5(32'h38b76bc9),
	.w6(32'hbb83748f),
	.w7(32'hbad41331),
	.w8(32'h3b80f292),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99e0d8),
	.w1(32'h3c1d90e3),
	.w2(32'h3c028f94),
	.w3(32'h3c93cd5c),
	.w4(32'hbb513046),
	.w5(32'hbb9eb85b),
	.w6(32'h3c1e2652),
	.w7(32'h3b9628a9),
	.w8(32'hba4f69d7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b2e9),
	.w1(32'hba637c40),
	.w2(32'h3bf7d827),
	.w3(32'h3babeb6d),
	.w4(32'hba96c1bc),
	.w5(32'h38d032a1),
	.w6(32'hbab27a02),
	.w7(32'h3b9cb0fc),
	.w8(32'h3c1f8980),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d530b26),
	.w1(32'h3ca116b7),
	.w2(32'h3c121f19),
	.w3(32'h3cb96909),
	.w4(32'hbb4ab861),
	.w5(32'h3a622220),
	.w6(32'hbbd5a976),
	.w7(32'hbcc3d459),
	.w8(32'hbcbb4686),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa798b5),
	.w1(32'h3b325479),
	.w2(32'hbb9e6ae4),
	.w3(32'h398f8407),
	.w4(32'hba067f6b),
	.w5(32'hbbfd4265),
	.w6(32'h3b0de95d),
	.w7(32'hbbb7783b),
	.w8(32'h3b3da18b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc23f4a),
	.w1(32'hbb433324),
	.w2(32'hbc22e4a0),
	.w3(32'h3b7caa63),
	.w4(32'hbc3a29ab),
	.w5(32'hbc8e3304),
	.w6(32'hbb4119d9),
	.w7(32'hbc19c21c),
	.w8(32'h3c1c7026),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c163c4f),
	.w1(32'h3b6f3d8b),
	.w2(32'h3ab7d8b5),
	.w3(32'h3acb479b),
	.w4(32'h390ec77c),
	.w5(32'hba11849f),
	.w6(32'h3b86640e),
	.w7(32'h3a1f2141),
	.w8(32'h3b5b9965),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf63a8f),
	.w1(32'h3c1865d3),
	.w2(32'h3b492034),
	.w3(32'h3b85481c),
	.w4(32'h3c2c6471),
	.w5(32'h3ae2cf7d),
	.w6(32'h3c329fdf),
	.w7(32'h383c1825),
	.w8(32'hbc1e264e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d3601),
	.w1(32'h3be33c3f),
	.w2(32'h3bf0eda5),
	.w3(32'hbb60df5d),
	.w4(32'h3b6a810b),
	.w5(32'h3a577834),
	.w6(32'h3b81a1e0),
	.w7(32'h3b224d83),
	.w8(32'h3b7d3fcc),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc51d19),
	.w1(32'h3b350bb0),
	.w2(32'h395adcd6),
	.w3(32'h3bd175af),
	.w4(32'h3aed7100),
	.w5(32'h3b00e1af),
	.w6(32'h3a6b25db),
	.w7(32'hb96c8d39),
	.w8(32'hbb3cbda7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb883f2),
	.w1(32'hb9a15760),
	.w2(32'hbb6007ea),
	.w3(32'hbb41d4b4),
	.w4(32'hbb1a1049),
	.w5(32'hbb9738c7),
	.w6(32'h3b3bd1ed),
	.w7(32'hbba40e94),
	.w8(32'hbaec1e62),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae98cdd),
	.w1(32'h3b81fa27),
	.w2(32'hba44caa0),
	.w3(32'h3ada3e39),
	.w4(32'h3b26b199),
	.w5(32'hbbda483c),
	.w6(32'h3af422e1),
	.w7(32'hbb48fca6),
	.w8(32'hbac9dd48),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb409bbd),
	.w1(32'hbac54fb8),
	.w2(32'h3ac7f9b4),
	.w3(32'hbb231892),
	.w4(32'hbb735fb2),
	.w5(32'h3a1f3e8a),
	.w6(32'hb9c6bf56),
	.w7(32'hba936775),
	.w8(32'hbad7327a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81d290),
	.w1(32'h3bb3a69b),
	.w2(32'hbbb87447),
	.w3(32'h3b99689a),
	.w4(32'h3b9bc9da),
	.w5(32'hbb8d68ac),
	.w6(32'h3b02e691),
	.w7(32'hbbd05ae9),
	.w8(32'hbc15eda4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdfe3a),
	.w1(32'h3b847a75),
	.w2(32'h3be31131),
	.w3(32'hbbcd24a6),
	.w4(32'hbb391f0b),
	.w5(32'h3beb9ff2),
	.w6(32'h3985f527),
	.w7(32'h3b5dc9dd),
	.w8(32'hbb74fd90),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b850815),
	.w1(32'h3b3eac51),
	.w2(32'hbbd9828b),
	.w3(32'h3b860f59),
	.w4(32'h3bd9f889),
	.w5(32'h3aa9a714),
	.w6(32'hbb51cbc5),
	.w7(32'hbbd01591),
	.w8(32'h3ad1924f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d4c76),
	.w1(32'h39e6f3aa),
	.w2(32'hbacbf629),
	.w3(32'h3c258526),
	.w4(32'hbbb3d45d),
	.w5(32'hbc1870d5),
	.w6(32'h3abe84c9),
	.w7(32'hbc5632e1),
	.w8(32'hbc08f848),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810ea5),
	.w1(32'hbb0779b0),
	.w2(32'h3bff8ee2),
	.w3(32'hbbc1a4f7),
	.w4(32'hbaa6a6f2),
	.w5(32'h3c464c89),
	.w6(32'hba796683),
	.w7(32'h3b1817db),
	.w8(32'h3b211475),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf511d),
	.w1(32'hbbe53078),
	.w2(32'h3aa99c7c),
	.w3(32'h3bdd6e2d),
	.w4(32'hbc0bdb22),
	.w5(32'h39a21408),
	.w6(32'hbb6dfa41),
	.w7(32'hbb91fcde),
	.w8(32'h3b9ec841),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4c050),
	.w1(32'h3ad35cbe),
	.w2(32'h3c336fd3),
	.w3(32'h3b637dc5),
	.w4(32'hbb13cd2d),
	.w5(32'h3bb57b63),
	.w6(32'h3a72fe60),
	.w7(32'h3bbd05bc),
	.w8(32'h3bb5c422),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca755a8),
	.w1(32'h3c474d2a),
	.w2(32'hb962bc0f),
	.w3(32'h3c10ba36),
	.w4(32'h3c207d39),
	.w5(32'h3ab306a5),
	.w6(32'h3c273391),
	.w7(32'hbb71fdcc),
	.w8(32'hbbeba976),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb281c3e),
	.w1(32'h3b666b4b),
	.w2(32'h3b54cd8e),
	.w3(32'h3ba52715),
	.w4(32'h3911c03e),
	.w5(32'h3b2c462f),
	.w6(32'h3b20c800),
	.w7(32'hb9fe53e8),
	.w8(32'h3aeebe55),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38a7a7),
	.w1(32'hbb3ed776),
	.w2(32'hbb532e08),
	.w3(32'h3b8b7135),
	.w4(32'hbaafe803),
	.w5(32'hb84f9890),
	.w6(32'h3add3fff),
	.w7(32'hb9ffaf4a),
	.w8(32'hba1e22ba),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e8c78),
	.w1(32'h3a1f38db),
	.w2(32'hba7ef7ae),
	.w3(32'h3bc950d0),
	.w4(32'hba74801c),
	.w5(32'hba9695c1),
	.w6(32'hbbc7376d),
	.w7(32'hbbba6827),
	.w8(32'hba85accd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde3887),
	.w1(32'h3aab2cf2),
	.w2(32'h3bf59a1a),
	.w3(32'h3c040a6d),
	.w4(32'h3b7a1cdc),
	.w5(32'hba92c223),
	.w6(32'h3a225acd),
	.w7(32'h3bb89400),
	.w8(32'hbba8f425),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd936ad),
	.w1(32'h3bb2645a),
	.w2(32'h3caeb040),
	.w3(32'h3c528ad4),
	.w4(32'h3a0052e5),
	.w5(32'h3be1b3bd),
	.w6(32'h384fc50e),
	.w7(32'h3beb15f5),
	.w8(32'h3b7bb62f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb6991d),
	.w1(32'hbb741e91),
	.w2(32'hbba32f44),
	.w3(32'h3c2da525),
	.w4(32'hbb97fe52),
	.w5(32'hbbeaf58c),
	.w6(32'hb973c0dd),
	.w7(32'hbba50334),
	.w8(32'hbbcb17e4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d8ce3),
	.w1(32'hbb35b7ce),
	.w2(32'h3b58b506),
	.w3(32'h3c39f572),
	.w4(32'h3a92fe0b),
	.w5(32'h3b8157fa),
	.w6(32'h3b94668c),
	.w7(32'hbb9c9d0d),
	.w8(32'h39b1e6d6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c208346),
	.w1(32'hbb437a9e),
	.w2(32'hbb8da21b),
	.w3(32'h3c2ada3c),
	.w4(32'hbb8a7451),
	.w5(32'hbbe620ab),
	.w6(32'hbafdd3e4),
	.w7(32'hbbeed8cd),
	.w8(32'hbb778ae9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5964e),
	.w1(32'h395b65c2),
	.w2(32'h377076ee),
	.w3(32'hbab261a9),
	.w4(32'hbc03a41c),
	.w5(32'hbbfc0a19),
	.w6(32'hbc2803da),
	.w7(32'hbc0b593c),
	.w8(32'h3b780688),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d924f),
	.w1(32'hbbae5e6c),
	.w2(32'hbae241ff),
	.w3(32'h3c0881e7),
	.w4(32'hbad5f790),
	.w5(32'hbbb734a4),
	.w6(32'h3b82cf51),
	.w7(32'hbba7fe0f),
	.w8(32'h3c0ec334),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b6c29),
	.w1(32'h3c394022),
	.w2(32'h3c9ce497),
	.w3(32'h3c3ce31e),
	.w4(32'hba50d6d0),
	.w5(32'h3b866b49),
	.w6(32'hbbf6567c),
	.w7(32'hbc39015a),
	.w8(32'h3b560b53),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c510cd6),
	.w1(32'h3af51996),
	.w2(32'h3bfe0eaa),
	.w3(32'hbb1e7f45),
	.w4(32'hbbd71b0d),
	.w5(32'hbb425aae),
	.w6(32'hb915dede),
	.w7(32'h3b84b44c),
	.w8(32'hbb9a8f8f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15e875),
	.w1(32'hbbbf0d74),
	.w2(32'hbb94d16f),
	.w3(32'h3b48a355),
	.w4(32'hbc288db9),
	.w5(32'hbc0a22d1),
	.w6(32'hbb67942e),
	.w7(32'hbc29917c),
	.w8(32'hbbabb30f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bfb44),
	.w1(32'h3baa1486),
	.w2(32'h3c04aebf),
	.w3(32'hba952251),
	.w4(32'h3ad7d361),
	.w5(32'h3bc21a54),
	.w6(32'h3b01917a),
	.w7(32'h3b8c522f),
	.w8(32'h3b671606),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34ea6a),
	.w1(32'h3c450407),
	.w2(32'h3ba3ebc8),
	.w3(32'h3be4f977),
	.w4(32'h3c28ca66),
	.w5(32'h3b452fad),
	.w6(32'h3be4291e),
	.w7(32'h3b386557),
	.w8(32'h386b1bb8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39980e),
	.w1(32'hbbbd62b7),
	.w2(32'h3c0e84ab),
	.w3(32'h3b8d4419),
	.w4(32'hbc14e152),
	.w5(32'hbbb406c4),
	.w6(32'hba9c61a7),
	.w7(32'h3bfe0e45),
	.w8(32'h3be333e1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c233cfb),
	.w1(32'h3b6d5f01),
	.w2(32'hbbb030e5),
	.w3(32'h3b90b6b4),
	.w4(32'h3bb14faf),
	.w5(32'hbb9baa50),
	.w6(32'h3b7e5529),
	.w7(32'hbb91989e),
	.w8(32'hbad4be8e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c257ac5),
	.w1(32'h3c87f7e6),
	.w2(32'hbb64965f),
	.w3(32'h3c3f94d3),
	.w4(32'h3bf2f9e3),
	.w5(32'hbc32a6cb),
	.w6(32'h3c3598d0),
	.w7(32'hbc4deae3),
	.w8(32'hbc3b7dc6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50388b),
	.w1(32'hbb27a563),
	.w2(32'h35581bb8),
	.w3(32'hbc786b2e),
	.w4(32'hbb07fc66),
	.w5(32'hbb3a4382),
	.w6(32'hba8f83d8),
	.w7(32'hbaa68850),
	.w8(32'hbae09456),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d057e),
	.w1(32'h3bcd51cf),
	.w2(32'h3b71b61d),
	.w3(32'hbb1fe159),
	.w4(32'h3ba46c3b),
	.w5(32'h3b09cad1),
	.w6(32'h3b801a68),
	.w7(32'h3a7f443f),
	.w8(32'hbb17bb49),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc3374),
	.w1(32'h3b3ca9dc),
	.w2(32'h3b0f6381),
	.w3(32'h3a31f0b2),
	.w4(32'hbaf6ef6e),
	.w5(32'hbb9052ad),
	.w6(32'hbad4c24f),
	.w7(32'hbb391269),
	.w8(32'hbb858b72),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f6f48),
	.w1(32'h3bd1a617),
	.w2(32'h3c206003),
	.w3(32'h3b1b4344),
	.w4(32'h3bcfca1d),
	.w5(32'h3ad72625),
	.w6(32'hbbb6b991),
	.w7(32'hbb00b3c0),
	.w8(32'h3c19b961),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4185),
	.w1(32'h3b7457f1),
	.w2(32'hbaaac389),
	.w3(32'h3bd3b885),
	.w4(32'hbb0c3bb6),
	.w5(32'hbb3958ba),
	.w6(32'h3b5c0a68),
	.w7(32'hba4b023d),
	.w8(32'h39231a6d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a419c4d),
	.w1(32'h3c1b2b4c),
	.w2(32'h3c02f7a0),
	.w3(32'h3b9ecf77),
	.w4(32'h3c16a1ff),
	.w5(32'h3bc4302d),
	.w6(32'h3b29b1e8),
	.w7(32'hb9791efa),
	.w8(32'hbbcb0348),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf673c3),
	.w1(32'h3c465871),
	.w2(32'h3c038a88),
	.w3(32'h3c0c4799),
	.w4(32'hbae441cd),
	.w5(32'hbb7bb8ca),
	.w6(32'hbb6bcddc),
	.w7(32'hbc0ec23b),
	.w8(32'h3b012b9b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82992a),
	.w1(32'h3b02de1a),
	.w2(32'hbbb5ef75),
	.w3(32'h3c21a15c),
	.w4(32'h3bb2a987),
	.w5(32'hbb3083df),
	.w6(32'h3b9cd671),
	.w7(32'hbb703826),
	.w8(32'h3bb82d77),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25ffd1),
	.w1(32'h3b47a8e6),
	.w2(32'h3a356f13),
	.w3(32'h3bc5ecf2),
	.w4(32'h3b2984c2),
	.w5(32'hbb5e4caf),
	.w6(32'h3bf13e9e),
	.w7(32'h3b53a59b),
	.w8(32'hbaac7aab),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc2483),
	.w1(32'h3875e630),
	.w2(32'h3ba0d8f0),
	.w3(32'h3a8d8d35),
	.w4(32'hbb85c446),
	.w5(32'hbb54bdb0),
	.w6(32'h3b6bd2a3),
	.w7(32'h3b05f9a2),
	.w8(32'h3bd57e72),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba1055),
	.w1(32'hbbedbfa7),
	.w2(32'hbb1399d2),
	.w3(32'h3b6d46a1),
	.w4(32'hbc2c8829),
	.w5(32'hbba42b69),
	.w6(32'hbad2f2a5),
	.w7(32'hba7e0ea1),
	.w8(32'h3b9a6c1e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae83a60),
	.w1(32'hbc18b1de),
	.w2(32'hbaacea40),
	.w3(32'h3ba1ad72),
	.w4(32'hbbecf7d8),
	.w5(32'h3bbff25a),
	.w6(32'hbc18bc5a),
	.w7(32'hbba32f75),
	.w8(32'h3aef595b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51fdd4),
	.w1(32'hbb27885b),
	.w2(32'hbb1ef27c),
	.w3(32'h3c9537e6),
	.w4(32'hbc21d71f),
	.w5(32'hba937bde),
	.w6(32'hbbac66e7),
	.w7(32'hbb8f845f),
	.w8(32'h3b090564),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adae71d),
	.w1(32'hbba74404),
	.w2(32'h3b8d555d),
	.w3(32'h3c14bdc1),
	.w4(32'hbc0124cf),
	.w5(32'hba8bea8c),
	.w6(32'hbb99d9cd),
	.w7(32'h39d339c5),
	.w8(32'h3b610808),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c185d30),
	.w1(32'hbb10920c),
	.w2(32'h3bf666fa),
	.w3(32'h3bf3eae4),
	.w4(32'hbc054f5a),
	.w5(32'h3b54a353),
	.w6(32'hbb8dd3f8),
	.w7(32'hbaf66efa),
	.w8(32'h3b92ce95),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95e89d),
	.w1(32'hbbcc3486),
	.w2(32'h38d345ea),
	.w3(32'h3c829370),
	.w4(32'hbbed486e),
	.w5(32'hbb3fd8c5),
	.w6(32'h3914b8e1),
	.w7(32'hbacaf222),
	.w8(32'h3c40b778),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21fc6c),
	.w1(32'h3c018b75),
	.w2(32'h3b86f3a8),
	.w3(32'h3ba15897),
	.w4(32'h38ae6e9f),
	.w5(32'hbb98e8fd),
	.w6(32'h3b69aef5),
	.w7(32'hbb34e9fd),
	.w8(32'h3b004694),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd6a33),
	.w1(32'h3b8c54fd),
	.w2(32'h3c268d73),
	.w3(32'hbbbd311e),
	.w4(32'h3b766e4d),
	.w5(32'h3bf12655),
	.w6(32'h3b51c0b1),
	.w7(32'h3bef3dcc),
	.w8(32'hb98ae99c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c152e5d),
	.w1(32'h3c0e984e),
	.w2(32'h3c28563b),
	.w3(32'h3c3036ac),
	.w4(32'h3b519cfc),
	.w5(32'h3c15ec13),
	.w6(32'h3b86884a),
	.w7(32'h3ba3258a),
	.w8(32'hbb0e6a7f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d7d38),
	.w1(32'h3c091df7),
	.w2(32'h3b1d782e),
	.w3(32'h3c2986c5),
	.w4(32'h3b8a99ff),
	.w5(32'h3abcb823),
	.w6(32'hbae5c9ab),
	.w7(32'hbc0f5259),
	.w8(32'hba95a98e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd3d73b),
	.w1(32'h3aa6b107),
	.w2(32'h3b6521ff),
	.w3(32'h3cc19a27),
	.w4(32'h3bd01830),
	.w5(32'hb98cee2b),
	.w6(32'h3c368b66),
	.w7(32'hba92bd8b),
	.w8(32'h3b459490),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f5316),
	.w1(32'h3acb3284),
	.w2(32'h3bdc4ced),
	.w3(32'h3c86cff5),
	.w4(32'hbb857628),
	.w5(32'h3b5caa88),
	.w6(32'h3baf46c0),
	.w7(32'hbbaa679e),
	.w8(32'hbb502fe8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c170acf),
	.w1(32'h3b36cdea),
	.w2(32'h3bcfa500),
	.w3(32'h3c4ad291),
	.w4(32'h3ba0e094),
	.w5(32'h3afdf599),
	.w6(32'hba8122b4),
	.w7(32'hbae3751b),
	.w8(32'h3bf6c89d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0b490),
	.w1(32'hba8bb2ca),
	.w2(32'h398ecbe4),
	.w3(32'hba0d3864),
	.w4(32'h3abceb6f),
	.w5(32'h3a9d44e0),
	.w6(32'hbaba34d9),
	.w7(32'hb916d361),
	.w8(32'h3bf65e4d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9fd42),
	.w1(32'h3bb8a0b5),
	.w2(32'h3ba881fb),
	.w3(32'h3b0baa0f),
	.w4(32'h3bc64b19),
	.w5(32'h3ae6c398),
	.w6(32'h3bc98997),
	.w7(32'h3abb76b0),
	.w8(32'h3b4d6a28),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51e860),
	.w1(32'hbb7f5518),
	.w2(32'hbacfe11d),
	.w3(32'h3c026d67),
	.w4(32'hbb95c568),
	.w5(32'hba754f92),
	.w6(32'hbb9675f6),
	.w7(32'hba9f8b8b),
	.w8(32'h3bb6c642),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b627d27),
	.w1(32'hbb9fed8d),
	.w2(32'h3bf2045b),
	.w3(32'h3b84c1ed),
	.w4(32'hbbd12925),
	.w5(32'hbba32099),
	.w6(32'h3a93b41a),
	.w7(32'h3b2794c0),
	.w8(32'hba572aa7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18c91b),
	.w1(32'hbb5ce6de),
	.w2(32'hbb32e9aa),
	.w3(32'h3aa4032c),
	.w4(32'hbbd10c60),
	.w5(32'hbb779869),
	.w6(32'h3c307464),
	.w7(32'h3b3f8196),
	.w8(32'h3ae6d337),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89bc251),
	.w1(32'h3ab0b1a1),
	.w2(32'h39c63554),
	.w3(32'hbb3847bc),
	.w4(32'h3ba2b98f),
	.w5(32'h39c918a2),
	.w6(32'hba3ae0bd),
	.w7(32'hba8bd6eb),
	.w8(32'hbb37abd6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba978c37),
	.w1(32'h3b2022e2),
	.w2(32'h3bc3c715),
	.w3(32'hbbb1fee4),
	.w4(32'h3adcd252),
	.w5(32'h3b5047f5),
	.w6(32'h3b9107dc),
	.w7(32'h3b7e9111),
	.w8(32'h3a7b597b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f77a4),
	.w1(32'h383157a0),
	.w2(32'h3bff2495),
	.w3(32'h3b442000),
	.w4(32'h3a4fd61d),
	.w5(32'h3bb1b076),
	.w6(32'h3acede6f),
	.w7(32'h3b38cb03),
	.w8(32'h3b57228a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb319c),
	.w1(32'hbc141f14),
	.w2(32'hbbe8c77d),
	.w3(32'h3bf5a191),
	.w4(32'hbb9f27ba),
	.w5(32'hbc2edc5a),
	.w6(32'hbb043148),
	.w7(32'hbba3ef75),
	.w8(32'h3c0cda88),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c809d3e),
	.w1(32'hbb0ad7f2),
	.w2(32'h3b86d740),
	.w3(32'h3cac8ba9),
	.w4(32'hbbd4d60f),
	.w5(32'hbae5f71a),
	.w6(32'hbabaf0f9),
	.w7(32'hbac5138e),
	.w8(32'h399fc7c0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c261004),
	.w1(32'hbbc24a8d),
	.w2(32'hbb421f61),
	.w3(32'h3b583993),
	.w4(32'hbb5b029e),
	.w5(32'hbae4f4cd),
	.w6(32'h3bb0148d),
	.w7(32'hba6eb651),
	.w8(32'hbb31cb86),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe442c),
	.w1(32'h3af94e95),
	.w2(32'h3c82e2e5),
	.w3(32'h3c354b3a),
	.w4(32'hbacce506),
	.w5(32'h3c1b3170),
	.w6(32'hbb1945a2),
	.w7(32'h3c08cdaa),
	.w8(32'h3c286570),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2de19b),
	.w1(32'h3a0ef1bb),
	.w2(32'h3c1d961b),
	.w3(32'h3c31cc61),
	.w4(32'h3a9ee6a0),
	.w5(32'h3c2628f0),
	.w6(32'h39175c68),
	.w7(32'h3c06e0ca),
	.w8(32'h3c3da55a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1acf1),
	.w1(32'hbc32506c),
	.w2(32'h3ac25d71),
	.w3(32'h3c0c8aec),
	.w4(32'hbc0d4725),
	.w5(32'hbba8703e),
	.w6(32'hbba8452c),
	.w7(32'h3ac6b064),
	.w8(32'h3b8b18dd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025702),
	.w1(32'hbba68bda),
	.w2(32'hbafd4c75),
	.w3(32'h3a4f5e9a),
	.w4(32'h3ae49e48),
	.w5(32'hbaf8024d),
	.w6(32'hbc12dba1),
	.w7(32'hbbad6c3d),
	.w8(32'hb83646de),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2599c),
	.w1(32'hba1a4d94),
	.w2(32'h3aed59f6),
	.w3(32'hbc194de8),
	.w4(32'hbaf1ff66),
	.w5(32'h3ac8f746),
	.w6(32'h3af7b9ee),
	.w7(32'h3b704d91),
	.w8(32'hbbe9e820),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1154e5),
	.w1(32'hbbd2d8cd),
	.w2(32'hbb35676c),
	.w3(32'hbb8db69f),
	.w4(32'h3b651d78),
	.w5(32'hba98a4d3),
	.w6(32'h3bdffe4d),
	.w7(32'hbb2a30b3),
	.w8(32'hbb6f7e66),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd90322),
	.w1(32'h3b9b9f4e),
	.w2(32'h3adb722a),
	.w3(32'h399ebe32),
	.w4(32'hbb621e37),
	.w5(32'hba76bed2),
	.w6(32'h3b839c2b),
	.w7(32'h3c3530c0),
	.w8(32'h3bcb2768),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38547e8f),
	.w1(32'h3a46ab9a),
	.w2(32'h3ba8891f),
	.w3(32'h3b5b8e6b),
	.w4(32'hbaee77da),
	.w5(32'h3bf38be9),
	.w6(32'h3b14ed86),
	.w7(32'h3bdc4c2f),
	.w8(32'h3c0f8eba),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9fce6f),
	.w1(32'h3bef4f6c),
	.w2(32'h3a9d13b5),
	.w3(32'h3c7e6df4),
	.w4(32'h3b4f7e96),
	.w5(32'hbb2996d7),
	.w6(32'h3b85fde3),
	.w7(32'hbbba8b8b),
	.w8(32'hbb4c0158),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac805ea),
	.w1(32'hbbbbc8db),
	.w2(32'h3a6b3a88),
	.w3(32'hbab6e9c5),
	.w4(32'hba82a71c),
	.w5(32'h3b69635f),
	.w6(32'hbb82eab0),
	.w7(32'h3b8ef88a),
	.w8(32'h3c2d8f5f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c660807),
	.w1(32'hbbb6afb1),
	.w2(32'h3ba447f7),
	.w3(32'h3c64a89e),
	.w4(32'hbc3865a6),
	.w5(32'hbac610d3),
	.w6(32'h39122dbd),
	.w7(32'h37c0b048),
	.w8(32'h3bf9c2ab),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a656c),
	.w1(32'hbb81d328),
	.w2(32'hbc900f29),
	.w3(32'h3bbcda2a),
	.w4(32'hbb78f348),
	.w5(32'hbc5ed11c),
	.w6(32'h39f1917a),
	.w7(32'hbc145ab0),
	.w8(32'hbbe17ddd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63843f),
	.w1(32'h3b313a8c),
	.w2(32'h38e037fd),
	.w3(32'hbc7db4a5),
	.w4(32'h3ba9bcdf),
	.w5(32'h3a561897),
	.w6(32'h3b55093b),
	.w7(32'h3ade6d3f),
	.w8(32'h3ab579fd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd35f53),
	.w1(32'h3b84a86f),
	.w2(32'h3b30be53),
	.w3(32'h3b6c47b6),
	.w4(32'hbb1223f1),
	.w5(32'hba2538d0),
	.w6(32'h3bff60a5),
	.w7(32'h3ad2898a),
	.w8(32'h3bfd68e2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57215b),
	.w1(32'h3b1a7859),
	.w2(32'h3b2d0245),
	.w3(32'h3ad78ac4),
	.w4(32'h3a420402),
	.w5(32'h3b2efd43),
	.w6(32'h3bf34bf0),
	.w7(32'h3a6b1d80),
	.w8(32'h3a8ce3ae),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e2123),
	.w1(32'h3c132002),
	.w2(32'h3c0fee87),
	.w3(32'h3b8671e5),
	.w4(32'h3926f925),
	.w5(32'h3b832ce8),
	.w6(32'h3bd813a1),
	.w7(32'h3b910d4b),
	.w8(32'h39a1bef9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bf276),
	.w1(32'hbbb03c90),
	.w2(32'hbb5e8b25),
	.w3(32'h3a592114),
	.w4(32'hbb3da94d),
	.w5(32'h3ab3049d),
	.w6(32'hbad073bf),
	.w7(32'hbac2375d),
	.w8(32'h39fe8c42),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f6a60),
	.w1(32'hba1533aa),
	.w2(32'hbab690f7),
	.w3(32'h3c73464e),
	.w4(32'hbb9a6800),
	.w5(32'hba4c8326),
	.w6(32'hbab71976),
	.w7(32'hbb807f7c),
	.w8(32'h3a644f8f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8e587),
	.w1(32'h3b1c5b33),
	.w2(32'h3b26d24f),
	.w3(32'hba11128e),
	.w4(32'h3b38cfd8),
	.w5(32'h3ae30fca),
	.w6(32'h39293ffc),
	.w7(32'hba6b550c),
	.w8(32'hb5d9a282),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b982d49),
	.w1(32'hb9720147),
	.w2(32'hbb37e8db),
	.w3(32'h3b3407c9),
	.w4(32'hbc01cf4f),
	.w5(32'hbc3923f6),
	.w6(32'h3a5fde41),
	.w7(32'hbb327327),
	.w8(32'h3c01267a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f868d),
	.w1(32'h3b22df82),
	.w2(32'h3bbee5b4),
	.w3(32'h3b80c185),
	.w4(32'h3b45f210),
	.w5(32'h3b0113b8),
	.w6(32'h3b319e97),
	.w7(32'h3ab1f6e7),
	.w8(32'h3b9e88ac),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cf6f9),
	.w1(32'hbb21e71e),
	.w2(32'h3bd45860),
	.w3(32'h3b22b63c),
	.w4(32'hba9d81a5),
	.w5(32'h3b85600a),
	.w6(32'h3b79863d),
	.w7(32'h3be880b9),
	.w8(32'h3bef6965),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c714e78),
	.w1(32'hbb75414b),
	.w2(32'hb910729c),
	.w3(32'h3c1e94e7),
	.w4(32'hbb5f71d2),
	.w5(32'h3a371b0f),
	.w6(32'hbb4352bf),
	.w7(32'hbb10f75a),
	.w8(32'h3a5a7d85),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b92c9),
	.w1(32'h3bad7223),
	.w2(32'h3bf82c96),
	.w3(32'h3c145b17),
	.w4(32'h3c0e7da0),
	.w5(32'hb9a719d7),
	.w6(32'h3c32eaf7),
	.w7(32'hbb09e8a4),
	.w8(32'hbb021352),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fc8a9),
	.w1(32'h3a34c6d6),
	.w2(32'h3b1fa934),
	.w3(32'hb9eec03c),
	.w4(32'h3b179f81),
	.w5(32'h3adad112),
	.w6(32'h3b1b41a3),
	.w7(32'h3bae8fd6),
	.w8(32'hb5fcce5b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a195d02),
	.w1(32'hbb93a3e9),
	.w2(32'hba03cfeb),
	.w3(32'h3b00b0da),
	.w4(32'hbb86405b),
	.w5(32'h3a9c7a3e),
	.w6(32'hbae59784),
	.w7(32'h3a27eca5),
	.w8(32'h3a1c10af),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac990af),
	.w1(32'h3b1ca7f9),
	.w2(32'h3bbfac14),
	.w3(32'hb95280fc),
	.w4(32'h3b7d75b5),
	.w5(32'h3a784adb),
	.w6(32'hba0d44b2),
	.w7(32'h3af11826),
	.w8(32'h3bcf45a2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcf42c),
	.w1(32'hbb44b68f),
	.w2(32'hbc19f0cf),
	.w3(32'h3b80bf9a),
	.w4(32'hbc04e1a8),
	.w5(32'hb9f7e1e8),
	.w6(32'hbc190008),
	.w7(32'h395c53ec),
	.w8(32'h3ae58e6e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8628e0),
	.w1(32'h3bbac683),
	.w2(32'h3bb9633f),
	.w3(32'h3bd118c1),
	.w4(32'h3bf62d3c),
	.w5(32'h3b480174),
	.w6(32'hbb38efc8),
	.w7(32'hb8f33922),
	.w8(32'hba29fdfb),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34b92),
	.w1(32'h3a253af8),
	.w2(32'h3b952d57),
	.w3(32'h3a37505a),
	.w4(32'hbad49d52),
	.w5(32'h3acc7506),
	.w6(32'h3983a30e),
	.w7(32'h3a668c69),
	.w8(32'h3987e731),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c2c16),
	.w1(32'hbb0a5563),
	.w2(32'hbb6a516b),
	.w3(32'h3a87a828),
	.w4(32'h3ac32df7),
	.w5(32'h3b583d3f),
	.w6(32'h3bace419),
	.w7(32'hbabb59e4),
	.w8(32'hbb2571b7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule