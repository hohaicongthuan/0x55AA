module layer_8_featuremap_85(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f01a9a),
	.w1(32'h39687ae4),
	.w2(32'h39e1c32d),
	.w3(32'h3a1468f0),
	.w4(32'h37995261),
	.w5(32'h38b135a3),
	.w6(32'h39af64dc),
	.w7(32'h3a70ef15),
	.w8(32'hb6256df3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b87102),
	.w1(32'h39dd90d6),
	.w2(32'h3957bf9f),
	.w3(32'h39d21a23),
	.w4(32'h396adffd),
	.w5(32'hb79955aa),
	.w6(32'h3926594b),
	.w7(32'h39d942cd),
	.w8(32'hb94d0012),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391bdb9b),
	.w1(32'h38a51717),
	.w2(32'h37cd9b1a),
	.w3(32'h396c88ee),
	.w4(32'hb85c30ed),
	.w5(32'hb97dfb96),
	.w6(32'hb89dd4ae),
	.w7(32'h39324e4a),
	.w8(32'hb9a857c5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ceb49),
	.w1(32'hbb27b94e),
	.w2(32'hbb31f0f6),
	.w3(32'hbab370cd),
	.w4(32'hb94f8453),
	.w5(32'hb9a477b2),
	.w6(32'hbabe449a),
	.w7(32'hbb3be960),
	.w8(32'h39c32a96),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a350833),
	.w1(32'h397fcbf0),
	.w2(32'h3a257904),
	.w3(32'h39ef5e52),
	.w4(32'h37cf725f),
	.w5(32'h39709f66),
	.w6(32'h39566d97),
	.w7(32'h3a371054),
	.w8(32'h3ae266db),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac09616),
	.w1(32'h3ad260b5),
	.w2(32'h3aaca151),
	.w3(32'h3ac2aabf),
	.w4(32'h3aa4fb77),
	.w5(32'h3a02e579),
	.w6(32'h3afaf050),
	.w7(32'h3afff014),
	.w8(32'hb8d5c30d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c9ace),
	.w1(32'h3a0991ff),
	.w2(32'h39d2e817),
	.w3(32'h3a0c1afd),
	.w4(32'h38f74931),
	.w5(32'hb9252937),
	.w6(32'h39abb3fe),
	.w7(32'h3a7f2c5b),
	.w8(32'h39c5155a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39bbde),
	.w1(32'hb8fd272d),
	.w2(32'h39f8d8b9),
	.w3(32'h39f8ede8),
	.w4(32'h381ddec4),
	.w5(32'h39be0a89),
	.w6(32'h37b368fa),
	.w7(32'h3a34d790),
	.w8(32'hb8aa7052),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d0348),
	.w1(32'h3a1b90cb),
	.w2(32'h3a150be2),
	.w3(32'h3a46454f),
	.w4(32'h3954b991),
	.w5(32'hb8df6748),
	.w6(32'h3941f88b),
	.w7(32'h3a91f269),
	.w8(32'hba61d722),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359319),
	.w1(32'hbb885f74),
	.w2(32'hbad50fc3),
	.w3(32'hbb3a075d),
	.w4(32'hbb0b91f4),
	.w5(32'hbb1a07d5),
	.w6(32'h39905ed4),
	.w7(32'hbaeacfe0),
	.w8(32'hb99799bb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ccfcdf),
	.w1(32'hb9a33ae1),
	.w2(32'hb989c837),
	.w3(32'hb9004521),
	.w4(32'hba1b26a0),
	.w5(32'hba2ac7a1),
	.w6(32'hb98218d7),
	.w7(32'hb93ae8aa),
	.w8(32'hb86a4178),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a15cd),
	.w1(32'h39b7ec01),
	.w2(32'h39738701),
	.w3(32'h39f43537),
	.w4(32'h3912ccc7),
	.w5(32'hb8ff2a8e),
	.w6(32'h39280645),
	.w7(32'h3a0e4f9c),
	.w8(32'hb7dd5307),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4a381),
	.w1(32'h39d4a31e),
	.w2(32'h39959408),
	.w3(32'h392bc79c),
	.w4(32'hb7510b6e),
	.w5(32'hb865c09c),
	.w6(32'h38b16dea),
	.w7(32'h3a0cb8b8),
	.w8(32'h3b099713),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3f37a),
	.w1(32'h3ae7523a),
	.w2(32'h3aca5f8d),
	.w3(32'h3ad8af0d),
	.w4(32'h3ab7c887),
	.w5(32'h3a2f9411),
	.w6(32'h3b1198d2),
	.w7(32'h3b1d97e2),
	.w8(32'h3a70f851),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9513dc),
	.w1(32'h3a786edc),
	.w2(32'h3a5c14c7),
	.w3(32'h3a9a629e),
	.w4(32'h3a524a22),
	.w5(32'h393126f6),
	.w6(32'h3a96046a),
	.w7(32'h3aa07bde),
	.w8(32'hb8714613),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a084c),
	.w1(32'hb90bd0aa),
	.w2(32'h39a08ffe),
	.w3(32'h375e48d3),
	.w4(32'hb9b839e7),
	.w5(32'hb8d92a64),
	.w6(32'hb8fd00e5),
	.w7(32'hb6f0904d),
	.w8(32'hba452fd8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fa432),
	.w1(32'hbab3b642),
	.w2(32'hbb8596f1),
	.w3(32'hba18cffd),
	.w4(32'h3b247f5b),
	.w5(32'h3b0f357c),
	.w6(32'hb99353eb),
	.w7(32'hba166751),
	.w8(32'hba26101b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b55b5),
	.w1(32'hb8fbf564),
	.w2(32'hb78d4fa6),
	.w3(32'hb942f0c9),
	.w4(32'hb9bbc3c5),
	.w5(32'hb973e7cd),
	.w6(32'hba01b813),
	.w7(32'hb725f50d),
	.w8(32'hb95fac99),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3806b0df),
	.w1(32'hba8f52e2),
	.w2(32'hb9d56036),
	.w3(32'hb9504f1a),
	.w4(32'hbaaa7f09),
	.w5(32'hba062c40),
	.w6(32'hba811769),
	.w7(32'h392a2fd7),
	.w8(32'h3b5ea916),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381e4425),
	.w1(32'h3b100e41),
	.w2(32'hbb0cda51),
	.w3(32'h39b9efea),
	.w4(32'h392f176c),
	.w5(32'h3af1e8e6),
	.w6(32'h38931e01),
	.w7(32'hb8cda59e),
	.w8(32'h382ce961),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c2715),
	.w1(32'hb9e27426),
	.w2(32'h3880f6f6),
	.w3(32'h39defcbd),
	.w4(32'hb9e18b68),
	.w5(32'hb85f91db),
	.w6(32'hb95f13bf),
	.w7(32'h3a022400),
	.w8(32'h3a088d03),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a813a90),
	.w1(32'h3a169368),
	.w2(32'h3a5a567b),
	.w3(32'h3a573bfc),
	.w4(32'h39a53d1f),
	.w5(32'h39b27637),
	.w6(32'h39d11df0),
	.w7(32'h3a8dcce7),
	.w8(32'h37b7af7f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8521b8),
	.w1(32'hbabf3b0e),
	.w2(32'hb9c3a1cb),
	.w3(32'hba8a2e44),
	.w4(32'hba90d81d),
	.w5(32'h39a7cd78),
	.w6(32'hba4c9387),
	.w7(32'h37e5a053),
	.w8(32'hb7f5e8ec),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c214f5),
	.w1(32'hba49c23b),
	.w2(32'h3996a422),
	.w3(32'hb984ec09),
	.w4(32'hb9f774bd),
	.w5(32'h3a02e329),
	.w6(32'hba0fd778),
	.w7(32'h39eacb85),
	.w8(32'hb9146b82),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d78d03),
	.w1(32'h395cc541),
	.w2(32'hba0f51d9),
	.w3(32'hba9f8120),
	.w4(32'hba728791),
	.w5(32'hb8e49302),
	.w6(32'hbaa74fd4),
	.w7(32'hbaa4489e),
	.w8(32'h37801a15),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c0805),
	.w1(32'hbab17652),
	.w2(32'hb9a7379c),
	.w3(32'hba7f72ff),
	.w4(32'hba8790db),
	.w5(32'h399cb504),
	.w6(32'hba3e851e),
	.w7(32'h38306d98),
	.w8(32'hb370d622),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62bf66),
	.w1(32'hba96e062),
	.w2(32'hb98551fd),
	.w3(32'hba6179b8),
	.w4(32'hba634434),
	.w5(32'h3998b2be),
	.w6(32'hba2d00d0),
	.w7(32'h3829259b),
	.w8(32'hb9ec97fa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f73b46),
	.w1(32'hb9fb0399),
	.w2(32'hb885257f),
	.w3(32'hb92dafe4),
	.w4(32'hba9d1879),
	.w5(32'hba1d48a7),
	.w6(32'hb999bee9),
	.w7(32'h39296e31),
	.w8(32'h3a7b641e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ad3e9),
	.w1(32'hbab545fe),
	.w2(32'h3b3ac2ef),
	.w3(32'h3a8cd0a1),
	.w4(32'hbab21abd),
	.w5(32'hb89d6624),
	.w6(32'h3b28943b),
	.w7(32'h3af1b953),
	.w8(32'hb934bb12),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388394ac),
	.w1(32'h3814bfea),
	.w2(32'hb64b5f28),
	.w3(32'h38d3d603),
	.w4(32'hb74ffc08),
	.w5(32'hb9149caf),
	.w6(32'hb8c46b54),
	.w7(32'h37fb5bf6),
	.w8(32'hba3e70a9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb340a49),
	.w1(32'hba401c1b),
	.w2(32'hbb993280),
	.w3(32'hbb724eab),
	.w4(32'hba74e30f),
	.w5(32'hb9c5556f),
	.w6(32'hbac878b0),
	.w7(32'hbb6b4d3f),
	.w8(32'h3984a2d9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe78e6),
	.w1(32'h3a6d6f62),
	.w2(32'h3ab8a7eb),
	.w3(32'h3b02204f),
	.w4(32'hb95f1469),
	.w5(32'h3a0f7dd0),
	.w6(32'hb8d753a8),
	.w7(32'h3ad99687),
	.w8(32'h3a23095a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62cebc),
	.w1(32'hb90016e4),
	.w2(32'hbaf35339),
	.w3(32'hbadccd96),
	.w4(32'hb8d8e319),
	.w5(32'hb9b5f6bd),
	.w6(32'h3aa71d22),
	.w7(32'hb9684687),
	.w8(32'hbaf69580),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed9b5),
	.w1(32'hb8d467ee),
	.w2(32'hbb2aba51),
	.w3(32'hbb25af42),
	.w4(32'hb9e007cc),
	.w5(32'h38ba6429),
	.w6(32'hbb5f287e),
	.w7(32'hbbb026d9),
	.w8(32'h3af16d40),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba669c),
	.w1(32'h3aca9c01),
	.w2(32'h3ab3ad15),
	.w3(32'h3abfc110),
	.w4(32'h3aa24bd3),
	.w5(32'h3a214881),
	.w6(32'h3b013750),
	.w7(32'h3b0a49ff),
	.w8(32'h39103fa9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399878e1),
	.w1(32'hb968f553),
	.w2(32'h39099883),
	.w3(32'h381f4b44),
	.w4(32'hba15ca8e),
	.w5(32'h38af2526),
	.w6(32'hb9c41c35),
	.w7(32'h3a010d12),
	.w8(32'hba5103fa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e02a71),
	.w1(32'hb9fdab54),
	.w2(32'hba929671),
	.w3(32'hba8a016d),
	.w4(32'hba247f1c),
	.w5(32'hb9e3f240),
	.w6(32'hbabba8b8),
	.w7(32'hbac48e25),
	.w8(32'hba04354e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6a955),
	.w1(32'hb9a80c51),
	.w2(32'hb9782fd8),
	.w3(32'h38189613),
	.w4(32'hb9c6f75d),
	.w5(32'hba0a7965),
	.w6(32'hb9baa25a),
	.w7(32'hb6d60e60),
	.w8(32'h3ac7ff6a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c8723),
	.w1(32'h3ac5c523),
	.w2(32'h3aac3c3f),
	.w3(32'h3b061c3d),
	.w4(32'h3aa7c3dc),
	.w5(32'h3452910c),
	.w6(32'h3affd36a),
	.w7(32'h3af2b799),
	.w8(32'hb97c8736),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f4f2fd),
	.w1(32'h39916469),
	.w2(32'h388f1482),
	.w3(32'hb706a498),
	.w4(32'hba27b6da),
	.w5(32'hb9a5b76b),
	.w6(32'hb9302b7f),
	.w7(32'h39bf6c89),
	.w8(32'hb851d2c4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98537bf),
	.w1(32'hba1e3fb8),
	.w2(32'hb957b429),
	.w3(32'hb98b0439),
	.w4(32'hb9f067ca),
	.w5(32'h38619c9f),
	.w6(32'hb94205a3),
	.w7(32'hb8dc287a),
	.w8(32'hbf460d1c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf684620),
	.w1(32'hbe284486),
	.w2(32'hbf10822f),
	.w3(32'hbf386990),
	.w4(32'hbf3b2be0),
	.w5(32'h3e517f56),
	.w6(32'hbedf4ed7),
	.w7(32'hbee487b4),
	.w8(32'hbeff9ba2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9fde44),
	.w1(32'h3ea46589),
	.w2(32'hbf6c9596),
	.w3(32'hbf67beb6),
	.w4(32'hbf0db506),
	.w5(32'h3e38a4d2),
	.w6(32'hbf51774f),
	.w7(32'h3cdf95db),
	.w8(32'hbf7c3441),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d90b2dc),
	.w1(32'hbef72402),
	.w2(32'hbf2aa4ab),
	.w3(32'hbd5da755),
	.w4(32'hbd6172a8),
	.w5(32'hbdfb7e06),
	.w6(32'hbcb9ee35),
	.w7(32'hbeb77e5a),
	.w8(32'hbf9137d5),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf61f893),
	.w1(32'hbf641a81),
	.w2(32'hbf076185),
	.w3(32'hbc64c399),
	.w4(32'hbee36bea),
	.w5(32'hbf266a60),
	.w6(32'h3e73096b),
	.w7(32'h3dcf0f60),
	.w8(32'h3d1faaf2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3efeff8b),
	.w1(32'hbf2ee021),
	.w2(32'h3dabfe7e),
	.w3(32'h3e927d2f),
	.w4(32'hbf5712fd),
	.w5(32'hbf326235),
	.w6(32'hbd545574),
	.w7(32'hbed73eda),
	.w8(32'hbd1c6bc8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf74aa8b),
	.w1(32'hbf0e3147),
	.w2(32'hbf40d589),
	.w3(32'h3e26a1e4),
	.w4(32'hbf13ef6d),
	.w5(32'hbf5178e5),
	.w6(32'h3e8219de),
	.w7(32'hbf97811f),
	.w8(32'hbf2fbc67),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe577760),
	.w1(32'hbf361f79),
	.w2(32'h3f128e78),
	.w3(32'hbed7496d),
	.w4(32'hbf0cb9e3),
	.w5(32'hbdb2e8b7),
	.w6(32'hbea15a13),
	.w7(32'hbf25612d),
	.w8(32'hbebd5f06),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ee6a7f7),
	.w1(32'h3f0e4e8d),
	.w2(32'h3f373696),
	.w3(32'h3ef3198f),
	.w4(32'h3f341b3c),
	.w5(32'h3f879a49),
	.w6(32'h3ec2e6ff),
	.w7(32'h3f604f4c),
	.w8(32'h3fa0fc8f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f824c0e),
	.w1(32'h3f114262),
	.w2(32'h3f8244fb),
	.w3(32'h3f1df001),
	.w4(32'h3f9c9f1f),
	.w5(32'h3f9e0120),
	.w6(32'h3f18541b),
	.w7(32'h3f4ef41b),
	.w8(32'h3fd64140),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f01654b),
	.w1(32'h3f73b3d1),
	.w2(32'h3f4d99aa),
	.w3(32'h3f29a126),
	.w4(32'h3f278609),
	.w5(32'h3f51f008),
	.w6(32'h3fa0eb59),
	.w7(32'h3f98dd65),
	.w8(32'h3f331c8d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f30b63d),
	.w1(32'h3fb542e6),
	.w2(32'h3fb1dab7),
	.w3(32'h3f68be54),
	.w4(32'h3ef7e2de),
	.w5(32'h3f7c107a),
	.w6(32'h3f82b358),
	.w7(32'h3f3c50b9),
	.w8(32'h3fa10723),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f240a53),
	.w1(32'h3f89fcd0),
	.w2(32'h3f90916f),
	.w3(32'h3ed95d5b),
	.w4(32'h3f6a8789),
	.w5(32'h3eea0727),
	.w6(32'h3f9de7d9),
	.w7(32'h3ed4b740),
	.w8(32'h3f1663e6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f8a9db2),
	.w1(32'h3f8dcf2e),
	.w2(32'h3f625fa5),
	.w3(32'h3eecf702),
	.w4(32'h3efee374),
	.w5(32'h3f6e1f50),
	.w6(32'h3fbba14b),
	.w7(32'h3f54a283),
	.w8(32'h3f85fb65),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f94bcaa),
	.w1(32'h3f748968),
	.w2(32'h3f384b90),
	.w3(32'h3f902490),
	.w4(32'h3f80c594),
	.w5(32'h3f8d70bd),
	.w6(32'h3f3d82d6),
	.w7(32'h3f634cee),
	.w8(32'h3f452b58),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f28f80f),
	.w1(32'hbe33afb0),
	.w2(32'hbde0f102),
	.w3(32'h3d8671a8),
	.w4(32'h3d8663c4),
	.w5(32'h3da8a655),
	.w6(32'hbdda0d0d),
	.w7(32'hbdb0ea6b),
	.w8(32'h3d072e0d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e7bd100),
	.w1(32'h3d8eb218),
	.w2(32'hbe9fab2e),
	.w3(32'hbe556553),
	.w4(32'h3eaff448),
	.w5(32'hbe362e15),
	.w6(32'h3e427458),
	.w7(32'h3e9542f0),
	.w8(32'hbef13f8c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbea97b84),
	.w1(32'hbf09ccbe),
	.w2(32'hbeef0d84),
	.w3(32'hbe8aa4c2),
	.w4(32'hbf02d6fe),
	.w5(32'hbe473197),
	.w6(32'hbe3f43af),
	.w7(32'hbe2e543b),
	.w8(32'hbe98aa45),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc045708),
	.w1(32'hbe1034a0),
	.w2(32'hbd87139b),
	.w3(32'hbcc9c495),
	.w4(32'h3df294d9),
	.w5(32'h3e9af905),
	.w6(32'hbebdd969),
	.w7(32'hbd5a60df),
	.w8(32'hbdb2280e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe926863),
	.w1(32'h3d56e7fc),
	.w2(32'hbdfc3c61),
	.w3(32'h3e61bc14),
	.w4(32'hbe324af4),
	.w5(32'h3e83d1d0),
	.w6(32'hbdd874bb),
	.w7(32'hbe914f35),
	.w8(32'h3def06da),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d988753),
	.w1(32'h3f60fef7),
	.w2(32'hbea6f2d6),
	.w3(32'hbeca59c1),
	.w4(32'hbec080c0),
	.w5(32'h3cc52393),
	.w6(32'hbdf207cc),
	.w7(32'h3e0761b0),
	.w8(32'hbe0fad3f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbedd24a5),
	.w1(32'hbd98c3fa),
	.w2(32'hbe438560),
	.w3(32'h3d195a41),
	.w4(32'hbe3ddadf),
	.w5(32'hbe5030ff),
	.w6(32'hbeaab9c0),
	.w7(32'hbf124ac2),
	.w8(32'h3eacec1e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec3db49),
	.w1(32'h3b82956f),
	.w2(32'h3d400448),
	.w3(32'h3de5d2d3),
	.w4(32'h3b779951),
	.w5(32'h3cd0311c),
	.w6(32'h3b764fc8),
	.w7(32'h3c2af5d3),
	.w8(32'h3cd4142d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d126c18),
	.w1(32'h3d0a2d0c),
	.w2(32'h3e058d9d),
	.w3(32'h3dd2919d),
	.w4(32'h3c81bd21),
	.w5(32'h3cbe92a2),
	.w6(32'h3d1d41f5),
	.w7(32'h3cb288fc),
	.w8(32'h3dea96e6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d36b5aa),
	.w1(32'h3d87253b),
	.w2(32'h3d009d8b),
	.w3(32'h3e22bdf6),
	.w4(32'h3e2bcab4),
	.w5(32'h3e2f7d7f),
	.w6(32'h3c5f056f),
	.w7(32'h3da368a9),
	.w8(32'h3d1bb7c1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d394524),
	.w1(32'h3cd1aa39),
	.w2(32'h3b46d961),
	.w3(32'h3d3625ff),
	.w4(32'h3daaeef3),
	.w5(32'h3c8d5b22),
	.w6(32'h3cafc3ef),
	.w7(32'h3e21db5c),
	.w8(32'h3dfd0e34),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1fc667),
	.w1(32'h3e600230),
	.w2(32'h3ce23ab9),
	.w3(32'h3d73d363),
	.w4(32'h3e043d4e),
	.w5(32'h3b20ff1c),
	.w6(32'h3d5bf49f),
	.w7(32'h3e2df395),
	.w8(32'h3d4c6f81),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceb088f),
	.w1(32'h3b271b39),
	.w2(32'h3cabb5a6),
	.w3(32'h3cc445fb),
	.w4(32'h3df6c358),
	.w5(32'h3d0896a8),
	.w6(32'h3e0ea7d7),
	.w7(32'h3db5ad14),
	.w8(32'h3c6e6081),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3a1671),
	.w1(32'h3db55587),
	.w2(32'h3d712846),
	.w3(32'h3d85acf7),
	.w4(32'h3d3bcb06),
	.w5(32'h3d06a6b2),
	.w6(32'h3d35ca91),
	.w7(32'h3d30f3c6),
	.w8(32'h3cd72c79),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dc7caf6),
	.w1(32'h3ba9de23),
	.w2(32'hbb69a09d),
	.w3(32'h3d56313a),
	.w4(32'hbb9d3b4a),
	.w5(32'hbbb779ab),
	.w6(32'h3cdc0af7),
	.w7(32'h3b318176),
	.w8(32'hbaf1a04e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7109bd),
	.w1(32'h3ae6b4db),
	.w2(32'h3c83cba9),
	.w3(32'h3b47b179),
	.w4(32'hba8e896b),
	.w5(32'h3a7ac3f7),
	.w6(32'hba1419ed),
	.w7(32'h3c495250),
	.w8(32'hbc0f0498),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51d6c7),
	.w1(32'hbb1b7d68),
	.w2(32'h3b5d71be),
	.w3(32'h3941a45b),
	.w4(32'h3b4594fe),
	.w5(32'hb9a09a3e),
	.w6(32'h3b353df5),
	.w7(32'h3986bbc0),
	.w8(32'hbb8b7f46),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc188f66),
	.w1(32'h3a934e9a),
	.w2(32'hbba0e1fe),
	.w3(32'h3b854e11),
	.w4(32'h3bcfad77),
	.w5(32'h3d3b521c),
	.w6(32'hba7db75d),
	.w7(32'h3bac22ea),
	.w8(32'h3b8aa3dd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c122c59),
	.w1(32'h3cd93a28),
	.w2(32'hbbd3e358),
	.w3(32'hbc3ea539),
	.w4(32'hbb9dbb94),
	.w5(32'h3b1cf232),
	.w6(32'hbb6d9d60),
	.w7(32'hbaa5c2fb),
	.w8(32'hbba972d6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cdf34),
	.w1(32'hbbed2613),
	.w2(32'hba07627c),
	.w3(32'h3c2fe020),
	.w4(32'h3bed5b85),
	.w5(32'h3b93cd35),
	.w6(32'hbb98f615),
	.w7(32'hbbd4a5ed),
	.w8(32'h3c2f7dfe),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af84a40),
	.w1(32'hbaac91d2),
	.w2(32'h3b38c7d0),
	.w3(32'h3c5ab6db),
	.w4(32'h3b0c066c),
	.w5(32'h3c0ec286),
	.w6(32'h3af5ac87),
	.w7(32'hba01e65f),
	.w8(32'h3b152746),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e8655),
	.w1(32'hb8f4feff),
	.w2(32'h3a914143),
	.w3(32'hbbe1d3a5),
	.w4(32'h3c64f485),
	.w5(32'hbbc21db5),
	.w6(32'hbc64e526),
	.w7(32'h3c28a17c),
	.w8(32'hbac18f3e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c99c5c),
	.w1(32'h3a899798),
	.w2(32'hba717fef),
	.w3(32'h3b0454e4),
	.w4(32'h3a80992e),
	.w5(32'hba3a97b3),
	.w6(32'h3bd33c73),
	.w7(32'h3b4e0248),
	.w8(32'h3c181edc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d094),
	.w1(32'hbb675a4c),
	.w2(32'hbb332df0),
	.w3(32'h3b829844),
	.w4(32'hbb42fa3e),
	.w5(32'h3b2b4126),
	.w6(32'h3b1eb464),
	.w7(32'h3af1996e),
	.w8(32'h3c11a647),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1de8a),
	.w1(32'hbb35e8af),
	.w2(32'hbb194b67),
	.w3(32'hbb3484c7),
	.w4(32'h3ba226b5),
	.w5(32'hbbf5487e),
	.w6(32'hbad53542),
	.w7(32'h3a1b4972),
	.w8(32'hb902fc14),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be82f73),
	.w1(32'hbc0771ff),
	.w2(32'h3c2382c8),
	.w3(32'hb9910047),
	.w4(32'hbbd1ebdc),
	.w5(32'hbbf09942),
	.w6(32'h3b83b4ae),
	.w7(32'hbb933cac),
	.w8(32'h3bcd440b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba8f03),
	.w1(32'hbb6bd007),
	.w2(32'hbaed27bb),
	.w3(32'h3b04f844),
	.w4(32'h3b4e0d4d),
	.w5(32'h3b5463f5),
	.w6(32'hbc01a5ae),
	.w7(32'hba88d82e),
	.w8(32'h3a787a9b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42e57c),
	.w1(32'h3a894384),
	.w2(32'h39d76bd3),
	.w3(32'hbbed7d8c),
	.w4(32'hbd05bd6b),
	.w5(32'hbbbbb636),
	.w6(32'hbb25702d),
	.w7(32'hb857dca2),
	.w8(32'hbafe1a59),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cf4d4),
	.w1(32'hbb1629a8),
	.w2(32'hbb7e8419),
	.w3(32'h3ad039ed),
	.w4(32'h3b3a72ef),
	.w5(32'hbba2b3c6),
	.w6(32'h3a34abe2),
	.w7(32'hbacf96f1),
	.w8(32'hbaee1099),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabadd31),
	.w1(32'h3c2fa854),
	.w2(32'hbb91230d),
	.w3(32'hbba755ad),
	.w4(32'h3b4fa707),
	.w5(32'h3b898d95),
	.w6(32'h3bef4701),
	.w7(32'hbc012480),
	.w8(32'h3c8374fe),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c207d7f),
	.w1(32'h3b325d90),
	.w2(32'h3c13aa83),
	.w3(32'hbbde39dd),
	.w4(32'hbb18f3c3),
	.w5(32'hbbe35cc9),
	.w6(32'h3c0f2706),
	.w7(32'h3bd81eba),
	.w8(32'hbbe8a742),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8726c),
	.w1(32'h3bd0c8b1),
	.w2(32'h3b569a16),
	.w3(32'h3bcdee10),
	.w4(32'hbbc910cb),
	.w5(32'h3d183a99),
	.w6(32'hbb7b9e0c),
	.w7(32'h3c27ef0f),
	.w8(32'hbc327c89),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbafb5),
	.w1(32'h3c11d5bd),
	.w2(32'hbc0ca4de),
	.w3(32'hbb9bddf2),
	.w4(32'hbc3dae17),
	.w5(32'hbb510d02),
	.w6(32'hbb554abe),
	.w7(32'hbbc98393),
	.w8(32'hbb8c3678),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b23cf),
	.w1(32'h36858ec2),
	.w2(32'h3b923259),
	.w3(32'hbc46fe23),
	.w4(32'h3af78550),
	.w5(32'h3b9b5d26),
	.w6(32'h3b0a253e),
	.w7(32'hbc15a889),
	.w8(32'hbc1b8287),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aa1f5),
	.w1(32'h3b9a2eca),
	.w2(32'hbbd86ddc),
	.w3(32'h3c0cb73e),
	.w4(32'hbbd6f9f0),
	.w5(32'hbb5afa41),
	.w6(32'h3b6545f5),
	.w7(32'hbb2ba5ba),
	.w8(32'hbc3c8dde),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc9d34d),
	.w1(32'hba9f57c8),
	.w2(32'h3bdb415c),
	.w3(32'hbbf3b138),
	.w4(32'hbc05ecb1),
	.w5(32'h3c3a0369),
	.w6(32'h3b0ba1b4),
	.w7(32'hbbcf10e0),
	.w8(32'hba913fd2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86d783),
	.w1(32'h3bb92b4e),
	.w2(32'h3b36b6f0),
	.w3(32'h3acb8991),
	.w4(32'h37153772),
	.w5(32'hbbda490d),
	.w6(32'h3bffc48d),
	.w7(32'hbc0e2411),
	.w8(32'h3b9859cf),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9864231),
	.w1(32'hbc0aba2e),
	.w2(32'h3c1a4f71),
	.w3(32'h3c884227),
	.w4(32'h3a41ef0a),
	.w5(32'h3b5c97eb),
	.w6(32'h3c0cba69),
	.w7(32'hbbc9ddd8),
	.w8(32'h3cbab6f9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08cee7),
	.w1(32'hbb3e73cd),
	.w2(32'h3c1888e9),
	.w3(32'h3bc89dc2),
	.w4(32'h3b4b360b),
	.w5(32'hbbb886ca),
	.w6(32'h3ab55452),
	.w7(32'hbbb9cec0),
	.w8(32'hbc25e6de),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0d53d),
	.w1(32'hbc385a90),
	.w2(32'hbb61e4c9),
	.w3(32'hbb553769),
	.w4(32'h3c00507f),
	.w5(32'h3b108a95),
	.w6(32'hbb875f70),
	.w7(32'hbc21ee70),
	.w8(32'h3b4333cb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ba210),
	.w1(32'h3d343ef2),
	.w2(32'h3b6855a7),
	.w3(32'hbbb7c162),
	.w4(32'hb93e4d28),
	.w5(32'h3b994fe6),
	.w6(32'h3c5815dc),
	.w7(32'hbac7672e),
	.w8(32'hbb08ad50),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa0488),
	.w1(32'h3ba8b0e0),
	.w2(32'hbc6954e4),
	.w3(32'hbb457196),
	.w4(32'h3b2a5d43),
	.w5(32'hbafff153),
	.w6(32'hbba641e8),
	.w7(32'hbb8db446),
	.w8(32'hba84f559),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c5fed),
	.w1(32'h3a77ffd9),
	.w2(32'hba7c5440),
	.w3(32'h3992f494),
	.w4(32'hbb36b68f),
	.w5(32'h3af6aa02),
	.w6(32'hbc1e92ad),
	.w7(32'h3c41d320),
	.w8(32'hbc620a85),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab06b5e),
	.w1(32'hbb343536),
	.w2(32'hbb538ab6),
	.w3(32'hba971b08),
	.w4(32'h390bd025),
	.w5(32'hbb3d329a),
	.w6(32'h3aa834fa),
	.w7(32'h3b5333cb),
	.w8(32'hbc2fe6a9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5de9eb),
	.w1(32'hbc60642c),
	.w2(32'hbab85e40),
	.w3(32'h3c440fb0),
	.w4(32'h3b3fdae5),
	.w5(32'hbb2e580d),
	.w6(32'h3bf2e8ed),
	.w7(32'hb9a4674f),
	.w8(32'h3c7f7eb9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb902ae8),
	.w1(32'h3ad3e8b0),
	.w2(32'hbbc112d5),
	.w3(32'hbbe68099),
	.w4(32'h3b4136ab),
	.w5(32'h3b1482ba),
	.w6(32'h3b0f2993),
	.w7(32'h3b65b680),
	.w8(32'hba6463e5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f28cc),
	.w1(32'hbba3bfe4),
	.w2(32'hbc26e29c),
	.w3(32'hbaebb493),
	.w4(32'hbbd7124e),
	.w5(32'hbb0fcf63),
	.w6(32'h3b870953),
	.w7(32'h3bc9ebd7),
	.w8(32'hbb7ba3e8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b38bc),
	.w1(32'hbc1a05ac),
	.w2(32'hba97ad20),
	.w3(32'hbbda3706),
	.w4(32'h3bc36ed0),
	.w5(32'hb9d5749f),
	.w6(32'hb9c62216),
	.w7(32'hbbdf1d00),
	.w8(32'h3c1b1b54),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08e8ab),
	.w1(32'h3b2a495b),
	.w2(32'hb9a0eb92),
	.w3(32'hbc85b90f),
	.w4(32'h3b28b30f),
	.w5(32'hbb1da10d),
	.w6(32'hbafa0fde),
	.w7(32'h3c48c0f0),
	.w8(32'hbc3e6936),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2be94c),
	.w1(32'hbb9be969),
	.w2(32'hbc6ca9cc),
	.w3(32'hbb9b8a08),
	.w4(32'hbae13b1c),
	.w5(32'hbb94ca38),
	.w6(32'h3ba4265b),
	.w7(32'hb93f0d2c),
	.w8(32'hb99b24aa),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6acd86),
	.w1(32'h3ada5ca5),
	.w2(32'hbb9d5768),
	.w3(32'h3a687618),
	.w4(32'h3beadc94),
	.w5(32'hbc1f63eb),
	.w6(32'hbc6d5abf),
	.w7(32'h3b829ef7),
	.w8(32'hbb45e51f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b9fac),
	.w1(32'h3b240696),
	.w2(32'h3ad60e59),
	.w3(32'hba56c51f),
	.w4(32'h3ba4e528),
	.w5(32'hbb8261e2),
	.w6(32'h3b9817f3),
	.w7(32'hbadd963b),
	.w8(32'h3820eefc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0574ce),
	.w1(32'hba22973a),
	.w2(32'hbadc1b60),
	.w3(32'h3caa94f9),
	.w4(32'hbaa1f4ba),
	.w5(32'hbb4081f3),
	.w6(32'h3c8fa2fc),
	.w7(32'h3acdb0af),
	.w8(32'h3ac67a10),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4f2f8),
	.w1(32'hbb60b7b6),
	.w2(32'h3c9e9114),
	.w3(32'hbc2a9c23),
	.w4(32'h3c5e29e0),
	.w5(32'h3b35807e),
	.w6(32'h3b370f87),
	.w7(32'hbbc92b64),
	.w8(32'hbc19fe82),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2af6bd),
	.w1(32'hbbad091f),
	.w2(32'hbafc36d0),
	.w3(32'h3bff6da1),
	.w4(32'h3b6bd12c),
	.w5(32'h3ad6b83b),
	.w6(32'h3bfd85fd),
	.w7(32'h3d6811cb),
	.w8(32'h3a6e5ff6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd038e9),
	.w1(32'hba449fc5),
	.w2(32'h3b84435d),
	.w3(32'hb8edeb86),
	.w4(32'hbc021a4e),
	.w5(32'hbb773ec4),
	.w6(32'hbb8bd6a8),
	.w7(32'h3bd0df58),
	.w8(32'hbc1e5843),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb918029),
	.w1(32'h3ae4404b),
	.w2(32'hbba5a57c),
	.w3(32'h3b079349),
	.w4(32'hbb038a0a),
	.w5(32'h3b2bc409),
	.w6(32'h3aee080f),
	.w7(32'hba8295c9),
	.w8(32'hba1c2f8e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0b2e0),
	.w1(32'h3a8e8b48),
	.w2(32'hbb8b7a04),
	.w3(32'h3c03e693),
	.w4(32'h3b1f9e1f),
	.w5(32'h3cc05cf0),
	.w6(32'h3d48d3f4),
	.w7(32'hbbc5754c),
	.w8(32'h3ab18394),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dc232b7),
	.w1(32'h3ae64c3c),
	.w2(32'hb92a356a),
	.w3(32'hbbd9d2e0),
	.w4(32'h3c6f1b5f),
	.w5(32'h3b8dbe09),
	.w6(32'hbcad608f),
	.w7(32'hba39a5ff),
	.w8(32'hbcc35b0c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1f9480),
	.w1(32'h3a8ae4ad),
	.w2(32'hbc856702),
	.w3(32'hba9436da),
	.w4(32'hbcc32f0b),
	.w5(32'h3c6e3ad2),
	.w6(32'hb87df32e),
	.w7(32'h3c811289),
	.w8(32'h3c827fe8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbbf6f9),
	.w1(32'hbc32d635),
	.w2(32'h3a9ff995),
	.w3(32'h3d486314),
	.w4(32'hbb95e1bc),
	.w5(32'h3bd470f1),
	.w6(32'hbbc907f7),
	.w7(32'h3c09b9a0),
	.w8(32'hbab2577d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de5d5a),
	.w1(32'h3bcae661),
	.w2(32'hbc1deca2),
	.w3(32'h3cdaa958),
	.w4(32'h3b7fda28),
	.w5(32'h3b228d09),
	.w6(32'h3a851597),
	.w7(32'h3b03322c),
	.w8(32'h3bcb11a1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bf680),
	.w1(32'hbb9117da),
	.w2(32'hbc8384e4),
	.w3(32'hbd0b8f42),
	.w4(32'h3c5af075),
	.w5(32'h3bdcddfe),
	.w6(32'hbbcfffcd),
	.w7(32'h374d7995),
	.w8(32'hbac323c7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4b468),
	.w1(32'hbbeca8c3),
	.w2(32'h3b260394),
	.w3(32'hbc8dadd8),
	.w4(32'hbcd98570),
	.w5(32'h3b392544),
	.w6(32'hbc167f95),
	.w7(32'h3bb89fbd),
	.w8(32'hbc747aa3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98bfbb),
	.w1(32'h3bda0b5a),
	.w2(32'h3c116230),
	.w3(32'hbbfd2c7d),
	.w4(32'h3bdc986b),
	.w5(32'h39f1f29e),
	.w6(32'hba314aac),
	.w7(32'hbcd20274),
	.w8(32'h3c65dda4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c375d90),
	.w1(32'h3cd05909),
	.w2(32'h3c4f5f58),
	.w3(32'hbc3b758e),
	.w4(32'h3c5bfbac),
	.w5(32'hbb65ea8b),
	.w6(32'h3cc746a3),
	.w7(32'hbb95322e),
	.w8(32'hbc80c15a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d00c7),
	.w1(32'h3c29993f),
	.w2(32'h3d4bdaf5),
	.w3(32'h3c88d0df),
	.w4(32'hbc08d3c9),
	.w5(32'h3c2964ad),
	.w6(32'h3b4983f2),
	.w7(32'h3c38266f),
	.w8(32'h3b71e03f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e3070),
	.w1(32'hbc5ab2e2),
	.w2(32'hbaf6a601),
	.w3(32'h3cd7645b),
	.w4(32'hbbdb9dcb),
	.w5(32'h3b14eef3),
	.w6(32'h3cbf3f3e),
	.w7(32'h3b21d191),
	.w8(32'h3adead1f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82eda7),
	.w1(32'hbc8f6f31),
	.w2(32'hbca693bb),
	.w3(32'hba9bb7cb),
	.w4(32'h3c6bad6b),
	.w5(32'h3c7b72e9),
	.w6(32'hbb04a533),
	.w7(32'hbbebc044),
	.w8(32'hbc340c02),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72724e),
	.w1(32'hbba36e21),
	.w2(32'h3badf841),
	.w3(32'h3a3e33a1),
	.w4(32'hbbb77562),
	.w5(32'hbd3d2f80),
	.w6(32'hb79dec58),
	.w7(32'h3b46c748),
	.w8(32'hb995a200),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad746f),
	.w1(32'h3bf75e4b),
	.w2(32'h3ae78f07),
	.w3(32'h3b405005),
	.w4(32'h3c08d883),
	.w5(32'h3a96c32d),
	.w6(32'hba9165db),
	.w7(32'h3bb3fdc1),
	.w8(32'h3c37cc60),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc9e5e0),
	.w1(32'hbd2375a2),
	.w2(32'hbcfa3bbb),
	.w3(32'h3b6b363e),
	.w4(32'h3c07d115),
	.w5(32'h3ba250fd),
	.w6(32'hba939a3c),
	.w7(32'h3933780f),
	.w8(32'hbc7462a9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c080696),
	.w1(32'h3b7d463c),
	.w2(32'h3c5f4d43),
	.w3(32'hbc667f53),
	.w4(32'h3cb2d270),
	.w5(32'h3b37265a),
	.w6(32'hbbde2544),
	.w7(32'h3c1255ee),
	.w8(32'hbc06e2a0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule