module layer_10_featuremap_181(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c1a22b),
	.w1(32'hb755b215),
	.w2(32'hb6e8d641),
	.w3(32'hb7ce1188),
	.w4(32'hb6d3f3c7),
	.w5(32'hb67d658c),
	.w6(32'hb7cdf287),
	.w7(32'h36a57fd8),
	.w8(32'hb686e63e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ababc39),
	.w1(32'h3a1fc2c3),
	.w2(32'h3a598ebc),
	.w3(32'h3a834ae5),
	.w4(32'h39cc4eb9),
	.w5(32'h39d9f5d6),
	.w6(32'h39aa58d5),
	.w7(32'hb9556b0d),
	.w8(32'h39b3b6ff),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72b3e3e),
	.w1(32'hb6aaac94),
	.w2(32'hb7427737),
	.w3(32'hb6b4fa73),
	.w4(32'hb50db5a4),
	.w5(32'hb6ed8613),
	.w6(32'h35d21c79),
	.w7(32'h366d234d),
	.w8(32'hb655683c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fc4a47),
	.w1(32'hb7e33535),
	.w2(32'hb81ad9ee),
	.w3(32'h379c4ee8),
	.w4(32'hb7ca2384),
	.w5(32'hb84888ea),
	.w6(32'h37f375dd),
	.w7(32'hb4b60c7a),
	.w8(32'hb7845b6f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82c85a4),
	.w1(32'h38b7385b),
	.w2(32'h39560d6d),
	.w3(32'hb8ddd079),
	.w4(32'h37cf1bbc),
	.w5(32'h391bfbca),
	.w6(32'hb8ced0b5),
	.w7(32'hb7f74ce9),
	.w8(32'h382f8525),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387714fb),
	.w1(32'h385d52a6),
	.w2(32'hb74e8da6),
	.w3(32'h382d480f),
	.w4(32'h386827be),
	.w5(32'h375c8249),
	.w6(32'hb5bd8dde),
	.w7(32'h369a4f72),
	.w8(32'h359ccc86),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eff8a),
	.w1(32'h3a442460),
	.w2(32'h3b3d3e50),
	.w3(32'hb8533bca),
	.w4(32'h3901ed26),
	.w5(32'h3ac80257),
	.w6(32'hb985f461),
	.w7(32'hba1b9942),
	.w8(32'h3a34c8c0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2123cd),
	.w1(32'h3aed1be5),
	.w2(32'h3b69758d),
	.w3(32'hba59dc0e),
	.w4(32'hbae6b3ba),
	.w5(32'hba64ca33),
	.w6(32'hbad5f41d),
	.w7(32'hbad41976),
	.w8(32'hb9e9a524),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911773b),
	.w1(32'hba201207),
	.w2(32'hb9d98c64),
	.w3(32'h381f22e7),
	.w4(32'hba2d7932),
	.w5(32'hba1b700d),
	.w6(32'h382a4095),
	.w7(32'hb9cf6978),
	.w8(32'hb906e5d7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0fc50),
	.w1(32'h3b6ae55c),
	.w2(32'h3bcc889f),
	.w3(32'h397dfe39),
	.w4(32'hb972dc96),
	.w5(32'h3b05e6b9),
	.w6(32'hbafcaf65),
	.w7(32'hbb46e69c),
	.w8(32'hb9e85054),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93dd922),
	.w1(32'h383d524a),
	.w2(32'h39fc2bdc),
	.w3(32'hb9a3a7af),
	.w4(32'hb88b0e0d),
	.w5(32'h39b578b7),
	.w6(32'hb93b80c6),
	.w7(32'h3682b818),
	.w8(32'h39997f99),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4626f9),
	.w1(32'hba028459),
	.w2(32'h3aca5542),
	.w3(32'h3b0a6bc5),
	.w4(32'hbb6115ba),
	.w5(32'hb9b5cdd7),
	.w6(32'h3b3731a2),
	.w7(32'hbb62f0bf),
	.w8(32'h391c377e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6d641),
	.w1(32'h3bb7922d),
	.w2(32'h3bfeb978),
	.w3(32'hba3a2dff),
	.w4(32'hba52282c),
	.w5(32'h3a5ebb09),
	.w6(32'hbb121f44),
	.w7(32'hbb85ad90),
	.w8(32'hba77438e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afaab67),
	.w1(32'h3b5d1c07),
	.w2(32'h3b6a3ea7),
	.w3(32'h3aad12d1),
	.w4(32'h3b487601),
	.w5(32'h3b6445a8),
	.w6(32'h39526d87),
	.w7(32'h3b160dcc),
	.w8(32'h3b5c6c29),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2da4bf),
	.w1(32'h3b091be7),
	.w2(32'h3b375850),
	.w3(32'h39c8ecd7),
	.w4(32'hba3cfccb),
	.w5(32'h3a14b1af),
	.w6(32'hb9c70819),
	.w7(32'hba8a41f1),
	.w8(32'h3aa816c5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b615b72),
	.w1(32'h3b658c87),
	.w2(32'h3b80deda),
	.w3(32'h39870089),
	.w4(32'hb89eaa62),
	.w5(32'hb9a9522b),
	.w6(32'hba080691),
	.w7(32'hba95415c),
	.w8(32'hbac667bc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb773bbda),
	.w1(32'hb981a7d1),
	.w2(32'h374441f4),
	.w3(32'hb90db785),
	.w4(32'hb884ffca),
	.w5(32'h394475c4),
	.w6(32'hb8b1242d),
	.w7(32'hb8d0092d),
	.w8(32'h39a0e1a5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f7c27),
	.w1(32'h3b9d3a78),
	.w2(32'h3bbd222f),
	.w3(32'h3a17dbbb),
	.w4(32'h39f2ca3c),
	.w5(32'h3afcdfa8),
	.w6(32'hbb20036b),
	.w7(32'hbb31809a),
	.w8(32'h39a019ab),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b900b31),
	.w1(32'h3b85f2d3),
	.w2(32'h3b1c6343),
	.w3(32'h3ab5a968),
	.w4(32'h3a9b967d),
	.w5(32'h3a13f87a),
	.w6(32'hba5b9821),
	.w7(32'hba15bf02),
	.w8(32'hba0dd4e8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78fb5a7),
	.w1(32'hb50c894f),
	.w2(32'hb724535f),
	.w3(32'hb72bfa95),
	.w4(32'h33ab7dc6),
	.w5(32'h3599b84b),
	.w6(32'hb71e24af),
	.w7(32'h3637e430),
	.w8(32'h36a243de),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82fe9a4),
	.w1(32'hb7f40e24),
	.w2(32'hb86797c9),
	.w3(32'hb789714c),
	.w4(32'h3591d678),
	.w5(32'hb7fcd256),
	.w6(32'hb7710b26),
	.w7(32'h34c34202),
	.w8(32'hb7efe4eb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9940666),
	.w1(32'hb9c65e6c),
	.w2(32'h3aaf8fbb),
	.w3(32'hb9e505fc),
	.w4(32'hba60151b),
	.w5(32'h3a49fbfa),
	.w6(32'h39a21c32),
	.w7(32'hba1397b3),
	.w8(32'h39f10626),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bb824),
	.w1(32'h3c1fa7d5),
	.w2(32'h3c23d5ad),
	.w3(32'h3bcc8dc5),
	.w4(32'h3b833ec6),
	.w5(32'h3bcf8a01),
	.w6(32'h3a6ad52f),
	.w7(32'hb9be9865),
	.w8(32'h3bb6edf8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e8a7a),
	.w1(32'h3b6e8e0b),
	.w2(32'h3bda607b),
	.w3(32'h39b5615d),
	.w4(32'hb88c9402),
	.w5(32'h3b11ab21),
	.w6(32'hbabfa442),
	.w7(32'hbb1ec254),
	.w8(32'hb8c7b192),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc1cd1),
	.w1(32'h3b6fadca),
	.w2(32'h3bad072f),
	.w3(32'h3b2359a7),
	.w4(32'hb9e0da8d),
	.w5(32'h3af97ee8),
	.w6(32'h3ac0a446),
	.w7(32'hbb0b0977),
	.w8(32'h3a24232b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8252300),
	.w1(32'hb9255dce),
	.w2(32'hb9ea92ec),
	.w3(32'h390bb193),
	.w4(32'h399e8bbc),
	.w5(32'hb996159c),
	.w6(32'h38b9c9c8),
	.w7(32'h3a204d9a),
	.w8(32'h393901d3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ee559),
	.w1(32'hb8389aed),
	.w2(32'hb81b36a5),
	.w3(32'hb7c94ce0),
	.w4(32'h36f713a8),
	.w5(32'h383acc38),
	.w6(32'h36942ece),
	.w7(32'h3755c7db),
	.w8(32'h382b79fd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a955650),
	.w1(32'h3a099022),
	.w2(32'h3a8d1f74),
	.w3(32'hb9b5f569),
	.w4(32'hba8cb5f1),
	.w5(32'hba38d83c),
	.w6(32'h3a3ff5e6),
	.w7(32'hba7f795f),
	.w8(32'hba737c9f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe9583),
	.w1(32'hba085fe5),
	.w2(32'h39e87434),
	.w3(32'h3aa6a66c),
	.w4(32'hba1ede4e),
	.w5(32'h38cb1548),
	.w6(32'h3b26b6df),
	.w7(32'hb92fae56),
	.w8(32'h3a0a977e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23d059),
	.w1(32'h3a9db2d1),
	.w2(32'h3af6b65d),
	.w3(32'h3a251278),
	.w4(32'h3975027c),
	.w5(32'hb8619564),
	.w6(32'hb93a8dc8),
	.w7(32'hb81603d8),
	.w8(32'hb9c18511),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6551da8),
	.w1(32'hb7b28413),
	.w2(32'h36155625),
	.w3(32'h3721891c),
	.w4(32'hb6d86a3a),
	.w5(32'h37713005),
	.w6(32'h381f9812),
	.w7(32'h37efb417),
	.w8(32'h381b1ae0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93677f8),
	.w1(32'hb8f9eb2e),
	.w2(32'h37066190),
	.w3(32'hb95aeafa),
	.w4(32'hb90cfc27),
	.w5(32'h3900a457),
	.w6(32'hb9506629),
	.w7(32'hb85643c4),
	.w8(32'h398733d6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3ce51),
	.w1(32'h3b092e2d),
	.w2(32'h3b6dd17a),
	.w3(32'hb9b69130),
	.w4(32'h38cfca38),
	.w5(32'h3a9b93c9),
	.w6(32'hbaa89202),
	.w7(32'hba42d795),
	.w8(32'h39d8c246),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8556fa),
	.w1(32'h3985e406),
	.w2(32'h3a2bc8d7),
	.w3(32'h3a9a7577),
	.w4(32'hb829da16),
	.w5(32'hb99c3fde),
	.w6(32'h3a8642e7),
	.w7(32'h39888e8f),
	.w8(32'h3943fd68),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a28bc7),
	.w1(32'hb9e4374f),
	.w2(32'hb9bb2e8a),
	.w3(32'h395259b3),
	.w4(32'hb9a10ed6),
	.w5(32'hb9ae380b),
	.w6(32'h39f52bd8),
	.w7(32'hb87ca3f3),
	.w8(32'hb98f129d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1da05),
	.w1(32'h3a13c515),
	.w2(32'h3aef6a9a),
	.w3(32'h38b84d4f),
	.w4(32'hba5aa992),
	.w5(32'hb795cf87),
	.w6(32'hb7a7475f),
	.w7(32'hba8d0b8b),
	.w8(32'hb8e0f8e3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe0579),
	.w1(32'h3b822b3a),
	.w2(32'h3c00f866),
	.w3(32'hbb3b874f),
	.w4(32'h3a8418ab),
	.w5(32'h3b75a263),
	.w6(32'hbb89cb3c),
	.w7(32'hbacf30fb),
	.w8(32'h3b1bb896),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2423b),
	.w1(32'h3a49431c),
	.w2(32'h3bbfe086),
	.w3(32'h3b4e2e44),
	.w4(32'hb8d09bc8),
	.w5(32'h3bcba27f),
	.w6(32'h3b97b664),
	.w7(32'h3a940696),
	.w8(32'h3b464f31),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd44ce6),
	.w1(32'h3a56920f),
	.w2(32'h3badb822),
	.w3(32'h3ba7a077),
	.w4(32'hb69c7f1d),
	.w5(32'h3b870ee4),
	.w6(32'h3be90672),
	.w7(32'h3b2cfc90),
	.w8(32'h3b75c239),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2df52),
	.w1(32'h39a178bc),
	.w2(32'h384f53d9),
	.w3(32'h3a05c141),
	.w4(32'hba350333),
	.w5(32'h38fb7bc8),
	.w6(32'h3960384a),
	.w7(32'hba861511),
	.w8(32'hb9bf7661),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec43a6),
	.w1(32'hb99c92cc),
	.w2(32'hb980415d),
	.w3(32'hb9de7ab0),
	.w4(32'hb8f7aa87),
	.w5(32'hb9764d80),
	.w6(32'hb9828a48),
	.w7(32'hb93592fc),
	.w8(32'hb985d695),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e36e3f),
	.w1(32'hb8ebdd21),
	.w2(32'hb91e37cd),
	.w3(32'h389e61fa),
	.w4(32'h3871099d),
	.w5(32'hb87d854a),
	.w6(32'h393d4702),
	.w7(32'h38959818),
	.w8(32'hb913c1a7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae81bf3),
	.w1(32'h3a514079),
	.w2(32'h3a5ea107),
	.w3(32'h3b10eb68),
	.w4(32'h3af16f89),
	.w5(32'h3ac5b58b),
	.w6(32'h3b2268aa),
	.w7(32'h3af02e9f),
	.w8(32'h3ab1b3b1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaf969),
	.w1(32'h3b812225),
	.w2(32'h3b3daded),
	.w3(32'h3ad78739),
	.w4(32'h3aafe8a4),
	.w5(32'h3a47268a),
	.w6(32'h3a293932),
	.w7(32'hba165a2d),
	.w8(32'hba646994),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68bc52),
	.w1(32'h3b38bce1),
	.w2(32'h3baff9dc),
	.w3(32'h39e5efac),
	.w4(32'hb7c365db),
	.w5(32'h3ac9e255),
	.w6(32'hba213ce7),
	.w7(32'hba8ac498),
	.w8(32'h398656c4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96113e),
	.w1(32'h3b829280),
	.w2(32'h3c0377a9),
	.w3(32'h3a1eb3f2),
	.w4(32'h394cd13d),
	.w5(32'h3b1e665c),
	.w6(32'hba9dc8dd),
	.w7(32'hbb40d581),
	.w8(32'hb9fc578f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83df8d),
	.w1(32'h3b1ac179),
	.w2(32'h3b501924),
	.w3(32'h3b36c488),
	.w4(32'h3ab39219),
	.w5(32'h3abf0ffe),
	.w6(32'h3ae73bd5),
	.w7(32'h3a3cfb17),
	.w8(32'h39e13eef),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0e798),
	.w1(32'h3bdc4d1b),
	.w2(32'h3b1fe082),
	.w3(32'h3b0641c5),
	.w4(32'h3b0d89bb),
	.w5(32'hba85bb4d),
	.w6(32'hba96012c),
	.w7(32'h3a670df5),
	.w8(32'h38d61b61),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a0b1e),
	.w1(32'hb95f8e00),
	.w2(32'hb97e5fc0),
	.w3(32'hb900c071),
	.w4(32'h395fdaef),
	.w5(32'hb933d6a2),
	.w6(32'h372af365),
	.w7(32'h3992d6b0),
	.w8(32'hb9db17ef),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81fc834),
	.w1(32'hb97eeeeb),
	.w2(32'hba339b0b),
	.w3(32'h3a1f9d2a),
	.w4(32'h3900b42a),
	.w5(32'hba80ae74),
	.w6(32'h3a2ac987),
	.w7(32'h385abb88),
	.w8(32'hba8fe2fd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79c16f5),
	.w1(32'h376922e9),
	.w2(32'hb9783178),
	.w3(32'h39befb77),
	.w4(32'h39caa3ea),
	.w5(32'hb96d9b1d),
	.w6(32'h399350b2),
	.w7(32'h3989505a),
	.w8(32'hb95f0734),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b744022),
	.w1(32'h3b5582da),
	.w2(32'h3baa566a),
	.w3(32'h3ad3f438),
	.w4(32'h3ab8ba0b),
	.w5(32'h3b115811),
	.w6(32'hb94197fd),
	.w7(32'hb9fe26f7),
	.w8(32'hb9dabf22),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41fde0),
	.w1(32'h3a3f7102),
	.w2(32'h3adb6146),
	.w3(32'h3984772e),
	.w4(32'h39897044),
	.w5(32'h3a54d6d2),
	.w6(32'hb980f13a),
	.w7(32'hb9f08a15),
	.w8(32'h39e98ca4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf0dad),
	.w1(32'h3b7b4609),
	.w2(32'h3bc7d1ce),
	.w3(32'h38370fca),
	.w4(32'hb8a6b712),
	.w5(32'h3b19da5f),
	.w6(32'hbb1128d6),
	.w7(32'hbb3b8c04),
	.w8(32'hb91e2abe),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f11c91),
	.w1(32'h390d6fa7),
	.w2(32'h3a1d0575),
	.w3(32'h39bb0961),
	.w4(32'hb8e25bfc),
	.w5(32'h39b7f42e),
	.w6(32'h3a160b73),
	.w7(32'h3726a43d),
	.w8(32'h3a0bb50d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375ac116),
	.w1(32'hb88e8198),
	.w2(32'hb92bbcf0),
	.w3(32'h37bf5bbd),
	.w4(32'hb79dfe74),
	.w5(32'hb92b309f),
	.w6(32'h38593aff),
	.w7(32'h38df9129),
	.w8(32'hb8a0c76b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c22404),
	.w1(32'h37f5a13a),
	.w2(32'h3759a7dc),
	.w3(32'h37b3cce5),
	.w4(32'h373a6749),
	.w5(32'h342b696b),
	.w6(32'h370c2c4c),
	.w7(32'h368ac043),
	.w8(32'hb71db941),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f55da),
	.w1(32'h382f5144),
	.w2(32'h382868ab),
	.w3(32'h3795e4f0),
	.w4(32'h3824235b),
	.w5(32'h36f58220),
	.w6(32'h378bdfd3),
	.w7(32'h37fb54f6),
	.w8(32'h369d7a72),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5df2b),
	.w1(32'hb9ba6933),
	.w2(32'h39a9fc1a),
	.w3(32'h39868e4c),
	.w4(32'hb9d1882b),
	.w5(32'h3908ad9c),
	.w6(32'h3a7d4a18),
	.w7(32'h397c3f08),
	.w8(32'h3a026bbe),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3873e16a),
	.w1(32'h39cb5f51),
	.w2(32'h399ed001),
	.w3(32'hb9c70f61),
	.w4(32'h3978a656),
	.w5(32'h38c15efe),
	.w6(32'hb9baaec6),
	.w7(32'h393df591),
	.w8(32'h37b3311d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00b075),
	.w1(32'h3a536244),
	.w2(32'h3b091110),
	.w3(32'h3aa4414a),
	.w4(32'hba6f022b),
	.w5(32'hb9c10af6),
	.w6(32'h3ab923a8),
	.w7(32'hbaf12378),
	.w8(32'hba5b5284),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ef365),
	.w1(32'h39ea85dd),
	.w2(32'h3a565e9c),
	.w3(32'h39dad0ac),
	.w4(32'h3a3ffcf9),
	.w5(32'h39dc301e),
	.w6(32'hba0c7f5c),
	.w7(32'h39e5f271),
	.w8(32'h3a7d4b24),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8db4a12),
	.w1(32'hb8875581),
	.w2(32'hb86ccb0a),
	.w3(32'hb7c99a8a),
	.w4(32'h379040ce),
	.w5(32'hb8209173),
	.w6(32'h345eb702),
	.w7(32'h379384ee),
	.w8(32'hb728c6e5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80be815),
	.w1(32'hb7e69b0d),
	.w2(32'hb8676bd1),
	.w3(32'hb784c7d0),
	.w4(32'hb684a396),
	.w5(32'hb7fd2ddf),
	.w6(32'hb7fa3feb),
	.w7(32'hb58e8b2d),
	.w8(32'hb7a9b5f7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886cdaf),
	.w1(32'h352023b7),
	.w2(32'h390ce62f),
	.w3(32'h372a37a1),
	.w4(32'hb802cc74),
	.w5(32'h390cd9b0),
	.w6(32'hb70163ff),
	.w7(32'hb8384fc2),
	.w8(32'h38eb2fdc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b8c051),
	.w1(32'hb829b209),
	.w2(32'hb7ed388b),
	.w3(32'hb8223a66),
	.w4(32'h3715d70c),
	.w5(32'h372d1ab1),
	.w6(32'hb769bde9),
	.w7(32'h3797c78c),
	.w8(32'h372beec1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae89f91),
	.w1(32'h3a926259),
	.w2(32'h3aec3276),
	.w3(32'h38b3ce19),
	.w4(32'hb9d0ad79),
	.w5(32'h374ce78a),
	.w6(32'h3843b9b7),
	.w7(32'hb9e5b6fc),
	.w8(32'hba5764ec),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cc917),
	.w1(32'h3b847c6f),
	.w2(32'h3c2239cb),
	.w3(32'h39c14737),
	.w4(32'h3a4ed95a),
	.w5(32'h3badf5b5),
	.w6(32'hba81cbf4),
	.w7(32'hbb12bfd8),
	.w8(32'h3aaa39a8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae071c3),
	.w1(32'h3ae76dbc),
	.w2(32'h3bcc5cdf),
	.w3(32'hba2fbc3f),
	.w4(32'hbaf6ed56),
	.w5(32'h3b06682d),
	.w6(32'hba8ba558),
	.w7(32'hbb4f463c),
	.w8(32'h39a9a7a1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb40482),
	.w1(32'h3b3f61ed),
	.w2(32'h3be1607e),
	.w3(32'h3a22c20a),
	.w4(32'hbb571a09),
	.w5(32'hbad072cb),
	.w6(32'hba4756a0),
	.w7(32'hbb690705),
	.w8(32'h3aa99d43),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89bcde1),
	.w1(32'hb7cdc369),
	.w2(32'hb89331d8),
	.w3(32'hb815f8cb),
	.w4(32'h36a36f2b),
	.w5(32'hb80ff714),
	.w6(32'hb7ef09a1),
	.w7(32'h37344cbe),
	.w8(32'hb80325ab),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901c9d8),
	.w1(32'hb87db31b),
	.w2(32'hb8ed2e14),
	.w3(32'hb87a5476),
	.w4(32'h36c72c89),
	.w5(32'hb85d83b0),
	.w6(32'hb86d8746),
	.w7(32'h3722386e),
	.w8(32'hb81d2c82),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8736862),
	.w1(32'hb582bd88),
	.w2(32'hb8fe5ea4),
	.w3(32'hb885612f),
	.w4(32'h37aaf5ab),
	.w5(32'hb8a97215),
	.w6(32'hb707da02),
	.w7(32'h38a4466c),
	.w8(32'hb87020ac),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f2cd7),
	.w1(32'h39889b2e),
	.w2(32'h3aaf81c8),
	.w3(32'h39ca125d),
	.w4(32'hb96d50f8),
	.w5(32'h3a635f01),
	.w6(32'h3a01001a),
	.w7(32'hb9804360),
	.w8(32'h39740b66),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a944e9),
	.w1(32'hb8e2f935),
	.w2(32'hb9212c6d),
	.w3(32'h38bfbcb0),
	.w4(32'h38a98b9b),
	.w5(32'hb8c869c3),
	.w6(32'h3903a414),
	.w7(32'h38cf46ac),
	.w8(32'hb8cdbc63),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adda7e4),
	.w1(32'h3acf7599),
	.w2(32'h3b26e954),
	.w3(32'h38ee9b57),
	.w4(32'hb90b6cce),
	.w5(32'h3a477f2c),
	.w6(32'hba2bdb03),
	.w7(32'hbace222d),
	.w8(32'hba3aa5f4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ac568),
	.w1(32'h3b00a860),
	.w2(32'h3ab8fd37),
	.w3(32'h3a1b9aac),
	.w4(32'hbb2d7dd5),
	.w5(32'hbb4cac78),
	.w6(32'h3aed5880),
	.w7(32'hbac50628),
	.w8(32'hbb358c4a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98fc93),
	.w1(32'h3b572ce2),
	.w2(32'h3b3269c0),
	.w3(32'h3ae61c1a),
	.w4(32'h38ab747b),
	.w5(32'hba93aefc),
	.w6(32'h3853d286),
	.w7(32'hbacbe445),
	.w8(32'hba9ddb47),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34ac76),
	.w1(32'h3b1a5fb4),
	.w2(32'h3b725a5d),
	.w3(32'h39fff2f3),
	.w4(32'h39a98587),
	.w5(32'h3af5b878),
	.w6(32'hb95f4f7e),
	.w7(32'hba4a1144),
	.w8(32'h3a434974),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5ddd3),
	.w1(32'h3ab77ca2),
	.w2(32'h3b0b6647),
	.w3(32'h3a153d2b),
	.w4(32'h3968de73),
	.w5(32'h3a774c5e),
	.w6(32'hba455ed5),
	.w7(32'hbaa08fb4),
	.w8(32'hba1b5d26),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971afce),
	.w1(32'h3849024b),
	.w2(32'h3af283c7),
	.w3(32'hb9c1bb96),
	.w4(32'hba1d4bae),
	.w5(32'h399800ff),
	.w6(32'hba07b0ba),
	.w7(32'hba3d7528),
	.w8(32'hb847d489),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b141d3d),
	.w1(32'h3b0e0615),
	.w2(32'h3b61039e),
	.w3(32'h39a6202c),
	.w4(32'h3a3f4c02),
	.w5(32'h3acd2627),
	.w6(32'hba24cd1e),
	.w7(32'hba63f9a8),
	.w8(32'h39c9cfae),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74257ef),
	.w1(32'hb6e14c7c),
	.w2(32'hb7916ab1),
	.w3(32'hb69e241f),
	.w4(32'h3681cf28),
	.w5(32'hb64169f7),
	.w6(32'hb60a7286),
	.w7(32'h36b9ed2c),
	.w8(32'h34b28d02),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7864e49),
	.w1(32'hb7a8d567),
	.w2(32'hb7eb84c6),
	.w3(32'hb71ccce8),
	.w4(32'hb68c433e),
	.w5(32'hb63366f3),
	.w6(32'hb75a75cd),
	.w7(32'h36143e5b),
	.w8(32'hb7252a8f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75acb5c),
	.w1(32'hb50f5b4d),
	.w2(32'hb7ed2689),
	.w3(32'hb5021b82),
	.w4(32'h36ff8b72),
	.w5(32'hb8005055),
	.w6(32'h37f56b92),
	.w7(32'h36c09a30),
	.w8(32'hb7388ede),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a84478),
	.w1(32'hb643e6ef),
	.w2(32'hb7b240f2),
	.w3(32'hb794d8b1),
	.w4(32'h36b02c04),
	.w5(32'hb6eabbf4),
	.w6(32'h36d07283),
	.w7(32'h375421c1),
	.w8(32'h35e2235f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e4083),
	.w1(32'h3a8f12c8),
	.w2(32'h3abf61d7),
	.w3(32'h3b27554c),
	.w4(32'h3a14e1d8),
	.w5(32'h3b1d57b2),
	.w6(32'h3a7894f1),
	.w7(32'hb849bc91),
	.w8(32'h3a93e746),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b5517),
	.w1(32'hb9ac07ec),
	.w2(32'h398313ba),
	.w3(32'hba16a4ca),
	.w4(32'hba56f0cd),
	.w5(32'hb97abf0f),
	.w6(32'h39e0cb71),
	.w7(32'hba2e5273),
	.w8(32'hb97f84af),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c9d16),
	.w1(32'h3b80b8c1),
	.w2(32'h3ba15053),
	.w3(32'h3a983901),
	.w4(32'h3a60a957),
	.w5(32'h3b1586ab),
	.w6(32'hbaaa0d52),
	.w7(32'hbab7bb75),
	.w8(32'h3a6bb5e5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7b6ff),
	.w1(32'h3bade569),
	.w2(32'h3bad4638),
	.w3(32'h3bd1289c),
	.w4(32'h3b8f3495),
	.w5(32'h3b7b2373),
	.w6(32'h3b981485),
	.w7(32'h3b1b493f),
	.w8(32'h3b4a5181),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7a2a5),
	.w1(32'h3a44abcd),
	.w2(32'h3b685c56),
	.w3(32'h3a8ab6cb),
	.w4(32'h38dbaeb4),
	.w5(32'h3b3f33cb),
	.w6(32'h3b1dc121),
	.w7(32'h3a1c1c65),
	.w8(32'h3b301047),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b227696),
	.w1(32'h3b3b3fc7),
	.w2(32'h3b8aebae),
	.w3(32'h3a5c0416),
	.w4(32'h3a7e8028),
	.w5(32'h3b4c388b),
	.w6(32'h3a52a693),
	.w7(32'hb991d624),
	.w8(32'h3acf7ac5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fa813),
	.w1(32'hb950480d),
	.w2(32'h3b0184fe),
	.w3(32'hbb1805c8),
	.w4(32'hbae940ef),
	.w5(32'h3ab75362),
	.w6(32'hbb4c6ca5),
	.w7(32'hbb5f8289),
	.w8(32'hba954514),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1000b),
	.w1(32'h3b996ed9),
	.w2(32'h3b8f51ba),
	.w3(32'h3b7cc932),
	.w4(32'h3b1779d4),
	.w5(32'h3b6407d8),
	.w6(32'h3aab29b7),
	.w7(32'h3a15bd23),
	.w8(32'h3b3a40c5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45f5d5),
	.w1(32'h3b19ff8a),
	.w2(32'h3b604e65),
	.w3(32'h3aa91a19),
	.w4(32'h3a610f72),
	.w5(32'h3b13250d),
	.w6(32'hba58a2b3),
	.w7(32'hba95d79f),
	.w8(32'h3a8e1b3d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6ee2f),
	.w1(32'h3b0d1a7a),
	.w2(32'h3b3ef1b2),
	.w3(32'h3a2c7429),
	.w4(32'hba79e432),
	.w5(32'h3a23e717),
	.w6(32'hb9591696),
	.w7(32'hbb0a8e02),
	.w8(32'hba3fce67),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fea94c),
	.w1(32'h3a02ab0b),
	.w2(32'hb9c5223f),
	.w3(32'h39e1fe95),
	.w4(32'h3a1356d1),
	.w5(32'hb9b2d35f),
	.w6(32'h39e99f43),
	.w7(32'h39748e02),
	.w8(32'hb9e306bb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8c054),
	.w1(32'h3b9f3a4d),
	.w2(32'h3ba0ad36),
	.w3(32'h3abf1b86),
	.w4(32'h3a1e19f6),
	.w5(32'h38d76ef5),
	.w6(32'hba951869),
	.w7(32'hbac9c70f),
	.w8(32'hba379030),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1b701),
	.w1(32'h3b81bbbb),
	.w2(32'h3bfda15d),
	.w3(32'hbb0c2f07),
	.w4(32'hbb05fb25),
	.w5(32'h3b154b31),
	.w6(32'hbb564c64),
	.w7(32'hbb86554c),
	.w8(32'hbab29b09),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad187e1),
	.w1(32'h3b4c7382),
	.w2(32'h3be6a5a3),
	.w3(32'hbb1ce348),
	.w4(32'hbae78669),
	.w5(32'h3b4b3db4),
	.w6(32'hbaf25a7a),
	.w7(32'hbb7bd4f1),
	.w8(32'h3a79a9fb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb15ba2),
	.w1(32'h3b9039ab),
	.w2(32'h3c061cfc),
	.w3(32'h3bbafc35),
	.w4(32'h3b188c16),
	.w5(32'h3c189ea3),
	.w6(32'h3b71dc58),
	.w7(32'h3b4b650c),
	.w8(32'h3bdd36ae),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f06b1),
	.w1(32'h3b84e392),
	.w2(32'h3b975da2),
	.w3(32'h3a940c47),
	.w4(32'h398a2aa5),
	.w5(32'h39057c7e),
	.w6(32'hbab31622),
	.w7(32'hbaff09f4),
	.w8(32'hba74055c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b41b3),
	.w1(32'h3bbfcf64),
	.w2(32'h3bc9226c),
	.w3(32'h3a8237d0),
	.w4(32'h3b737a49),
	.w5(32'h3b87f82b),
	.w6(32'hbb0abfde),
	.w7(32'h3a0a8423),
	.w8(32'h3b3adf1a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36634f),
	.w1(32'hb92b46ff),
	.w2(32'hba722984),
	.w3(32'h39f5a7ce),
	.w4(32'h3a5c1b5a),
	.w5(32'hba03a8bc),
	.w6(32'h3a0a4b29),
	.w7(32'h3a3fd177),
	.w8(32'hba48cc66),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a5ea8),
	.w1(32'h3bbb66d3),
	.w2(32'h3c07745d),
	.w3(32'h39a82f83),
	.w4(32'hb9e482fc),
	.w5(32'h3b6043d5),
	.w6(32'hba15f67b),
	.w7(32'hbaf90661),
	.w8(32'hb9e8df04),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7f782),
	.w1(32'h3a8e3317),
	.w2(32'h3a996e30),
	.w3(32'h39d9d5aa),
	.w4(32'hbaa87e78),
	.w5(32'hba705506),
	.w6(32'h3a6035ca),
	.w7(32'hbb0d4faf),
	.w8(32'hbae737d7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68b9757),
	.w1(32'h37bb2db8),
	.w2(32'h38adb5fa),
	.w3(32'h372571b5),
	.w4(32'h3729ea46),
	.w5(32'h381cd2ba),
	.w6(32'hb86ac098),
	.w7(32'hb801d645),
	.w8(32'h37b88958),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4a8dd),
	.w1(32'h39ee3167),
	.w2(32'h3a86ad83),
	.w3(32'h3a03233a),
	.w4(32'h39b629db),
	.w5(32'h3a40bb1d),
	.w6(32'h39b7885c),
	.w7(32'h39869d13),
	.w8(32'h39c00bee),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba17d99),
	.w1(32'h3b6b7f92),
	.w2(32'hb702b340),
	.w3(32'h3b18f0bf),
	.w4(32'h3abaf53f),
	.w5(32'hba947f60),
	.w6(32'h3a40a553),
	.w7(32'h3a8d0fac),
	.w8(32'hba14715d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed9dbb),
	.w1(32'h3aebebc1),
	.w2(32'h3b112472),
	.w3(32'hb8ce9213),
	.w4(32'h39ebe5ff),
	.w5(32'hba316a75),
	.w6(32'hba0f83aa),
	.w7(32'hba51b875),
	.w8(32'hbb058874),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fd24d),
	.w1(32'h3b5200e0),
	.w2(32'h3b0dd057),
	.w3(32'h3b025d61),
	.w4(32'h3b00ed47),
	.w5(32'h3b1c833e),
	.w6(32'h398814f2),
	.w7(32'h3abfb8ea),
	.w8(32'h3b469bf8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af599f6),
	.w1(32'h3b45adf6),
	.w2(32'h3b2a8df3),
	.w3(32'h38b25d48),
	.w4(32'h3a2a37ad),
	.w5(32'h3a8e2bf3),
	.w6(32'hba725df2),
	.w7(32'h396259fb),
	.w8(32'h39f8623a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6938c7),
	.w1(32'hb95018a1),
	.w2(32'h3ac3efa4),
	.w3(32'hb81c1479),
	.w4(32'hba61c429),
	.w5(32'h3a78b9da),
	.w6(32'h3a596f27),
	.w7(32'hb9ca3bbc),
	.w8(32'h3a9e2ca4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe4be0),
	.w1(32'h3af089d5),
	.w2(32'h3b47520a),
	.w3(32'hb9106c68),
	.w4(32'h39dcaffa),
	.w5(32'h3ac32d94),
	.w6(32'hba9308de),
	.w7(32'hba86d91f),
	.w8(32'hba06d6f4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00ec66),
	.w1(32'h3a965904),
	.w2(32'h3adf2ce1),
	.w3(32'h3a56817e),
	.w4(32'h3977d43a),
	.w5(32'h399d7838),
	.w6(32'h39840c2d),
	.w7(32'hb9293750),
	.w8(32'hb84e927d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c76a0d),
	.w1(32'hb81b3c4a),
	.w2(32'hb7a81810),
	.w3(32'hb87b440e),
	.w4(32'h36b59206),
	.w5(32'hb799f173),
	.w6(32'hb8bbce7b),
	.w7(32'hb7e549bf),
	.w8(32'hb82ff1e2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b32f68),
	.w1(32'hb72334a4),
	.w2(32'hb7fdb088),
	.w3(32'hb7304bbc),
	.w4(32'h3727a2a2),
	.w5(32'hb69fb954),
	.w6(32'hb7625e66),
	.w7(32'h37227e3c),
	.w8(32'hb6c6e3e7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37212aeb),
	.w1(32'hb8cf95fb),
	.w2(32'h36efff4d),
	.w3(32'hb908eac0),
	.w4(32'hb8fa9fa5),
	.w5(32'h38cf0958),
	.w6(32'hb8bd6976),
	.w7(32'hb9071eac),
	.w8(32'hb8634f64),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fce255),
	.w1(32'hb8b0fa0d),
	.w2(32'h38a7676e),
	.w3(32'h38320d2c),
	.w4(32'h388e0a6e),
	.w5(32'h38f671bf),
	.w6(32'hb7cc27b7),
	.w7(32'hb88ec82c),
	.w8(32'hb808299e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e78c0),
	.w1(32'h3ab8108a),
	.w2(32'h3b7055ae),
	.w3(32'h39b7a3a1),
	.w4(32'hb99261ca),
	.w5(32'h3a1faffe),
	.w6(32'hba25257b),
	.w7(32'hbad31a34),
	.w8(32'hb9ec379c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd7f59),
	.w1(32'h396abd7e),
	.w2(32'h3a26d82a),
	.w3(32'hb9617a42),
	.w4(32'h39737f91),
	.w5(32'h3a3fa651),
	.w6(32'hb8fd063e),
	.w7(32'h3917f5ba),
	.w8(32'h39e5d431),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbb121),
	.w1(32'h3acc6025),
	.w2(32'h3acc2785),
	.w3(32'h39a04c64),
	.w4(32'hb911ec6f),
	.w5(32'h38f3cc82),
	.w6(32'hb8b2d9be),
	.w7(32'hba0965e2),
	.w8(32'h39a3f966),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb85a8),
	.w1(32'h3b748045),
	.w2(32'h3b02a815),
	.w3(32'h3b632abd),
	.w4(32'h3a32744d),
	.w5(32'h3915b116),
	.w6(32'h3b397535),
	.w7(32'h39fabd68),
	.w8(32'h3a882590),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b1d197),
	.w1(32'hb7d6b91c),
	.w2(32'hb8ca839c),
	.w3(32'hb8ca082e),
	.w4(32'hb90bac7b),
	.w5(32'hb8d40594),
	.w6(32'hb92a5e81),
	.w7(32'hb951ce7f),
	.w8(32'hb93bba71),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1a8f2),
	.w1(32'hb8fde402),
	.w2(32'h386d1918),
	.w3(32'hb9b2a123),
	.w4(32'hb94caaa6),
	.w5(32'hb855e416),
	.w6(32'hb906bf04),
	.w7(32'hb90ebd35),
	.w8(32'h38be995d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7969a31),
	.w1(32'hb70811d1),
	.w2(32'h375d9e96),
	.w3(32'h35f09a8f),
	.w4(32'h370bb1df),
	.w5(32'h3807e3bd),
	.w6(32'h37700526),
	.w7(32'h376145a1),
	.w8(32'h38003613),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4935d),
	.w1(32'h3ad29b36),
	.w2(32'h39e708a7),
	.w3(32'h3a650502),
	.w4(32'h3a896ea5),
	.w5(32'h39227bbd),
	.w6(32'hb8846044),
	.w7(32'h3a09547c),
	.w8(32'h3939df00),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a239120),
	.w1(32'hb8e94244),
	.w2(32'h3b44030d),
	.w3(32'hbaa97a1a),
	.w4(32'hbaaf691c),
	.w5(32'h3a9efc0f),
	.w6(32'hbafb8abc),
	.w7(32'hbb1fedb8),
	.w8(32'hba58647b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6feda0),
	.w1(32'h3b381f0e),
	.w2(32'h3b9c79e6),
	.w3(32'h3824ef94),
	.w4(32'hb921a24a),
	.w5(32'h3aef7e10),
	.w6(32'hbb145c65),
	.w7(32'hbab6d2ea),
	.w8(32'h3a93dd19),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79044ad),
	.w1(32'hb7969c30),
	.w2(32'hb7625f8d),
	.w3(32'hb6be11ef),
	.w4(32'hb695913d),
	.w5(32'hb5e31e89),
	.w6(32'hb6594ce1),
	.w7(32'h36c2d47e),
	.w8(32'h36b1c5c3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0ed62),
	.w1(32'hb9156245),
	.w2(32'h3a9e966c),
	.w3(32'hba20e4a4),
	.w4(32'hba8aa803),
	.w5(32'h38bca0c7),
	.w6(32'hb8c39beb),
	.w7(32'hb93a614d),
	.w8(32'h3a370a0b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3c0d7),
	.w1(32'h3a7fe03d),
	.w2(32'h3b023031),
	.w3(32'h3a9ed7b9),
	.w4(32'h39deff39),
	.w5(32'h3ab00d1d),
	.w6(32'h3a8112e2),
	.w7(32'hba2926ba),
	.w8(32'h395c223f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b50ac),
	.w1(32'h3a3cb550),
	.w2(32'h3aadab4f),
	.w3(32'hb8366c79),
	.w4(32'hb9808bdf),
	.w5(32'h39d1e6a0),
	.w6(32'hb8823fa1),
	.w7(32'hb9a41434),
	.w8(32'h399926f0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03aa9b),
	.w1(32'h3a5e32d6),
	.w2(32'h3b72cc14),
	.w3(32'h39f6df09),
	.w4(32'h38ad5c76),
	.w5(32'h3b2c1c94),
	.w6(32'h396edae6),
	.w7(32'hb9cc3e9d),
	.w8(32'h3b1aac09),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b982bf8),
	.w1(32'h3b8bd9f9),
	.w2(32'h3bc33e3b),
	.w3(32'h393aab8c),
	.w4(32'h39008b23),
	.w5(32'h3b01c8d2),
	.w6(32'hbacddb44),
	.w7(32'hbb6a1988),
	.w8(32'hba89ab64),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c6797),
	.w1(32'h3b1a7fed),
	.w2(32'h398e35dd),
	.w3(32'h3ac1df91),
	.w4(32'h3ab527a3),
	.w5(32'h3a05bb63),
	.w6(32'h3a27124a),
	.w7(32'h3aa9b206),
	.w8(32'h3a651866),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b90a2),
	.w1(32'h3b9c0e25),
	.w2(32'h3ba4dbe4),
	.w3(32'h3add0b68),
	.w4(32'h3a369973),
	.w5(32'h3951c186),
	.w6(32'hbb08620c),
	.w7(32'hba85977b),
	.w8(32'h39bb3861),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badb064),
	.w1(32'h3b9c7bc1),
	.w2(32'h3be0844b),
	.w3(32'h3b143ca3),
	.w4(32'h3afabb8c),
	.w5(32'h3ba891ef),
	.w6(32'h39e455b4),
	.w7(32'hb9a28ba7),
	.w8(32'h3b492988),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41b310),
	.w1(32'h3ad43818),
	.w2(32'h3ac288da),
	.w3(32'h3addcc88),
	.w4(32'h3a8104b5),
	.w5(32'h3a3b5ab1),
	.w6(32'h3a4ca1b3),
	.w7(32'h3a088188),
	.w8(32'h3a55f016),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50720d),
	.w1(32'h3b2f166e),
	.w2(32'h3ab051ac),
	.w3(32'h3af1aa3e),
	.w4(32'h3abe0a69),
	.w5(32'h39ed8804),
	.w6(32'hb9efe67e),
	.w7(32'h3909c593),
	.w8(32'h3a3794c6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bf89b),
	.w1(32'h3a0b5bd1),
	.w2(32'h3a951b05),
	.w3(32'hb99956eb),
	.w4(32'hb9be225b),
	.w5(32'h38e69186),
	.w6(32'hba12352f),
	.w7(32'hba241c89),
	.w8(32'hb9316143),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdafdd7),
	.w1(32'h3b9085be),
	.w2(32'h3b07c828),
	.w3(32'h3b64ae97),
	.w4(32'h3ad89f32),
	.w5(32'h3a588cbc),
	.w6(32'h3992ad4e),
	.w7(32'hb99f5209),
	.w8(32'h3aaa7b99),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7e411),
	.w1(32'h3ab72671),
	.w2(32'h3b1424ea),
	.w3(32'h39fbc0d4),
	.w4(32'h3a032c92),
	.w5(32'h3b13a378),
	.w6(32'hb9edab0a),
	.w7(32'hba709971),
	.w8(32'h3a7bceb2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75fed0f),
	.w1(32'hb7051b4e),
	.w2(32'hb6b29ab8),
	.w3(32'hb59a0ff1),
	.w4(32'h377074ef),
	.w5(32'h375be1bd),
	.w6(32'h35f4127c),
	.w7(32'h372a9d6d),
	.w8(32'h3781e65a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6da82a9),
	.w1(32'hb77c1475),
	.w2(32'hb705eece),
	.w3(32'hb6c58c38),
	.w4(32'hb78d6231),
	.w5(32'hb7a74c60),
	.w6(32'hb717ec66),
	.w7(32'hb7073fd6),
	.w8(32'hb463bc9f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac32ce9),
	.w1(32'h39f88389),
	.w2(32'h37d24687),
	.w3(32'h3a710305),
	.w4(32'hba2fda01),
	.w5(32'hba9b3540),
	.w6(32'h3a09b7bb),
	.w7(32'hb9edfba5),
	.w8(32'hba74f7df),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baecd71),
	.w1(32'h3b89d272),
	.w2(32'h3afcf14c),
	.w3(32'h3ae4aca1),
	.w4(32'h3a4a61fa),
	.w5(32'h3ab56c23),
	.w6(32'h3a3d7be0),
	.w7(32'hb9f8ed28),
	.w8(32'h38caaf80),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb2ad5),
	.w1(32'h3b56d083),
	.w2(32'h3bb9b47a),
	.w3(32'h39e42cb3),
	.w4(32'hbaf4baa2),
	.w5(32'h3984dfed),
	.w6(32'h3930b817),
	.w7(32'hbb3dc43f),
	.w8(32'hba6fc0e7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82680db),
	.w1(32'hb7c0a85c),
	.w2(32'hb7b08deb),
	.w3(32'hb79b9156),
	.w4(32'hb78ebe85),
	.w5(32'hb804db31),
	.w6(32'hb6142dd2),
	.w7(32'hb7a5f3a1),
	.w8(32'hb7f2136b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b862c5a),
	.w1(32'h3b4367f7),
	.w2(32'h3b8470e4),
	.w3(32'h3a9db216),
	.w4(32'h3959c9e2),
	.w5(32'h3ab03b5a),
	.w6(32'hba602905),
	.w7(32'hbaa97738),
	.w8(32'hb9a9a9ff),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e7740),
	.w1(32'h3b2b2eec),
	.w2(32'h3acf47dc),
	.w3(32'h3b025d6b),
	.w4(32'h39a87545),
	.w5(32'hba198553),
	.w6(32'h39835770),
	.w7(32'hba361a9f),
	.w8(32'hba8183fd),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d6332),
	.w1(32'h3b6b7ad5),
	.w2(32'h3b52d497),
	.w3(32'h3af49fa7),
	.w4(32'h3a8c2312),
	.w5(32'h3956223c),
	.w6(32'hb9d53658),
	.w7(32'hba6fe457),
	.w8(32'hb9c7132f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c14d16),
	.w1(32'h3a34f08b),
	.w2(32'h3b63dcd7),
	.w3(32'hbab63a7e),
	.w4(32'hbb2c83f7),
	.w5(32'h3a88988d),
	.w6(32'hbb1dff39),
	.w7(32'hbb8d1ff1),
	.w8(32'hbabcf7aa),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d13c6),
	.w1(32'h39379b65),
	.w2(32'h3ae3d9d1),
	.w3(32'h3ac7bbca),
	.w4(32'h39ac5733),
	.w5(32'h3ada929d),
	.w6(32'h3ad67c6e),
	.w7(32'h397295d3),
	.w8(32'h39b0c75d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9374052),
	.w1(32'hba18c12e),
	.w2(32'hba21500f),
	.w3(32'h39c782a4),
	.w4(32'h3a13f2ae),
	.w5(32'h3981cff7),
	.w6(32'h3a3d845c),
	.w7(32'h39e428c3),
	.w8(32'h39446cca),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5f8e3),
	.w1(32'hb906a865),
	.w2(32'hba67f089),
	.w3(32'h3ab278ca),
	.w4(32'hb95afd86),
	.w5(32'hba9b34fa),
	.w6(32'h3aef05a0),
	.w7(32'h3a53e27b),
	.w8(32'hba648da9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51de20),
	.w1(32'h3ac61e99),
	.w2(32'h3b951295),
	.w3(32'h3aca1745),
	.w4(32'h39b30eaf),
	.w5(32'h3bb15bac),
	.w6(32'h3a94236f),
	.w7(32'hb928ed78),
	.w8(32'h3b5e5a7d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993100d),
	.w1(32'hbab64d80),
	.w2(32'h3a62b813),
	.w3(32'hb908b77f),
	.w4(32'hbad1ceef),
	.w5(32'h3a07767c),
	.w6(32'h3a9d0adb),
	.w7(32'hb9dcb773),
	.w8(32'h3a1c9b5c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3c15d),
	.w1(32'h39eedcfd),
	.w2(32'h3a495822),
	.w3(32'h381dfd42),
	.w4(32'h39ac2690),
	.w5(32'h3a2f7fa5),
	.w6(32'hb8f7955e),
	.w7(32'hb99b974d),
	.w8(32'hb8c9d272),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a997f),
	.w1(32'h398e98f6),
	.w2(32'h3909e9f1),
	.w3(32'h395cc74a),
	.w4(32'h39ddef0c),
	.w5(32'h396264fe),
	.w6(32'h394c6725),
	.w7(32'h39e5a37a),
	.w8(32'h39bfa860),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b254726),
	.w1(32'h3b1939e0),
	.w2(32'h3b11836b),
	.w3(32'h3a24703c),
	.w4(32'h38981b7d),
	.w5(32'h3a959f18),
	.w6(32'hba7b7129),
	.w7(32'hba9a1ecb),
	.w8(32'h3a111def),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74fa5a3),
	.w1(32'h378f272f),
	.w2(32'h382476b5),
	.w3(32'h35b8d958),
	.w4(32'h37f7759f),
	.w5(32'h3891461c),
	.w6(32'h373a6189),
	.w7(32'h37d33bc5),
	.w8(32'h38838d34),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac151cc),
	.w1(32'h3a8f5a3a),
	.w2(32'h3abb365d),
	.w3(32'hb9332470),
	.w4(32'h39afed9e),
	.w5(32'h3a031c68),
	.w6(32'hba127ea4),
	.w7(32'hba133416),
	.w8(32'hb96c5901),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9405d51),
	.w1(32'hb9059b39),
	.w2(32'h3977abbf),
	.w3(32'hb9e22d9a),
	.w4(32'hb9976241),
	.w5(32'h39321495),
	.w6(32'hb996a079),
	.w7(32'h38180834),
	.w8(32'h39010bf9),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cd829),
	.w1(32'hbb774990),
	.w2(32'h393706ce),
	.w3(32'hbb1763ec),
	.w4(32'hbbb3c5a1),
	.w5(32'hbb5c274f),
	.w6(32'h388e7eab),
	.w7(32'hbb7acd88),
	.w8(32'hbb21ebf9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907625f),
	.w1(32'h37000ca3),
	.w2(32'hb55e2b12),
	.w3(32'hb8d23256),
	.w4(32'h38a360c0),
	.w5(32'h37bfe0b7),
	.w6(32'hb908958e),
	.w7(32'h38281b52),
	.w8(32'hb7f442e5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3585aeba),
	.w1(32'hb91becd4),
	.w2(32'hb93d95a3),
	.w3(32'h384c500c),
	.w4(32'hb8a5106f),
	.w5(32'h38429711),
	.w6(32'h38e43b44),
	.w7(32'h36ddb632),
	.w8(32'h3968432d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46d366),
	.w1(32'h3b4586b6),
	.w2(32'h3a209ee4),
	.w3(32'h3accf42c),
	.w4(32'h3b6770bc),
	.w5(32'h3b26f770),
	.w6(32'hba11c5b9),
	.w7(32'h3b3cabb6),
	.w8(32'h3b005cb6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b817ba1),
	.w1(32'h3b4abe72),
	.w2(32'h3bec020f),
	.w3(32'h3afec410),
	.w4(32'h3ae4bb9b),
	.w5(32'h3b9548e4),
	.w6(32'hb98d24cd),
	.w7(32'hb9399abb),
	.w8(32'h3a3e4998),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18541d),
	.w1(32'hba34aaae),
	.w2(32'h3a7d46e5),
	.w3(32'h3a4b26cd),
	.w4(32'hba333d78),
	.w5(32'h3a016024),
	.w6(32'h3b0df700),
	.w7(32'h37f4d6c2),
	.w8(32'h3a2b1e9e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b6545),
	.w1(32'h3b2c606a),
	.w2(32'h3b289b96),
	.w3(32'h3acd72d9),
	.w4(32'h3a2f362b),
	.w5(32'h39ccb26e),
	.w6(32'h39f72103),
	.w7(32'h3a49334b),
	.w8(32'h3a9585b5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86d749),
	.w1(32'h3a366fe4),
	.w2(32'h39c5c5ec),
	.w3(32'h39de2778),
	.w4(32'h391a14b9),
	.w5(32'h3955ab79),
	.w6(32'h391b1c0b),
	.w7(32'h39177e20),
	.w8(32'h39dd4d1e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcf241),
	.w1(32'h3bd02ccf),
	.w2(32'h3c22acb4),
	.w3(32'h39ce93bb),
	.w4(32'hbae286ac),
	.w5(32'h3b6a9e5d),
	.w6(32'hbb3f79b1),
	.w7(32'hbbd88810),
	.w8(32'hb980bb87),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b437f67),
	.w1(32'h3abe1f4e),
	.w2(32'h3b69d74c),
	.w3(32'h3a8359bf),
	.w4(32'hba72e325),
	.w5(32'h3ab461a4),
	.w6(32'h3a0fc8dc),
	.w7(32'hbb067202),
	.w8(32'h398e37fb),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081912),
	.w1(32'h3b464529),
	.w2(32'h3bd3693c),
	.w3(32'hb9c6d265),
	.w4(32'h3a4b8dd7),
	.w5(32'h3b0b885a),
	.w6(32'hbadd826c),
	.w7(32'hba791243),
	.w8(32'h397742f8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e8bc8a),
	.w1(32'hb8cebf10),
	.w2(32'h37c726ff),
	.w3(32'hb885306d),
	.w4(32'h3907f0e9),
	.w5(32'h39692e22),
	.w6(32'hb7c1c9dd),
	.w7(32'h399ce027),
	.w8(32'h39cd8f6b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36aabe),
	.w1(32'h3b4da2ad),
	.w2(32'h3b7ae351),
	.w3(32'h3a3ee3dc),
	.w4(32'h3aa387cb),
	.w5(32'h3b309558),
	.w6(32'hbafcc99d),
	.w7(32'hb9c729f4),
	.w8(32'h3ade4ea1),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cdd841),
	.w1(32'hb811b866),
	.w2(32'hb842ea9c),
	.w3(32'hb7e8d3c9),
	.w4(32'hb7ff5de0),
	.w5(32'hb80ea07b),
	.w6(32'hb7fb5489),
	.w7(32'hb7b1736f),
	.w8(32'hb7c71998),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba593c6a),
	.w1(32'h39c4314c),
	.w2(32'h3ab852b5),
	.w3(32'hba2d88e5),
	.w4(32'h393921a2),
	.w5(32'h37ad0714),
	.w6(32'hba848c94),
	.w7(32'hb90eb925),
	.w8(32'hb89c0fc0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39918b97),
	.w1(32'hba140187),
	.w2(32'hb9455ef3),
	.w3(32'hb8c0eb2e),
	.w4(32'hba00df85),
	.w5(32'hb79b9bfc),
	.w6(32'h3743fb18),
	.w7(32'hb9a79e05),
	.w8(32'hb9098583),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37129d),
	.w1(32'h3b244aac),
	.w2(32'h3b518b03),
	.w3(32'h3ad46a79),
	.w4(32'h39d23541),
	.w5(32'h3a9eb222),
	.w6(32'h3a540ada),
	.w7(32'hba973a13),
	.w8(32'h393a1ec3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80d6c45),
	.w1(32'hb71e0902),
	.w2(32'hb7239a01),
	.w3(32'hb7c31db9),
	.w4(32'hb5a7fb31),
	.w5(32'hb6c3767b),
	.w6(32'hb7c0ca51),
	.w7(32'hb60c1aa4),
	.w8(32'hb767d16a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ea3ed3),
	.w1(32'hb8821e86),
	.w2(32'hb7da596f),
	.w3(32'hb7fbf489),
	.w4(32'h38368645),
	.w5(32'hb7c48aff),
	.w6(32'h37f481fb),
	.w7(32'h3889c8bc),
	.w8(32'hb7e1b8dd),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a87b7e),
	.w1(32'hba0b68de),
	.w2(32'hb90b7508),
	.w3(32'h3988ea9a),
	.w4(32'hba32a946),
	.w5(32'hb99c06c8),
	.w6(32'h3a4f9438),
	.w7(32'hb9734952),
	.w8(32'hb9676b02),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11d320),
	.w1(32'h3b912166),
	.w2(32'h3b8c4043),
	.w3(32'h399c8085),
	.w4(32'h3ac084a6),
	.w5(32'h3b1a4d3f),
	.w6(32'hba30db2e),
	.w7(32'hba4a03bf),
	.w8(32'h3a65312b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc1e54),
	.w1(32'hb88d214e),
	.w2(32'h381aa60c),
	.w3(32'hb9062d24),
	.w4(32'hb891d019),
	.w5(32'h3888ad4f),
	.w6(32'hb8adad3d),
	.w7(32'hb8420fcf),
	.w8(32'h37ed8e8d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39166d38),
	.w1(32'h399ef069),
	.w2(32'h3a974b39),
	.w3(32'h3825e713),
	.w4(32'hb8ea0f09),
	.w5(32'h3a2f2015),
	.w6(32'h38b753be),
	.w7(32'hb9ad6e52),
	.w8(32'h3988d1e8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d0870),
	.w1(32'h3be6cf9d),
	.w2(32'h3be16949),
	.w3(32'h3b7e9567),
	.w4(32'hbb040ff9),
	.w5(32'hbba94aa7),
	.w6(32'h3a86c255),
	.w7(32'hbbd972dd),
	.w8(32'hbbcb021e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2d718),
	.w1(32'h3aa1206d),
	.w2(32'h3b70ca3c),
	.w3(32'h3b83d3e5),
	.w4(32'h3af529f5),
	.w5(32'h3ba8a73d),
	.w6(32'h3aa32b9b),
	.w7(32'h3afce42a),
	.w8(32'h3b8b82d3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37de65c9),
	.w1(32'h38601a73),
	.w2(32'hb6b2f39f),
	.w3(32'hb857b930),
	.w4(32'h38930fad),
	.w5(32'h37a0025d),
	.w6(32'hb7097f94),
	.w7(32'h39441ecb),
	.w8(32'h391ba29e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d3d89),
	.w1(32'hb8154005),
	.w2(32'hb55f8445),
	.w3(32'hb78788e6),
	.w4(32'hb708f51f),
	.w5(32'h379102b0),
	.w6(32'hb7116a68),
	.w7(32'hb6e1b035),
	.w8(32'h3795f08c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9104b56),
	.w1(32'hb7bf21d9),
	.w2(32'h37905a4e),
	.w3(32'h375f97f1),
	.w4(32'h39aa4cc2),
	.w5(32'h38c04c9e),
	.w6(32'h394af73c),
	.w7(32'h39c05b8e),
	.w8(32'h389b6ca9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a4c431),
	.w1(32'h35148f1a),
	.w2(32'hb7bce741),
	.w3(32'h36c73080),
	.w4(32'hb513ee85),
	.w5(32'hb754ce55),
	.w6(32'hb6869dae),
	.w7(32'hb7624838),
	.w8(32'hb6c698d5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9617b2),
	.w1(32'h3accdbbe),
	.w2(32'h3a854a23),
	.w3(32'h38bc2425),
	.w4(32'h3a5a01f2),
	.w5(32'h3a201ebd),
	.w6(32'hba017754),
	.w7(32'h399f4902),
	.w8(32'h3a088456),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c8e17),
	.w1(32'h3b6a6c4f),
	.w2(32'h3bba35e0),
	.w3(32'h3a21cb73),
	.w4(32'h39b02f88),
	.w5(32'h3b9b22a3),
	.w6(32'hba0f4d72),
	.w7(32'hbb1be97a),
	.w8(32'h3a46493c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89eea8),
	.w1(32'h3b21cfad),
	.w2(32'h3b372c25),
	.w3(32'h39bcd86e),
	.w4(32'hbab2190f),
	.w5(32'h3a548f11),
	.w6(32'hb8b1e46b),
	.w7(32'hbb0eca73),
	.w8(32'hb9395e16),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22ef45),
	.w1(32'h39e212e3),
	.w2(32'h3a0fa880),
	.w3(32'h39c5afcc),
	.w4(32'h398b5a8e),
	.w5(32'h399a7023),
	.w6(32'h39b6f800),
	.w7(32'h39118f6c),
	.w8(32'h390b0ce5),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbb294),
	.w1(32'h3bb966b2),
	.w2(32'h3b8c71dc),
	.w3(32'h3b0b5f2b),
	.w4(32'h3b0c002e),
	.w5(32'h3a858d51),
	.w6(32'h39711022),
	.w7(32'hb9c4eddc),
	.w8(32'h3a48dd24),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a4a11),
	.w1(32'h39e17ad0),
	.w2(32'h3a87d80d),
	.w3(32'hb9e236c6),
	.w4(32'hba8063bb),
	.w5(32'hb9a9df7d),
	.w6(32'h3841506e),
	.w7(32'hbaa9eb04),
	.w8(32'hba84f549),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ed588),
	.w1(32'hb7ff79d0),
	.w2(32'hb827b7d4),
	.w3(32'hb838998a),
	.w4(32'hb4c14a35),
	.w5(32'hb73ff667),
	.w6(32'hb81d3386),
	.w7(32'h360dba1a),
	.w8(32'hb72e4eae),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f03928),
	.w1(32'hb85f58de),
	.w2(32'hb806157c),
	.w3(32'hb8edd49a),
	.w4(32'hb8bbd6fb),
	.w5(32'hb8f9cb20),
	.w6(32'hb8b94fe8),
	.w7(32'hb90aee9a),
	.w8(32'hb92d4123),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90cd183),
	.w1(32'hb8d0b700),
	.w2(32'hb8fd1718),
	.w3(32'hb815ff82),
	.w4(32'h36b39902),
	.w5(32'hb822bcd4),
	.w6(32'hb822f687),
	.w7(32'h373b983a),
	.w8(32'hb7f9344b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b816ba8),
	.w1(32'h3a522c48),
	.w2(32'h3956326e),
	.w3(32'hba0514c1),
	.w4(32'hbac8d165),
	.w5(32'hbb0adf1b),
	.w6(32'hba3ad2f4),
	.w7(32'hbb122e1e),
	.w8(32'hbb976c93),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6624ea),
	.w1(32'hbb1eb0b1),
	.w2(32'h3b488646),
	.w3(32'h3aa5f01e),
	.w4(32'hbb1b3cc3),
	.w5(32'h3b54588b),
	.w6(32'h3a788970),
	.w7(32'hbb033c6d),
	.w8(32'h3a4ec7dd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7522f9),
	.w1(32'h3b1cbe18),
	.w2(32'h3af658b4),
	.w3(32'h3b001013),
	.w4(32'h3a742950),
	.w5(32'h3a38f602),
	.w6(32'h3a379c0e),
	.w7(32'h3a34a33f),
	.w8(32'h3a95b1eb),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbba0e),
	.w1(32'h392b2aca),
	.w2(32'h3a1b0d2c),
	.w3(32'h3a3d1170),
	.w4(32'h391d416d),
	.w5(32'h3a3e031c),
	.w6(32'h3aadee68),
	.w7(32'h3a2373ef),
	.w8(32'h39bf2731),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc79260),
	.w1(32'h3b88f790),
	.w2(32'h3b159ffd),
	.w3(32'h3b39bf56),
	.w4(32'h3b145d63),
	.w5(32'h3ae5ebca),
	.w6(32'h3aee6f6c),
	.w7(32'h3aa2ae52),
	.w8(32'h3adba552),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b098804),
	.w1(32'h3acb6e3a),
	.w2(32'h3aefb349),
	.w3(32'h3922c610),
	.w4(32'hb8309141),
	.w5(32'h3998866c),
	.w6(32'hb9c969f9),
	.w7(32'hba53b68d),
	.w8(32'hb9e12f9d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74dcc1),
	.w1(32'h3add86c1),
	.w2(32'h3be52d68),
	.w3(32'hb9e3fad5),
	.w4(32'hbbb493d7),
	.w5(32'hba8f74ba),
	.w6(32'hba7953c0),
	.w7(32'hbbf8690d),
	.w8(32'hbb41f9ba),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c9e2ed),
	.w1(32'h37a0be6a),
	.w2(32'h369bd661),
	.w3(32'h37d41f62),
	.w4(32'h37c86307),
	.w5(32'h37e21030),
	.w6(32'h37aa285d),
	.w7(32'h37dccf67),
	.w8(32'h383e4d87),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7df2c25),
	.w1(32'hb7f3b699),
	.w2(32'hb7b62e03),
	.w3(32'hb80cc0c7),
	.w4(32'hb80bc7c9),
	.w5(32'hb75711ab),
	.w6(32'hb697025a),
	.w7(32'hb787a703),
	.w8(32'hb70685f9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71b3fa),
	.w1(32'h3ab5156c),
	.w2(32'h3bb4a467),
	.w3(32'hba00a8a3),
	.w4(32'hba42684b),
	.w5(32'h3b1d66dd),
	.w6(32'hbab85ce5),
	.w7(32'hbb28e7c7),
	.w8(32'h3a84a810),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b530948),
	.w1(32'h3b3183e6),
	.w2(32'h3bf0f20a),
	.w3(32'h3a66e71e),
	.w4(32'h3a97e558),
	.w5(32'h3b83451b),
	.w6(32'hbab37d63),
	.w7(32'hbadc8292),
	.w8(32'h3a44c489),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b884e2d),
	.w1(32'h3b4ea1f6),
	.w2(32'h3b79b1db),
	.w3(32'h3a8a0f84),
	.w4(32'hb9c0cb06),
	.w5(32'h3a820c65),
	.w6(32'hb9e18aaf),
	.w7(32'hbad52f93),
	.w8(32'hb87aa078),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8992436),
	.w1(32'hb889a1e7),
	.w2(32'hb7dd831b),
	.w3(32'hb8dd4b2c),
	.w4(32'hb8a1c81d),
	.w5(32'hb83ccbd8),
	.w6(32'hb7d6be3a),
	.w7(32'hb770c949),
	.w8(32'h35bcf9c3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83890c3),
	.w1(32'hb87132b8),
	.w2(32'hb875ec3e),
	.w3(32'hb8905fcf),
	.w4(32'hb6cfd652),
	.w5(32'hb81c85ad),
	.w6(32'hb831e03c),
	.w7(32'hb77cd80a),
	.w8(32'hb7be6df1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c88e1),
	.w1(32'hb8eba382),
	.w2(32'hb91d41ad),
	.w3(32'hb7b5197e),
	.w4(32'hb91737cd),
	.w5(32'hb954f4e1),
	.w6(32'hb7fbada7),
	.w7(32'hb8bb4ee3),
	.w8(32'hb9162f67),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e7261),
	.w1(32'hb929dc0f),
	.w2(32'h3997d4ff),
	.w3(32'hba04a42a),
	.w4(32'hba36f200),
	.w5(32'hb9aa4649),
	.w6(32'h3937908c),
	.w7(32'hba31a8cb),
	.w8(32'hba171cf8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c3c61),
	.w1(32'h3af6b90a),
	.w2(32'h3b45bb69),
	.w3(32'hba31b9f6),
	.w4(32'hbbb9f23b),
	.w5(32'hbb33a873),
	.w6(32'hb93ad157),
	.w7(32'hbc00610e),
	.w8(32'hbb90e9db),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bd256),
	.w1(32'h3b9a6ba7),
	.w2(32'h3b57368c),
	.w3(32'h3af337ff),
	.w4(32'h3b40659d),
	.w5(32'h3afed717),
	.w6(32'hba5dd0aa),
	.w7(32'h38ab7e5f),
	.w8(32'h3abc46c2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d44da),
	.w1(32'h3a102bcf),
	.w2(32'h3b4c4e69),
	.w3(32'hb9e4fe8e),
	.w4(32'hba17af81),
	.w5(32'h3b17e30e),
	.w6(32'h38d12b45),
	.w7(32'hbaa01776),
	.w8(32'h3ab6db36),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b186de0),
	.w1(32'h3b43bdf1),
	.w2(32'h3b5c8774),
	.w3(32'h3b10e9b3),
	.w4(32'h3af8053e),
	.w5(32'h3ae2571c),
	.w6(32'h3af1630e),
	.w7(32'h3ace6ae7),
	.w8(32'h3b0bba6f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb786fe05),
	.w1(32'hb6f07577),
	.w2(32'hb66a35d2),
	.w3(32'hb73fef52),
	.w4(32'hb53bbd38),
	.w5(32'h36411623),
	.w6(32'hb6ffd8b3),
	.w7(32'h36802543),
	.w8(32'h36e39c84),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81cb5da),
	.w1(32'hb7f1ce55),
	.w2(32'hb820f5f5),
	.w3(32'hb78e0d27),
	.w4(32'hb72338a6),
	.w5(32'hb7e26867),
	.w6(32'hb7014abf),
	.w7(32'hb69fb5fd),
	.w8(32'hb7c05dd8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf6fb5),
	.w1(32'hb832f9dd),
	.w2(32'hb84297b4),
	.w3(32'hb88f011d),
	.w4(32'h38b8dfcb),
	.w5(32'hb6e65029),
	.w6(32'hb8c4fb6f),
	.w7(32'h37f12529),
	.w8(32'h376d9e7a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb828187c),
	.w1(32'hb5c54cb3),
	.w2(32'hb82ad1e1),
	.w3(32'hb7b7dfdd),
	.w4(32'h37ce3277),
	.w5(32'hb809c37a),
	.w6(32'hb7b751bf),
	.w7(32'h3798eccc),
	.w8(32'hb741f41d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e7616),
	.w1(32'hb98209b8),
	.w2(32'h3a094536),
	.w3(32'h38d8853d),
	.w4(32'hb9b1c220),
	.w5(32'h3954a77c),
	.w6(32'h3796a5db),
	.w7(32'hb9ef9814),
	.w8(32'h38aa4a94),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b598a1b),
	.w1(32'h3b2f9543),
	.w2(32'h3b7bc29d),
	.w3(32'h3aa7797b),
	.w4(32'h3aaf7b1b),
	.w5(32'h3afbbfb6),
	.w6(32'hb9cd6396),
	.w7(32'hba271ab0),
	.w8(32'h38f0c0c4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bc2f4),
	.w1(32'h3b26a182),
	.w2(32'h3ab34aa5),
	.w3(32'h3ae4bb85),
	.w4(32'hb8cfe4e0),
	.w5(32'hba63f2f6),
	.w6(32'h3a232e73),
	.w7(32'h397122da),
	.w8(32'h39f5aa5a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8282c73),
	.w1(32'hb7887872),
	.w2(32'h37a74e54),
	.w3(32'hb83e7bc9),
	.w4(32'hb6e6bc30),
	.w5(32'h37dc2526),
	.w6(32'hb812d40c),
	.w7(32'hb7a0fd1a),
	.w8(32'hb48084d3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a78d9),
	.w1(32'h3b6eafa8),
	.w2(32'h3bb4f72e),
	.w3(32'h3a45b66a),
	.w4(32'h3a903155),
	.w5(32'h3b2422ad),
	.w6(32'hbab36610),
	.w7(32'hbac2b7d3),
	.w8(32'h3a2fcead),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399dd48d),
	.w1(32'h39bf6901),
	.w2(32'h3ad51a17),
	.w3(32'hba3e9e2b),
	.w4(32'hba90e721),
	.w5(32'hb9593da2),
	.w6(32'hbac61ac1),
	.w7(32'hbaf8848e),
	.w8(32'hba81dafe),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2f687),
	.w1(32'hb84bcd64),
	.w2(32'hb92834b4),
	.w3(32'h390a77a9),
	.w4(32'hb7e8ffbb),
	.w5(32'hb928e923),
	.w6(32'h39350b0f),
	.w7(32'h38e02a2f),
	.w8(32'h37e91096),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2be68),
	.w1(32'h3aa8bbb1),
	.w2(32'h3aead2a0),
	.w3(32'h37112b23),
	.w4(32'h39aed7cf),
	.w5(32'h3a40a77a),
	.w6(32'hb9f57f6b),
	.w7(32'hba0a6692),
	.w8(32'h39024238),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dff37b),
	.w1(32'h391cc2ac),
	.w2(32'h376555ec),
	.w3(32'h393602b9),
	.w4(32'h3955dd9a),
	.w5(32'h380f3e6d),
	.w6(32'h3950bb61),
	.w7(32'h3965eae6),
	.w8(32'h3837d985),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9236422),
	.w1(32'hb8f1c1ec),
	.w2(32'hb78f4a2f),
	.w3(32'hb842c899),
	.w4(32'hb5cbebf0),
	.w5(32'hb82be4c3),
	.w6(32'h379ea594),
	.w7(32'h38b00e04),
	.w8(32'hb92b468d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87f5e5f),
	.w1(32'hb828bc5a),
	.w2(32'hb764a5bc),
	.w3(32'hb879cb23),
	.w4(32'hb7a36906),
	.w5(32'hb6c0fbee),
	.w6(32'hb87b232f),
	.w7(32'hb7276096),
	.w8(32'h372daad5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f5a358),
	.w1(32'h368811d8),
	.w2(32'h37460ed3),
	.w3(32'hb4456a03),
	.w4(32'h34ecdd90),
	.w5(32'h366f47da),
	.w6(32'hb4479d35),
	.w7(32'h3695709b),
	.w8(32'h3791f486),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60ec73),
	.w1(32'h3a22ea77),
	.w2(32'h3a9de85b),
	.w3(32'h39cb9aa9),
	.w4(32'hb8fabdf7),
	.w5(32'h3a7f0b37),
	.w6(32'h39f95689),
	.w7(32'hb7a122b1),
	.w8(32'h3a765574),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b451d),
	.w1(32'h3b82519f),
	.w2(32'h3be3e81b),
	.w3(32'h3a536c79),
	.w4(32'h3a2034f5),
	.w5(32'h3b3bc758),
	.w6(32'hbacace86),
	.w7(32'hbb036905),
	.w8(32'h3a1f32fb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35d2c8),
	.w1(32'h3ade52a5),
	.w2(32'h3b32282d),
	.w3(32'h39a418ad),
	.w4(32'hb98af1d4),
	.w5(32'h3a242105),
	.w6(32'hba802d90),
	.w7(32'hbaa2117e),
	.w8(32'hb870a0db),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b848904),
	.w1(32'h3b380042),
	.w2(32'h3b483dca),
	.w3(32'h3a9e9e8b),
	.w4(32'h3a0e9c99),
	.w5(32'h3aeb02d4),
	.w6(32'hb853db8e),
	.w7(32'hbad0a30c),
	.w8(32'hba764127),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81f97fd),
	.w1(32'h38a2bf48),
	.w2(32'h39982b1f),
	.w3(32'hb91b225f),
	.w4(32'hb8620d8e),
	.w5(32'h3940f12c),
	.w6(32'hb907f5e2),
	.w7(32'hb8e73f01),
	.w8(32'h390f2a36),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a99c23),
	.w1(32'hb5702f7c),
	.w2(32'hb6fddc54),
	.w3(32'hb7809898),
	.w4(32'h361f985f),
	.w5(32'h36893da1),
	.w6(32'hb790b9d9),
	.w7(32'hb67a4fea),
	.w8(32'h35faa75a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d3b964),
	.w1(32'hb85aeafd),
	.w2(32'hb86240f7),
	.w3(32'hb803f4a5),
	.w4(32'hb7e41215),
	.w5(32'hb812c973),
	.w6(32'hb795d17e),
	.w7(32'hb86a7425),
	.w8(32'hb80045b1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80db93c),
	.w1(32'hb8128f92),
	.w2(32'hb7c48b71),
	.w3(32'hb77d5d87),
	.w4(32'h37165611),
	.w5(32'hb64545c0),
	.w6(32'hb782eec3),
	.w7(32'h37e59450),
	.w8(32'h37a5437e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cb017),
	.w1(32'h3b70fef5),
	.w2(32'h3b467dbe),
	.w3(32'h3af4af7d),
	.w4(32'h3aa89c7b),
	.w5(32'h3ac05fb1),
	.w6(32'h38a5f525),
	.w7(32'hba11b31b),
	.w8(32'h398e18d5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e78b0a),
	.w1(32'hb91ef93c),
	.w2(32'hb88ab36f),
	.w3(32'hb9380c71),
	.w4(32'h38448320),
	.w5(32'hb8ecff9e),
	.w6(32'hb88df53a),
	.w7(32'hb8e86f6d),
	.w8(32'hb9c1302c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7e7f2),
	.w1(32'hb9c76697),
	.w2(32'h3a8b6248),
	.w3(32'h39ab3496),
	.w4(32'hb9aa1603),
	.w5(32'h3a8d8ab2),
	.w6(32'h3a6506d8),
	.w7(32'h390c9713),
	.w8(32'h3a83e1dd),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39800b42),
	.w1(32'hb903f22e),
	.w2(32'h39ca906d),
	.w3(32'h39a126cf),
	.w4(32'hb8afdfcd),
	.w5(32'h3989c270),
	.w6(32'h39fd8f57),
	.w7(32'h381e4e42),
	.w8(32'h39fb03ad),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8341f2b),
	.w1(32'h38b3c53b),
	.w2(32'h36e97945),
	.w3(32'h38f01ca1),
	.w4(32'h390b2052),
	.w5(32'hb8c69d00),
	.w6(32'h3921bb6c),
	.w7(32'h38ee9be8),
	.w8(32'hb8d68042),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adea16b),
	.w1(32'h3a8e31c4),
	.w2(32'h3a00ca94),
	.w3(32'h39c88c91),
	.w4(32'h38e2a468),
	.w5(32'hb91bc66d),
	.w6(32'h394230dd),
	.w7(32'hba0fc048),
	.w8(32'hb913ac0c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70b85de),
	.w1(32'hb79d8b20),
	.w2(32'hb753daea),
	.w3(32'h370f39e2),
	.w4(32'h37812379),
	.w5(32'h369ce527),
	.w6(32'hb5016248),
	.w7(32'h36f4a488),
	.w8(32'h36cc7c74),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58789d),
	.w1(32'h3b27904b),
	.w2(32'h3b8ecd4f),
	.w3(32'h3aee20a1),
	.w4(32'h3908cfa0),
	.w5(32'h3ac3fc2b),
	.w6(32'hb9b7d699),
	.w7(32'hba65fb5a),
	.w8(32'h3a3af7c9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f2d228),
	.w1(32'h390a5b8c),
	.w2(32'hb9c59e5a),
	.w3(32'hb752f99e),
	.w4(32'h391002f1),
	.w5(32'hb9d4b849),
	.w6(32'h399bc25e),
	.w7(32'hb8aceab8),
	.w8(32'h37a36b05),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa82f04),
	.w1(32'hbadde15f),
	.w2(32'h39d54c52),
	.w3(32'h3a8c665c),
	.w4(32'hbadbd304),
	.w5(32'h3a22ce59),
	.w6(32'h3af568a0),
	.w7(32'hba4bd14b),
	.w8(32'h3ab9a56e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule