module layer_10_featuremap_371(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdc848),
	.w1(32'h3b3b5cf8),
	.w2(32'h3ac6f8b1),
	.w3(32'hbc0635a4),
	.w4(32'h3a37b654),
	.w5(32'h3b1990ef),
	.w6(32'hbbfc4769),
	.w7(32'h3c08a1b6),
	.w8(32'hbb896e1c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc8ea6e),
	.w1(32'h3c152234),
	.w2(32'hbc879995),
	.w3(32'hbb34eb16),
	.w4(32'hbbdaceb5),
	.w5(32'hbaa993ab),
	.w6(32'hbcd4bedc),
	.w7(32'hbc5a9ac7),
	.w8(32'h3bc1cec9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b350b78),
	.w1(32'h3990c4e8),
	.w2(32'h3c6b0a48),
	.w3(32'hbbd60433),
	.w4(32'h3bbab615),
	.w5(32'h3c006f5c),
	.w6(32'h3d0fee44),
	.w7(32'h3ba483ff),
	.w8(32'hbc029266),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ffac),
	.w1(32'h3c68ccdd),
	.w2(32'h3bd32bfd),
	.w3(32'h3b7f662b),
	.w4(32'h376a9cbc),
	.w5(32'h3c8e7313),
	.w6(32'hbb93a5cd),
	.w7(32'h3ba8f420),
	.w8(32'h3a4b19fb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6da00),
	.w1(32'h3c361265),
	.w2(32'hba9aa972),
	.w3(32'hbd5ddaf2),
	.w4(32'hbb4be305),
	.w5(32'h3aa8aeec),
	.w6(32'h3b8513f3),
	.w7(32'hba8427b3),
	.w8(32'hbd0be2e5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd376f5),
	.w1(32'h3a016405),
	.w2(32'hbbdf72f1),
	.w3(32'h3b38864f),
	.w4(32'h3ba29993),
	.w5(32'h3c2ced24),
	.w6(32'hba7f2698),
	.w7(32'hbc230d09),
	.w8(32'h3c421447),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40a9fd),
	.w1(32'h3aa23a48),
	.w2(32'hbc24542e),
	.w3(32'hbc9e97b5),
	.w4(32'h3d0fc0de),
	.w5(32'hbd10a768),
	.w6(32'hbae2efde),
	.w7(32'hbb1e7a87),
	.w8(32'hbc138d56),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b80e2),
	.w1(32'h3c1f5407),
	.w2(32'hbc82d8f0),
	.w3(32'hbc4522a6),
	.w4(32'hbc03776d),
	.w5(32'h3bce10e4),
	.w6(32'hbc0c87ff),
	.w7(32'hbc85daa5),
	.w8(32'h3c4a73af),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca313d8),
	.w1(32'h3c063759),
	.w2(32'hbc23396b),
	.w3(32'hba2cb745),
	.w4(32'hbc20fbfd),
	.w5(32'hbc056800),
	.w6(32'hbb44c836),
	.w7(32'h3ab75c81),
	.w8(32'hbb5aec02),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd89253),
	.w1(32'hbc6b05a4),
	.w2(32'hbbea9e4b),
	.w3(32'h3aa1d335),
	.w4(32'h3c832eba),
	.w5(32'hbae9357d),
	.w6(32'hbb96a6bb),
	.w7(32'hba64b14f),
	.w8(32'hbc4bcb3e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a707b71),
	.w1(32'hbb8010de),
	.w2(32'h3ae23c5c),
	.w3(32'h3b6f0e32),
	.w4(32'h3b9fdfbf),
	.w5(32'hbcee3bc1),
	.w6(32'hbb59d430),
	.w7(32'hbbe0e91e),
	.w8(32'h3ae8be81),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ca06f),
	.w1(32'hbc87d281),
	.w2(32'hbd55b51e),
	.w3(32'hbc3a1e5c),
	.w4(32'hbc799b82),
	.w5(32'h3c0c7292),
	.w6(32'h39dd5ef8),
	.w7(32'h3bcf5654),
	.w8(32'hbc89e962),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66cd59),
	.w1(32'h3bd9b8fa),
	.w2(32'hbc935f6f),
	.w3(32'hbb262380),
	.w4(32'h3b8bbf43),
	.w5(32'h3c6b116e),
	.w6(32'h3bff3b0d),
	.w7(32'h3ba22b6c),
	.w8(32'hbd09ae5b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf3ca6),
	.w1(32'hbc82a7c4),
	.w2(32'hbc7af1a1),
	.w3(32'hbc24220c),
	.w4(32'h3d308976),
	.w5(32'hbc2d2e8e),
	.w6(32'h3c182c7c),
	.w7(32'h3c8d1fa0),
	.w8(32'hbb96d246),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc535e76),
	.w1(32'h3c096c0c),
	.w2(32'h3beda0c8),
	.w3(32'hb9672d17),
	.w4(32'hbc4edfe2),
	.w5(32'hb9cf6c63),
	.w6(32'h3b74e3af),
	.w7(32'h3c521bb1),
	.w8(32'h3bb8945f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1db74),
	.w1(32'hbc3f18ba),
	.w2(32'hbc67c16d),
	.w3(32'hbc10d52b),
	.w4(32'h3c08a45a),
	.w5(32'hbc71bd8b),
	.w6(32'h3c3589cb),
	.w7(32'h3967511e),
	.w8(32'hbce0830e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda1eed),
	.w1(32'h3c3d29ee),
	.w2(32'hbc1d4679),
	.w3(32'hbb35d86b),
	.w4(32'h3a7d5752),
	.w5(32'hbc5786d3),
	.w6(32'hbaf8a0f5),
	.w7(32'hbb0e1b16),
	.w8(32'hba7a74f2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9243fa5),
	.w1(32'h3aa54368),
	.w2(32'hbd2cec99),
	.w3(32'h3a47896b),
	.w4(32'h3bf7ce0b),
	.w5(32'hbc63314f),
	.w6(32'hbb2a589f),
	.w7(32'hbd8f5f7a),
	.w8(32'hbcdaaa0a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70120e),
	.w1(32'hbb60145d),
	.w2(32'hbca0a1dd),
	.w3(32'hbb7587bc),
	.w4(32'hba8472da),
	.w5(32'h3b190b04),
	.w6(32'h3b6b2cd3),
	.w7(32'h3c54c40a),
	.w8(32'hbc961e34),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c468fc8),
	.w1(32'h3cc2312d),
	.w2(32'h3c3e42ea),
	.w3(32'hbc4269de),
	.w4(32'h3d61cd8d),
	.w5(32'h3c04fbac),
	.w6(32'h3c71a6a4),
	.w7(32'hba437d15),
	.w8(32'hbc205bee),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bb020),
	.w1(32'h3ac33725),
	.w2(32'h3cf71413),
	.w3(32'h39799bb5),
	.w4(32'hbb21d78a),
	.w5(32'hbad0b31d),
	.w6(32'h3b0f99a3),
	.w7(32'h3b161eca),
	.w8(32'hbbf794e6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc901a15),
	.w1(32'h3c9f4e5b),
	.w2(32'h3b15676d),
	.w3(32'hba595366),
	.w4(32'hbb7d99df),
	.w5(32'hbba065be),
	.w6(32'hbd241156),
	.w7(32'h3aad152d),
	.w8(32'h3bd76626),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9352fa),
	.w1(32'hbc9295fd),
	.w2(32'hbd2d0b4d),
	.w3(32'hb934d8b5),
	.w4(32'h3cba8911),
	.w5(32'h3c955e6e),
	.w6(32'h3cd359bd),
	.w7(32'hbab24426),
	.w8(32'hbcebf0f8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb82cd7),
	.w1(32'hbc04010d),
	.w2(32'hb9b390e8),
	.w3(32'h3c71c441),
	.w4(32'h3c038d6e),
	.w5(32'hbabe2cb4),
	.w6(32'hbb64d1cd),
	.w7(32'hbb96eff8),
	.w8(32'h3adef3ed),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badec80),
	.w1(32'h3d04ba86),
	.w2(32'h3d0048aa),
	.w3(32'h3c0360c7),
	.w4(32'hbd6d87d8),
	.w5(32'hbb12e8f4),
	.w6(32'h3b76c09a),
	.w7(32'hbbc03a09),
	.w8(32'hbc528a23),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc6079),
	.w1(32'hb9a24cbb),
	.w2(32'hbb8846a3),
	.w3(32'h3c1d9b8b),
	.w4(32'h3b19dc09),
	.w5(32'hbc1a083c),
	.w6(32'h3c4ffc13),
	.w7(32'h3c5eb47e),
	.w8(32'hbbcdb221),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37d0bc),
	.w1(32'h3c076bd0),
	.w2(32'hbaee3635),
	.w3(32'h3c3121b2),
	.w4(32'hbb754179),
	.w5(32'h3adefd1f),
	.w6(32'h3a9a4609),
	.w7(32'hbba5d4b1),
	.w8(32'hbbdb3df9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13b7cf),
	.w1(32'hbcc2b2ff),
	.w2(32'hbac85ae3),
	.w3(32'h3c8d3bb8),
	.w4(32'hbc147adb),
	.w5(32'hbc59a396),
	.w6(32'hbcaec1d2),
	.w7(32'hbc8571e6),
	.w8(32'h3b404b99),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2ebec),
	.w1(32'h3c4de4ef),
	.w2(32'hbbd75c2b),
	.w3(32'h3c311dc2),
	.w4(32'hb8d31f99),
	.w5(32'h3bf7ee85),
	.w6(32'hb90bb9eb),
	.w7(32'hbaf374d2),
	.w8(32'h3b93fb04),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72a941),
	.w1(32'h3c91c6da),
	.w2(32'h3c4a934d),
	.w3(32'h38dfa2be),
	.w4(32'hbc597d75),
	.w5(32'hbc3c19b9),
	.w6(32'h3c5b6171),
	.w7(32'h3a40a1c8),
	.w8(32'h3c15340d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a80dc0),
	.w1(32'h3ae19153),
	.w2(32'h3c8b8b0f),
	.w3(32'h3b734b06),
	.w4(32'hbc05388a),
	.w5(32'hbbfbd066),
	.w6(32'h3a979d25),
	.w7(32'hbb81ab22),
	.w8(32'h3c2c58a1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19edf6),
	.w1(32'hba79c900),
	.w2(32'h3ca2aaf9),
	.w3(32'hbc1ac002),
	.w4(32'hbb9760f3),
	.w5(32'h3b3fec31),
	.w6(32'hba9b7bc2),
	.w7(32'h3b6e795d),
	.w8(32'hbbaa676d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44e3eb),
	.w1(32'hbb984d19),
	.w2(32'h3b02b387),
	.w3(32'hbc006ba5),
	.w4(32'hb8a34380),
	.w5(32'hbc25b15a),
	.w6(32'hbaade66d),
	.w7(32'hbb8335ec),
	.w8(32'hb85cd5d7),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5abcef),
	.w1(32'h3d3a1b1f),
	.w2(32'h3ad57142),
	.w3(32'hba82d135),
	.w4(32'hbb0a6967),
	.w5(32'h3a024f47),
	.w6(32'hba8f212e),
	.w7(32'hbbae4d1d),
	.w8(32'hbb3ba864),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30ecb8),
	.w1(32'hbb426d34),
	.w2(32'hbc8ddedc),
	.w3(32'h3ba4b37d),
	.w4(32'h3c92fa69),
	.w5(32'h3b0f45ed),
	.w6(32'h39ab382f),
	.w7(32'h3c2fa410),
	.w8(32'hbc01623e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c267458),
	.w1(32'h3c316809),
	.w2(32'hbc19ade8),
	.w3(32'hbbb69e9b),
	.w4(32'hbb62bc29),
	.w5(32'h3c6cd1eb),
	.w6(32'hbc3b853d),
	.w7(32'hbb0b7310),
	.w8(32'h3b92394f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfd8419),
	.w1(32'h39b8065a),
	.w2(32'hba9a4f50),
	.w3(32'hbcd0d3b4),
	.w4(32'hbc4f9e3a),
	.w5(32'h3cb93373),
	.w6(32'hbac48b87),
	.w7(32'h3d060c00),
	.w8(32'h3cfd23ac),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89bdda),
	.w1(32'h3b845c9a),
	.w2(32'h3ca408e2),
	.w3(32'hbcaf2d60),
	.w4(32'hbc8b9f13),
	.w5(32'hbc184d81),
	.w6(32'hbc4a599a),
	.w7(32'hbc149e5a),
	.w8(32'hbc506aff),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bf100),
	.w1(32'hbc982295),
	.w2(32'h3c4f3466),
	.w3(32'h3bfad171),
	.w4(32'hbcf774e4),
	.w5(32'h3c03374f),
	.w6(32'hbc2153cb),
	.w7(32'hbc1b889f),
	.w8(32'hbbd9b53e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65d805),
	.w1(32'h3b732605),
	.w2(32'h3ba52cc4),
	.w3(32'h3b1b4a69),
	.w4(32'hbc21c3ae),
	.w5(32'hbb1cc04a),
	.w6(32'hbbf6ea72),
	.w7(32'h3bb2da48),
	.w8(32'h3b8ad2a2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4671b),
	.w1(32'h3bb2ab4d),
	.w2(32'h3c0b6ae0),
	.w3(32'hbbd4c742),
	.w4(32'hbbf9a30e),
	.w5(32'hbbc12405),
	.w6(32'hb924bf6f),
	.w7(32'h3abfbf0f),
	.w8(32'h3b669ec5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2decf9),
	.w1(32'hb9fac5ba),
	.w2(32'h3b12350d),
	.w3(32'hbb5f7d8d),
	.w4(32'h38312eec),
	.w5(32'h3b894be3),
	.w6(32'h3b9be4b5),
	.w7(32'h3a91db1b),
	.w8(32'h3be97890),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b643928),
	.w1(32'h3bd39d00),
	.w2(32'hbc07d945),
	.w3(32'h3c0aeff5),
	.w4(32'h39186b7a),
	.w5(32'h3c5d1962),
	.w6(32'hbc421282),
	.w7(32'h3bd93e20),
	.w8(32'h3ab0dd60),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa1d8d),
	.w1(32'hbc4ea0c8),
	.w2(32'hbcce728e),
	.w3(32'h3a496e1e),
	.w4(32'h3be38044),
	.w5(32'hbc9f09ad),
	.w6(32'h3be48dff),
	.w7(32'hbbe7389c),
	.w8(32'hbc52dad1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc218e11),
	.w1(32'hbaaed70f),
	.w2(32'h3bfe68cc),
	.w3(32'h3b22a376),
	.w4(32'h3abff155),
	.w5(32'h3b97b2e2),
	.w6(32'h3a1d7825),
	.w7(32'h3c200d6f),
	.w8(32'h3bb81df1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a904b8c),
	.w1(32'h3bfc6531),
	.w2(32'h3cec516c),
	.w3(32'hba4502f2),
	.w4(32'hbc013bb7),
	.w5(32'hbcc7688d),
	.w6(32'h3b6828a6),
	.w7(32'hbb5e5e8a),
	.w8(32'hbb45cb09),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7310a0),
	.w1(32'hba2ee1e5),
	.w2(32'h3b324d97),
	.w3(32'hbacfe6f4),
	.w4(32'hba21d1fe),
	.w5(32'hbbd0f200),
	.w6(32'h3b5daf3c),
	.w7(32'h3c0071aa),
	.w8(32'h3b77d680),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc7fa7),
	.w1(32'hbb157b0e),
	.w2(32'hbcffc561),
	.w3(32'h3c87f630),
	.w4(32'h3c4e4a39),
	.w5(32'hbbe22aa1),
	.w6(32'h3c2667e4),
	.w7(32'hbbf97f9c),
	.w8(32'hbd0b659b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cdf6b),
	.w1(32'h3b0f525a),
	.w2(32'hbb653af0),
	.w3(32'hbaba5156),
	.w4(32'hba23ca8e),
	.w5(32'hba820884),
	.w6(32'hbac429ab),
	.w7(32'hbb83c66d),
	.w8(32'h3b19efe0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3871557a),
	.w1(32'hbaa7b42e),
	.w2(32'h3ac9093c),
	.w3(32'h3b5bf615),
	.w4(32'hbc80c9f7),
	.w5(32'h3be3c50d),
	.w6(32'hbb8dfdaa),
	.w7(32'h3bc72229),
	.w8(32'h3b008b2f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b706c3f),
	.w1(32'h3c36649b),
	.w2(32'h3b252178),
	.w3(32'hbac7ad78),
	.w4(32'hbade0050),
	.w5(32'hb896f6a6),
	.w6(32'hbb2801e4),
	.w7(32'hbba5f483),
	.w8(32'h391e859a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd83c0a),
	.w1(32'hbbf3b6bd),
	.w2(32'h3b6d29c8),
	.w3(32'h3c2d7037),
	.w4(32'h3c1182d5),
	.w5(32'hbb510e00),
	.w6(32'h3c5fbf3c),
	.w7(32'hbb685a26),
	.w8(32'h3882fa6a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b767878),
	.w1(32'h3b230d44),
	.w2(32'hbc035097),
	.w3(32'hbc14300e),
	.w4(32'h3b5731a6),
	.w5(32'h3c2a251f),
	.w6(32'hba07128d),
	.w7(32'h3c02d64f),
	.w8(32'h3aa0a368),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d9bf8),
	.w1(32'hbc302737),
	.w2(32'hbcf24504),
	.w3(32'hba2beeef),
	.w4(32'h3b6b85ad),
	.w5(32'hbc6b642e),
	.w6(32'h3c4ab395),
	.w7(32'hba2d9ece),
	.w8(32'hba2434bf),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b72c6),
	.w1(32'hb96e7ba6),
	.w2(32'h3c05fc6d),
	.w3(32'h3c8fdc7b),
	.w4(32'h3b895e66),
	.w5(32'hbc463707),
	.w6(32'hbbf6bbe5),
	.w7(32'hba7cf1d9),
	.w8(32'hba999844),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb88a4d),
	.w1(32'h3c5995bc),
	.w2(32'h3c15647b),
	.w3(32'hbc9a0eff),
	.w4(32'h3b16e93d),
	.w5(32'h3a824c1e),
	.w6(32'hb954427e),
	.w7(32'hbbeb07e1),
	.w8(32'h398d7a58),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fa8a9),
	.w1(32'h3aedd4f5),
	.w2(32'h3b815184),
	.w3(32'hba956f18),
	.w4(32'hbaccb99e),
	.w5(32'h3b23a121),
	.w6(32'h3c9076e1),
	.w7(32'hba5e8383),
	.w8(32'h3903a92f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f424b),
	.w1(32'h3a7cd3d7),
	.w2(32'h3c3eea0a),
	.w3(32'h3c39502e),
	.w4(32'h3c20c5d1),
	.w5(32'h3b516fae),
	.w6(32'hbc09ad54),
	.w7(32'h3d057bf3),
	.w8(32'h3bf8fbe2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cb249),
	.w1(32'h3baf3edf),
	.w2(32'hbc32a083),
	.w3(32'h3cb44ae0),
	.w4(32'hbac9e6bf),
	.w5(32'h3a5d4600),
	.w6(32'h39856328),
	.w7(32'hbb88df2a),
	.w8(32'h3bf8ee59),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1567c),
	.w1(32'h3c3cb246),
	.w2(32'hbbea3f43),
	.w3(32'hbc92cf8d),
	.w4(32'hbc3b5c60),
	.w5(32'hbc0fe55b),
	.w6(32'hb9d2310c),
	.w7(32'hbc18921a),
	.w8(32'hbc0c2bdc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ae80a),
	.w1(32'h3c2d533b),
	.w2(32'hbce55d09),
	.w3(32'hbb81c474),
	.w4(32'h3a9c609f),
	.w5(32'h3b1148ce),
	.w6(32'hbc86547a),
	.w7(32'hbc5134ea),
	.w8(32'hbc9d785b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6aab96),
	.w1(32'hbb1cbc5c),
	.w2(32'hbb67a8c8),
	.w3(32'hbaa9b76f),
	.w4(32'h3c58242a),
	.w5(32'hbc84a5dc),
	.w6(32'hbc9deb99),
	.w7(32'hbc6c647e),
	.w8(32'h3bbed87c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42e796),
	.w1(32'hbb930e67),
	.w2(32'h3a86715a),
	.w3(32'h3c531660),
	.w4(32'hbb83b8e2),
	.w5(32'hbc0d0f64),
	.w6(32'hbc4bda7d),
	.w7(32'h3bf83be7),
	.w8(32'h3aef927a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ad03e),
	.w1(32'h3c3c6216),
	.w2(32'hbc8f15fd),
	.w3(32'h3c790c02),
	.w4(32'hbbb86653),
	.w5(32'h3c11211a),
	.w6(32'h3b8077a9),
	.w7(32'hbabf0971),
	.w8(32'h3bb3dd28),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56313e),
	.w1(32'hbc1dc1c9),
	.w2(32'h3bc34175),
	.w3(32'hba28da27),
	.w4(32'hbb64dc45),
	.w5(32'hbb567370),
	.w6(32'h3bd7a261),
	.w7(32'h3c1550ad),
	.w8(32'hba1929a7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7252cd),
	.w1(32'hbb7ff200),
	.w2(32'hbc1db372),
	.w3(32'hbb6d88da),
	.w4(32'hba5fa6aa),
	.w5(32'h3b31f21b),
	.w6(32'h396895bd),
	.w7(32'h3c1bcb1f),
	.w8(32'h3aeb2057),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bc1cc),
	.w1(32'hbcf0204e),
	.w2(32'hbdc23508),
	.w3(32'h3b4a4356),
	.w4(32'h3ca00ff1),
	.w5(32'hbc6c6ea2),
	.w6(32'hbb2306cf),
	.w7(32'h3c803d5f),
	.w8(32'h3b07aaeb),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80764f),
	.w1(32'h3b8acacf),
	.w2(32'hbbe1cfba),
	.w3(32'h3c2ff812),
	.w4(32'hbba08c03),
	.w5(32'hbc3d5cad),
	.w6(32'hbb43baf2),
	.w7(32'hbbce0c52),
	.w8(32'hbc5b72f5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefdcd7),
	.w1(32'h3c277033),
	.w2(32'hbc0cf512),
	.w3(32'hbbeb53ad),
	.w4(32'h3bd93dbd),
	.w5(32'hbd062aa9),
	.w6(32'h3cbc3491),
	.w7(32'hbc137209),
	.w8(32'hbc87e54c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f5fc2),
	.w1(32'h3cb64d5c),
	.w2(32'h3d7a639a),
	.w3(32'h3c1e7476),
	.w4(32'hbc887f22),
	.w5(32'hbc14e214),
	.w6(32'hbb9d4e53),
	.w7(32'hba8076e9),
	.w8(32'h3c97995c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf19fb0),
	.w1(32'h3bbb7c1a),
	.w2(32'hbc00141b),
	.w3(32'h3b9217ee),
	.w4(32'h3b725542),
	.w5(32'h3b35f471),
	.w6(32'hbbf4ca47),
	.w7(32'hbc697e99),
	.w8(32'hbc7fba8a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e8142),
	.w1(32'h3c261d3f),
	.w2(32'h3c2d31fa),
	.w3(32'h3bf21077),
	.w4(32'h392e3072),
	.w5(32'h3a71cffe),
	.w6(32'h3c070883),
	.w7(32'hbb27c790),
	.w8(32'hbc0049a5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18721a),
	.w1(32'h3ab46fb4),
	.w2(32'h3cdbce19),
	.w3(32'hbc0d360c),
	.w4(32'hbc761654),
	.w5(32'hbc8b89ea),
	.w6(32'hba27db50),
	.w7(32'h3c3a9e91),
	.w8(32'h3c69c736),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb928c5f),
	.w1(32'h38fbc9bb),
	.w2(32'hbc2f7620),
	.w3(32'h3b2fdb86),
	.w4(32'h3b21e800),
	.w5(32'hbbd9c708),
	.w6(32'hbb810951),
	.w7(32'h3a572202),
	.w8(32'hbbec92c2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66c968),
	.w1(32'h3bdcb13d),
	.w2(32'hbbdf48cb),
	.w3(32'h3b600481),
	.w4(32'h3a4f787f),
	.w5(32'hbc3611f2),
	.w6(32'h3b903125),
	.w7(32'hba571301),
	.w8(32'h3b31614b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b762ab8),
	.w1(32'h3b389b35),
	.w2(32'hbd1345e9),
	.w3(32'h3c09720a),
	.w4(32'h3a879970),
	.w5(32'hbadd4170),
	.w6(32'hbc1760b7),
	.w7(32'h3bba33b5),
	.w8(32'hbc07a047),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf53edf),
	.w1(32'h3b9deeb4),
	.w2(32'hbc1326be),
	.w3(32'hbbd93a73),
	.w4(32'h3be860ce),
	.w5(32'hbb0e4fde),
	.w6(32'h3c1a5e42),
	.w7(32'hbab5b53e),
	.w8(32'hbc129a7e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e589a),
	.w1(32'h3c033ebc),
	.w2(32'h3c1489fb),
	.w3(32'h3be8b89c),
	.w4(32'hbc0db684),
	.w5(32'h3b25a07c),
	.w6(32'h3c4d175b),
	.w7(32'h3b1f4e05),
	.w8(32'hba6a4d90),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e54f),
	.w1(32'hbba2fb8d),
	.w2(32'hbb51571d),
	.w3(32'hbcafd1fe),
	.w4(32'h3bbc7c88),
	.w5(32'h3cce486d),
	.w6(32'h3b9e7dec),
	.w7(32'h3a5313a9),
	.w8(32'hbb916847),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c484945),
	.w1(32'hbc4387d0),
	.w2(32'hbd0f12b0),
	.w3(32'h3c059f9f),
	.w4(32'h3ce3c6d7),
	.w5(32'hbc9057ae),
	.w6(32'h382f034c),
	.w7(32'h3c02600d),
	.w8(32'h3a8d4b01),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc397a48),
	.w1(32'hbaba7755),
	.w2(32'hbb0aad8e),
	.w3(32'h3b6541e3),
	.w4(32'hbbb627da),
	.w5(32'hbad6a4c1),
	.w6(32'h3b8cdd9e),
	.w7(32'h3c3e5005),
	.w8(32'h3b1a4dab),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cb56a),
	.w1(32'hbbe1230a),
	.w2(32'h3bf552f0),
	.w3(32'hbc3c1fdd),
	.w4(32'h3c0213fc),
	.w5(32'hbc853833),
	.w6(32'hbb7f0fa0),
	.w7(32'h3b540163),
	.w8(32'hbb8a6902),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0878cf),
	.w1(32'hbc5933b7),
	.w2(32'hbc01a948),
	.w3(32'hbad4b762),
	.w4(32'hbb8fd963),
	.w5(32'hbbb4e435),
	.w6(32'hbc368add),
	.w7(32'hbc6958b1),
	.w8(32'hbbe4888e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71f786),
	.w1(32'h3c8943c3),
	.w2(32'hba511bfd),
	.w3(32'h3c2494fc),
	.w4(32'hbb95f0ae),
	.w5(32'hbb981a6d),
	.w6(32'hbc2dba76),
	.w7(32'hbc8cc86e),
	.w8(32'h3b894c5b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfb78d),
	.w1(32'hbb9ebf6c),
	.w2(32'hbb4688e7),
	.w3(32'hba618dd1),
	.w4(32'h3c14d2a3),
	.w5(32'hbb34b4cf),
	.w6(32'hbb33cf76),
	.w7(32'hbb427024),
	.w8(32'hbbb44a69),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66d7fa),
	.w1(32'h3c09b6a2),
	.w2(32'hbb829542),
	.w3(32'hbbe403b5),
	.w4(32'hbbcb4f4a),
	.w5(32'hbb2c59f9),
	.w6(32'hbb4e8990),
	.w7(32'hbbd528d1),
	.w8(32'h3b05753d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e03e3),
	.w1(32'h3d4be1a1),
	.w2(32'h3c8086bb),
	.w3(32'h3c4dcdd8),
	.w4(32'hbc0c2d71),
	.w5(32'hb9695175),
	.w6(32'hbba6c49c),
	.w7(32'hbc1c1b99),
	.w8(32'h3b5e8127),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf6ba8),
	.w1(32'hba852d7a),
	.w2(32'hbbb60808),
	.w3(32'h3b87546f),
	.w4(32'h3b9af05e),
	.w5(32'h3c7d3390),
	.w6(32'h3bafd90b),
	.w7(32'hbd5547fd),
	.w8(32'h3a5a7136),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34165b),
	.w1(32'h3c4bffc0),
	.w2(32'h3c9f0d3e),
	.w3(32'h3abad25a),
	.w4(32'h3bfdd1de),
	.w5(32'h3c766598),
	.w6(32'h3bc6fc4f),
	.w7(32'h3b827886),
	.w8(32'h3c8e37a3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18a61e),
	.w1(32'h3ab6d6e3),
	.w2(32'hbc5b856a),
	.w3(32'h3c246f97),
	.w4(32'h3a0576a6),
	.w5(32'hbbcc8b10),
	.w6(32'hbbca69ff),
	.w7(32'hbb4c97ba),
	.w8(32'hbc8ebd1b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91185c),
	.w1(32'hbaf84073),
	.w2(32'h3c0ab6b2),
	.w3(32'hbc1d8bba),
	.w4(32'hbc09b801),
	.w5(32'hbc276f48),
	.w6(32'h3b3c38f9),
	.w7(32'h3ba1bca2),
	.w8(32'hbafc8a90),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b1eee),
	.w1(32'hbcc00d79),
	.w2(32'hbcae6155),
	.w3(32'h3c2d0d13),
	.w4(32'h3be8ed18),
	.w5(32'hbc137acb),
	.w6(32'h3cc27ac2),
	.w7(32'h3b95929d),
	.w8(32'hbc6a3292),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0f7bc),
	.w1(32'hb9803aeb),
	.w2(32'h3c289ff8),
	.w3(32'hbc0063de),
	.w4(32'hbc86af23),
	.w5(32'hbbc30a4c),
	.w6(32'hbc220184),
	.w7(32'hbc51828b),
	.w8(32'h3b7c5da6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab34baf),
	.w1(32'hba53fd50),
	.w2(32'hbd15e236),
	.w3(32'h3c5c331e),
	.w4(32'h3c3d4bc4),
	.w5(32'hbbc7a009),
	.w6(32'h3c0be4ce),
	.w7(32'hbb24b471),
	.w8(32'hbbdfe292),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32f5af),
	.w1(32'h3bfd0015),
	.w2(32'hbcbff285),
	.w3(32'h3c1d30aa),
	.w4(32'hbba7e87c),
	.w5(32'h39c21774),
	.w6(32'h3a8f12f2),
	.w7(32'h3bb7e223),
	.w8(32'h3b4f225a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c009957),
	.w1(32'h3c06bf4f),
	.w2(32'h3bce2696),
	.w3(32'hbbdf65b8),
	.w4(32'hbae5c821),
	.w5(32'h3bf9ffc9),
	.w6(32'hba61d862),
	.w7(32'h3bfddee4),
	.w8(32'h3bc765e2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa896c4),
	.w1(32'hbb52db03),
	.w2(32'hbc04d71e),
	.w3(32'hbc369f4a),
	.w4(32'h3b60cebb),
	.w5(32'h3c873186),
	.w6(32'hba9d5f8c),
	.w7(32'hba7f25e0),
	.w8(32'hb91bfb6e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d57f311),
	.w1(32'hbcaece8e),
	.w2(32'hbc18e4f9),
	.w3(32'h3b56b0ca),
	.w4(32'h3c5252fe),
	.w5(32'hbb898a90),
	.w6(32'h39b4c377),
	.w7(32'h3b8c8782),
	.w8(32'hbc2b586b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d727b),
	.w1(32'hbcfab906),
	.w2(32'h3bc3266b),
	.w3(32'hbc3e55db),
	.w4(32'h3b434ab4),
	.w5(32'hbd73061b),
	.w6(32'hbca83e86),
	.w7(32'h3d005c3d),
	.w8(32'h3b1f3e32),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31a17d),
	.w1(32'hba97e516),
	.w2(32'h3ce0cd7f),
	.w3(32'hbcacd316),
	.w4(32'hbbf54849),
	.w5(32'h3c9aaba0),
	.w6(32'h3c451261),
	.w7(32'h3c9c064e),
	.w8(32'h3cafd5a0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefd218),
	.w1(32'h3c2430e8),
	.w2(32'h3cbd1ca8),
	.w3(32'hbc246a9c),
	.w4(32'h3bc10b33),
	.w5(32'h3bd8584c),
	.w6(32'hbb456d73),
	.w7(32'hbb502f70),
	.w8(32'h3b94f6bd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea7dba),
	.w1(32'h3c28fe9a),
	.w2(32'h3c4230db),
	.w3(32'hbb361cb7),
	.w4(32'hbb023749),
	.w5(32'h3b45e482),
	.w6(32'hbc4dd90c),
	.w7(32'h3b031017),
	.w8(32'h3bfa269a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5fb18),
	.w1(32'h3a86d3be),
	.w2(32'hba8fdeb4),
	.w3(32'hbae9aaa0),
	.w4(32'h3c01c14a),
	.w5(32'h3cb0bddb),
	.w6(32'h3c32ea85),
	.w7(32'h3ca266a1),
	.w8(32'h3c8919ac),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbf0dd),
	.w1(32'h3b904d42),
	.w2(32'hbc5e192e),
	.w3(32'hbb061f18),
	.w4(32'hbbc14b74),
	.w5(32'hba109b92),
	.w6(32'hbadc9fd9),
	.w7(32'h3b0dc234),
	.w8(32'h3c82bcf2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0860cc),
	.w1(32'hbcddde60),
	.w2(32'h3cd2b4df),
	.w3(32'hbd198d16),
	.w4(32'hbc2bab32),
	.w5(32'h3a92d328),
	.w6(32'h3c9048ff),
	.w7(32'h3cca64fc),
	.w8(32'h3ce7aa48),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47def4),
	.w1(32'hbca6dbc2),
	.w2(32'hbc209d06),
	.w3(32'h3b5fd8b9),
	.w4(32'hbc82e59a),
	.w5(32'hbb86e6bb),
	.w6(32'hbb918751),
	.w7(32'h3bebf7ce),
	.w8(32'hbca303be),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb94698),
	.w1(32'hbc861ad0),
	.w2(32'h3bccefe7),
	.w3(32'h3c4e7443),
	.w4(32'h3be9015a),
	.w5(32'hb927c0ca),
	.w6(32'h3b0f1121),
	.w7(32'hbb48d8e3),
	.w8(32'h3b7c0fac),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8485bb),
	.w1(32'hbc007e73),
	.w2(32'hbb39900e),
	.w3(32'hbc5493e2),
	.w4(32'hb9c19016),
	.w5(32'hbb49ef9d),
	.w6(32'hbc20442f),
	.w7(32'h3b06085d),
	.w8(32'hbc191360),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcef403),
	.w1(32'hbc9458e7),
	.w2(32'hbb9d3ae6),
	.w3(32'h3c9813ef),
	.w4(32'h3b723f96),
	.w5(32'hbb18e0a7),
	.w6(32'hbbd44048),
	.w7(32'hbb2de7bf),
	.w8(32'hbac98ff1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c42a35),
	.w1(32'hbb7fb8d0),
	.w2(32'h3c4c17af),
	.w3(32'hbb82bb47),
	.w4(32'hbb2b162c),
	.w5(32'hbc8ce050),
	.w6(32'h3bef4f86),
	.w7(32'h3bf2a104),
	.w8(32'h3c1db284),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec3dc),
	.w1(32'hbc9a6202),
	.w2(32'hbc5bbbc6),
	.w3(32'h3bc08fb7),
	.w4(32'hbc906a33),
	.w5(32'hbcf8a1a0),
	.w6(32'hbbc67fa8),
	.w7(32'hbb4b840f),
	.w8(32'hbc9080a7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066a9a),
	.w1(32'hbba25aa8),
	.w2(32'h3bc3f2fb),
	.w3(32'h3b70ebaa),
	.w4(32'hbbf3961d),
	.w5(32'h3a7a6d0c),
	.w6(32'h3b25e301),
	.w7(32'h3c2705eb),
	.w8(32'hb9751cbf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e3f8d),
	.w1(32'h3cc42b7b),
	.w2(32'h3c6f82bb),
	.w3(32'hbbdefc92),
	.w4(32'hbb87e5f8),
	.w5(32'hb9a0ce5c),
	.w6(32'h3be2aabf),
	.w7(32'h3b90768f),
	.w8(32'hbbd8ea85),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd4a2d),
	.w1(32'hbcaf78c1),
	.w2(32'hbc7ba8ab),
	.w3(32'hbc9cce0f),
	.w4(32'hbb6d72e7),
	.w5(32'hbc8104f0),
	.w6(32'h3ba5e8a2),
	.w7(32'h3bb04197),
	.w8(32'h3b4d0cb7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2c39bb),
	.w1(32'h3b57bba4),
	.w2(32'h3bc410e8),
	.w3(32'h3bcca63b),
	.w4(32'h3bc7f070),
	.w5(32'h3c34a071),
	.w6(32'hbb9433ce),
	.w7(32'hbb64aa0d),
	.w8(32'h3c55800e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0267d5),
	.w1(32'hbbc46fb3),
	.w2(32'h3b5b14a9),
	.w3(32'hbbb15550),
	.w4(32'hbdb51458),
	.w5(32'h3b613963),
	.w6(32'hb96425e0),
	.w7(32'h3b24f7be),
	.w8(32'h3c089bc2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5b3670),
	.w1(32'h3b62d360),
	.w2(32'hbbae88f7),
	.w3(32'hbb008018),
	.w4(32'hbb14afe9),
	.w5(32'h3c8f454e),
	.w6(32'hbbc5ad4f),
	.w7(32'hb9624d91),
	.w8(32'hbd10a81d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7e7a3),
	.w1(32'hbbda79c0),
	.w2(32'hbb161d41),
	.w3(32'h3c694882),
	.w4(32'hb9270416),
	.w5(32'hbb1f76d6),
	.w6(32'hbc2586a7),
	.w7(32'hbbbda6d0),
	.w8(32'h3c861e29),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e56b9),
	.w1(32'h3b713293),
	.w2(32'hbc7658f1),
	.w3(32'h3b5b065a),
	.w4(32'hba024a43),
	.w5(32'hbb3ca6ae),
	.w6(32'hbb47e1d7),
	.w7(32'h3b78c3c6),
	.w8(32'h3b5db34f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54a6f4),
	.w1(32'hbb37e4b5),
	.w2(32'h3c26d36c),
	.w3(32'hbc9dd7df),
	.w4(32'h3b3eb28e),
	.w5(32'hbc9003f5),
	.w6(32'h3b4b85be),
	.w7(32'hbb30deae),
	.w8(32'h3c232771),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82fe5f),
	.w1(32'hb99d9ccd),
	.w2(32'hbc44f126),
	.w3(32'h3b0a851e),
	.w4(32'hbb9892f0),
	.w5(32'hb9f2a5d8),
	.w6(32'h3c250eb2),
	.w7(32'hbc22bc76),
	.w8(32'hbb174ade),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb29aba),
	.w1(32'h3bf3a14b),
	.w2(32'hbc9515e7),
	.w3(32'h3c0bdeba),
	.w4(32'h3c929b19),
	.w5(32'hbc64c9e8),
	.w6(32'hb9c91be3),
	.w7(32'h3aea9f44),
	.w8(32'hb9aa49e9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18d7c1),
	.w1(32'h3a21d0a1),
	.w2(32'h3cce8aca),
	.w3(32'hbbff4231),
	.w4(32'h3a330a82),
	.w5(32'h3bb7d35f),
	.w6(32'h37a3e93f),
	.w7(32'h3bdd36a3),
	.w8(32'h3c17ba00),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af83516),
	.w1(32'h3c17d37b),
	.w2(32'h3c3bf433),
	.w3(32'hb9fdf07b),
	.w4(32'hbb5526c5),
	.w5(32'h3b2ded7c),
	.w6(32'hbb9c6757),
	.w7(32'h3c1ae908),
	.w8(32'h3ad053b5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba957340),
	.w1(32'h3bcd5af7),
	.w2(32'hbc67579e),
	.w3(32'h3bbe9b44),
	.w4(32'hb9b80000),
	.w5(32'h3cce57e3),
	.w6(32'hbc9c7889),
	.w7(32'h3923db2a),
	.w8(32'h3ba173d7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee8b13),
	.w1(32'hb953ef04),
	.w2(32'h3c023df6),
	.w3(32'h3b947909),
	.w4(32'h3880d427),
	.w5(32'h3c12eb54),
	.w6(32'hbcba490e),
	.w7(32'hba4ee83d),
	.w8(32'h3bdaed8d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc143fbd),
	.w1(32'h3add9766),
	.w2(32'hbcc54c31),
	.w3(32'h3c1280d3),
	.w4(32'hb9d86828),
	.w5(32'hbd95def3),
	.w6(32'h3aa283f4),
	.w7(32'h3b095f3f),
	.w8(32'hbc895e7b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09f09f),
	.w1(32'h3d008ab7),
	.w2(32'hbc12955e),
	.w3(32'hbbaf3d83),
	.w4(32'hbc228b14),
	.w5(32'hbda8e816),
	.w6(32'h3b74c3b4),
	.w7(32'hbc202b19),
	.w8(32'hbc895f7d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a2628),
	.w1(32'hbc46bf63),
	.w2(32'hbcb778bf),
	.w3(32'h3bcb00d3),
	.w4(32'hb9965b8e),
	.w5(32'h3c122500),
	.w6(32'h3ba91839),
	.w7(32'hb9f40cd8),
	.w8(32'hbc53cb92),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1d2ea),
	.w1(32'hbc096169),
	.w2(32'h3c3eeafb),
	.w3(32'h3af92777),
	.w4(32'h3c5520a9),
	.w5(32'hbbd8e2d8),
	.w6(32'h3abcbf66),
	.w7(32'h3bac51b1),
	.w8(32'hbadcdbc9),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5306e1),
	.w1(32'h3c1a595c),
	.w2(32'h3c0e3e46),
	.w3(32'h3c5118cd),
	.w4(32'hbc44b7b9),
	.w5(32'h3b13204c),
	.w6(32'hbab719fe),
	.w7(32'h3ba8f51e),
	.w8(32'h3905f38d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0bcc9),
	.w1(32'h3b0fb2fc),
	.w2(32'h39aac746),
	.w3(32'h3bd57552),
	.w4(32'h3d028549),
	.w5(32'h3c7ebdd2),
	.w6(32'h3ba9aa88),
	.w7(32'h3a99a32e),
	.w8(32'hbb68d14f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba575f0),
	.w1(32'h3b18a4c9),
	.w2(32'hbb514de4),
	.w3(32'h3c118b4b),
	.w4(32'h3bb5e780),
	.w5(32'hbe158712),
	.w6(32'h3b793b50),
	.w7(32'hbd319204),
	.w8(32'hb9cfdf4e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc233a61),
	.w1(32'hbbf4b843),
	.w2(32'hbbc7b825),
	.w3(32'hb8837afd),
	.w4(32'hbc9f69b8),
	.w5(32'hbb166edc),
	.w6(32'h3bed5258),
	.w7(32'h3bb185ce),
	.w8(32'h3a826f64),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a3799),
	.w1(32'hbcbae9b1),
	.w2(32'hbcf61cec),
	.w3(32'h3c2d7890),
	.w4(32'h3c3e8ea3),
	.w5(32'hba008896),
	.w6(32'h3a3fe40f),
	.w7(32'h3ab197b7),
	.w8(32'hbc8c159f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4a7b0),
	.w1(32'h3b47e6c0),
	.w2(32'h3cc8d7c9),
	.w3(32'hbc2c6169),
	.w4(32'h3b9816dd),
	.w5(32'hb9bdc194),
	.w6(32'h3ae88f43),
	.w7(32'h3b7c8569),
	.w8(32'h3c16c7d4),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f22a4),
	.w1(32'hbc062c3a),
	.w2(32'hbcb0a18c),
	.w3(32'h3b67894e),
	.w4(32'h3c98ab0f),
	.w5(32'hbce297dd),
	.w6(32'h3b9b7d9b),
	.w7(32'h3c08d009),
	.w8(32'hba96d51c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb56a77),
	.w1(32'hbda012dd),
	.w2(32'hbcba0181),
	.w3(32'hbb23b790),
	.w4(32'h3c3ab0b4),
	.w5(32'hbc3823a5),
	.w6(32'h3c63dfd7),
	.w7(32'hb83498dc),
	.w8(32'hbb68604b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b363f2e),
	.w1(32'h3b888c62),
	.w2(32'h3c203245),
	.w3(32'h3c474943),
	.w4(32'h3c0d739b),
	.w5(32'h3bd1ec60),
	.w6(32'h3c0b4491),
	.w7(32'h3c8c75df),
	.w8(32'h3c0d9b93),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb875088),
	.w1(32'hbc0e69fb),
	.w2(32'hbc9dae89),
	.w3(32'hbba62d30),
	.w4(32'h3c0cd6e1),
	.w5(32'hbc6a3110),
	.w6(32'h3c238188),
	.w7(32'h3af13c28),
	.w8(32'h3c1bbfe8),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921e03d),
	.w1(32'h3bbcb5df),
	.w2(32'hbb8c9e15),
	.w3(32'h3d3a9317),
	.w4(32'h3b70bebc),
	.w5(32'hbbcbab94),
	.w6(32'h3af647ec),
	.w7(32'hbbae2ad3),
	.w8(32'h3a2b9923),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc176f0),
	.w1(32'hbbe967bd),
	.w2(32'h3cad47bd),
	.w3(32'h3c91ddb4),
	.w4(32'hbc8ab357),
	.w5(32'hbbccd231),
	.w6(32'h3b8700f1),
	.w7(32'h3d9c45b1),
	.w8(32'hba95e594),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f60cc5),
	.w1(32'hbbf2756d),
	.w2(32'hbc514384),
	.w3(32'hbbee7b6a),
	.w4(32'hbdcd7d8b),
	.w5(32'hbbc005ec),
	.w6(32'hb9ed8de5),
	.w7(32'hbbeed93e),
	.w8(32'h3b40fbae),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41197a),
	.w1(32'hbc336387),
	.w2(32'hbc227d89),
	.w3(32'hbb0f2e3a),
	.w4(32'h3adfc9ce),
	.w5(32'hbb5a161b),
	.w6(32'h3cfed500),
	.w7(32'hbbf72a11),
	.w8(32'hbcfe83d5),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e83a),
	.w1(32'hbad08467),
	.w2(32'h3ad202af),
	.w3(32'h3b89888e),
	.w4(32'h3bfa7f92),
	.w5(32'hbba492f5),
	.w6(32'hbb316b6f),
	.w7(32'h3b8a835e),
	.w8(32'h3b61dbfa),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a3416),
	.w1(32'h3ae256a5),
	.w2(32'hbc17315c),
	.w3(32'hbc6c1850),
	.w4(32'hbb1ea92e),
	.w5(32'h3c917f8e),
	.w6(32'hbbd67a2a),
	.w7(32'hbd1c8485),
	.w8(32'h3c20d743),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bbad5),
	.w1(32'hbd4bb711),
	.w2(32'h3b3e5608),
	.w3(32'h3bb721ae),
	.w4(32'hbcc48e6e),
	.w5(32'h3bacb2b4),
	.w6(32'hbcad2bda),
	.w7(32'h3ba2f283),
	.w8(32'h3c010bd6),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf58204),
	.w1(32'hba3e01f6),
	.w2(32'hbba967ed),
	.w3(32'h3cb1fcaa),
	.w4(32'h3ab55f14),
	.w5(32'h3bfbf013),
	.w6(32'h3b12237c),
	.w7(32'hbc83d8f0),
	.w8(32'hbbcc6c93),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5c89b),
	.w1(32'hbbd3924b),
	.w2(32'hbd1e856d),
	.w3(32'hbb7a42a8),
	.w4(32'hb949aae5),
	.w5(32'hb8bd33df),
	.w6(32'h3c4da6d3),
	.w7(32'h3b90e5eb),
	.w8(32'h3c1d68b1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc92d3),
	.w1(32'h3ac64632),
	.w2(32'hbc272bc3),
	.w3(32'h3afb122b),
	.w4(32'hbc6e57b8),
	.w5(32'hbc133d9a),
	.w6(32'hbcb42770),
	.w7(32'hbb633ab0),
	.w8(32'hbc85895d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558ccd),
	.w1(32'h3be9d787),
	.w2(32'hbaf225bc),
	.w3(32'h3c3fced5),
	.w4(32'hbcb73a34),
	.w5(32'h3bec2cf5),
	.w6(32'h3d771259),
	.w7(32'hbc824abb),
	.w8(32'h3d511258),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8102a6),
	.w1(32'hbb3cff17),
	.w2(32'hbc8f464a),
	.w3(32'hba05f7b3),
	.w4(32'h3c88a256),
	.w5(32'h3be5401c),
	.w6(32'h3c619932),
	.w7(32'h3bb7c8b7),
	.w8(32'hbb6285b8),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2472fe),
	.w1(32'hbb21a28f),
	.w2(32'hbcdb8588),
	.w3(32'hbb223df5),
	.w4(32'h3c161471),
	.w5(32'hbcc08a44),
	.w6(32'hbcb27e23),
	.w7(32'hbca202fc),
	.w8(32'hbc29aed4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77043c),
	.w1(32'h3c10caf9),
	.w2(32'h3c84ba0d),
	.w3(32'h3bf78088),
	.w4(32'hbba9dcb0),
	.w5(32'hbb871f0c),
	.w6(32'hbac7c6de),
	.w7(32'hbbfa59b7),
	.w8(32'h3b8fc7f7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08aa5c),
	.w1(32'hbc2c7026),
	.w2(32'h39dfa410),
	.w3(32'hbbc80b10),
	.w4(32'hbbe93cf1),
	.w5(32'h3b622ab7),
	.w6(32'hbb78e6cd),
	.w7(32'h3b8e70c1),
	.w8(32'h3b5d014c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d1b2b),
	.w1(32'hbb01cbca),
	.w2(32'h3d09aac0),
	.w3(32'hba512f82),
	.w4(32'h3bf3ff50),
	.w5(32'hbc94a0de),
	.w6(32'hbdba8f11),
	.w7(32'h3b85cfa9),
	.w8(32'hbb800188),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd064e6a),
	.w1(32'hbc110d63),
	.w2(32'h3a13be47),
	.w3(32'hba3fbb19),
	.w4(32'hbca5e542),
	.w5(32'h3b6c55ca),
	.w6(32'h3be6cf55),
	.w7(32'hbb3e4daa),
	.w8(32'h3b95e0ab),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6c72),
	.w1(32'h3cacd296),
	.w2(32'h3bc2b66f),
	.w3(32'h3a90a320),
	.w4(32'hbb9c79d5),
	.w5(32'h3a6ea414),
	.w6(32'h3973f241),
	.w7(32'h3be89dc1),
	.w8(32'hbb54906c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23a1d6),
	.w1(32'hbb30dd04),
	.w2(32'hbb32fc5c),
	.w3(32'hbdebcc1e),
	.w4(32'hb8c3014e),
	.w5(32'h3b1bb913),
	.w6(32'hbbefa509),
	.w7(32'h3b937e5e),
	.w8(32'h397e6854),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc801115),
	.w1(32'h3a5e6b2b),
	.w2(32'h3cb36f1a),
	.w3(32'hbbba7e23),
	.w4(32'h3c180284),
	.w5(32'hbc967352),
	.w6(32'h3b80823e),
	.w7(32'h3d17e938),
	.w8(32'hbc84c95b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd54a0f),
	.w1(32'hb90d283e),
	.w2(32'hbcc30073),
	.w3(32'hbb549cd0),
	.w4(32'hbc7918f4),
	.w5(32'h3bcf269f),
	.w6(32'h3c32a62f),
	.w7(32'h3b978dcc),
	.w8(32'hbc16c141),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d02005f),
	.w1(32'hbbf5944a),
	.w2(32'hbcaf03ac),
	.w3(32'h3ac388cd),
	.w4(32'h39a04fe1),
	.w5(32'hbb8b7710),
	.w6(32'h3c3dd214),
	.w7(32'hbb4794ef),
	.w8(32'h3ba24f1d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89403b),
	.w1(32'hb8a33188),
	.w2(32'h3b7357e9),
	.w3(32'hbbb105ca),
	.w4(32'h3bced21a),
	.w5(32'hbab13dab),
	.w6(32'hbac08091),
	.w7(32'hbb6a62ce),
	.w8(32'hbcacfd02),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3377dd),
	.w1(32'hbbaa6a3b),
	.w2(32'hba3aa64c),
	.w3(32'hbc540045),
	.w4(32'hbd63456c),
	.w5(32'h3bf19d4d),
	.w6(32'hbc14ebef),
	.w7(32'h3b3559d4),
	.w8(32'hbb90d997),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4feab6),
	.w1(32'h3c26453c),
	.w2(32'h3b5b7b41),
	.w3(32'h3c0fbc72),
	.w4(32'h3b3ff63d),
	.w5(32'hbc23d1c0),
	.w6(32'hbc01c217),
	.w7(32'hbbbb68bd),
	.w8(32'hbd61eee1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c890dde),
	.w1(32'h3bb8f4a8),
	.w2(32'hbc17f858),
	.w3(32'hbc962857),
	.w4(32'hbb965d5e),
	.w5(32'h3bdee51e),
	.w6(32'hbc0d2781),
	.w7(32'hbbeb82d8),
	.w8(32'hbc027358),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32d88d),
	.w1(32'h3a631827),
	.w2(32'hbcfea33a),
	.w3(32'hbba0a57b),
	.w4(32'hb9f768fe),
	.w5(32'h3c0765a9),
	.w6(32'hbc162320),
	.w7(32'hbc6ee063),
	.w8(32'h3c492789),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd50a),
	.w1(32'hbbb71869),
	.w2(32'hbc188395),
	.w3(32'hbd947260),
	.w4(32'hbb4bd54e),
	.w5(32'h3bc81498),
	.w6(32'h3c29e9b7),
	.w7(32'hbbb9bfb8),
	.w8(32'h3c78d95d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bcae0),
	.w1(32'h3c645642),
	.w2(32'hbc24ed63),
	.w3(32'h3b9620e3),
	.w4(32'hbbb271a2),
	.w5(32'hbb1dd8cf),
	.w6(32'h3ac24ca2),
	.w7(32'hbd2297b4),
	.w8(32'hbcac40e5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba180d5a),
	.w1(32'hb956fbc4),
	.w2(32'h3b0851e5),
	.w3(32'h3ad96b7c),
	.w4(32'hba21215a),
	.w5(32'hbb840605),
	.w6(32'hbc2224cd),
	.w7(32'h3c034ead),
	.w8(32'hbc38192e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b852e53),
	.w1(32'h3b094921),
	.w2(32'hbb8168d2),
	.w3(32'h3bc2e189),
	.w4(32'hbc6f1fc9),
	.w5(32'hbb81c585),
	.w6(32'h3a858a94),
	.w7(32'hba19ecbc),
	.w8(32'h3c4fab7f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82a915),
	.w1(32'hbae9e395),
	.w2(32'hbc6881bd),
	.w3(32'hbbb762e2),
	.w4(32'h3b68fe62),
	.w5(32'hbc77a675),
	.w6(32'hba4f53d8),
	.w7(32'hbc0c278e),
	.w8(32'hba447cc6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0001e8),
	.w1(32'hbc84b7ba),
	.w2(32'hbb725ff5),
	.w3(32'h3c753f86),
	.w4(32'h3c36b419),
	.w5(32'h3c73a0a3),
	.w6(32'hbb57321e),
	.w7(32'h3b3adf6e),
	.w8(32'h3c97a71e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e7046),
	.w1(32'hbd21609e),
	.w2(32'hbd39504b),
	.w3(32'h3c5e7e95),
	.w4(32'h3bf56344),
	.w5(32'h3c898806),
	.w6(32'hb8b5d638),
	.w7(32'hbb672c4b),
	.w8(32'h3d4acc24),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbf991),
	.w1(32'hbbdf99d4),
	.w2(32'hbca6ac70),
	.w3(32'h3c1d7773),
	.w4(32'hbb965320),
	.w5(32'hbc743ac5),
	.w6(32'h3c01c56d),
	.w7(32'hbc20130d),
	.w8(32'hbc810345),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f0d32),
	.w1(32'hbbaf0e1f),
	.w2(32'hbbc1dd76),
	.w3(32'hbc284cd7),
	.w4(32'hba009590),
	.w5(32'hbc19039b),
	.w6(32'hba98907e),
	.w7(32'hbc9a7178),
	.w8(32'h3ade18eb),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe83c9a),
	.w1(32'hbb653217),
	.w2(32'hbba12577),
	.w3(32'h3ab9cd98),
	.w4(32'h3b8ef140),
	.w5(32'h3ace80f3),
	.w6(32'h3b1b9226),
	.w7(32'h3bba1938),
	.w8(32'hbbe4f9c2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9084e),
	.w1(32'h3bf35289),
	.w2(32'hbb0a11cf),
	.w3(32'h3c6923b5),
	.w4(32'h3cabf297),
	.w5(32'hbb9b46da),
	.w6(32'hbbd24921),
	.w7(32'hbb8c835f),
	.w8(32'hbb81e3fc),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c319401),
	.w1(32'h3b77cb3b),
	.w2(32'hbc23f1c0),
	.w3(32'h3aa6e47c),
	.w4(32'hbb2ee0f5),
	.w5(32'h3af5cd21),
	.w6(32'hbbdae363),
	.w7(32'h3a4a93ba),
	.w8(32'h3a4cd457),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6759d2),
	.w1(32'hbbc1d125),
	.w2(32'hbcdae179),
	.w3(32'h3b2754cb),
	.w4(32'hbaa295d9),
	.w5(32'h3b5ca695),
	.w6(32'hbc092aaf),
	.w7(32'hbb34698f),
	.w8(32'h3bbf6ea2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8bf5f),
	.w1(32'hbd6bafa5),
	.w2(32'hbc67ffa5),
	.w3(32'h3c03977b),
	.w4(32'h3b46baa0),
	.w5(32'hbac7b771),
	.w6(32'h3aff486a),
	.w7(32'h3c6e5252),
	.w8(32'h3ad17620),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d1b45),
	.w1(32'h3b02ca0d),
	.w2(32'h3b926cc0),
	.w3(32'hbb97296e),
	.w4(32'hbca21b24),
	.w5(32'h3b2e6207),
	.w6(32'hbbae7e90),
	.w7(32'h3c7d65dc),
	.w8(32'h3a309d6d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cb59f),
	.w1(32'hbd11a7d0),
	.w2(32'h3d003d0e),
	.w3(32'hbc6e2b11),
	.w4(32'hbb054943),
	.w5(32'h3b83f538),
	.w6(32'hb94e9fd3),
	.w7(32'hbb7d427c),
	.w8(32'hbc195fbe),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a91c0),
	.w1(32'hbc659627),
	.w2(32'h3ac2b356),
	.w3(32'h3a0a9d5e),
	.w4(32'h3ba8e96c),
	.w5(32'hbc8004e3),
	.w6(32'h3b82848b),
	.w7(32'hbc161a1f),
	.w8(32'hbc83d843),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3df29),
	.w1(32'hbc92a2a4),
	.w2(32'hbc2119f8),
	.w3(32'h3c203481),
	.w4(32'hbb9bf3fe),
	.w5(32'hba870e8f),
	.w6(32'hbc24142e),
	.w7(32'h3b462f4f),
	.w8(32'hbc5eb280),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30dd29),
	.w1(32'hbb5397a5),
	.w2(32'h3ba66ebc),
	.w3(32'hbc6508cc),
	.w4(32'hbc89ce38),
	.w5(32'h3ca87d83),
	.w6(32'hbb6ad67b),
	.w7(32'h3b0607e6),
	.w8(32'h3c9dd56d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02a7c7),
	.w1(32'h3a8eec09),
	.w2(32'h3aedfdd7),
	.w3(32'hbaf2f2d0),
	.w4(32'hbb8db4c6),
	.w5(32'h3aba9882),
	.w6(32'hbc0b9612),
	.w7(32'hbaac07b5),
	.w8(32'h3ae40459),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44210f),
	.w1(32'hbba50dd2),
	.w2(32'hbc89d507),
	.w3(32'h3a3a829c),
	.w4(32'h3bf72588),
	.w5(32'hbb57163a),
	.w6(32'h3a1b0e67),
	.w7(32'h3c0561fb),
	.w8(32'hbc827e22),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd2c8b),
	.w1(32'hbc8152f3),
	.w2(32'hbc801716),
	.w3(32'h3cdbb614),
	.w4(32'hbbce4382),
	.w5(32'hbccdacda),
	.w6(32'hbcb1793c),
	.w7(32'hbb1708fd),
	.w8(32'h3c5c91f9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17c22c),
	.w1(32'h3af0aae6),
	.w2(32'hbba3b96d),
	.w3(32'h3b4f3541),
	.w4(32'hbc2431dd),
	.w5(32'hbc15dfcd),
	.w6(32'h3c0235d9),
	.w7(32'hbbd58735),
	.w8(32'h3bc5c74a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17f1e9),
	.w1(32'h3bdf1b93),
	.w2(32'hbba75e5f),
	.w3(32'h3bc38853),
	.w4(32'h3a244db6),
	.w5(32'h3ac7e98c),
	.w6(32'h3b5a803d),
	.w7(32'h3b382a5b),
	.w8(32'h3b5b4208),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01a8bc),
	.w1(32'h3bbd658c),
	.w2(32'hbbfbda04),
	.w3(32'h3bf96d81),
	.w4(32'hba57646d),
	.w5(32'h3afda09a),
	.w6(32'hbb43d0a2),
	.w7(32'hbc20904a),
	.w8(32'hbc8802f9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1e451),
	.w1(32'hbb05e4c5),
	.w2(32'hbaa09504),
	.w3(32'h3b5126fc),
	.w4(32'hbc026e57),
	.w5(32'h3af17b9b),
	.w6(32'hba1eaf96),
	.w7(32'h3c643d01),
	.w8(32'hba3815a1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd41ac8),
	.w1(32'h3b99f62f),
	.w2(32'hba3a845b),
	.w3(32'hbba1f4b8),
	.w4(32'h3bff08e4),
	.w5(32'hb8f35366),
	.w6(32'h3b4558ef),
	.w7(32'hbab96285),
	.w8(32'h3b74ccfe),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d5434),
	.w1(32'hbb293283),
	.w2(32'hbbaf7a2c),
	.w3(32'h3b7f3162),
	.w4(32'hbbeec52f),
	.w5(32'h3c09d576),
	.w6(32'h3c210c90),
	.w7(32'h389b99ec),
	.w8(32'hbc283e7f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb413f3),
	.w1(32'h3cad0558),
	.w2(32'h3cb61f64),
	.w3(32'hbcd5d6f4),
	.w4(32'h3bc7d19f),
	.w5(32'h3c48639d),
	.w6(32'hba9ce8ee),
	.w7(32'hbbcac37c),
	.w8(32'h3b9680d0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf09ef),
	.w1(32'h3c9b7448),
	.w2(32'h3be1edbe),
	.w3(32'hbb213d23),
	.w4(32'hb98157c4),
	.w5(32'hbb87184b),
	.w6(32'h3b6d4843),
	.w7(32'h3b44532d),
	.w8(32'h3c805b71),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cf0d9),
	.w1(32'hbc8733fe),
	.w2(32'hbc08bd55),
	.w3(32'h3bb69ea0),
	.w4(32'h3c1163e4),
	.w5(32'h3bbf9988),
	.w6(32'h3c6ac814),
	.w7(32'h3b5c607e),
	.w8(32'hbc7ad46e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ffc4f),
	.w1(32'h3b83c141),
	.w2(32'hbb6c4827),
	.w3(32'h3a851f20),
	.w4(32'hbd144f5a),
	.w5(32'hbbacb0e1),
	.w6(32'hbafa4788),
	.w7(32'hba9b4e25),
	.w8(32'h3c2d7fcc),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d9320),
	.w1(32'hbb82a180),
	.w2(32'hbad169dd),
	.w3(32'hbb212c0e),
	.w4(32'hbac37b8b),
	.w5(32'h3b89444d),
	.w6(32'h3b2f8300),
	.w7(32'hba876df0),
	.w8(32'hbc7b8d30),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcead9f),
	.w1(32'hbc17c106),
	.w2(32'hbb25093c),
	.w3(32'hbcf8adb6),
	.w4(32'hbc5736cd),
	.w5(32'h3d57a47f),
	.w6(32'h3b01cee6),
	.w7(32'h3b29ffe2),
	.w8(32'h3bbf8b64),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09960e),
	.w1(32'h3cd5f883),
	.w2(32'h3ab49dad),
	.w3(32'h3c35f410),
	.w4(32'hbc0151b8),
	.w5(32'h3c0b9f77),
	.w6(32'hbbac5ca9),
	.w7(32'h3c4d3b57),
	.w8(32'h3a9e7fb6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0090cf),
	.w1(32'h3cdf3e71),
	.w2(32'h3b950e8d),
	.w3(32'hbc45f362),
	.w4(32'hbb7fc3e0),
	.w5(32'hbb6984ca),
	.w6(32'hbc5400f3),
	.w7(32'hbbf8218d),
	.w8(32'hbbb6b79f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc226682),
	.w1(32'h3b58b61e),
	.w2(32'h3c0361d3),
	.w3(32'hbbb0e61d),
	.w4(32'hba997576),
	.w5(32'hbbc3ae62),
	.w6(32'h3b4cf715),
	.w7(32'h3cdb103a),
	.w8(32'hbb62d535),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c550df9),
	.w1(32'hb950eac6),
	.w2(32'h3bc00d07),
	.w3(32'hbb5ea561),
	.w4(32'hbb2dad94),
	.w5(32'h3b62ee1f),
	.w6(32'h3b2dbb9c),
	.w7(32'h3b9969e2),
	.w8(32'h3b4fc649),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e324e),
	.w1(32'h3bc00b52),
	.w2(32'h3bba6ae5),
	.w3(32'h3bb117cd),
	.w4(32'hbba6f083),
	.w5(32'h3c778076),
	.w6(32'h3b52c9bc),
	.w7(32'hbc5298e8),
	.w8(32'h3d839466),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9fc12e),
	.w1(32'h3b80c474),
	.w2(32'h3bb04d86),
	.w3(32'h3b495aef),
	.w4(32'hbb68879e),
	.w5(32'hbbd08169),
	.w6(32'h3b0f363d),
	.w7(32'h3ab9075d),
	.w8(32'h3b3fc810),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa79e),
	.w1(32'hb9d0aab9),
	.w2(32'hbc1e7b07),
	.w3(32'h3b472774),
	.w4(32'h3c337c93),
	.w5(32'hbbc60a1c),
	.w6(32'hba6241df),
	.w7(32'hbaeb2b47),
	.w8(32'h3b872c73),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4c03b),
	.w1(32'hbc3b9958),
	.w2(32'hbc25b56a),
	.w3(32'h3b143880),
	.w4(32'h3bab728f),
	.w5(32'h3bd68c3a),
	.w6(32'h3b2b87c9),
	.w7(32'h3bb87aee),
	.w8(32'h3ae51640),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad10d6c),
	.w1(32'hbb92d5d7),
	.w2(32'h3b4b2829),
	.w3(32'hb9e21d73),
	.w4(32'h3c75db11),
	.w5(32'hbb681b65),
	.w6(32'hbbbf7941),
	.w7(32'h3a1a37f4),
	.w8(32'h3cfe939b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba34d7e),
	.w1(32'hbb1f75e1),
	.w2(32'hb98bf08a),
	.w3(32'hbbeb1c31),
	.w4(32'hbbd9ef18),
	.w5(32'hbab4f4ed),
	.w6(32'h3b1d4876),
	.w7(32'hbd1e9117),
	.w8(32'hbabbf443),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1812f),
	.w1(32'h3bc0213e),
	.w2(32'h3b831849),
	.w3(32'h3b93d649),
	.w4(32'hbbf3dbd9),
	.w5(32'hbcb23df1),
	.w6(32'h3c8301ad),
	.w7(32'hbb4e1916),
	.w8(32'hbc38b1e3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c960663),
	.w1(32'h3bda7126),
	.w2(32'hbc425998),
	.w3(32'hbd0a488b),
	.w4(32'h3af8b7e9),
	.w5(32'hbc30ede8),
	.w6(32'h3c151637),
	.w7(32'hbbc8db7c),
	.w8(32'hbc88004f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde502a),
	.w1(32'h3cc53fc9),
	.w2(32'h3b87e6b5),
	.w3(32'h3c1ae67d),
	.w4(32'h3bc0ea7b),
	.w5(32'hbbfee5bd),
	.w6(32'h3c35a47b),
	.w7(32'hbbb61a15),
	.w8(32'hba663d20),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf79f99),
	.w1(32'hbb93de70),
	.w2(32'hbd4ef993),
	.w3(32'hbb5b6431),
	.w4(32'h3cd48232),
	.w5(32'h3b480f83),
	.w6(32'hbaefb4d7),
	.w7(32'h3c868cf5),
	.w8(32'hbb2ee12d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb332b6),
	.w1(32'h39b7fc8f),
	.w2(32'hba18b5ce),
	.w3(32'h3bb4c4bc),
	.w4(32'hbc23badb),
	.w5(32'h3b6fc765),
	.w6(32'h3bbfa755),
	.w7(32'hbad2275c),
	.w8(32'h3c49fc2d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad058c8),
	.w1(32'hbc4eeb89),
	.w2(32'h3be0cc45),
	.w3(32'h3c06c701),
	.w4(32'h3c829732),
	.w5(32'hbc769142),
	.w6(32'hbb893e64),
	.w7(32'hbbc36f78),
	.w8(32'hb9dd2416),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a967b0c),
	.w1(32'h3b82a901),
	.w2(32'hbc32ecf5),
	.w3(32'hbc9eb370),
	.w4(32'hbb2728bb),
	.w5(32'h3bc908fa),
	.w6(32'h3c2d9cc2),
	.w7(32'h3c0941fb),
	.w8(32'hbccc57a7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dbed6),
	.w1(32'h3c0e6f20),
	.w2(32'hbc7d452e),
	.w3(32'h3cf42017),
	.w4(32'h3a494c82),
	.w5(32'hbc916975),
	.w6(32'h3c201784),
	.w7(32'hbaa1ed52),
	.w8(32'hbc7499ec),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c945dbc),
	.w1(32'h3c03e5e7),
	.w2(32'hbb94ee5e),
	.w3(32'hbba147a8),
	.w4(32'h3c2c33b9),
	.w5(32'h3c6ef18d),
	.w6(32'h3c6f514d),
	.w7(32'h3c35a748),
	.w8(32'h3b139e12),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b101c3d),
	.w1(32'h3c0ea31c),
	.w2(32'h3c47324e),
	.w3(32'hbcd80ca1),
	.w4(32'hbcaaf80f),
	.w5(32'hbc4777c5),
	.w6(32'hbb2e5f97),
	.w7(32'hbb1c2aa2),
	.w8(32'hbbf40a64),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe0082),
	.w1(32'hba740467),
	.w2(32'h3be81d82),
	.w3(32'hbc6a765b),
	.w4(32'hbbe75c96),
	.w5(32'hbba88201),
	.w6(32'hbbf24a30),
	.w7(32'h3aac5f3c),
	.w8(32'h3cca2ed1),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be52360),
	.w1(32'h3b06505a),
	.w2(32'h3c09ba80),
	.w3(32'h3c9bb037),
	.w4(32'h3bc1779e),
	.w5(32'hbb2c10c5),
	.w6(32'h3a884a0e),
	.w7(32'h3c60a5b1),
	.w8(32'h3aa9600c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad38366),
	.w1(32'h3b7443a1),
	.w2(32'hbbbc86e2),
	.w3(32'h3a547338),
	.w4(32'h39a8f973),
	.w5(32'hbb3ff1e9),
	.w6(32'hbacb3032),
	.w7(32'hbb24c8b5),
	.w8(32'hba7f2661),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c800b37),
	.w1(32'hbadeaa7d),
	.w2(32'hbc0a737e),
	.w3(32'hbb8fe30b),
	.w4(32'h39da719e),
	.w5(32'hba7e234f),
	.w6(32'hbb15e063),
	.w7(32'hbc0421e0),
	.w8(32'h3ac95171),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb153a24),
	.w1(32'hba782876),
	.w2(32'h3a25a8aa),
	.w3(32'h3aed4a38),
	.w4(32'h3d206631),
	.w5(32'hbbeb5c0e),
	.w6(32'hbb8396f0),
	.w7(32'h3b5304ad),
	.w8(32'h3b11a635),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33668c),
	.w1(32'hb916994f),
	.w2(32'hbb284da7),
	.w3(32'hbb804e47),
	.w4(32'hbca14ec5),
	.w5(32'h3c75cca0),
	.w6(32'hbb4ce9ec),
	.w7(32'hbbdf9ef4),
	.w8(32'hbc29004b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d02f2),
	.w1(32'h3c08f35f),
	.w2(32'hbb914371),
	.w3(32'h3bcb3e8c),
	.w4(32'h3c758b8b),
	.w5(32'hbc551733),
	.w6(32'hbaa610f3),
	.w7(32'hba392e89),
	.w8(32'h3ae14969),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87d4c1),
	.w1(32'h3c838d98),
	.w2(32'h3c15ebe4),
	.w3(32'h38afe8ed),
	.w4(32'hbb28da5e),
	.w5(32'hbba66b92),
	.w6(32'hbc3a643f),
	.w7(32'h3b2179cc),
	.w8(32'hbc869254),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4afd7),
	.w1(32'h3c1cfdbb),
	.w2(32'hbaa93c1d),
	.w3(32'h3be3a17c),
	.w4(32'hbaf46e07),
	.w5(32'hbba6c46d),
	.w6(32'h3c1268a3),
	.w7(32'hbc50a685),
	.w8(32'h3c3527e4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caad382),
	.w1(32'h3c1d4cff),
	.w2(32'hbc9efde1),
	.w3(32'hbbd7a80a),
	.w4(32'h3c087433),
	.w5(32'h3c828308),
	.w6(32'h3c3c4ace),
	.w7(32'hbc6fee07),
	.w8(32'hbd55d23e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9fc4aa),
	.w1(32'h3c1695d8),
	.w2(32'hbc9bb9be),
	.w3(32'hba8a9512),
	.w4(32'h3c59e452),
	.w5(32'hbc3b9bd1),
	.w6(32'hbb9ab2bb),
	.w7(32'h3c540dac),
	.w8(32'hbc8d69b0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc36a46),
	.w1(32'hba770d9f),
	.w2(32'h3becaf72),
	.w3(32'h3bded635),
	.w4(32'h3c8aeba5),
	.w5(32'h3b3cd49f),
	.w6(32'h3b38e427),
	.w7(32'h3b1ab391),
	.w8(32'hbc429b48),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0b26b),
	.w1(32'h3bd1e57a),
	.w2(32'hbd3fe15a),
	.w3(32'h3b9a7f9d),
	.w4(32'hbbad2401),
	.w5(32'hbc199fec),
	.w6(32'h3b480438),
	.w7(32'hbb9861e5),
	.w8(32'hbca2231f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc07ed7),
	.w1(32'h3b526ad8),
	.w2(32'hbc259ed3),
	.w3(32'hbb311557),
	.w4(32'h3c25ff55),
	.w5(32'hbbf6fb24),
	.w6(32'hbb49108d),
	.w7(32'h3c1fdd0f),
	.w8(32'h3c6cb52c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f5f88),
	.w1(32'hbae82d97),
	.w2(32'h3c5346be),
	.w3(32'h3b3558b2),
	.w4(32'hba0bab82),
	.w5(32'hbc78c806),
	.w6(32'hbbe3e003),
	.w7(32'h3c3b4236),
	.w8(32'hbbea47cd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbde76f),
	.w1(32'h3c195e69),
	.w2(32'h3c24b135),
	.w3(32'hbb83fc9b),
	.w4(32'h3bc19f0c),
	.w5(32'hbca9c364),
	.w6(32'h3bf628e2),
	.w7(32'hbc8a6778),
	.w8(32'h3b9aba2c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40b7d2),
	.w1(32'hbc0a501c),
	.w2(32'h3ad4b1a9),
	.w3(32'h3b7a80d3),
	.w4(32'hb9a3563a),
	.w5(32'hbc02ca4f),
	.w6(32'hbc58188f),
	.w7(32'h3984083a),
	.w8(32'hbaa35ff5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b225b92),
	.w1(32'h3c230028),
	.w2(32'h3cca322f),
	.w3(32'hba93b7eb),
	.w4(32'hbc5a0c29),
	.w5(32'h3baba896),
	.w6(32'h3a4c469a),
	.w7(32'hb9c14b63),
	.w8(32'hb98263dc),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43a04c),
	.w1(32'hbc97c09a),
	.w2(32'hbcff6550),
	.w3(32'h3ba8daef),
	.w4(32'hbb99679d),
	.w5(32'hbc045634),
	.w6(32'hbbd168b4),
	.w7(32'hba4d48a6),
	.w8(32'hbc047362),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae23870),
	.w1(32'hbd038b4f),
	.w2(32'hbcdcdc1c),
	.w3(32'h3b38b9ff),
	.w4(32'h3c4d17fe),
	.w5(32'hbc79b7b7),
	.w6(32'h3c258f2d),
	.w7(32'h3ab7b1a9),
	.w8(32'h3c344429),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca4cf6),
	.w1(32'hbc693bbf),
	.w2(32'hbd1f42db),
	.w3(32'hba6c0dbc),
	.w4(32'h38b5f617),
	.w5(32'hbbc54983),
	.w6(32'h3c94f013),
	.w7(32'h3aa4a511),
	.w8(32'hbb17d9db),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b4163),
	.w1(32'h3bdb43d7),
	.w2(32'h3ba6a5fd),
	.w3(32'h3baba973),
	.w4(32'h3b4fdacf),
	.w5(32'hbc3650b8),
	.w6(32'h3be9e213),
	.w7(32'hbc062771),
	.w8(32'hbb0d7967),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bcea1),
	.w1(32'hbc2fef28),
	.w2(32'h3c81d46b),
	.w3(32'h3ba9f925),
	.w4(32'h3b5ae3fe),
	.w5(32'h3baf6d05),
	.w6(32'hbb5ff176),
	.w7(32'hbb270791),
	.w8(32'hbc029d68),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39740afe),
	.w1(32'h3a748452),
	.w2(32'h3c7c10f5),
	.w3(32'h39e7b978),
	.w4(32'hbba769c9),
	.w5(32'h3c1f8dcb),
	.w6(32'hbb11ba35),
	.w7(32'h3c3f91f2),
	.w8(32'hbc815a0c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79179e),
	.w1(32'h3b0e13bc),
	.w2(32'h3cffa861),
	.w3(32'h39fa6520),
	.w4(32'h3c67fe79),
	.w5(32'hbba87a1a),
	.w6(32'h3c321133),
	.w7(32'h3c36b4dc),
	.w8(32'hbbbbdffb),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66ab15),
	.w1(32'hbc0ae48a),
	.w2(32'hb9af137f),
	.w3(32'hbbc9112f),
	.w4(32'h3b7d4dae),
	.w5(32'hbb89ea5c),
	.w6(32'hbc5062d6),
	.w7(32'h3a076d0a),
	.w8(32'hbccfb125),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003779),
	.w1(32'hbb9595b8),
	.w2(32'hbc6d82e8),
	.w3(32'hbbc19a46),
	.w4(32'hbc80f357),
	.w5(32'h3bb7d668),
	.w6(32'h3b8a1973),
	.w7(32'h3bbeebe8),
	.w8(32'hbba08904),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4141b8),
	.w1(32'h3c8851f8),
	.w2(32'h3a9e9f1f),
	.w3(32'hbc38d29c),
	.w4(32'hbc9c5fc2),
	.w5(32'hbc8ed4e5),
	.w6(32'hbbc07857),
	.w7(32'h3aa3c351),
	.w8(32'hbbe2bcd8),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e2170),
	.w1(32'hbb104108),
	.w2(32'hba63cef3),
	.w3(32'hbb0eeada),
	.w4(32'hbcda51f5),
	.w5(32'hbad75fd1),
	.w6(32'h3994a5ad),
	.w7(32'h3a82638f),
	.w8(32'h3a040db6),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb824d4b),
	.w1(32'h3cb2a3b0),
	.w2(32'hbbc98225),
	.w3(32'h3b3daaf5),
	.w4(32'hbc416fd0),
	.w5(32'h3bdbd397),
	.w6(32'h3b36e458),
	.w7(32'hbb0c01d0),
	.w8(32'h3b53cb82),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44d8cb),
	.w1(32'hbc0e4b9b),
	.w2(32'hbc03c43c),
	.w3(32'hbc095f3d),
	.w4(32'h3bc7c57c),
	.w5(32'h3bbf867a),
	.w6(32'hbb7cedd2),
	.w7(32'h3a5c1efb),
	.w8(32'hbc41f211),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47cbbf),
	.w1(32'hbc7d310e),
	.w2(32'h3b2c63f8),
	.w3(32'h3a8253a1),
	.w4(32'hbcb42206),
	.w5(32'hbb702e39),
	.w6(32'h3b45a2d6),
	.w7(32'hbc80f522),
	.w8(32'h3c293068),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cc5b1),
	.w1(32'hbc9a510b),
	.w2(32'hbcd544fd),
	.w3(32'hb9cbd30f),
	.w4(32'h3ce21dd6),
	.w5(32'hbc267225),
	.w6(32'h3c09e3d0),
	.w7(32'h3c9c09c9),
	.w8(32'hbba3b478),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaa3cd),
	.w1(32'hbc01688e),
	.w2(32'h3af5d3c3),
	.w3(32'h3b0a1a27),
	.w4(32'hbb863ac8),
	.w5(32'h3be4b248),
	.w6(32'h3c0cf018),
	.w7(32'hbbb89049),
	.w8(32'hbba49bd7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3195b),
	.w1(32'hbbae5a52),
	.w2(32'h3c4e3b36),
	.w3(32'h3afee9ca),
	.w4(32'hbbe744b0),
	.w5(32'hbc02d82e),
	.w6(32'h3c05321d),
	.w7(32'hbb29cb24),
	.w8(32'hbbed013d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule