module layer_10_featuremap_194(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4a445),
	.w1(32'h3bb2dd19),
	.w2(32'h3bef46fb),
	.w3(32'hbb62ff14),
	.w4(32'hbb7c6187),
	.w5(32'h3c36feb0),
	.w6(32'h3ca62160),
	.w7(32'h3c42072f),
	.w8(32'h39948952),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1fb5e),
	.w1(32'h3c072708),
	.w2(32'hbb590a9b),
	.w3(32'h3d0a9682),
	.w4(32'h3ba1967e),
	.w5(32'hbbb66e33),
	.w6(32'h3c650283),
	.w7(32'h3b2755f3),
	.w8(32'hbb0137ad),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b319a6d),
	.w1(32'h3b9f1b2e),
	.w2(32'h3b3e4349),
	.w3(32'h3b2502d3),
	.w4(32'hbab6fcdc),
	.w5(32'hbb150d96),
	.w6(32'h39cce917),
	.w7(32'hba37d85d),
	.w8(32'hbaeba421),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa41902),
	.w1(32'h3c19f405),
	.w2(32'hbc4b0fa9),
	.w3(32'hb998b181),
	.w4(32'hbc05f4cd),
	.w5(32'hbc994759),
	.w6(32'h3bd9cb76),
	.w7(32'hbc5abade),
	.w8(32'hbc1e6929),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0162e3),
	.w1(32'h3c00b43a),
	.w2(32'hbad5f4cc),
	.w3(32'hbc27f767),
	.w4(32'h3ab97b41),
	.w5(32'hbbc04c48),
	.w6(32'h39c01577),
	.w7(32'hbc2eb269),
	.w8(32'h3b4aced6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c5da5),
	.w1(32'h3a834e8c),
	.w2(32'hbb9720ec),
	.w3(32'h3abcb084),
	.w4(32'hbb1d06c3),
	.w5(32'hbb891315),
	.w6(32'hbb13011a),
	.w7(32'hbb3a25ad),
	.w8(32'hb86ec7fa),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8274dc),
	.w1(32'h3c11917f),
	.w2(32'h3d0b32ce),
	.w3(32'hbc863789),
	.w4(32'h3b5e01c7),
	.w5(32'h3d1d5342),
	.w6(32'hbcc513ec),
	.w7(32'hbbb534af),
	.w8(32'h3cd43fc9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06c1c8),
	.w1(32'h3c9bff77),
	.w2(32'h3d5b86d5),
	.w3(32'h3cdbc5bb),
	.w4(32'h3bdbae95),
	.w5(32'h3bd7c65c),
	.w6(32'h3cadfffa),
	.w7(32'h3c903a9a),
	.w8(32'h3c70f62c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba836ca1),
	.w1(32'hbb0773b5),
	.w2(32'h3ba72c16),
	.w3(32'hbb1188e5),
	.w4(32'hbacf81e0),
	.w5(32'h3bd393a6),
	.w6(32'h3b180066),
	.w7(32'h3b7ff30d),
	.w8(32'h3bcf394b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d260373),
	.w1(32'h3bc84728),
	.w2(32'h3d81c182),
	.w3(32'h3c960b52),
	.w4(32'hbcde42f0),
	.w5(32'h3ce9d9b0),
	.w6(32'hbba3dea4),
	.w7(32'hbcf65faa),
	.w8(32'h3c1b84bd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05b38a),
	.w1(32'h3c154bc2),
	.w2(32'h3bb52f35),
	.w3(32'h3b910745),
	.w4(32'h39c4e243),
	.w5(32'h3aac38dd),
	.w6(32'h3b9d2bd6),
	.w7(32'hbb934b31),
	.w8(32'hbac9b7c2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf674bf),
	.w1(32'hbcb3149a),
	.w2(32'h3d318ad8),
	.w3(32'h3c08bcba),
	.w4(32'hbcf8564d),
	.w5(32'h3cdd7976),
	.w6(32'hbc38e748),
	.w7(32'hbd2e2366),
	.w8(32'h3d00b309),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf1afb6),
	.w1(32'h3a4b13c3),
	.w2(32'h3d86507b),
	.w3(32'hbc142492),
	.w4(32'hbccdb3b0),
	.w5(32'h3d20a9df),
	.w6(32'hbca5c985),
	.w7(32'hbd15a858),
	.w8(32'h3c5dfa2b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ed449),
	.w1(32'h3c328369),
	.w2(32'h3c72a2c2),
	.w3(32'h3c26e3e8),
	.w4(32'h3bfad25a),
	.w5(32'h3c03a9c5),
	.w6(32'h3c5bda17),
	.w7(32'h3c34377d),
	.w8(32'h3b8c127e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67d008),
	.w1(32'h3bb4045e),
	.w2(32'hbbe583e8),
	.w3(32'h3bca6c5c),
	.w4(32'hbc65f73e),
	.w5(32'hbc9e0a4e),
	.w6(32'h3cac7b74),
	.w7(32'hbcce10a3),
	.w8(32'hbc494343),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d06fa79),
	.w1(32'h3ca17557),
	.w2(32'h3d477e29),
	.w3(32'hbc5f4f9a),
	.w4(32'hbc494368),
	.w5(32'h3cd21e7a),
	.w6(32'h3b05935c),
	.w7(32'hbb98c26c),
	.w8(32'h3cc2145c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc1c0c),
	.w1(32'h3b11a3a9),
	.w2(32'h3b7324a2),
	.w3(32'h3b89eab4),
	.w4(32'h3aa1ec75),
	.w5(32'h3a88c9c7),
	.w6(32'hbb897a77),
	.w7(32'hbb93f7d5),
	.w8(32'hbbc449ca),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99762c),
	.w1(32'h3be5638d),
	.w2(32'h3d902f5d),
	.w3(32'hbb87c8de),
	.w4(32'hbca2a1f3),
	.w5(32'h3d363f5b),
	.w6(32'hbb2ba14f),
	.w7(32'hbc0429cd),
	.w8(32'h3d05ff23),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8610bb),
	.w1(32'h3b64299a),
	.w2(32'h3d1d44b8),
	.w3(32'hbb730347),
	.w4(32'hbc82b3fb),
	.w5(32'h3cccf427),
	.w6(32'hbb8d8bd0),
	.w7(32'hbc804b3e),
	.w8(32'h3c58f3fb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b199b81),
	.w1(32'hbaf5ad5a),
	.w2(32'h3b574b08),
	.w3(32'hbb1686c2),
	.w4(32'hba812521),
	.w5(32'h3b3bd9a9),
	.w6(32'hb88f0da7),
	.w7(32'h3b4d35af),
	.w8(32'h3b34eb40),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35a969),
	.w1(32'hbb85bfd5),
	.w2(32'hbb630fb9),
	.w3(32'h3b06649f),
	.w4(32'hbb84ba94),
	.w5(32'hbb527200),
	.w6(32'hbb88b52d),
	.w7(32'hbb0c7f2c),
	.w8(32'hbb5f5fd1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e56bd),
	.w1(32'hbc6f50e0),
	.w2(32'h3c0817e0),
	.w3(32'hbb9dae6a),
	.w4(32'hbcc4f0d5),
	.w5(32'hbc6245ff),
	.w6(32'h3c1ca753),
	.w7(32'hbc104a70),
	.w8(32'hbc4a2a31),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd0f3b2),
	.w1(32'h3d033108),
	.w2(32'h3d849c4a),
	.w3(32'h3d9806bb),
	.w4(32'hbc95f41f),
	.w5(32'h3d5dbe44),
	.w6(32'h3d4a007d),
	.w7(32'h3b872a35),
	.w8(32'h3d61000c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1295ae),
	.w1(32'h3bb795e1),
	.w2(32'h3cfab175),
	.w3(32'h3c1f0d68),
	.w4(32'hbcbbcc89),
	.w5(32'h3be3bfbb),
	.w6(32'h3c4bf50b),
	.w7(32'hbd112520),
	.w8(32'hbc4e056e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d30a0f3),
	.w1(32'hbc670d7e),
	.w2(32'hbba4fbf2),
	.w3(32'h3cee0faf),
	.w4(32'hbc9508bf),
	.w5(32'hbc87bdf4),
	.w6(32'h3d09e86d),
	.w7(32'hbceb12af),
	.w8(32'hbd06cd2c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385f1dc5),
	.w1(32'h3bbc3e1e),
	.w2(32'h3c4f8237),
	.w3(32'h3af0960e),
	.w4(32'h3b130786),
	.w5(32'hbb349f1f),
	.w6(32'hbbc95bc1),
	.w7(32'h3b50949a),
	.w8(32'hbb163982),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb100aab),
	.w1(32'h39b419f0),
	.w2(32'hb755568a),
	.w3(32'hbba3384a),
	.w4(32'h39c150d7),
	.w5(32'hba1ed5e5),
	.w6(32'h3a08267e),
	.w7(32'h3a2d144e),
	.w8(32'h3aaceb41),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bdbc7),
	.w1(32'hbc89fab3),
	.w2(32'h3c436655),
	.w3(32'h3cd66cf6),
	.w4(32'hbb2834f5),
	.w5(32'hbc5ae14b),
	.w6(32'h3cd9a1be),
	.w7(32'hbc88e090),
	.w8(32'hbcc7cf3f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5aa35b),
	.w1(32'hbb0c4f39),
	.w2(32'h3c0c1789),
	.w3(32'h3be17add),
	.w4(32'hbb852fea),
	.w5(32'h3b9d5627),
	.w6(32'h3c8aa19e),
	.w7(32'h3c59cc63),
	.w8(32'h3b6e84d7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9edbbc),
	.w1(32'hbcf5c76d),
	.w2(32'hbc093e4f),
	.w3(32'h3a4aa0be),
	.w4(32'hbc83c1f8),
	.w5(32'hbc99eea0),
	.w6(32'h3b9a2a02),
	.w7(32'hbc819b90),
	.w8(32'hbd04c206),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e1528),
	.w1(32'hb9887c09),
	.w2(32'hbace6e56),
	.w3(32'h3b4ae681),
	.w4(32'h39c2ab92),
	.w5(32'hba5bed3b),
	.w6(32'hb7f8ccd6),
	.w7(32'h3a3331fa),
	.w8(32'hba82b60a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39dd31),
	.w1(32'h3aa5d648),
	.w2(32'h3824b5bc),
	.w3(32'hba9355b7),
	.w4(32'hba3c5098),
	.w5(32'hba37a97f),
	.w6(32'h3ac63083),
	.w7(32'h3a1cb3d0),
	.w8(32'hbab835c3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0bf97),
	.w1(32'h3bf2b28c),
	.w2(32'h3d1d0795),
	.w3(32'hbc1a169e),
	.w4(32'hbc1451dc),
	.w5(32'h3c800b7a),
	.w6(32'h3baa4d5c),
	.w7(32'hbb894159),
	.w8(32'h3ba76f92),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e25b4),
	.w1(32'h3c275c8c),
	.w2(32'h3c92a21d),
	.w3(32'h3c4d01be),
	.w4(32'h3bee40d9),
	.w5(32'h3b888f91),
	.w6(32'h3caba1a8),
	.w7(32'h3bf56a02),
	.w8(32'hba3fa4ba),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388e2d9c),
	.w1(32'hbb14a340),
	.w2(32'h3ba945d6),
	.w3(32'hbbb144bf),
	.w4(32'hbc2a226e),
	.w5(32'h3b431326),
	.w6(32'hbbb5c98e),
	.w7(32'h3aab15e9),
	.w8(32'h3b85790b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7a364),
	.w1(32'hbb75831c),
	.w2(32'h3cab6f8b),
	.w3(32'hba07eacf),
	.w4(32'hbc169a28),
	.w5(32'h3c532738),
	.w6(32'hbbda3b5d),
	.w7(32'hbbb1f685),
	.w8(32'h3c4a1f17),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d99a5d1),
	.w1(32'hbd00afe1),
	.w2(32'h3d82773a),
	.w3(32'h3da266e8),
	.w4(32'hbd48841e),
	.w5(32'h3d129100),
	.w6(32'h3cca98cf),
	.w7(32'hbda351ad),
	.w8(32'h3ccf6054),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3da81a5d),
	.w1(32'hbcef08b6),
	.w2(32'hbda7ccd7),
	.w3(32'h3d82b539),
	.w4(32'hbd01ee7d),
	.w5(32'hbdbc784a),
	.w6(32'h3ddc1a3a),
	.w7(32'hbc812b00),
	.w8(32'hbd80b453),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d329626),
	.w1(32'hbc557f8e),
	.w2(32'hbd4c89e2),
	.w3(32'h3d843894),
	.w4(32'h3ba77896),
	.w5(32'hbd21653c),
	.w6(32'h3dbd18a9),
	.w7(32'h3c825167),
	.w8(32'hbcabc835),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c9843),
	.w1(32'hbc0dfa1b),
	.w2(32'hbccf756c),
	.w3(32'h3c2861eb),
	.w4(32'hbc3ee712),
	.w5(32'hbcdfa025),
	.w6(32'h3c869d6f),
	.w7(32'hbc6881d5),
	.w8(32'hbcadeea0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6a45a),
	.w1(32'hbb3aae07),
	.w2(32'h3b190fbc),
	.w3(32'hbaedccb7),
	.w4(32'h3a16f508),
	.w5(32'h3b06a309),
	.w6(32'h3aed80f5),
	.w7(32'h3b273466),
	.w8(32'hba0834cd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dcf51a),
	.w1(32'hbb9f73b4),
	.w2(32'hbad3f691),
	.w3(32'h3ad6a252),
	.w4(32'h3b3afaee),
	.w5(32'h39e0de31),
	.w6(32'hbb61b14f),
	.w7(32'hbc2d203f),
	.w8(32'hbb2f866e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc06299),
	.w1(32'hbbbcef2f),
	.w2(32'hb9f85544),
	.w3(32'h3ca52601),
	.w4(32'hbbb5319e),
	.w5(32'h3a3bb956),
	.w6(32'h3cbb1700),
	.w7(32'hbacc554e),
	.w8(32'h3b6f366f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cead29d),
	.w1(32'hbaac994a),
	.w2(32'h3d85b4c4),
	.w3(32'h3c751606),
	.w4(32'hbcdadf1e),
	.w5(32'h3d0fb446),
	.w6(32'hbbe6a6bf),
	.w7(32'hbbf902ad),
	.w8(32'h3d22a344),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d370db4),
	.w1(32'hbb8d2b04),
	.w2(32'h3cea95f8),
	.w3(32'h3ca64b22),
	.w4(32'hbcb84c50),
	.w5(32'h3bd60047),
	.w6(32'h3cd2c350),
	.w7(32'hbcf7abf1),
	.w8(32'hbca1cbe7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d30106e),
	.w1(32'h3bd4ef70),
	.w2(32'h3d1b3f8c),
	.w3(32'h3c3b8e20),
	.w4(32'hbd2aab45),
	.w5(32'h3b5a563d),
	.w6(32'h3c876a4c),
	.w7(32'hbd256723),
	.w8(32'hbc77f2fe),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d31e92a),
	.w1(32'h3cd0dc5a),
	.w2(32'h3c93765c),
	.w3(32'h3cde4ec9),
	.w4(32'h3bf24675),
	.w5(32'hbba1250a),
	.w6(32'h3d246d34),
	.w7(32'hbc86712d),
	.w8(32'h3b8b28f4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca214c3),
	.w1(32'h3b2f2f2f),
	.w2(32'h3db5ac13),
	.w3(32'hbbe0eb5c),
	.w4(32'hbc621254),
	.w5(32'h3d8e9a21),
	.w6(32'hbccca067),
	.w7(32'hbc08da91),
	.w8(32'h3d1ba509),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf6d9a),
	.w1(32'h3ae9ca46),
	.w2(32'h3b94c663),
	.w3(32'h3a918dcd),
	.w4(32'h38f374ac),
	.w5(32'hb68d5f04),
	.w6(32'h3b8723e3),
	.w7(32'h3acf8108),
	.w8(32'hbac6f087),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1956a7),
	.w1(32'hbb9787f5),
	.w2(32'hbc108aa9),
	.w3(32'h3ab164c3),
	.w4(32'hba4328e4),
	.w5(32'hbb86d9bd),
	.w6(32'h3a9c6a82),
	.w7(32'hbb60d076),
	.w8(32'hbb495b5a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86dfcf),
	.w1(32'hbb885d26),
	.w2(32'h3aff7b41),
	.w3(32'hbb882fef),
	.w4(32'hbaa068d6),
	.w5(32'hbb11e0d3),
	.w6(32'hba5971c7),
	.w7(32'h3a800774),
	.w8(32'h3aae57e6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfd1d4b),
	.w1(32'h3c2019aa),
	.w2(32'h3cee4b11),
	.w3(32'h3b0a6dd9),
	.w4(32'h394038a6),
	.w5(32'h3cbf238c),
	.w6(32'hba5d733b),
	.w7(32'h3a890cb4),
	.w8(32'h3c57b1ed),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f79af),
	.w1(32'h39a31744),
	.w2(32'h3b9a9e2c),
	.w3(32'h3c38ac25),
	.w4(32'hbb89fd77),
	.w5(32'h3c4a278e),
	.w6(32'h3a21c17f),
	.w7(32'hbb907580),
	.w8(32'h3c6cae10),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccb73fd),
	.w1(32'h3cb73815),
	.w2(32'h3da9e1ec),
	.w3(32'hbbe26f85),
	.w4(32'hbcc0cdab),
	.w5(32'h3d33c64b),
	.w6(32'hbcd2b547),
	.w7(32'hbd0d29cd),
	.w8(32'h3cc9dc99),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0e378),
	.w1(32'h3ab14cb4),
	.w2(32'h3c1610ba),
	.w3(32'hba40d11e),
	.w4(32'hbae86cde),
	.w5(32'h3bccdc31),
	.w6(32'h3b8b9328),
	.w7(32'h3a1ef806),
	.w8(32'h3bea5fe0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13ffc7),
	.w1(32'h375851f6),
	.w2(32'hbb2eea39),
	.w3(32'hbb282944),
	.w4(32'h3b93dd7e),
	.w5(32'hbb838f8a),
	.w6(32'h3ba56494),
	.w7(32'hba2929c6),
	.w8(32'h3baba8e5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adef4bd),
	.w1(32'hbb78bc3a),
	.w2(32'hbba360f7),
	.w3(32'h3b6dc8e9),
	.w4(32'hb95b4d1e),
	.w5(32'h3a6e124c),
	.w6(32'h3b5eedc3),
	.w7(32'h3aabcb0a),
	.w8(32'h3aa358a8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2048fa),
	.w1(32'h3c202719),
	.w2(32'hbc6fa946),
	.w3(32'h3bb60a46),
	.w4(32'hbb0a9627),
	.w5(32'hbc0c36bf),
	.w6(32'h3afdca34),
	.w7(32'hbbf1d5a2),
	.w8(32'h39febee0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86569b),
	.w1(32'hbbf37e20),
	.w2(32'hbb870292),
	.w3(32'h3bb71c77),
	.w4(32'hbbfee5ee),
	.w5(32'hbb78bc3d),
	.w6(32'h3bc575c1),
	.w7(32'hbb011829),
	.w8(32'hbb8bcc7b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b507f5c),
	.w1(32'h3b960629),
	.w2(32'h3a9bf274),
	.w3(32'h3aa9eeec),
	.w4(32'h39b6e557),
	.w5(32'h3b04b655),
	.w6(32'h3af90c67),
	.w7(32'hb91a46d4),
	.w8(32'hba9457b3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d07a5),
	.w1(32'h3b129926),
	.w2(32'h3cfc548b),
	.w3(32'h3a5361b1),
	.w4(32'hbc10eccc),
	.w5(32'h3c917d7a),
	.w6(32'hbbba42fb),
	.w7(32'hbc4b5d0f),
	.w8(32'h3c393996),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0c445),
	.w1(32'h3bd59e3b),
	.w2(32'h3d0c3c68),
	.w3(32'hbb71453f),
	.w4(32'hbb1ebd46),
	.w5(32'h3ce9e97e),
	.w6(32'h3bbf7c43),
	.w7(32'h3afce708),
	.w8(32'h3c89d0f4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb816a15),
	.w1(32'hbb6c726c),
	.w2(32'h3c5b0f53),
	.w3(32'h3a570b69),
	.w4(32'h3a7d6436),
	.w5(32'h3ba7db16),
	.w6(32'h3ba889ea),
	.w7(32'h3b2b01fa),
	.w8(32'hba1b7d5e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe74eab),
	.w1(32'hbc228a5c),
	.w2(32'h3a09a489),
	.w3(32'h3c03b4b3),
	.w4(32'hbc23db8f),
	.w5(32'hbaa36f8a),
	.w6(32'hbc225ddc),
	.w7(32'hba3ada8b),
	.w8(32'h3bc1d17e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf38312),
	.w1(32'h3b6bffd1),
	.w2(32'hbb2bad5e),
	.w3(32'h3b9174b7),
	.w4(32'h3a5debdc),
	.w5(32'h3a4024fd),
	.w6(32'h3a046bc9),
	.w7(32'hbb188399),
	.w8(32'h39b0a158),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998eea8),
	.w1(32'h3b144d6e),
	.w2(32'hbc0d1a93),
	.w3(32'hbb5f6bef),
	.w4(32'hbb93d611),
	.w5(32'hbba5aac8),
	.w6(32'h3ac80663),
	.w7(32'hbbc869bf),
	.w8(32'h3a3698c8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc599b47),
	.w1(32'h3cd5f731),
	.w2(32'h3d9975c0),
	.w3(32'hbca21d3c),
	.w4(32'hbc39612c),
	.w5(32'h3d1cd5ea),
	.w6(32'hbd0c45a0),
	.w7(32'hbcd6bffa),
	.w8(32'h3c96fad8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10a491),
	.w1(32'h3b307b5e),
	.w2(32'h3d545b95),
	.w3(32'hbcff913e),
	.w4(32'hbd3b3b53),
	.w5(32'h3d054627),
	.w6(32'h3bf5ad28),
	.w7(32'hbc788693),
	.w8(32'h3cfb6135),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0fe53e),
	.w1(32'h3c53ef08),
	.w2(32'h3d1ce602),
	.w3(32'hbae21a46),
	.w4(32'hbca7e7af),
	.w5(32'h3c82d0e4),
	.w6(32'h3bdf6981),
	.w7(32'hbbc37e20),
	.w8(32'h3ce9fd6f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d63cb3c),
	.w1(32'hbd4707c5),
	.w2(32'hbcb9a967),
	.w3(32'h3c8c5b7d),
	.w4(32'hbdada716),
	.w5(32'hbd9ebeee),
	.w6(32'h3d31e7e4),
	.w7(32'hbdab4f11),
	.w8(32'hbd6a720d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c460b68),
	.w1(32'hbb6c524e),
	.w2(32'h3a8ed0bb),
	.w3(32'hbb37ea5a),
	.w4(32'hbb435012),
	.w5(32'h3b43b731),
	.w6(32'hbb485c2a),
	.w7(32'h3a94f21a),
	.w8(32'h3af73ffd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814a9b),
	.w1(32'h3adbf6fa),
	.w2(32'hbb1735b3),
	.w3(32'h3aeb5cb4),
	.w4(32'h3a37781f),
	.w5(32'hba6ce277),
	.w6(32'h38c18d7d),
	.w7(32'hbaebacb2),
	.w8(32'hbb1fd265),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba862f5c),
	.w1(32'h3b885a96),
	.w2(32'hbab2c44f),
	.w3(32'hbb1930f5),
	.w4(32'h3b18ccf7),
	.w5(32'h39df07d7),
	.w6(32'h3a937266),
	.w7(32'hb9d46e18),
	.w8(32'hbb1f0a5c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a824f0f),
	.w1(32'hbb14d846),
	.w2(32'h3c1b3ad4),
	.w3(32'hbb7b308c),
	.w4(32'hbbe51b0e),
	.w5(32'h3be96b17),
	.w6(32'hbba2727d),
	.w7(32'hbbfa55ea),
	.w8(32'h3bc9248f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba800ff2),
	.w1(32'hbb90d908),
	.w2(32'hbb0cbcd4),
	.w3(32'hbb7d6747),
	.w4(32'h3a90e3b8),
	.w5(32'h3ba6b264),
	.w6(32'hbb9998c7),
	.w7(32'hbb480cab),
	.w8(32'h3b358d54),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24fd3e),
	.w1(32'h3c4477b7),
	.w2(32'h3d713352),
	.w3(32'h3bb8435a),
	.w4(32'h3c15973c),
	.w5(32'h3c5fc68a),
	.w6(32'hbc8a3ece),
	.w7(32'hbc280256),
	.w8(32'h3c744650),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2cb6a6),
	.w1(32'hbc3a20d6),
	.w2(32'h3cf25592),
	.w3(32'h3bfe0f51),
	.w4(32'hbd0e3679),
	.w5(32'hbb9d849c),
	.w6(32'h3bbe3070),
	.w7(32'hbc85899a),
	.w8(32'h3c28179c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce9d2b0),
	.w1(32'hbb90e59e),
	.w2(32'h3d17480d),
	.w3(32'h3c20dcee),
	.w4(32'hbc8c9889),
	.w5(32'h3c0572f3),
	.w6(32'h3c34829f),
	.w7(32'hbc5d163e),
	.w8(32'hbc943642),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38bca3),
	.w1(32'h3c6f9c01),
	.w2(32'h3d29ad1a),
	.w3(32'h3bc2b909),
	.w4(32'hbb8cfb27),
	.w5(32'h3ca01417),
	.w6(32'h3b8e01e6),
	.w7(32'hbb26bc4c),
	.w8(32'h3c610867),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb392c2d),
	.w1(32'h3bae8992),
	.w2(32'h3ce43fd3),
	.w3(32'hbc82c5e8),
	.w4(32'hbcb9117b),
	.w5(32'h3c611abc),
	.w6(32'hbc074722),
	.w7(32'hbcb8792a),
	.w8(32'hbb4429aa),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fd3db),
	.w1(32'hbae15ee2),
	.w2(32'h3c31d4a0),
	.w3(32'h3aaf0eae),
	.w4(32'hb9ec492c),
	.w5(32'h3bd75269),
	.w6(32'h3c2fb04d),
	.w7(32'hbbe5a012),
	.w8(32'h3acfdb4c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a507345),
	.w1(32'h3ada541f),
	.w2(32'h3cc2c466),
	.w3(32'hbb861225),
	.w4(32'hbba4bd7f),
	.w5(32'h3cb75a1e),
	.w6(32'hbbe75c0c),
	.w7(32'hbca26c7f),
	.w8(32'h3c01922c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc8665),
	.w1(32'hbbb8fe75),
	.w2(32'h3b879172),
	.w3(32'hba40bf5b),
	.w4(32'hb95081e6),
	.w5(32'h3c24fa0f),
	.w6(32'hbb729bfb),
	.w7(32'h3af26f49),
	.w8(32'h3ba94f3b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3d09c),
	.w1(32'hbaed8f8c),
	.w2(32'hb9d5f7b4),
	.w3(32'h3bb2b0d6),
	.w4(32'hbb2e059c),
	.w5(32'hbac947f1),
	.w6(32'h3aaf17e3),
	.w7(32'h3a8b76f7),
	.w8(32'h3a2b9bad),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a977ea3),
	.w1(32'h3b0a3b01),
	.w2(32'h3a87cfa0),
	.w3(32'h3af85d16),
	.w4(32'h3b391a24),
	.w5(32'h3aeb14ba),
	.w6(32'h3aed0d31),
	.w7(32'hbb24b8b7),
	.w8(32'hbaf739f1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e72cf),
	.w1(32'hbba39847),
	.w2(32'hbc5673a7),
	.w3(32'hbaf07eff),
	.w4(32'hbaec10ad),
	.w5(32'hbc31a227),
	.w6(32'h3b971e8c),
	.w7(32'hbba9d64f),
	.w8(32'hbbfc9157),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4c7676),
	.w1(32'hbb0e50cd),
	.w2(32'hbbf80e89),
	.w3(32'h3d1982ad),
	.w4(32'hbba616f9),
	.w5(32'hbcb6a276),
	.w6(32'h3d0cb2f1),
	.w7(32'h3b99b5e4),
	.w8(32'hbc64c3b5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50234c),
	.w1(32'hbbd8994a),
	.w2(32'hbba4e419),
	.w3(32'hbb6f7305),
	.w4(32'hbc1632e7),
	.w5(32'hbbf2e734),
	.w6(32'hba88dc88),
	.w7(32'hbbcdb1fc),
	.w8(32'hbb73a9b7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd80618),
	.w1(32'h3c24f310),
	.w2(32'h3ca868f2),
	.w3(32'h3bc1dd41),
	.w4(32'hbc5ae8a6),
	.w5(32'h3c563736),
	.w6(32'h3c2815d3),
	.w7(32'hbc43ef60),
	.w8(32'h3a9673b1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced84ac),
	.w1(32'h3ca02af0),
	.w2(32'h3d467e3f),
	.w3(32'h3ce9060c),
	.w4(32'h3c01940a),
	.w5(32'h3cf676ba),
	.w6(32'h3cc42b43),
	.w7(32'h3c859708),
	.w8(32'h3cd89449),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca015aa),
	.w1(32'hbc3b0d00),
	.w2(32'hbcb1a394),
	.w3(32'h3cdb311e),
	.w4(32'hbbda8ddb),
	.w5(32'hbd02fd8f),
	.w6(32'h3d09ddd5),
	.w7(32'hbbfdd55c),
	.w8(32'hbcbf340d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad4586),
	.w1(32'h3a1b1393),
	.w2(32'h3d51f051),
	.w3(32'h3ac39323),
	.w4(32'hbce1764b),
	.w5(32'h3d08a49b),
	.w6(32'hbd1910f0),
	.w7(32'hbd3a9508),
	.w8(32'h3c895748),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60ef29),
	.w1(32'hbcf82b01),
	.w2(32'hbd0ae05f),
	.w3(32'h3c0c41da),
	.w4(32'hbd2f5f7f),
	.w5(32'hbd2a5e8f),
	.w6(32'hbac0d13d),
	.w7(32'hbd42794b),
	.w8(32'hbd39dbb6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0c89df),
	.w1(32'h3cb3f3c8),
	.w2(32'h3d364b2c),
	.w3(32'h3c85d973),
	.w4(32'h3b80126b),
	.w5(32'h3cce7aad),
	.w6(32'h3ccf1154),
	.w7(32'h3c42cef9),
	.w8(32'h3d057ecd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce9d51a),
	.w1(32'h3c8ba4f7),
	.w2(32'h3cb5e1f9),
	.w3(32'h3c21bc10),
	.w4(32'hbb0157a5),
	.w5(32'h3af338dd),
	.w6(32'h3c2112da),
	.w7(32'hbc389cd1),
	.w8(32'hbbad0802),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccbf62e),
	.w1(32'hbc523fa5),
	.w2(32'hbd0b6f31),
	.w3(32'h3c9398cd),
	.w4(32'hbcd5cb93),
	.w5(32'hbd411c48),
	.w6(32'h3d1ffcfe),
	.w7(32'hbca50ba5),
	.w8(32'hbd4ea9f7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb961001),
	.w1(32'h3b09ada2),
	.w2(32'h3b21f4f7),
	.w3(32'hbb73e584),
	.w4(32'h3a6fe4e7),
	.w5(32'h3abafced),
	.w6(32'h3aba3809),
	.w7(32'hb819caf8),
	.w8(32'hbaf03ee8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6644d),
	.w1(32'h3bbc52ea),
	.w2(32'h3d5ab93c),
	.w3(32'h3b3e52d6),
	.w4(32'hbcbec4cb),
	.w5(32'h3cb8e14f),
	.w6(32'h3c652a4d),
	.w7(32'hbc37d280),
	.w8(32'h3bff3d20),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76a5c5),
	.w1(32'h3c6463f6),
	.w2(32'h3d3dd28f),
	.w3(32'hbbe4f401),
	.w4(32'hbc9683e8),
	.w5(32'h3c84c1aa),
	.w6(32'hbcb44a6d),
	.w7(32'hbd2920d2),
	.w8(32'hb780c360),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8a6316),
	.w1(32'hbcd30672),
	.w2(32'h3d651648),
	.w3(32'h3d62d4d2),
	.w4(32'hbd8897de),
	.w5(32'h3d0cf702),
	.w6(32'h3c0fd22d),
	.w7(32'hbd33d0ed),
	.w8(32'h3d2d4f3b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd94c5f),
	.w1(32'hbc5e0191),
	.w2(32'hbde58c3e),
	.w3(32'h3dd5c6a4),
	.w4(32'hbccf588d),
	.w5(32'hbdc35bbf),
	.w6(32'h3ddf9219),
	.w7(32'hbc927b7c),
	.w8(32'hbd755032),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d210d60),
	.w1(32'hb9c0d03f),
	.w2(32'h3c148877),
	.w3(32'h3be3737b),
	.w4(32'hbca189b9),
	.w5(32'hb884d96e),
	.w6(32'h3c173f06),
	.w7(32'hbd28b128),
	.w8(32'hbcaa4d4f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4d7dc1),
	.w1(32'hbc17723f),
	.w2(32'h3d2e7696),
	.w3(32'h3d3a4651),
	.w4(32'hbd114ef7),
	.w5(32'h3c9b915d),
	.w6(32'hbca5bf5c),
	.w7(32'hbd45d3d2),
	.w8(32'h3bba1125),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb500c78),
	.w1(32'h3b14fcd8),
	.w2(32'hbb9a4fba),
	.w3(32'hbb9e6b9c),
	.w4(32'hbb44d7be),
	.w5(32'hbbbdd294),
	.w6(32'h3a1610a2),
	.w7(32'hbbb680ec),
	.w8(32'hbbcb25dd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9014be),
	.w1(32'h3c309e4a),
	.w2(32'h3d88c3b8),
	.w3(32'h3d31ca93),
	.w4(32'hbd547b1b),
	.w5(32'h3baf25dc),
	.w6(32'h3c935545),
	.w7(32'hbce88371),
	.w8(32'h3cf35527),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d164e26),
	.w1(32'hbcbfc230),
	.w2(32'h3c5a468e),
	.w3(32'h3c628234),
	.w4(32'hbc8a8c7f),
	.w5(32'h3b225604),
	.w6(32'hbbedc51b),
	.w7(32'hbcd192dd),
	.w8(32'hbc085d68),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5c6d8),
	.w1(32'hb8f00e49),
	.w2(32'h3bd9502a),
	.w3(32'h3a94da1e),
	.w4(32'hbba489bc),
	.w5(32'hbb5c7a20),
	.w6(32'hba0facb3),
	.w7(32'hbbba2717),
	.w8(32'hbb98dffb),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c263428),
	.w1(32'h3b819746),
	.w2(32'h3b8d737a),
	.w3(32'hbbb62c62),
	.w4(32'hbc0fda4d),
	.w5(32'h389a0e0a),
	.w6(32'h38a0b24d),
	.w7(32'h3b5805de),
	.w8(32'h3b2e10ee),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c911391),
	.w1(32'h3b9c1a4e),
	.w2(32'h3cde36b6),
	.w3(32'h3c069632),
	.w4(32'hbbdcf600),
	.w5(32'h3c91ad17),
	.w6(32'h3c171fe3),
	.w7(32'hbb8a5ae2),
	.w8(32'h3c406b40),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be56030),
	.w1(32'hbc16a733),
	.w2(32'h3c1d464e),
	.w3(32'hba49f26e),
	.w4(32'hbc8a79a2),
	.w5(32'hbbdd4e65),
	.w6(32'h3c1539ac),
	.w7(32'hbc94d274),
	.w8(32'hbca86bc9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c526a44),
	.w1(32'h3aaa1b38),
	.w2(32'hbc927186),
	.w3(32'h3c8b7abf),
	.w4(32'h3c28125c),
	.w5(32'hbcaaeccd),
	.w6(32'h3d0e9cea),
	.w7(32'h3c2b55bf),
	.w8(32'hbc83c7d1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b851d),
	.w1(32'hbc20b535),
	.w2(32'h3c6e7971),
	.w3(32'h3c03084d),
	.w4(32'hbc387f68),
	.w5(32'h3c604011),
	.w6(32'h3c87a4ec),
	.w7(32'h3c3e1efc),
	.w8(32'hbb3b6cb9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24f639),
	.w1(32'hbc6077fd),
	.w2(32'hbc06e7f8),
	.w3(32'h3c67f103),
	.w4(32'hbcd19ffa),
	.w5(32'hbba57eee),
	.w6(32'h3b7e3f11),
	.w7(32'hbc703c02),
	.w8(32'h3b8cb2eb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8d4d9),
	.w1(32'h3c98976a),
	.w2(32'h3d3abd6a),
	.w3(32'h3a5dd2c4),
	.w4(32'hbba5114c),
	.w5(32'h3cdc6c70),
	.w6(32'hbc354b42),
	.w7(32'hbc09448d),
	.w8(32'h3cba403e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d1879),
	.w1(32'hbba0fa36),
	.w2(32'h3c565a5c),
	.w3(32'h3b558b7d),
	.w4(32'hbbfa4d78),
	.w5(32'h3b916e80),
	.w6(32'h3c80e435),
	.w7(32'hbc0364e1),
	.w8(32'hbace4807),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b1902),
	.w1(32'h3a1c51dc),
	.w2(32'hbac8ce3a),
	.w3(32'h3a9e2de5),
	.w4(32'hbb454683),
	.w5(32'hbb485cc8),
	.w6(32'h3a53a24e),
	.w7(32'hb89419c9),
	.w8(32'hbb5ac494),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f87d29),
	.w1(32'h3b50ada3),
	.w2(32'h3ad7b57f),
	.w3(32'hbb79203b),
	.w4(32'h39fcab2b),
	.w5(32'h3a4f8710),
	.w6(32'h398a53cb),
	.w7(32'hb8844f45),
	.w8(32'h3b38efcd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb050f44),
	.w1(32'h397eee75),
	.w2(32'hbb51c98b),
	.w3(32'hbad324f0),
	.w4(32'hbb155975),
	.w5(32'hbb200f4f),
	.w6(32'hbad74b69),
	.w7(32'hbb4c0ff0),
	.w8(32'hbb13e89c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa43ddc),
	.w1(32'h3c08a819),
	.w2(32'h3b8356bc),
	.w3(32'hba95078f),
	.w4(32'h3a4cc8a8),
	.w5(32'h3b95cd78),
	.w6(32'h3b6f6949),
	.w7(32'hbbcf5b31),
	.w8(32'hbbbcaaf3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1680e),
	.w1(32'hb98ffa20),
	.w2(32'h3b9bfa93),
	.w3(32'h3c21fc3c),
	.w4(32'hbc99d6af),
	.w5(32'hbbd8948d),
	.w6(32'h3be181ff),
	.w7(32'hbcd35b79),
	.w8(32'hbc885435),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be793a8),
	.w1(32'h3c0cff4f),
	.w2(32'h3ac51a0e),
	.w3(32'hbbb35dad),
	.w4(32'h3ad7e58a),
	.w5(32'hba940bde),
	.w6(32'h3b425cf2),
	.w7(32'hbaa7d591),
	.w8(32'hbb8595e9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d852c),
	.w1(32'hbc43fe85),
	.w2(32'h3c67f9b5),
	.w3(32'hbad6bf12),
	.w4(32'hbc816800),
	.w5(32'h3bd1eb41),
	.w6(32'hbc300704),
	.w7(32'hbc333af4),
	.w8(32'h3baf9596),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1eef96),
	.w1(32'h3b785989),
	.w2(32'hbcb1c2bf),
	.w3(32'h3cee3c2f),
	.w4(32'h393ccea2),
	.w5(32'hbceb411a),
	.w6(32'h3d188fdd),
	.w7(32'h3bd8dd47),
	.w8(32'hbccdd491),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80f356),
	.w1(32'h3c226813),
	.w2(32'h3c81c1cb),
	.w3(32'hbb82b3a1),
	.w4(32'h3b84ee41),
	.w5(32'h3a2cacc7),
	.w6(32'h3b9a0ee6),
	.w7(32'hbbc8c2cc),
	.w8(32'hbb851790),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab9f9e),
	.w1(32'hbaedb3d4),
	.w2(32'hbc420c34),
	.w3(32'h3c19f119),
	.w4(32'hbbfb41f9),
	.w5(32'hbbfa42e5),
	.w6(32'h3a8afc78),
	.w7(32'hbacb860a),
	.w8(32'h3c02f71e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15894a),
	.w1(32'hbb19f2b5),
	.w2(32'hbac5406e),
	.w3(32'h3c0b1e6d),
	.w4(32'hbb2293f2),
	.w5(32'h3a563710),
	.w6(32'hba631301),
	.w7(32'h3a89651e),
	.w8(32'hb9f19853),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0739bd),
	.w1(32'h3b1aef46),
	.w2(32'h3ab2bf97),
	.w3(32'h3be990f9),
	.w4(32'h3b36d2a9),
	.w5(32'h3a7b5f1c),
	.w6(32'h3c1cc0a0),
	.w7(32'h3b7bea1a),
	.w8(32'h3b3a7e62),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbf7a3),
	.w1(32'h3b2fedc7),
	.w2(32'h3d2f6d05),
	.w3(32'hbd1a1afc),
	.w4(32'hbcce1af6),
	.w5(32'h3d34ffd1),
	.w6(32'hbcbb51ae),
	.w7(32'h3a742126),
	.w8(32'h3cdc6ccb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c250e27),
	.w1(32'h3c032082),
	.w2(32'h3d652da7),
	.w3(32'hbc33a7af),
	.w4(32'hbcb64cf4),
	.w5(32'h3d026fa2),
	.w6(32'hbc108acd),
	.w7(32'hbca10b18),
	.w8(32'h3c870807),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb65cc),
	.w1(32'h3afac606),
	.w2(32'h3bcec5a4),
	.w3(32'hbada37f0),
	.w4(32'hba7fd3f8),
	.w5(32'h3b2e20d2),
	.w6(32'hbbafbb00),
	.w7(32'hbb38aa96),
	.w8(32'h3a7c58e4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ae5e9),
	.w1(32'h3b266148),
	.w2(32'h3c33a28e),
	.w3(32'h3b89683d),
	.w4(32'hbb6fbecb),
	.w5(32'h3b81e822),
	.w6(32'h3b7ca3c3),
	.w7(32'h3c00950b),
	.w8(32'h3c582bc8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c600fbe),
	.w1(32'hb8138aae),
	.w2(32'h3b933fc3),
	.w3(32'h3c39efce),
	.w4(32'hbb4f7412),
	.w5(32'hbabf954f),
	.w6(32'h3c10e80d),
	.w7(32'hbc04d90b),
	.w8(32'hbb9ca112),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83f90c),
	.w1(32'h3b8a49e3),
	.w2(32'h3c934a04),
	.w3(32'h39019915),
	.w4(32'hbb98f717),
	.w5(32'h3be50f0a),
	.w6(32'h3b7f0729),
	.w7(32'hba8824b6),
	.w8(32'h3bcd54ac),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92e689),
	.w1(32'h3c7dd4a5),
	.w2(32'h3cc7a4b3),
	.w3(32'h3aa5dec3),
	.w4(32'h3b33ace2),
	.w5(32'h3c54747c),
	.w6(32'hba536a88),
	.w7(32'hbb06f344),
	.w8(32'h3bb52c0e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c275225),
	.w1(32'h3c3c4095),
	.w2(32'h3d8a8b4e),
	.w3(32'hbc2a89ba),
	.w4(32'hbccca7b4),
	.w5(32'h3d2402ac),
	.w6(32'hbc421198),
	.w7(32'hbcc4bb5b),
	.w8(32'h3c8dfdbe),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf5088),
	.w1(32'hbbcefa57),
	.w2(32'hbc1a8b10),
	.w3(32'h3ca6be58),
	.w4(32'hbc129fc7),
	.w5(32'hbc810f06),
	.w6(32'h3ccc99fd),
	.w7(32'hbc4cf92c),
	.w8(32'hbc84cf4e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdfe7c5),
	.w1(32'h3c8b384b),
	.w2(32'h3ccfee65),
	.w3(32'h3a390074),
	.w4(32'hbc05cc8d),
	.w5(32'h3bcc81dd),
	.w6(32'hba738af1),
	.w7(32'hbc3ea4ae),
	.w8(32'h3c14bac9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b70fd),
	.w1(32'h3c7685e7),
	.w2(32'h3d4f0068),
	.w3(32'h3ab9ec40),
	.w4(32'hbc499a8f),
	.w5(32'h3d11d724),
	.w6(32'hbc6385ee),
	.w7(32'hbc804112),
	.w8(32'h3cb95bba),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf93f00),
	.w1(32'hbb607e8c),
	.w2(32'hbba648c8),
	.w3(32'h3c10ed25),
	.w4(32'hbc720939),
	.w5(32'hbc253dd5),
	.w6(32'h3c814ee4),
	.w7(32'hbc4bbc9d),
	.w8(32'hbc449f7f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7dad51),
	.w1(32'h3ae9ad5c),
	.w2(32'h3cbeb127),
	.w3(32'h3c1f2ff9),
	.w4(32'hbc428b64),
	.w5(32'h3c3c6f7f),
	.w6(32'h3aea5273),
	.w7(32'hbc5d432d),
	.w8(32'h3c1310c5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce2cf),
	.w1(32'hb84d83d5),
	.w2(32'h3bcb0ca4),
	.w3(32'h38d099d3),
	.w4(32'hbba7248e),
	.w5(32'h38228b6b),
	.w6(32'h3a8c016e),
	.w7(32'hbbeb8eb9),
	.w8(32'hbb387f93),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca02dd6),
	.w1(32'hbd16aa97),
	.w2(32'hbd63f980),
	.w3(32'h3cd5e309),
	.w4(32'hbcbea55d),
	.w5(32'hbd50a8ef),
	.w6(32'h3d4530ac),
	.w7(32'hbc387d08),
	.w8(32'hbd398eac),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca41cf6),
	.w1(32'h3b04643b),
	.w2(32'hbbb35adc),
	.w3(32'h3c66563d),
	.w4(32'hbb3875f1),
	.w5(32'hbc470761),
	.w6(32'h3c9e78f6),
	.w7(32'hba054d28),
	.w8(32'hbc245d6c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9838d),
	.w1(32'hb8f3f716),
	.w2(32'h390f4264),
	.w3(32'hb995d0bd),
	.w4(32'hb90aec34),
	.w5(32'h36996b85),
	.w6(32'hb75e2e18),
	.w7(32'hba01a0ff),
	.w8(32'hba447a09),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d081d),
	.w1(32'h3bbc82de),
	.w2(32'h3ba328dc),
	.w3(32'hba39298b),
	.w4(32'h3a9f90dd),
	.w5(32'hba341624),
	.w6(32'h3b77930c),
	.w7(32'h3b4f1a01),
	.w8(32'hbb07bef9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c583b),
	.w1(32'hbae8a827),
	.w2(32'h3b407acd),
	.w3(32'h3b1e8664),
	.w4(32'hbb94d783),
	.w5(32'hbc170012),
	.w6(32'h3b1d3940),
	.w7(32'hbbfc391f),
	.w8(32'hbc265785),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1b480c),
	.w1(32'hbae03ec8),
	.w2(32'hbc3f7823),
	.w3(32'h3cd443f0),
	.w4(32'hbc6a64b7),
	.w5(32'hbcbbf319),
	.w6(32'h3ce1f45a),
	.w7(32'hbcad1f27),
	.w8(32'hbcf42d29),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb35dce),
	.w1(32'h3bb76c24),
	.w2(32'h3d301dbd),
	.w3(32'h3bfeae8e),
	.w4(32'hbc79978c),
	.w5(32'h3c8906e1),
	.w6(32'hbb5c2f0e),
	.w7(32'hbcc4a659),
	.w8(32'hb93c95e5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afc60f),
	.w1(32'hba82d2c6),
	.w2(32'h3a63e594),
	.w3(32'hb9b20aaf),
	.w4(32'hbacae65d),
	.w5(32'hba632059),
	.w6(32'h39b82f9d),
	.w7(32'h3a75a304),
	.w8(32'h3a0fdb21),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63838f),
	.w1(32'h3c16f7c3),
	.w2(32'h3d38d301),
	.w3(32'h3be51796),
	.w4(32'hbc20598a),
	.w5(32'h3cce1102),
	.w6(32'hb98c79be),
	.w7(32'hbcb781de),
	.w8(32'h3c0b50b5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca94ff5),
	.w1(32'h3c0926f8),
	.w2(32'h3c84d665),
	.w3(32'h3c262dde),
	.w4(32'hbb13398f),
	.w5(32'h3b768e6f),
	.w6(32'h3c828636),
	.w7(32'hbc267363),
	.w8(32'hbb413fb9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d00be),
	.w1(32'h3ac4e15f),
	.w2(32'h3d24cd86),
	.w3(32'h3bca9344),
	.w4(32'hbc495b17),
	.w5(32'h3cc8be15),
	.w6(32'hbc833b80),
	.w7(32'hbd0b3389),
	.w8(32'h3c22d439),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdfecd),
	.w1(32'hbd01e332),
	.w2(32'h3c2d5a60),
	.w3(32'hbc4aafa3),
	.w4(32'hbd2b6585),
	.w5(32'hbc9e5638),
	.w6(32'h3c2735bf),
	.w7(32'hbd2e1e6f),
	.w8(32'hbd1af292),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2c638),
	.w1(32'h3c527a3a),
	.w2(32'h3b850049),
	.w3(32'h3c86d1d5),
	.w4(32'h3c43dbed),
	.w5(32'h3b877708),
	.w6(32'h3ca9a864),
	.w7(32'h3c6e72ac),
	.w8(32'h3c2f7d5d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b833a),
	.w1(32'hbb73256f),
	.w2(32'hbb86d81f),
	.w3(32'hbbea5bf5),
	.w4(32'hbb736413),
	.w5(32'hbb81768e),
	.w6(32'hbb0f66a2),
	.w7(32'hbb8b2b8e),
	.w8(32'hbb676392),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca428c6),
	.w1(32'hbc43a79d),
	.w2(32'hbc857778),
	.w3(32'h3c469d8b),
	.w4(32'hbc797edb),
	.w5(32'hbc93e436),
	.w6(32'h3cc35f12),
	.w7(32'hbc4e36fd),
	.w8(32'hbc79d91f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4aa61b),
	.w1(32'h3c81fd98),
	.w2(32'hbc1ce028),
	.w3(32'h3d052e47),
	.w4(32'h3c041c70),
	.w5(32'hbc4f566b),
	.w6(32'h3d3debe6),
	.w7(32'hbaf0f647),
	.w8(32'hba9bd576),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bb515),
	.w1(32'hbc5ae12f),
	.w2(32'hbc221aec),
	.w3(32'h3c046103),
	.w4(32'hbc8b4949),
	.w5(32'hbc98b548),
	.w6(32'h3c6f3545),
	.w7(32'hbc295f34),
	.w8(32'hbc8629c5),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c027805),
	.w1(32'h3b276d82),
	.w2(32'h3c485a1b),
	.w3(32'h3b304bf4),
	.w4(32'h3b371e38),
	.w5(32'h3c070311),
	.w6(32'hbb6d8df1),
	.w7(32'hbb6287a1),
	.w8(32'h3bca612a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b569c60),
	.w1(32'h3b7124e1),
	.w2(32'h3b9604cb),
	.w3(32'h3b2223c3),
	.w4(32'h3b8fd9aa),
	.w5(32'h3b93babf),
	.w6(32'h3adfc372),
	.w7(32'h3b8afb9c),
	.w8(32'h3b7ad661),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0d507),
	.w1(32'h3c205aa6),
	.w2(32'h3ccad0db),
	.w3(32'h3b660cd9),
	.w4(32'hbc23e539),
	.w5(32'h3c7248c4),
	.w6(32'h3be393ee),
	.w7(32'hbbba7aec),
	.w8(32'h3c10ec46),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb198271),
	.w1(32'hbbb9e32c),
	.w2(32'h39e79861),
	.w3(32'h3b54b9ef),
	.w4(32'hbb6867eb),
	.w5(32'hba3a1794),
	.w6(32'hbc24c2db),
	.w7(32'hbc3baca8),
	.w8(32'hbc0c59ca),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc52ac2),
	.w1(32'hbc1f1f74),
	.w2(32'h3a44eae7),
	.w3(32'hbc1b0f80),
	.w4(32'hbca19d33),
	.w5(32'hbbc25a97),
	.w6(32'h3c2df28d),
	.w7(32'hbc100be4),
	.w8(32'hbc198c6a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b43b62),
	.w1(32'h39be0e00),
	.w2(32'h3b153642),
	.w3(32'hb7c95e33),
	.w4(32'hb958052a),
	.w5(32'h3aa03657),
	.w6(32'h3a2f6e8a),
	.w7(32'h3a4b943c),
	.w8(32'h3a9cda9a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0a27f),
	.w1(32'hbc058e65),
	.w2(32'h3cb1597b),
	.w3(32'hbc812600),
	.w4(32'hbcb5adbb),
	.w5(32'h3be82c72),
	.w6(32'hb8888a4b),
	.w7(32'hbbf157c7),
	.w8(32'h3be8c883),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a350e94),
	.w1(32'h3a1d01d8),
	.w2(32'h3a869304),
	.w3(32'h3a4321e7),
	.w4(32'h39bf3c3d),
	.w5(32'h3a378035),
	.w6(32'hb7891460),
	.w7(32'h3a5283bd),
	.w8(32'h390fc6be),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace1f33),
	.w1(32'h3b0407eb),
	.w2(32'h3af03020),
	.w3(32'hb9d8acf2),
	.w4(32'h3aa23ec8),
	.w5(32'h3acac3fa),
	.w6(32'h3a7f70f2),
	.w7(32'h3aa1b688),
	.w8(32'h3b114053),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cea17e4),
	.w1(32'h3a9a7b1e),
	.w2(32'hbc1ce2f4),
	.w3(32'h3cc674da),
	.w4(32'hb9d4c6ea),
	.w5(32'hbc0ef93d),
	.w6(32'h3d01b4bf),
	.w7(32'hb886cf0a),
	.w8(32'hbc0f842e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d26af5c),
	.w1(32'hbb997a91),
	.w2(32'h3d268329),
	.w3(32'h3c9617ee),
	.w4(32'hbc9bdc0d),
	.w5(32'h3d25306c),
	.w6(32'h3c9389cd),
	.w7(32'hbc974b2d),
	.w8(32'h3c8c7f7e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c950774),
	.w1(32'hbb81f68d),
	.w2(32'hb8b1a4b0),
	.w3(32'h3bdf973f),
	.w4(32'hbbc765fc),
	.w5(32'hbb1bda07),
	.w6(32'h3c3637c7),
	.w7(32'hbb3c3473),
	.w8(32'h3ade7087),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb93adb),
	.w1(32'hbb655457),
	.w2(32'h3c24a78e),
	.w3(32'h3c3c49be),
	.w4(32'hbbcbfcac),
	.w5(32'h39f6978f),
	.w6(32'h3c355e48),
	.w7(32'hbc732108),
	.w8(32'hbbf0ff19),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61dee7),
	.w1(32'hba43e7c2),
	.w2(32'h3c38bf3a),
	.w3(32'hba13ce9d),
	.w4(32'hbba7caab),
	.w5(32'h3857dde1),
	.w6(32'h3acc3814),
	.w7(32'hbc1ed827),
	.w8(32'hba8cf02a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfa6bc1),
	.w1(32'h3bbbf767),
	.w2(32'h3d88898c),
	.w3(32'h3b3a629b),
	.w4(32'hbccefc19),
	.w5(32'h3d0ace8b),
	.w6(32'h3acfe6bb),
	.w7(32'hbc8a185b),
	.w8(32'h3cdb51ae),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccf650f),
	.w1(32'h3c071eec),
	.w2(32'h3cdb2397),
	.w3(32'h3c2f87e7),
	.w4(32'hbc339642),
	.w5(32'h3b9a614a),
	.w6(32'h399284b4),
	.w7(32'hbcb4eca2),
	.w8(32'h3a1adb92),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1639a7),
	.w1(32'h3b846a94),
	.w2(32'h3d512b60),
	.w3(32'hbc1b1583),
	.w4(32'hbc8aebf3),
	.w5(32'h3cffcea0),
	.w6(32'hbc31d8d6),
	.w7(32'hbcbeabbe),
	.w8(32'h3c5a1398),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc1866),
	.w1(32'h3bc1f083),
	.w2(32'hbae45e96),
	.w3(32'hba9c5fcc),
	.w4(32'h3bc5560a),
	.w5(32'hbb6761c4),
	.w6(32'h3bfeaf26),
	.w7(32'h3a5d91f3),
	.w8(32'hba702d4a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e55e),
	.w1(32'h3c0b9e9a),
	.w2(32'h3cbc8720),
	.w3(32'h3a60d93c),
	.w4(32'hbacefbfd),
	.w5(32'h3c93d3b0),
	.w6(32'hbb455336),
	.w7(32'hbbd13847),
	.w8(32'h3ba1322d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8ee30),
	.w1(32'h3a63eba8),
	.w2(32'h39bd931e),
	.w3(32'hbade8bb3),
	.w4(32'h3a756519),
	.w5(32'h392103b2),
	.w6(32'h3a05ecca),
	.w7(32'h399026d3),
	.w8(32'h3a06733f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb13a00),
	.w1(32'hbb2101dc),
	.w2(32'h3c40610e),
	.w3(32'hbbf1757f),
	.w4(32'hbbf9ce92),
	.w5(32'h3a64f18a),
	.w6(32'hbbb52818),
	.w7(32'hbbb80b8d),
	.w8(32'h3b68d08b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee95b1),
	.w1(32'hbc04fcf6),
	.w2(32'hbc091b9a),
	.w3(32'h3a25140a),
	.w4(32'hbbb8b11e),
	.w5(32'hbc015b0b),
	.w6(32'h3abfb2d4),
	.w7(32'hbb97dba4),
	.w8(32'hbbac9065),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c433135),
	.w1(32'h3c218062),
	.w2(32'h3ceace4e),
	.w3(32'hbb97f1e9),
	.w4(32'hbbf8387a),
	.w5(32'h3c411ae9),
	.w6(32'h3b80558a),
	.w7(32'hbb813534),
	.w8(32'h3c09bff9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f407f),
	.w1(32'h3aebeda2),
	.w2(32'h3a07a1cb),
	.w3(32'h399adaaf),
	.w4(32'h3b0b0c40),
	.w5(32'h3a980e35),
	.w6(32'h3abe0f50),
	.w7(32'h3a4ea55d),
	.w8(32'h39475b42),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba471e5b),
	.w1(32'h3b137596),
	.w2(32'h3af70e7e),
	.w3(32'h39ca066e),
	.w4(32'h3a29f822),
	.w5(32'hb9ceb639),
	.w6(32'h3a7a3b7f),
	.w7(32'hb7f805f4),
	.w8(32'hbb2403f3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38a4a0),
	.w1(32'h3bb0d119),
	.w2(32'h3bee3e03),
	.w3(32'hbbd73da7),
	.w4(32'hbbbf9aab),
	.w5(32'hbb5e3431),
	.w6(32'h3c262d55),
	.w7(32'h3b1f73d8),
	.w8(32'hbb0422b6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2daf2a),
	.w1(32'h3c96edad),
	.w2(32'h3d1ab1eb),
	.w3(32'h3c8f24f3),
	.w4(32'hbac3951d),
	.w5(32'h3cc494e2),
	.w6(32'h3baeea6c),
	.w7(32'h3b4e92f3),
	.w8(32'h3c8cefb8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ffdab),
	.w1(32'hbc8cf293),
	.w2(32'h3c5e716f),
	.w3(32'h3d1d5ed8),
	.w4(32'hbccb9c0d),
	.w5(32'hba89ae66),
	.w6(32'h3c8a4045),
	.w7(32'hbc9acf55),
	.w8(32'h3a9ccd71),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ee37e),
	.w1(32'h3b227526),
	.w2(32'h3b99807f),
	.w3(32'h3b4d2f81),
	.w4(32'h3a801699),
	.w5(32'h3b8fbb20),
	.w6(32'h3b75acb4),
	.w7(32'h39d32ecb),
	.w8(32'h3b71043a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c987a2a),
	.w1(32'hbbfce200),
	.w2(32'h3daa8ef8),
	.w3(32'hbcf0a229),
	.w4(32'hbd626fa1),
	.w5(32'h3d14e41f),
	.w6(32'hbd1f5589),
	.w7(32'hbd622b1b),
	.w8(32'h3cb2f3e1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6d0e66),
	.w1(32'h3bd7da15),
	.w2(32'h3bced3a2),
	.w3(32'h3d121092),
	.w4(32'h3b5e538b),
	.w5(32'hbc20ebba),
	.w6(32'h3d6864ba),
	.w7(32'hbcd707cc),
	.w8(32'hbcfed1ce),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3261a),
	.w1(32'hbb93bc71),
	.w2(32'h3c125ef6),
	.w3(32'hbb67ee8e),
	.w4(32'hbbf1f97a),
	.w5(32'h3b8f8b96),
	.w6(32'hbc46abcb),
	.w7(32'hbc6c17c0),
	.w8(32'h3b8a1dd3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b1527),
	.w1(32'h3b47a4ae),
	.w2(32'hbaac6359),
	.w3(32'hba18711d),
	.w4(32'h3b3a9356),
	.w5(32'hba40909b),
	.w6(32'h3b42f6db),
	.w7(32'hba911f8c),
	.w8(32'h393afd22),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba083a82),
	.w1(32'h3a874f44),
	.w2(32'h3a5518fe),
	.w3(32'hb968a333),
	.w4(32'hba450a9b),
	.w5(32'hba9fc8cd),
	.w6(32'hb9e31ebe),
	.w7(32'hba2aa604),
	.w8(32'hb9d83391),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6829820),
	.w1(32'h3a3597d8),
	.w2(32'hba9c1f70),
	.w3(32'hbac37202),
	.w4(32'h3a3913cf),
	.w5(32'hba4e091b),
	.w6(32'h39a2aa06),
	.w7(32'hba4c3a67),
	.w8(32'hb9c3ca9d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1c4eb),
	.w1(32'hbc222853),
	.w2(32'h3c65172c),
	.w3(32'h397362c5),
	.w4(32'hbc719c4f),
	.w5(32'h3c0d1622),
	.w6(32'hbacd3be1),
	.w7(32'hbbd261ad),
	.w8(32'h3c2fce49),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cee732d),
	.w1(32'h3c5b7b94),
	.w2(32'h3ce040fd),
	.w3(32'h3c179a3e),
	.w4(32'hbbc37d26),
	.w5(32'h3c811651),
	.w6(32'h3c4096a4),
	.w7(32'h3b3bd247),
	.w8(32'h3c7b6308),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2edffe),
	.w1(32'h3bff7e8c),
	.w2(32'h3d0b10ab),
	.w3(32'h3cdc671f),
	.w4(32'hbc921c89),
	.w5(32'hbac170d7),
	.w6(32'h3cbe5732),
	.w7(32'hbc912280),
	.w8(32'hbc3ec02c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f6cb2),
	.w1(32'hbb81e089),
	.w2(32'hba86ac9d),
	.w3(32'h3884d16b),
	.w4(32'hbbf47a84),
	.w5(32'hbbb74591),
	.w6(32'h3bd681c1),
	.w7(32'h3a8f2a3c),
	.w8(32'hb9ae8abf),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae671b),
	.w1(32'h3b919c51),
	.w2(32'h3d339a4e),
	.w3(32'hbb884286),
	.w4(32'hbcc79c64),
	.w5(32'h3c967caa),
	.w6(32'hbb8ea6f0),
	.w7(32'hbcc62168),
	.w8(32'h3c4415d8),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6465e1),
	.w1(32'hbaafb53f),
	.w2(32'h3c5e49f1),
	.w3(32'h3bde5e49),
	.w4(32'hbba698e4),
	.w5(32'h3b901740),
	.w6(32'hbb171c27),
	.w7(32'hbbf9ea08),
	.w8(32'h3bd210f5),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc7cab),
	.w1(32'h3a8a29b3),
	.w2(32'h3a24dbf0),
	.w3(32'h393ce01a),
	.w4(32'h3a91fe49),
	.w5(32'h39f4bda3),
	.w6(32'h3a1b70f9),
	.w7(32'h3a2c7ffd),
	.w8(32'hb90ca1e8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d6ee4),
	.w1(32'h3bc40398),
	.w2(32'h3c0ebce1),
	.w3(32'h3be9d836),
	.w4(32'h3b0ad5d4),
	.w5(32'h3b52478a),
	.w6(32'h3b9be309),
	.w7(32'h3b926b34),
	.w8(32'h3bfcd4f9),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99c40c),
	.w1(32'hba1ade52),
	.w2(32'h39bbc8b2),
	.w3(32'hbaaf47ce),
	.w4(32'hba3057b2),
	.w5(32'hb9df5e9d),
	.w6(32'hba23c51c),
	.w7(32'h3aaed42b),
	.w8(32'hb8a99a02),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4720c),
	.w1(32'hbade830f),
	.w2(32'h3bd70643),
	.w3(32'h3c106703),
	.w4(32'hbcab1ae4),
	.w5(32'hbc9a2fd7),
	.w6(32'h3bfaeb02),
	.w7(32'hbcb6db0b),
	.w8(32'hbc68babf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d291fca),
	.w1(32'h3a0fac14),
	.w2(32'hbc0af2a3),
	.w3(32'h3cbce81f),
	.w4(32'hbc2d3e13),
	.w5(32'hbcb53834),
	.w6(32'h3d27516e),
	.w7(32'hbb89f43b),
	.w8(32'hbbc03251),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d086427),
	.w1(32'h3b46fc5f),
	.w2(32'h3c022206),
	.w3(32'h3c8ec342),
	.w4(32'hbc082e3a),
	.w5(32'hbb4dedc0),
	.w6(32'h3cb715b5),
	.w7(32'hbc474cf9),
	.w8(32'hbaad22e8),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a7505),
	.w1(32'h3ba662ae),
	.w2(32'hbb48bff3),
	.w3(32'h3c347555),
	.w4(32'h3bc9c5ae),
	.w5(32'hba270e3a),
	.w6(32'h3c8451ff),
	.w7(32'h3bf6f3c3),
	.w8(32'h3ba8e0be),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2e85ba),
	.w1(32'h3c16095e),
	.w2(32'h3bf7c590),
	.w3(32'h3cbbf883),
	.w4(32'hbbb1ac8a),
	.w5(32'hbc8056b3),
	.w6(32'h3d2ab6a0),
	.w7(32'hbbcd9134),
	.w8(32'hbc437ba9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf372),
	.w1(32'h3af74981),
	.w2(32'h3cbbb97d),
	.w3(32'hbbac64e6),
	.w4(32'hbc214bf9),
	.w5(32'h3bf814ab),
	.w6(32'h3ae3ec2f),
	.w7(32'hbc2af2ce),
	.w8(32'h3b0b22bb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb93566),
	.w1(32'h397b7688),
	.w2(32'h3d459797),
	.w3(32'h3b159629),
	.w4(32'hbce02277),
	.w5(32'h3c5cdb83),
	.w6(32'hbc13e0b0),
	.w7(32'hbd006d1f),
	.w8(32'h3b2ae790),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15abd4),
	.w1(32'h3a0ef0f0),
	.w2(32'h3ab4710b),
	.w3(32'h3b956059),
	.w4(32'h3a5cf84b),
	.w5(32'h3ae3109c),
	.w6(32'hb9b8f37d),
	.w7(32'h3a6fc519),
	.w8(32'hb9ae9242),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba161800),
	.w1(32'h3b83a747),
	.w2(32'h3b88ec5a),
	.w3(32'h38dd813f),
	.w4(32'h3b0a8230),
	.w5(32'h3afb9daf),
	.w6(32'h3b8ea3c5),
	.w7(32'h3b54e46b),
	.w8(32'h3af335c5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08b895),
	.w1(32'hbb2f9b04),
	.w2(32'h3d0209e8),
	.w3(32'hbc29b1c7),
	.w4(32'hbd1dc417),
	.w5(32'h3bd72370),
	.w6(32'h3ba73460),
	.w7(32'hbc669456),
	.w8(32'h3c868e78),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4d083),
	.w1(32'hba5fda27),
	.w2(32'h3d0cf921),
	.w3(32'hba5e961a),
	.w4(32'hbcab84d4),
	.w5(32'h3cfc9c5c),
	.w6(32'h3b87786c),
	.w7(32'hbcc77d9f),
	.w8(32'h3c159835),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d2198),
	.w1(32'h3c444a9f),
	.w2(32'h3cd3c37d),
	.w3(32'h3c52761b),
	.w4(32'hbc8943b5),
	.w5(32'h3ae0ed9d),
	.w6(32'h3c879ffd),
	.w7(32'hbc743c80),
	.w8(32'hbc03db6d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aac02),
	.w1(32'h3c52c8d9),
	.w2(32'h3cf250ea),
	.w3(32'hbba40e9a),
	.w4(32'hbc6d9baa),
	.w5(32'h3cba1a9e),
	.w6(32'hbcce1abd),
	.w7(32'hbd003eb4),
	.w8(32'h3c27648f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75aaf6),
	.w1(32'h38ea0d7f),
	.w2(32'h39817fdb),
	.w3(32'hbb252203),
	.w4(32'hba8872be),
	.w5(32'hb896a15f),
	.w6(32'hba268e68),
	.w7(32'h3b6a25da),
	.w8(32'hb89a254f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabd2aa),
	.w1(32'h3b3f60e5),
	.w2(32'h3bc14018),
	.w3(32'hbb0ce5c6),
	.w4(32'hb8b5dcd3),
	.w5(32'h3b63c27b),
	.w6(32'hba084962),
	.w7(32'h395e42f6),
	.w8(32'h3b3f8958),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a1d63),
	.w1(32'hbd7aded7),
	.w2(32'h3d00ceca),
	.w3(32'h3cf5c8e2),
	.w4(32'hbd44e4a5),
	.w5(32'h3cf6f534),
	.w6(32'hbba4f7cf),
	.w7(32'hbd5a1b1e),
	.w8(32'h3c942450),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95ca47),
	.w1(32'h3bcd486b),
	.w2(32'h3d80c1ac),
	.w3(32'hbc4af716),
	.w4(32'hbd06c089),
	.w5(32'h3cf5e04b),
	.w6(32'hbca4d83d),
	.w7(32'hbcbe8a16),
	.w8(32'h3cea5ab4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4f6a1),
	.w1(32'hbc1267bb),
	.w2(32'h3c7f575e),
	.w3(32'h3c9fc203),
	.w4(32'hbc4c221c),
	.w5(32'h3c028f2a),
	.w6(32'hbc95c68b),
	.w7(32'hbcbae033),
	.w8(32'h3bb81600),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b8fe5),
	.w1(32'hbc4a4f7a),
	.w2(32'hbca76617),
	.w3(32'h3c8aba0d),
	.w4(32'hbc2c0258),
	.w5(32'hbcbd61ce),
	.w6(32'h3cebda4d),
	.w7(32'hbbeb2c9e),
	.w8(32'hbca15d2e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd4ae2d),
	.w1(32'h3c68824e),
	.w2(32'h3c95fff8),
	.w3(32'h3c9b103c),
	.w4(32'h3b7d29ee),
	.w5(32'hbbaf00f9),
	.w6(32'h3cf6718b),
	.w7(32'h3a9e3c12),
	.w8(32'hbc362aa1),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb93aa),
	.w1(32'hba10b8de),
	.w2(32'hba4622a3),
	.w3(32'h3add26fb),
	.w4(32'h3931ad30),
	.w5(32'h38657734),
	.w6(32'hb9abe865),
	.w7(32'hb9a35d90),
	.w8(32'hb8cb0175),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7358b8),
	.w1(32'h37e1c60d),
	.w2(32'hba69adc7),
	.w3(32'hba0e7afd),
	.w4(32'h3a0f663a),
	.w5(32'hba7a85bb),
	.w6(32'h38d5daa2),
	.w7(32'h399d69f9),
	.w8(32'hb918c911),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69f66),
	.w1(32'h3b934c03),
	.w2(32'h3be4ca86),
	.w3(32'hbc60f49d),
	.w4(32'hbb5a4a82),
	.w5(32'h3b832709),
	.w6(32'h3be132bf),
	.w7(32'h3bf43fa6),
	.w8(32'hb9f8abb6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99cb0c),
	.w1(32'hba80d17b),
	.w2(32'hbb402ad5),
	.w3(32'hbb659cf0),
	.w4(32'hba138f8e),
	.w5(32'hbb677755),
	.w6(32'hba6e23e6),
	.w7(32'hbb30e6ea),
	.w8(32'h38c0c4de),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07eb1a),
	.w1(32'h39b8c04c),
	.w2(32'h3c6086cc),
	.w3(32'hbb21b858),
	.w4(32'h3b17c8dc),
	.w5(32'h3c68f82b),
	.w6(32'hbc24901c),
	.w7(32'h3b1fef68),
	.w8(32'h3c26784c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3521b),
	.w1(32'hb8874111),
	.w2(32'h3cc18aad),
	.w3(32'h3acf5cb8),
	.w4(32'hbcaceeb0),
	.w5(32'h3c9d7bc7),
	.w6(32'h3b801b19),
	.w7(32'hbbf9d051),
	.w8(32'h3c65388d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cefc996),
	.w1(32'h3b272616),
	.w2(32'h3c0e4cd5),
	.w3(32'h3ca63a57),
	.w4(32'hbb516a4f),
	.w5(32'h3a7e7e92),
	.w6(32'h3c73bc34),
	.w7(32'hba38e2b5),
	.w8(32'h3a7eec85),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba883381),
	.w1(32'hba96abfe),
	.w2(32'h395470fb),
	.w3(32'hbac3d2b6),
	.w4(32'h38256b8e),
	.w5(32'h3a1e85d2),
	.w6(32'hbb49380e),
	.w7(32'hba4f460f),
	.w8(32'h39ad8f15),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1be6a5),
	.w1(32'hbcb21ce0),
	.w2(32'h3d4ab82f),
	.w3(32'h3cb5a768),
	.w4(32'hbcf8754d),
	.w5(32'h3cc111ed),
	.w6(32'hbc192548),
	.w7(32'hbd4a50dc),
	.w8(32'h3c8df71d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefdbee),
	.w1(32'h3b211480),
	.w2(32'h3cb7559e),
	.w3(32'hbc30a94b),
	.w4(32'hbc2bbd73),
	.w5(32'h3c46a86b),
	.w6(32'hbb9812e0),
	.w7(32'hbc1b0666),
	.w8(32'h3bcff038),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a2a34),
	.w1(32'h3ac25538),
	.w2(32'hb92e4848),
	.w3(32'h3a62dc87),
	.w4(32'h3a92cc81),
	.w5(32'hba87910f),
	.w6(32'h3a96751a),
	.w7(32'hb93fbe08),
	.w8(32'h3a8de519),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae127c6),
	.w1(32'hbbcf2680),
	.w2(32'h3c890a30),
	.w3(32'hbc33e631),
	.w4(32'hbc906e8e),
	.w5(32'h3c3e0fbe),
	.w6(32'hbc56ecf6),
	.w7(32'hbcb273b5),
	.w8(32'h3b6395b7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fbd36),
	.w1(32'hb9256797),
	.w2(32'hb9be1129),
	.w3(32'hba48f615),
	.w4(32'h3aaf53ad),
	.w5(32'h3a93b774),
	.w6(32'hb8bc60e1),
	.w7(32'hb887037d),
	.w8(32'hb9c7bb2b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b050e),
	.w1(32'hbb1905c2),
	.w2(32'h3984d7b8),
	.w3(32'h3aa17160),
	.w4(32'hbb2d9a64),
	.w5(32'hba355376),
	.w6(32'h3a729167),
	.w7(32'hb88adaeb),
	.w8(32'h3ace760b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96fc86f),
	.w1(32'hb7ec5042),
	.w2(32'hbaaeef0f),
	.w3(32'hba5d033c),
	.w4(32'hb844230a),
	.w5(32'hbb0dfebc),
	.w6(32'hb9714e72),
	.w7(32'hbac9640d),
	.w8(32'hb97df475),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ba167),
	.w1(32'hb92a4f39),
	.w2(32'hba7b6ddf),
	.w3(32'hbac4a314),
	.w4(32'hb8b23ebc),
	.w5(32'hb7fe37e0),
	.w6(32'hb996de9d),
	.w7(32'hb9b82bf6),
	.w8(32'hb836e64f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c025451),
	.w1(32'hbae10e74),
	.w2(32'hbbcbc677),
	.w3(32'h3c1784da),
	.w4(32'hbaed3f38),
	.w5(32'hbc129458),
	.w6(32'h3c409afd),
	.w7(32'hbb5ea186),
	.w8(32'hbc11ff0f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45dd9f),
	.w1(32'h3d04f08e),
	.w2(32'h3d8eb4d9),
	.w3(32'hbbea40eb),
	.w4(32'hbabed65b),
	.w5(32'h3d3f8c13),
	.w6(32'hbc9a04bb),
	.w7(32'hbca58149),
	.w8(32'h3c8e4aa5),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c013e27),
	.w1(32'hba5a7983),
	.w2(32'h3ce5aa9e),
	.w3(32'hbc0b283b),
	.w4(32'hbc83fd74),
	.w5(32'h3c795253),
	.w6(32'hbc0a4987),
	.w7(32'hbca3e9b6),
	.w8(32'h3b8fb039),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2703a7),
	.w1(32'h3c5a43e3),
	.w2(32'h3d493587),
	.w3(32'hbbbd98ce),
	.w4(32'hbc54ab0f),
	.w5(32'h3d118ded),
	.w6(32'hbc6bdc3d),
	.w7(32'hbc959bc9),
	.w8(32'h3c809940),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69ba8f),
	.w1(32'h3a350593),
	.w2(32'h3b3a8189),
	.w3(32'hb97eb2a2),
	.w4(32'hba01fdd2),
	.w5(32'h3a9e2b5b),
	.w6(32'h3a92579a),
	.w7(32'h39d92df1),
	.w8(32'h3aad9e8e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b5d88),
	.w1(32'h3b35f353),
	.w2(32'h3a2d5998),
	.w3(32'h380a76e5),
	.w4(32'h3a4464b6),
	.w5(32'hba4daa67),
	.w6(32'h3a35ae13),
	.w7(32'h3acc691c),
	.w8(32'h3b2366cf),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d2a2e),
	.w1(32'h3a01399d),
	.w2(32'hba3cec75),
	.w3(32'hba87fb57),
	.w4(32'h3a76cc32),
	.w5(32'hb9eecb78),
	.w6(32'h38a12847),
	.w7(32'hba43fe8c),
	.w8(32'h36a02755),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373c97f1),
	.w1(32'h3a79e167),
	.w2(32'hba4da8d7),
	.w3(32'hb9270dac),
	.w4(32'h3ab5769f),
	.w5(32'hb9fbb5a5),
	.w6(32'h3a5d75fd),
	.w7(32'hb9debf22),
	.w8(32'h39874df6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a4c45),
	.w1(32'h3c5d44f6),
	.w2(32'h3d125f4c),
	.w3(32'h3b656d1c),
	.w4(32'hbbef4694),
	.w5(32'h3c872259),
	.w6(32'hbc12359d),
	.w7(32'hbbebaccd),
	.w8(32'h3c80c0ae),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa26c56),
	.w1(32'hb945f915),
	.w2(32'hbaef5ffb),
	.w3(32'hb7b79146),
	.w4(32'hb93f4ef4),
	.w5(32'hbb1e634f),
	.w6(32'hba53451d),
	.w7(32'hbaf6ae89),
	.w8(32'hb9a4b90c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babd559),
	.w1(32'hba8b8cd4),
	.w2(32'h3aeac48d),
	.w3(32'h3bac3dbd),
	.w4(32'h3a5cdab1),
	.w5(32'h3b5fbfa5),
	.w6(32'h3c3c5c9d),
	.w7(32'h3b1f2f3b),
	.w8(32'h3bbff93d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066e2d),
	.w1(32'h3b5180e1),
	.w2(32'h3bada6d6),
	.w3(32'h3be24c32),
	.w4(32'h3a05f237),
	.w5(32'h3ac123e1),
	.w6(32'h3be4eea3),
	.w7(32'h3b272717),
	.w8(32'h3ac6cfc9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cbe82d),
	.w1(32'h3a38b82e),
	.w2(32'hb979b5a8),
	.w3(32'h3a812b4e),
	.w4(32'h3a059c67),
	.w5(32'hba028eba),
	.w6(32'h3a3d6e67),
	.w7(32'hb85448d7),
	.w8(32'h39c8cf9f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd468c3),
	.w1(32'hbaac680f),
	.w2(32'h3bdec995),
	.w3(32'h395c6ba5),
	.w4(32'hbbc3d673),
	.w5(32'h3b6634b0),
	.w6(32'hbba97d8b),
	.w7(32'hbc0b51aa),
	.w8(32'h3ad7170e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b1129),
	.w1(32'h3b958b61),
	.w2(32'h3bd68906),
	.w3(32'h3a31398f),
	.w4(32'h3b44bf52),
	.w5(32'h3ba3f474),
	.w6(32'h3ae7035a),
	.w7(32'h3ba37d2e),
	.w8(32'h3b7f3279),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd335ad),
	.w1(32'h3cf51797),
	.w2(32'h3d8de355),
	.w3(32'hbc641154),
	.w4(32'h3b857f42),
	.w5(32'h3d308ed1),
	.w6(32'hbc06cf8e),
	.w7(32'hbb842dd0),
	.w8(32'h3cce0f38),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b5b98),
	.w1(32'hbac4fefe),
	.w2(32'hbb988804),
	.w3(32'hba7fe136),
	.w4(32'hbaa91655),
	.w5(32'hbb5080b5),
	.w6(32'hbb37117f),
	.w7(32'hb9d0795f),
	.w8(32'h3b45689a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cced0bb),
	.w1(32'h3a7d4a8f),
	.w2(32'hbc2295c2),
	.w3(32'h3b5fc5be),
	.w4(32'hbcc035da),
	.w5(32'hbcf56a12),
	.w6(32'h3d1e1633),
	.w7(32'h3c38ba44),
	.w8(32'hbbe68952),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule