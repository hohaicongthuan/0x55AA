module layer_8_featuremap_131(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa7859),
	.w1(32'h3a761d99),
	.w2(32'h3b25cb78),
	.w3(32'hbbc00025),
	.w4(32'hbb71667f),
	.w5(32'hbb6afd7b),
	.w6(32'hbbccc0a0),
	.w7(32'h3b0bf246),
	.w8(32'h3ba8b2b3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb29f34),
	.w1(32'h3b9119db),
	.w2(32'h3acdd377),
	.w3(32'hbbaea3d0),
	.w4(32'h3ac70397),
	.w5(32'h3c765d0a),
	.w6(32'h3b69cadf),
	.w7(32'h3b39e896),
	.w8(32'h3c96ddf3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c962855),
	.w1(32'h3c6bb672),
	.w2(32'h3b39a243),
	.w3(32'h3c0df0cb),
	.w4(32'h3b1ba9b0),
	.w5(32'h39bb1577),
	.w6(32'h3c5979e6),
	.w7(32'h3b364271),
	.w8(32'h3963d0eb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb670a95),
	.w1(32'h3af24af0),
	.w2(32'hbb9ae1ae),
	.w3(32'hba5ba26c),
	.w4(32'h3b867c29),
	.w5(32'h3b9777a6),
	.w6(32'hbb76480a),
	.w7(32'hbb8dcbe9),
	.w8(32'hbb4bcb26),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c9ef0),
	.w1(32'h3b99559d),
	.w2(32'hb9b8c55f),
	.w3(32'h3b800554),
	.w4(32'h3b01346a),
	.w5(32'h3b379182),
	.w6(32'hba113b47),
	.w7(32'hb898efae),
	.w8(32'hbb5de1c8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47f491),
	.w1(32'h39445e30),
	.w2(32'h3be09fde),
	.w3(32'h3b9853e3),
	.w4(32'h3c248296),
	.w5(32'h3c55e5d2),
	.w6(32'h3bdaa75b),
	.w7(32'h3c3cb0ec),
	.w8(32'h3c0f072a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27a3f4),
	.w1(32'h3c36c482),
	.w2(32'h3a639b58),
	.w3(32'h3c659e5f),
	.w4(32'h3bd272ad),
	.w5(32'h3b922d70),
	.w6(32'h3c36a8ee),
	.w7(32'h3bec753b),
	.w8(32'h3c94b5cd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b1967),
	.w1(32'h3c8c4611),
	.w2(32'hb8c4f52c),
	.w3(32'h3b7e299b),
	.w4(32'h3b5fcedb),
	.w5(32'h3b8025bb),
	.w6(32'h3c9312b8),
	.w7(32'hbb0527ce),
	.w8(32'hbb7a32dd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1de363),
	.w1(32'h3bf06964),
	.w2(32'h3b3ce014),
	.w3(32'hbbeb5672),
	.w4(32'h3be59dc4),
	.w5(32'h3b1fac02),
	.w6(32'hbbb34b8f),
	.w7(32'hbb425447),
	.w8(32'hbb0d086a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86cf41),
	.w1(32'h3a8652e5),
	.w2(32'h3c2db74c),
	.w3(32'hbb9412fa),
	.w4(32'h3c22b476),
	.w5(32'h3a407147),
	.w6(32'hbbc5f403),
	.w7(32'h3c0d6e09),
	.w8(32'h3c922088),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c396f87),
	.w1(32'h3bd6eee6),
	.w2(32'hbbaf491b),
	.w3(32'hbc082735),
	.w4(32'hbc2fe322),
	.w5(32'hba9213a5),
	.w6(32'h3bd2eeec),
	.w7(32'hbc00547e),
	.w8(32'hbbccac70),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe88e5),
	.w1(32'h3ba5835a),
	.w2(32'h3b950465),
	.w3(32'h3b2c955d),
	.w4(32'h3b64219f),
	.w5(32'h3b74eb3a),
	.w6(32'hba2f7b41),
	.w7(32'h3c007034),
	.w8(32'h3aa91704),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff3c7),
	.w1(32'h3bb33aed),
	.w2(32'h3b41cbc8),
	.w3(32'hbb3da63a),
	.w4(32'hbb17385e),
	.w5(32'hba7193d8),
	.w6(32'hb94642f2),
	.w7(32'hba89f53b),
	.w8(32'hbb8f8219),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6b9ed),
	.w1(32'hbbb3cf58),
	.w2(32'h3b05f751),
	.w3(32'hbb3fec99),
	.w4(32'h3a85a7fc),
	.w5(32'h390a7aef),
	.w6(32'hbbd75abc),
	.w7(32'h3adc9dfa),
	.w8(32'h3afd2aa4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26501b),
	.w1(32'hba96e80d),
	.w2(32'h39d2c2d1),
	.w3(32'hba5bc762),
	.w4(32'hb82f30ca),
	.w5(32'hbac144ef),
	.w6(32'hbaef2b69),
	.w7(32'hb9087cf1),
	.w8(32'h3a51a379),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac86bee),
	.w1(32'hba2a1964),
	.w2(32'h3bc753d8),
	.w3(32'hba1074b8),
	.w4(32'hbac9997a),
	.w5(32'hba8573f0),
	.w6(32'h3980f8e9),
	.w7(32'h3bd4767b),
	.w8(32'h3c5584ca),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb4f74),
	.w1(32'h3adf8950),
	.w2(32'hbb24592e),
	.w3(32'h3ad5d14a),
	.w4(32'h38e97022),
	.w5(32'hbbb808b4),
	.w6(32'h3c89ce2d),
	.w7(32'hba385ded),
	.w8(32'hbb2d2929),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92ba0d),
	.w1(32'hbb88de38),
	.w2(32'hbb45abea),
	.w3(32'hbc3e804e),
	.w4(32'h3bdfe2e2),
	.w5(32'hbb81da1d),
	.w6(32'hbbb39c64),
	.w7(32'hb9c8ebeb),
	.w8(32'h3b047eae),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5e278),
	.w1(32'hbc7c302f),
	.w2(32'hbbe0e6e7),
	.w3(32'hbc806913),
	.w4(32'hbc05efa7),
	.w5(32'hbb311023),
	.w6(32'hbcac4eb0),
	.w7(32'hbc214d94),
	.w8(32'hbba05e5a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb679d08),
	.w1(32'hbbac95f1),
	.w2(32'hbc8265d4),
	.w3(32'hbc254ecf),
	.w4(32'hbb6ac24e),
	.w5(32'hbbbbb10d),
	.w6(32'hbc328e9f),
	.w7(32'h3a8b8bfa),
	.w8(32'hbb96a1e4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc784a3b),
	.w1(32'h3b1d7ce5),
	.w2(32'h3a0de014),
	.w3(32'h3ba440aa),
	.w4(32'h3b5026b5),
	.w5(32'hbb90af8f),
	.w6(32'hbba1ea2c),
	.w7(32'hba767099),
	.w8(32'hbc218b22),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62cced),
	.w1(32'h3c257c57),
	.w2(32'hbb768ce4),
	.w3(32'h3acab891),
	.w4(32'h3b64349b),
	.w5(32'h3abb10fd),
	.w6(32'h3bdb5165),
	.w7(32'hbb070195),
	.w8(32'hbba2d069),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18db6c),
	.w1(32'hbb32a150),
	.w2(32'hbb88971f),
	.w3(32'hbb2c0839),
	.w4(32'hbc074408),
	.w5(32'h3ab65d43),
	.w6(32'hbb983a2f),
	.w7(32'hbc199785),
	.w8(32'hbc07e86c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea772c),
	.w1(32'hbbb51d35),
	.w2(32'hbb96da64),
	.w3(32'hbba70cc0),
	.w4(32'hbc290336),
	.w5(32'hbc1c19d9),
	.w6(32'hbc08bc48),
	.w7(32'hbc0ebc26),
	.w8(32'hbbdb2511),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e915c),
	.w1(32'hbaf8ac48),
	.w2(32'h3c746a86),
	.w3(32'hbb301557),
	.w4(32'h3baa9a1d),
	.w5(32'h3cf1d9ff),
	.w6(32'hbadda133),
	.w7(32'h3cbc32fb),
	.w8(32'h3d36b099),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce04eb8),
	.w1(32'h3ba1a74e),
	.w2(32'hbc3c448a),
	.w3(32'h3bfb5db5),
	.w4(32'h39ebb852),
	.w5(32'hbae76cbc),
	.w6(32'h3c3a9136),
	.w7(32'hbc0047ee),
	.w8(32'hbcc9da0d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae32fd8),
	.w1(32'h3c831700),
	.w2(32'hbb952620),
	.w3(32'hbbc78702),
	.w4(32'hbba5bd2f),
	.w5(32'hbc549e2f),
	.w6(32'h3b401321),
	.w7(32'hbc30086d),
	.w8(32'hbbcd94d7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39fd27),
	.w1(32'h39461048),
	.w2(32'hbc723600),
	.w3(32'hbcd5902a),
	.w4(32'h3b1f725c),
	.w5(32'hbc88e2f7),
	.w6(32'hbcefa74e),
	.w7(32'hbcb72319),
	.w8(32'hbca8dfb9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb825994),
	.w1(32'h3c09ee41),
	.w2(32'h3b8edd92),
	.w3(32'hbb8ece42),
	.w4(32'h3bf5a642),
	.w5(32'h3bdc6508),
	.w6(32'h3b27056b),
	.w7(32'h3beb4ad5),
	.w8(32'hbb22149e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad70079),
	.w1(32'h3a60b9e6),
	.w2(32'h3c727695),
	.w3(32'h3c24ada5),
	.w4(32'h3cb9daae),
	.w5(32'h3c91b305),
	.w6(32'h39ceb685),
	.w7(32'h3cdb3b45),
	.w8(32'h3bee1ba7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21fdf9),
	.w1(32'hbc50e16a),
	.w2(32'h3b8d7220),
	.w3(32'hba01dae2),
	.w4(32'h3aa51830),
	.w5(32'h3b2f871e),
	.w6(32'hbca48a5f),
	.w7(32'h3b393316),
	.w8(32'h3b8aee41),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cc9ab),
	.w1(32'h3b63e55b),
	.w2(32'h3aba5f6b),
	.w3(32'h3a80297c),
	.w4(32'hbb980786),
	.w5(32'hbbd5d754),
	.w6(32'h3aa364a0),
	.w7(32'hba001e00),
	.w8(32'hbb8725dd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac054),
	.w1(32'hbb86517f),
	.w2(32'h3baac765),
	.w3(32'hbbc9f9e8),
	.w4(32'h3b9b924b),
	.w5(32'h3bebca6d),
	.w6(32'hbb5e6634),
	.w7(32'h3c4383bd),
	.w8(32'h3be4d901),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b480fa6),
	.w1(32'hba887f55),
	.w2(32'hbc1a3025),
	.w3(32'h3c163310),
	.w4(32'h3bc26f61),
	.w5(32'hbc55e69c),
	.w6(32'h3aa73ee2),
	.w7(32'hbb505667),
	.w8(32'hbbc30f9e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb3b92),
	.w1(32'h3b272d56),
	.w2(32'hbb9cba7a),
	.w3(32'hbb70cfb6),
	.w4(32'hbb7de6ef),
	.w5(32'hbac2042a),
	.w6(32'hbaf338fd),
	.w7(32'hbb272e47),
	.w8(32'hbba1bb73),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80a7a7),
	.w1(32'hb9119395),
	.w2(32'h3c6bee15),
	.w3(32'hbb105e2f),
	.w4(32'h3b896145),
	.w5(32'h3cbd37f2),
	.w6(32'hbb92ac89),
	.w7(32'h3c02c1c6),
	.w8(32'h3c9542dd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c849e99),
	.w1(32'h3bc9edaf),
	.w2(32'h3bb47477),
	.w3(32'h3ca20623),
	.w4(32'hbb19534a),
	.w5(32'h385bb879),
	.w6(32'h3c0edefd),
	.w7(32'h3b8b2c82),
	.w8(32'h3bb2c9f4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7bfd3),
	.w1(32'hbb4663ab),
	.w2(32'h3a52b4c9),
	.w3(32'hbb40d6d6),
	.w4(32'hbb9a153b),
	.w5(32'h3ca07101),
	.w6(32'h3c06a6a3),
	.w7(32'hbb56d8db),
	.w8(32'h3c9644c8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3bfe4),
	.w1(32'h3bee673c),
	.w2(32'hbbea7840),
	.w3(32'h3c209530),
	.w4(32'hbbe5721e),
	.w5(32'hba955f07),
	.w6(32'h3c0d7461),
	.w7(32'hbb95fe39),
	.w8(32'hbb449620),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fbcf9),
	.w1(32'h3af61392),
	.w2(32'hbabbff54),
	.w3(32'hbba3f994),
	.w4(32'hbb8dc57f),
	.w5(32'hbb8f053d),
	.w6(32'hbb9df2e8),
	.w7(32'hbbcb76f1),
	.w8(32'hbb9bdc11),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e06ab),
	.w1(32'hbb35ddaa),
	.w2(32'h3bd9586b),
	.w3(32'hbbaa3242),
	.w4(32'hbb96771e),
	.w5(32'h3b7b3fc3),
	.w6(32'hbbeb5608),
	.w7(32'hba32bdec),
	.w8(32'h3c5ea8be),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13a974),
	.w1(32'h3bd89cb4),
	.w2(32'hba919649),
	.w3(32'h3c052f0d),
	.w4(32'h3b08edda),
	.w5(32'hbbc69e4f),
	.w6(32'h3bb218e6),
	.w7(32'hba922118),
	.w8(32'h3ae858c0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e5f40),
	.w1(32'h3b3ae128),
	.w2(32'h3bcd64ac),
	.w3(32'hbad8505e),
	.w4(32'hbb4f4431),
	.w5(32'h3bd8d91d),
	.w6(32'h3b01f621),
	.w7(32'hbb8235d4),
	.w8(32'hb974c3fd),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b970fb9),
	.w1(32'hbc565d2f),
	.w2(32'h3a3c5792),
	.w3(32'hbb0a3bc4),
	.w4(32'hbb416424),
	.w5(32'hbb358c34),
	.w6(32'hbc0a6847),
	.w7(32'hbb2f4027),
	.w8(32'hbbf3a4cb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc064b49),
	.w1(32'hbc162619),
	.w2(32'hbb1a1e2c),
	.w3(32'hbba7f25a),
	.w4(32'hbbb9e643),
	.w5(32'hbb6b73d3),
	.w6(32'hbc51f482),
	.w7(32'hbb3fad14),
	.w8(32'hbb9ea270),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8476d),
	.w1(32'h38947a38),
	.w2(32'h3aaac846),
	.w3(32'hbb3ba8a1),
	.w4(32'hbb2fe8ec),
	.w5(32'hbb71685a),
	.w6(32'hbb6cde48),
	.w7(32'h3c37b25c),
	.w8(32'h3c36489a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed488e),
	.w1(32'hbbe72db5),
	.w2(32'hbbc2aba9),
	.w3(32'h3ae679e9),
	.w4(32'hba86b477),
	.w5(32'h3a40a2f9),
	.w6(32'h3c5de1db),
	.w7(32'hbb68e471),
	.w8(32'hbc287d84),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb622b99),
	.w1(32'hbbf7570c),
	.w2(32'h3ac03a15),
	.w3(32'hb9d67462),
	.w4(32'hbbd242ba),
	.w5(32'hbbcfac4b),
	.w6(32'hbc57d50a),
	.w7(32'hbb876dee),
	.w8(32'hbc04b8b9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b18ad),
	.w1(32'hbc2fc539),
	.w2(32'h3ad01db0),
	.w3(32'hbb8172d4),
	.w4(32'hbb419355),
	.w5(32'hbbb41659),
	.w6(32'hbc50be83),
	.w7(32'hbb8f6781),
	.w8(32'hba5d582e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e57f4),
	.w1(32'hbaf9dc0e),
	.w2(32'hb9707351),
	.w3(32'hbbc3013b),
	.w4(32'hbc2bd9a3),
	.w5(32'hbb3aff22),
	.w6(32'hbb99fa9e),
	.w7(32'hbb8221f3),
	.w8(32'h3bf9913d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88ed5d),
	.w1(32'hbb3ec965),
	.w2(32'h3c8b4001),
	.w3(32'hbae93fe5),
	.w4(32'h3c98edc8),
	.w5(32'h3c391999),
	.w6(32'hba85d754),
	.w7(32'h3c9c072e),
	.w8(32'h3ba0e2d3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf56a5),
	.w1(32'h39c8b7e0),
	.w2(32'h3b4b209b),
	.w3(32'h3b8a815a),
	.w4(32'h3b646749),
	.w5(32'hbbf17aa6),
	.w6(32'hbc6f1a44),
	.w7(32'hbc551ea4),
	.w8(32'hbc863c16),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2385d1),
	.w1(32'h3b7679bc),
	.w2(32'h3bb2fa51),
	.w3(32'hbba54524),
	.w4(32'hbbf237fe),
	.w5(32'h3b974a5e),
	.w6(32'hbc437f71),
	.w7(32'hbbcbcf4b),
	.w8(32'h3c065772),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15a806),
	.w1(32'h3ad48f96),
	.w2(32'h3b7ad882),
	.w3(32'h3c0f786c),
	.w4(32'hba1d505d),
	.w5(32'hb9ac71e8),
	.w6(32'hba1dd8db),
	.w7(32'h3af19de8),
	.w8(32'h3a16c6b5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27c816),
	.w1(32'hbb461260),
	.w2(32'hba95e757),
	.w3(32'h3a099f22),
	.w4(32'h3c12cec0),
	.w5(32'h3ba05be1),
	.w6(32'hbb3565d1),
	.w7(32'h3bafeee7),
	.w8(32'hbbe67783),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c20f5),
	.w1(32'hbaf58542),
	.w2(32'hbbd21462),
	.w3(32'hbb04470b),
	.w4(32'hbb9e3e22),
	.w5(32'hbbc2b689),
	.w6(32'h396d2c36),
	.w7(32'hbbee6905),
	.w8(32'hbb3c2385),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69aa0),
	.w1(32'h3b954992),
	.w2(32'hba2d21b0),
	.w3(32'hbb60fd91),
	.w4(32'h3a7e12ae),
	.w5(32'hbbd23d54),
	.w6(32'hbb3fd336),
	.w7(32'hbbc9444a),
	.w8(32'hbb961f21),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb6614),
	.w1(32'h3c15dbe9),
	.w2(32'h3b444f6e),
	.w3(32'hba8268a6),
	.w4(32'h3c65406c),
	.w5(32'h3bd63fbf),
	.w6(32'h39f5c59c),
	.w7(32'h3bb7d08d),
	.w8(32'hbaba7684),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b9886),
	.w1(32'hbb0acca9),
	.w2(32'h3b914d02),
	.w3(32'h3b90efbc),
	.w4(32'h3a9dc274),
	.w5(32'h3b103ed9),
	.w6(32'h3a174cf9),
	.w7(32'h3b2c6663),
	.w8(32'hba33f80f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8054f8),
	.w1(32'hbb9df96c),
	.w2(32'hbb39aff5),
	.w3(32'hb8f9c1f2),
	.w4(32'hbc4ca77d),
	.w5(32'hbb0d5055),
	.w6(32'hbb9fbb86),
	.w7(32'hbc879a51),
	.w8(32'hbb05d502),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c166015),
	.w1(32'h3ca84c37),
	.w2(32'h3bc30ce5),
	.w3(32'hbb944dd3),
	.w4(32'h3ac20d23),
	.w5(32'h3af01150),
	.w6(32'h3c3fce30),
	.w7(32'h3a2ba827),
	.w8(32'h3c5505fd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffb1c8),
	.w1(32'h3b9cbf34),
	.w2(32'hbb851eb5),
	.w3(32'h3a54c2b7),
	.w4(32'h39cb5b62),
	.w5(32'hb9fb1ccc),
	.w6(32'hbb9bfe5c),
	.w7(32'h3c38fc57),
	.w8(32'h3c21d87c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5b968),
	.w1(32'hbb4f6dc6),
	.w2(32'h3a4eb0c5),
	.w3(32'hbb07b822),
	.w4(32'h3a23d583),
	.w5(32'h3b016f24),
	.w6(32'h3b6fb12c),
	.w7(32'hba5c886f),
	.w8(32'hba5368f3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89fe18),
	.w1(32'h3b2d72ba),
	.w2(32'h3af4b748),
	.w3(32'hbb0d6e5a),
	.w4(32'hbc32fd3e),
	.w5(32'hbc058470),
	.w6(32'hbb95b156),
	.w7(32'hbb67b60f),
	.w8(32'hbb9c5f8a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e5124),
	.w1(32'h3abe8bb0),
	.w2(32'hbbb0d2b2),
	.w3(32'hbab97375),
	.w4(32'h3bb8d0d6),
	.w5(32'h3b55c300),
	.w6(32'hbab53bab),
	.w7(32'h3c3eb1c3),
	.w8(32'h3ac109b1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7be80),
	.w1(32'hbb841be5),
	.w2(32'hbb0a0c00),
	.w3(32'h3b2ce6be),
	.w4(32'h3ae95412),
	.w5(32'h3c7baa7a),
	.w6(32'h3b33ed94),
	.w7(32'h39f790a0),
	.w8(32'h3bff1482),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde3b5b),
	.w1(32'hbb65b376),
	.w2(32'hbc15e314),
	.w3(32'hb93a861b),
	.w4(32'h3b97215e),
	.w5(32'h3b6c3030),
	.w6(32'hbb83b5b1),
	.w7(32'h3a9af6df),
	.w8(32'hbb3e18a6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf0aff),
	.w1(32'hbb08b95a),
	.w2(32'h3c3a8f5a),
	.w3(32'hbb91d1ab),
	.w4(32'hbc04fb90),
	.w5(32'hbc066b71),
	.w6(32'hbb92a155),
	.w7(32'h3829330c),
	.w8(32'h3a4dd7a4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95ad09),
	.w1(32'hba9a5123),
	.w2(32'h3bc5f86d),
	.w3(32'h3bdfa5ea),
	.w4(32'hba75fcc8),
	.w5(32'h38d18ab7),
	.w6(32'h3c6feed3),
	.w7(32'h3bb3efc2),
	.w8(32'h3bd77d89),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af40089),
	.w1(32'hbc06d559),
	.w2(32'hba380105),
	.w3(32'hbc02fb3b),
	.w4(32'h3aa1183f),
	.w5(32'hbb8e541d),
	.w6(32'hbbd3053b),
	.w7(32'hbc2dc2f7),
	.w8(32'hbae8d4ec),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b516a23),
	.w1(32'h3b66097a),
	.w2(32'hbae197f8),
	.w3(32'h3c3d74ce),
	.w4(32'h3b963621),
	.w5(32'hbb73a8ba),
	.w6(32'h3aa31de0),
	.w7(32'hbc05f68a),
	.w8(32'hbc2c6fc9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34bcdb),
	.w1(32'hbb8c0fb8),
	.w2(32'hbc07e5b1),
	.w3(32'hbb1d77c2),
	.w4(32'hbc0d606d),
	.w5(32'hbc3b7a3e),
	.w6(32'hbc108bd7),
	.w7(32'hbbfcbb81),
	.w8(32'hbc00238b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7167e),
	.w1(32'hba37662b),
	.w2(32'h3c26224b),
	.w3(32'hbc012699),
	.w4(32'hbb0b6ffc),
	.w5(32'h39ef3de4),
	.w6(32'hbbfcb346),
	.w7(32'h3cba345d),
	.w8(32'h3cd5940c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30d447),
	.w1(32'h3b3c327f),
	.w2(32'h3c6515da),
	.w3(32'h3c0a9f6b),
	.w4(32'h3b46c12d),
	.w5(32'h3c4f7b87),
	.w6(32'h3cbf54fa),
	.w7(32'hba56ab3c),
	.w8(32'h3b374373),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ca821),
	.w1(32'h3b53f68e),
	.w2(32'hbb86d98c),
	.w3(32'h3c419abb),
	.w4(32'hbaf7d90d),
	.w5(32'hbaefc0ba),
	.w6(32'h3b98ed3e),
	.w7(32'hbb66c847),
	.w8(32'hbbdac2fc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7115bb),
	.w1(32'hbba85396),
	.w2(32'hbb7e130d),
	.w3(32'hbbca3e88),
	.w4(32'hbb578f0c),
	.w5(32'hbb579b2f),
	.w6(32'hbbfde76b),
	.w7(32'hbb243308),
	.w8(32'hba8f2879),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab831d1),
	.w1(32'hba3fd2fa),
	.w2(32'h3bc94e5d),
	.w3(32'hbb84215a),
	.w4(32'h3b469f21),
	.w5(32'hbb819bdc),
	.w6(32'hbbdbd51b),
	.w7(32'h3c3f4bb9),
	.w8(32'h3aed7206),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f724e3),
	.w1(32'h3b2324d6),
	.w2(32'hbb8109d9),
	.w3(32'hba69ce56),
	.w4(32'hbc1d594c),
	.w5(32'h3b0b848e),
	.w6(32'hbc004fb6),
	.w7(32'hbc59c488),
	.w8(32'hbb8998e6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec9dc4),
	.w1(32'h3bc7225f),
	.w2(32'h3b19ccd9),
	.w3(32'h3bd613be),
	.w4(32'hb9785895),
	.w5(32'h3ab87045),
	.w6(32'h3b9eefa0),
	.w7(32'hbb4497ec),
	.w8(32'hba50bebe),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e4403),
	.w1(32'h3c3eab52),
	.w2(32'hbc200063),
	.w3(32'h3c459c41),
	.w4(32'hbb70cd60),
	.w5(32'h3be2d61c),
	.w6(32'h3c245555),
	.w7(32'h3c079180),
	.w8(32'h3b7619f1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b31e8),
	.w1(32'h3c091a73),
	.w2(32'hbc31ab24),
	.w3(32'h3b7bd752),
	.w4(32'hbd245df6),
	.w5(32'hbb74da95),
	.w6(32'hbb358606),
	.w7(32'hbc535799),
	.w8(32'h3d62301c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbab07f),
	.w1(32'h3ad9ed84),
	.w2(32'h3c21aec0),
	.w3(32'h3ba129a9),
	.w4(32'h3c106b65),
	.w5(32'h3c2c7791),
	.w6(32'h3ca5256b),
	.w7(32'h3c1259c5),
	.w8(32'h3c9a6c04),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc44fa3),
	.w1(32'hbc403d52),
	.w2(32'hbc225dac),
	.w3(32'hbc632d8b),
	.w4(32'hbc6ed88b),
	.w5(32'hbc2f897b),
	.w6(32'hbce5ed38),
	.w7(32'hbc7b398c),
	.w8(32'hbb69dae5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5e23e),
	.w1(32'h3bffb147),
	.w2(32'h3a7fbb32),
	.w3(32'hbbf6dcf7),
	.w4(32'h3b09debd),
	.w5(32'h3c0ef49b),
	.w6(32'hbc979ba5),
	.w7(32'hbaacb2f5),
	.w8(32'hbb79bf23),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcda40),
	.w1(32'hbb25a260),
	.w2(32'hbcc220ea),
	.w3(32'hbc3dea04),
	.w4(32'hbcd943e2),
	.w5(32'h3b0258d8),
	.w6(32'hbc8401d9),
	.w7(32'hbd3b29e1),
	.w8(32'h39b3de26),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb80de3),
	.w1(32'h3c835d9c),
	.w2(32'hbbdeb45f),
	.w3(32'h3cde7ce6),
	.w4(32'hbb96fb6a),
	.w5(32'hbb99cb0c),
	.w6(32'h3d4ec990),
	.w7(32'hba713d0b),
	.w8(32'hbc646422),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca3631),
	.w1(32'hbbc586ca),
	.w2(32'h3c01a22a),
	.w3(32'h3c839e18),
	.w4(32'h3c1448f8),
	.w5(32'hba9502f9),
	.w6(32'h3cc7d825),
	.w7(32'h3c1530f7),
	.w8(32'hbc214950),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb914f27),
	.w1(32'hbca7a9a5),
	.w2(32'h3bd58c49),
	.w3(32'hbcb06dcb),
	.w4(32'h3c196b4a),
	.w5(32'h3c00ba07),
	.w6(32'hbccfa4d1),
	.w7(32'h3c240b05),
	.w8(32'h39e193ff),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd27f3),
	.w1(32'h3bfb9341),
	.w2(32'h3b45548b),
	.w3(32'h3c35da7f),
	.w4(32'h3c5d0c7b),
	.w5(32'h3b8384f6),
	.w6(32'h3c63f5ad),
	.w7(32'h3bd093f3),
	.w8(32'hbba7ab61),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc8dd3),
	.w1(32'h3b53caca),
	.w2(32'hbc3440e3),
	.w3(32'h3b202fed),
	.w4(32'hbc88f6a4),
	.w5(32'hbb3d28b6),
	.w6(32'hbab0720e),
	.w7(32'hbb546437),
	.w8(32'h3c586d71),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaf22b),
	.w1(32'h3bb704bb),
	.w2(32'h39103a95),
	.w3(32'hbb1a8c77),
	.w4(32'h3b4a8a59),
	.w5(32'h3b84c155),
	.w6(32'h3cf37ee6),
	.w7(32'hbbf4ba90),
	.w8(32'hbc9ee604),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c502c),
	.w1(32'h3ae5b655),
	.w2(32'hbb1ee869),
	.w3(32'h3aa37409),
	.w4(32'hbc4a908f),
	.w5(32'h3c88a0e1),
	.w6(32'h3b8792dc),
	.w7(32'hbc4da18d),
	.w8(32'h397568a9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf77171),
	.w1(32'h3c7a13e3),
	.w2(32'h3bf7304a),
	.w3(32'hba800b71),
	.w4(32'hbb9d683f),
	.w5(32'h3c0aff54),
	.w6(32'hbb79eab8),
	.w7(32'h3bb56349),
	.w8(32'hbc9b0d13),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e3769),
	.w1(32'hbab5f595),
	.w2(32'hbb73f1ab),
	.w3(32'h3b80043d),
	.w4(32'hbb851f67),
	.w5(32'hbccb621f),
	.w6(32'hbc6d84bc),
	.w7(32'hba7b04cf),
	.w8(32'hbd3100e9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc79006),
	.w1(32'h3c2c0df5),
	.w2(32'h3c335458),
	.w3(32'h3b54132d),
	.w4(32'h3b966418),
	.w5(32'h3c21fb02),
	.w6(32'h3d0b6eaa),
	.w7(32'h3c31dd9e),
	.w8(32'h3c7de354),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25da86),
	.w1(32'h3c16b9a4),
	.w2(32'hbb64312d),
	.w3(32'h3bc39a1a),
	.w4(32'hbc4df175),
	.w5(32'h3b57585d),
	.w6(32'h3c08222a),
	.w7(32'h3c26bd32),
	.w8(32'hbb4347a7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bd5e5),
	.w1(32'h3bb4ae71),
	.w2(32'h3cb929f9),
	.w3(32'hbbf96ddc),
	.w4(32'hbc8422fa),
	.w5(32'hbd1cd7c5),
	.w6(32'hbbf722b4),
	.w7(32'h3abf1b34),
	.w8(32'hbbc225cb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0c197f),
	.w1(32'hbc8103a1),
	.w2(32'hbcc53f40),
	.w3(32'h3bc5156a),
	.w4(32'hbcecb4d4),
	.w5(32'hbc8cc9c6),
	.w6(32'hbc2ba3d9),
	.w7(32'hbca7d5a2),
	.w8(32'h3c80840d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c022b9d),
	.w1(32'h3ba944d3),
	.w2(32'h3c4df3e9),
	.w3(32'hbbc0eafe),
	.w4(32'h3c604c61),
	.w5(32'h3c03686c),
	.w6(32'h3d2c82cd),
	.w7(32'h3c315a3f),
	.w8(32'h3b8e64aa),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aac5d),
	.w1(32'hbb3b202d),
	.w2(32'h3cb7c6e5),
	.w3(32'h3873575a),
	.w4(32'h3cc868bf),
	.w5(32'hbc540ac7),
	.w6(32'h3a03c3bd),
	.w7(32'h3cfe6189),
	.w8(32'hbd051806),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6850e),
	.w1(32'hbcea2c3e),
	.w2(32'hbc2d2182),
	.w3(32'hbd063345),
	.w4(32'hbac4beb2),
	.w5(32'h3ba112b4),
	.w6(32'hbd62c430),
	.w7(32'hbc0b2f29),
	.w8(32'hbbeea4cf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2279ae),
	.w1(32'hbc0f4348),
	.w2(32'hbb79007d),
	.w3(32'hba803d0a),
	.w4(32'hbb035b86),
	.w5(32'h3aace7bc),
	.w6(32'hbc3e492e),
	.w7(32'h3c711840),
	.w8(32'h3c533098),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b000681),
	.w1(32'hba2e2032),
	.w2(32'h3bb909ec),
	.w3(32'hbb9b49d4),
	.w4(32'hbbfa5bb2),
	.w5(32'h3b7dab34),
	.w6(32'hb954efd1),
	.w7(32'h3ac03178),
	.w8(32'h3b68bf7b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5cd5f),
	.w1(32'h3c845526),
	.w2(32'h3c8c3e89),
	.w3(32'hbc162831),
	.w4(32'h3c48025c),
	.w5(32'h3be2cd80),
	.w6(32'hbb31e854),
	.w7(32'h3c01086f),
	.w8(32'hbbbfb3ab),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0502c),
	.w1(32'h3b2fbef2),
	.w2(32'hbbbfe1a3),
	.w3(32'h3bc5ad39),
	.w4(32'h3b268e97),
	.w5(32'hbc34c134),
	.w6(32'hbc2ea023),
	.w7(32'h3b9da7ed),
	.w8(32'hbc646194),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb10892),
	.w1(32'h3cdd2dbe),
	.w2(32'h3c23281a),
	.w3(32'h3bf0acff),
	.w4(32'h3c72a97c),
	.w5(32'hbc82992a),
	.w6(32'h3cee68eb),
	.w7(32'h3c19ab23),
	.w8(32'hbc937834),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22d90b),
	.w1(32'hbc2b85f0),
	.w2(32'h3c1190be),
	.w3(32'hbc55d2b1),
	.w4(32'hbc41e45a),
	.w5(32'hbc8e23cd),
	.w6(32'hbce93a8f),
	.w7(32'h3b9b3cab),
	.w8(32'hbbe87137),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b402f3f),
	.w1(32'hbc48b403),
	.w2(32'h3c2eb5f3),
	.w3(32'hb909b650),
	.w4(32'h3b245985),
	.w5(32'hbc0427c0),
	.w6(32'hbcca5971),
	.w7(32'h3c614065),
	.w8(32'hba80ebc2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c1aef3),
	.w1(32'h3be69dac),
	.w2(32'h3b23d42e),
	.w3(32'h3b701dcf),
	.w4(32'hbc5f96c9),
	.w5(32'hbbb05c7c),
	.w6(32'h3a086841),
	.w7(32'hbc1489c7),
	.w8(32'h3a5f4b91),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c23aa),
	.w1(32'hba9c6304),
	.w2(32'h3c9a5729),
	.w3(32'h3bccd747),
	.w4(32'h3ccfd180),
	.w5(32'h3c484a76),
	.w6(32'hbb02b23c),
	.w7(32'h3d2a7c24),
	.w8(32'hb9f108fe),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49de0b),
	.w1(32'hbcc0d218),
	.w2(32'h3b9e538c),
	.w3(32'hbcc31001),
	.w4(32'hbb242cf4),
	.w5(32'hb98824ed),
	.w6(32'hbd83af0e),
	.w7(32'h3c33a7b0),
	.w8(32'hbbef8564),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30964c),
	.w1(32'hbbff50e2),
	.w2(32'hbc65ee05),
	.w3(32'h3bcb8e30),
	.w4(32'hbbb46e20),
	.w5(32'hbb07bf67),
	.w6(32'hbbcbb509),
	.w7(32'hbc88ab35),
	.w8(32'hbbe42077),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb50258),
	.w1(32'hbc3bc84a),
	.w2(32'hbc3deb4a),
	.w3(32'h3c3f4af1),
	.w4(32'hbb44c8d1),
	.w5(32'hbb6e6b12),
	.w6(32'hbb814495),
	.w7(32'hbc2c3ba1),
	.w8(32'h3c840571),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01c198),
	.w1(32'hbc062dc3),
	.w2(32'hbcb1925f),
	.w3(32'h3be1b9bb),
	.w4(32'hbca22603),
	.w5(32'hbcb08bca),
	.w6(32'h3a919133),
	.w7(32'hbc2cacf3),
	.w8(32'hbc722d12),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc840838),
	.w1(32'hba80a1a3),
	.w2(32'hbc343e72),
	.w3(32'hbbf18385),
	.w4(32'hbc085dfb),
	.w5(32'h3ba63b95),
	.w6(32'hbb21a14f),
	.w7(32'hbb4b8924),
	.w8(32'h3ca0f239),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ed53b),
	.w1(32'hba124a7b),
	.w2(32'hbccb9a65),
	.w3(32'h3aee13e0),
	.w4(32'hbd41334c),
	.w5(32'h3a79ebd7),
	.w6(32'hbc2443f4),
	.w7(32'hbd047087),
	.w8(32'h3d11b888),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac5315),
	.w1(32'h3c881d2e),
	.w2(32'hbb900868),
	.w3(32'h3bec9d80),
	.w4(32'hbc46eae3),
	.w5(32'hbb677b0a),
	.w6(32'h3d30bcec),
	.w7(32'hbc57e9f4),
	.w8(32'h3c1c723a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fecaf),
	.w1(32'h3ba44632),
	.w2(32'h3bc99fe1),
	.w3(32'h3b0fdb1d),
	.w4(32'hb9ddc28b),
	.w5(32'hbb0a81ab),
	.w6(32'h3af84f2a),
	.w7(32'h3b63d8fd),
	.w8(32'hbafbefb8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c434),
	.w1(32'h3bb1dfac),
	.w2(32'hbc5ff886),
	.w3(32'h3b8d2b60),
	.w4(32'hba5f492d),
	.w5(32'hbc6b0e27),
	.w6(32'h3a9ca6d2),
	.w7(32'hbc88a4a0),
	.w8(32'hbcce6ae5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7f0c3),
	.w1(32'h3bb2a71b),
	.w2(32'hbc7ec2d2),
	.w3(32'hbacfc812),
	.w4(32'hbb227ddb),
	.w5(32'hbbf687e2),
	.w6(32'hbb8ecf0a),
	.w7(32'hbbbea437),
	.w8(32'hbc0b6cb9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40cae5),
	.w1(32'hbbc2f670),
	.w2(32'h3b9760f7),
	.w3(32'hbbdb20bb),
	.w4(32'h3bec0f44),
	.w5(32'h3992e12a),
	.w6(32'hbc79bfec),
	.w7(32'h39711dc8),
	.w8(32'hbb2185e4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbabdbf),
	.w1(32'h3ba57c27),
	.w2(32'hbc10dd5b),
	.w3(32'hb9acf481),
	.w4(32'h3b90fcea),
	.w5(32'h3d1ea19d),
	.w6(32'h3a02ed8e),
	.w7(32'hbae3ab69),
	.w8(32'h3b642c21),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd20833),
	.w1(32'h3bb4f23f),
	.w2(32'h3bf45f05),
	.w3(32'hbb2cf4ec),
	.w4(32'hba4304b5),
	.w5(32'hbbf85531),
	.w6(32'hbc52f7ea),
	.w7(32'h3c0b92ee),
	.w8(32'hbb3258e1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7f7cc),
	.w1(32'h3c07277d),
	.w2(32'hbb116895),
	.w3(32'h3b92ebb2),
	.w4(32'hbb44dcbe),
	.w5(32'h3c979473),
	.w6(32'h3b20292e),
	.w7(32'hbc4b98f9),
	.w8(32'h3d0ffebf),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c264499),
	.w1(32'hbc5f2226),
	.w2(32'hbb459cf5),
	.w3(32'hbc6788ba),
	.w4(32'h3925bffe),
	.w5(32'hbc818dc7),
	.w6(32'hbccbc3aa),
	.w7(32'h3aeed21b),
	.w8(32'hbd0f4348),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fc29b),
	.w1(32'h3bdc29fa),
	.w2(32'h3b8b586f),
	.w3(32'hbc5e53d1),
	.w4(32'h3b2734ab),
	.w5(32'hbb432a0c),
	.w6(32'hbcabdfe3),
	.w7(32'h3b1049bc),
	.w8(32'hbc0528ad),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea8292),
	.w1(32'hbb01b470),
	.w2(32'hbc43308a),
	.w3(32'h3c17077d),
	.w4(32'hb9c899d9),
	.w5(32'hba887a87),
	.w6(32'h3b3353ab),
	.w7(32'hbc1b985f),
	.w8(32'hbc55afb6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fdadd),
	.w1(32'h3cf148a8),
	.w2(32'h3baac698),
	.w3(32'h3ce395e8),
	.w4(32'h3b575868),
	.w5(32'h3b36a91d),
	.w6(32'h3d1be327),
	.w7(32'h3aa98cca),
	.w8(32'h3b3f6d7f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule