module layer_8_featuremap_241(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda6a8b),
	.w1(32'hbc12e5d4),
	.w2(32'hbb8e92e4),
	.w3(32'h3b1fcd53),
	.w4(32'h3b3e265a),
	.w5(32'h3b747de6),
	.w6(32'h39e9d932),
	.w7(32'h3abd7984),
	.w8(32'hbbaacff2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c074b),
	.w1(32'h3bb728a0),
	.w2(32'h3b819123),
	.w3(32'h3c06a698),
	.w4(32'h3c1da678),
	.w5(32'h3bcf08d1),
	.w6(32'h3bab9873),
	.w7(32'h3a868cb1),
	.w8(32'h3ac20a8b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3e2a1),
	.w1(32'h3abdf0c7),
	.w2(32'h3b8c5667),
	.w3(32'h3babac08),
	.w4(32'h3b171afc),
	.w5(32'hbb2c757d),
	.w6(32'hbb811fe1),
	.w7(32'hbbb42baa),
	.w8(32'h3b2a4a94),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b875ebe),
	.w1(32'hbbd9802f),
	.w2(32'h3ac86835),
	.w3(32'hb9681c79),
	.w4(32'hbbcc71c4),
	.w5(32'hbb46f3fb),
	.w6(32'hba0aa027),
	.w7(32'hba8ddbc0),
	.w8(32'h3bdfa4e0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52e9ea),
	.w1(32'h3a3ecf9e),
	.w2(32'hbb9bd67f),
	.w3(32'h3c274f20),
	.w4(32'h3b6f47d6),
	.w5(32'hbadbb42f),
	.w6(32'h3bb4ebbf),
	.w7(32'h3b16272f),
	.w8(32'hbb3ec887),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0be4d),
	.w1(32'hbaf5af74),
	.w2(32'hbc348f5a),
	.w3(32'hba079c56),
	.w4(32'hbbfbbcb6),
	.w5(32'hbc28b2d4),
	.w6(32'hb95f3b2f),
	.w7(32'hbc0a7828),
	.w8(32'hbc513a55),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3df243),
	.w1(32'hbb05d650),
	.w2(32'hbb5d6671),
	.w3(32'hbbda7a5e),
	.w4(32'hbaf8829f),
	.w5(32'hbb45f930),
	.w6(32'hbb6303a4),
	.w7(32'hbb5e229d),
	.w8(32'hbba5aa68),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d4b1f),
	.w1(32'hbab37302),
	.w2(32'hbaeca59a),
	.w3(32'hbb9c291c),
	.w4(32'hbb09a158),
	.w5(32'hbba79e36),
	.w6(32'h39990666),
	.w7(32'hbb88c336),
	.w8(32'hbb8a9c45),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb83b1a),
	.w1(32'h3b9140e4),
	.w2(32'hbb75a25e),
	.w3(32'h3c0dbf74),
	.w4(32'h3bea327d),
	.w5(32'hbb655809),
	.w6(32'hb8958f5f),
	.w7(32'hbbe81c59),
	.w8(32'hbbc63270),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58432f),
	.w1(32'h3ad0f2ca),
	.w2(32'h3be8f549),
	.w3(32'h3bf504d4),
	.w4(32'h3c0530d7),
	.w5(32'h3c65fc48),
	.w6(32'h3a93fd4a),
	.w7(32'h3a89c65d),
	.w8(32'h3bc5b91c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9183d5),
	.w1(32'hbbd0f889),
	.w2(32'h3bf74196),
	.w3(32'h3cc2855d),
	.w4(32'hbb55b546),
	.w5(32'h3be47e04),
	.w6(32'hbaf7caed),
	.w7(32'h3bb60dee),
	.w8(32'h3b8156ee),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9aab5),
	.w1(32'hbb299baf),
	.w2(32'hbbfbadd2),
	.w3(32'h3bfe7c25),
	.w4(32'h3b24a5cb),
	.w5(32'hb9c174d6),
	.w6(32'h3af0c015),
	.w7(32'h3bafc7cd),
	.w8(32'hbb3062f4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9d0f4),
	.w1(32'h37d1db38),
	.w2(32'h3ba84db9),
	.w3(32'hba263690),
	.w4(32'h3c0532b6),
	.w5(32'h3c0bd199),
	.w6(32'hbb5c3e4b),
	.w7(32'hbbdcd974),
	.w8(32'hbb5835b7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34abd),
	.w1(32'h3b27a17b),
	.w2(32'hbb55a13e),
	.w3(32'h3b9d060d),
	.w4(32'hba98b9b0),
	.w5(32'h3b70391c),
	.w6(32'hbb87a86a),
	.w7(32'h3aa4a6b3),
	.w8(32'h3bc8185c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed3133),
	.w1(32'h3ad5285c),
	.w2(32'hbaf5b643),
	.w3(32'h3c35e85d),
	.w4(32'h39fc7642),
	.w5(32'hbb4d2c48),
	.w6(32'hb9216059),
	.w7(32'hbb12660e),
	.w8(32'hbaca95a2),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3249cf),
	.w1(32'h3bd35a36),
	.w2(32'h3af921a7),
	.w3(32'hbb06a846),
	.w4(32'h3bb96558),
	.w5(32'h3ba95bb4),
	.w6(32'h3adb8d03),
	.w7(32'h3ad38031),
	.w8(32'hbbce1616),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8207c9),
	.w1(32'hbc1a5781),
	.w2(32'hbc0735cd),
	.w3(32'hbae7f6a3),
	.w4(32'hbbd84045),
	.w5(32'hbc08b26e),
	.w6(32'hbc057c1f),
	.w7(32'hbc213926),
	.w8(32'hbc010e90),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdbf12),
	.w1(32'hbb37b399),
	.w2(32'hbc155c2a),
	.w3(32'hbb94c270),
	.w4(32'hbbf93664),
	.w5(32'h394cf085),
	.w6(32'hbb8193a7),
	.w7(32'hbb0dc0a4),
	.w8(32'h3b2721f7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d43ad),
	.w1(32'hbd2f732f),
	.w2(32'hbcf1c840),
	.w3(32'hb7b5ce16),
	.w4(32'hbcc3b8ec),
	.w5(32'hbc57f525),
	.w6(32'h3c48b3c5),
	.w7(32'hba42fbd5),
	.w8(32'h3b3b951f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8a3a7),
	.w1(32'hbc682d15),
	.w2(32'hbc826add),
	.w3(32'h3c70b575),
	.w4(32'hbb04c5d6),
	.w5(32'hbaf58415),
	.w6(32'h3bbcdd54),
	.w7(32'h3a32a241),
	.w8(32'hbab65808),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb913ea6),
	.w1(32'hbb420305),
	.w2(32'hbc161de8),
	.w3(32'h3b48ecbe),
	.w4(32'h3abad331),
	.w5(32'hbc2ccc2d),
	.w6(32'hbb523691),
	.w7(32'h3b6bceed),
	.w8(32'hbba65dc6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08a42b),
	.w1(32'h3c639f2a),
	.w2(32'h3a4d3fd8),
	.w3(32'hba28d7cc),
	.w4(32'h3ba95491),
	.w5(32'h3b1f8853),
	.w6(32'h3bc4fe05),
	.w7(32'hbb433c8e),
	.w8(32'hbb2c4224),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d120b3a),
	.w1(32'hbc3766b3),
	.w2(32'hbc3dd461),
	.w3(32'h3d28c9eb),
	.w4(32'hbbc58a2d),
	.w5(32'hbc0ac155),
	.w6(32'h3cb34542),
	.w7(32'h3b68d418),
	.w8(32'h3c542cb9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfca35d),
	.w1(32'hbb3833f0),
	.w2(32'hbb21db74),
	.w3(32'h3c841057),
	.w4(32'hb9e2f261),
	.w5(32'hba29e506),
	.w6(32'h3b34de0a),
	.w7(32'hbbf518ae),
	.w8(32'hba15df0c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b013699),
	.w1(32'hbbf5982d),
	.w2(32'hbc28ffe0),
	.w3(32'hb9f6714d),
	.w4(32'hbb91f111),
	.w5(32'hbc1cc321),
	.w6(32'hbbf3c5b2),
	.w7(32'hbc0da9e7),
	.w8(32'hbb7b5dbf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2d60f),
	.w1(32'hbb9f74b6),
	.w2(32'hbc7ea2df),
	.w3(32'h3b99d2e5),
	.w4(32'h3b10ff9f),
	.w5(32'hbc064c45),
	.w6(32'h3c788298),
	.w7(32'h3bfba3a8),
	.w8(32'hbbbd7735),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2200e4),
	.w1(32'h3be3d518),
	.w2(32'hb9e79a47),
	.w3(32'hbad54c3e),
	.w4(32'h3c06ff7a),
	.w5(32'hba48d5bb),
	.w6(32'h3b69d62c),
	.w7(32'h3c0a0e61),
	.w8(32'h3bd17f4a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d8642),
	.w1(32'hbcfe6e28),
	.w2(32'hbda54b32),
	.w3(32'h3bf5f5da),
	.w4(32'hbd84a53c),
	.w5(32'hbd8939da),
	.w6(32'hbc583d42),
	.w7(32'h3cc7b42b),
	.w8(32'hbcb4db48),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e674b),
	.w1(32'h3bc8ad93),
	.w2(32'h3a8680cc),
	.w3(32'h3ba25deb),
	.w4(32'h3bf2b12a),
	.w5(32'h3a362783),
	.w6(32'h3c71a454),
	.w7(32'h3bca4f87),
	.w8(32'hbb2c07c3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c5ed),
	.w1(32'h3aab67a1),
	.w2(32'hbb41cc64),
	.w3(32'hbbcc23b5),
	.w4(32'h3a945fed),
	.w5(32'hba1e6875),
	.w6(32'hbaaf431b),
	.w7(32'hbb1b7c68),
	.w8(32'h39dea92b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b353415),
	.w1(32'h3a43f11f),
	.w2(32'hbb11fb7a),
	.w3(32'h3bc39114),
	.w4(32'h3b0f67f9),
	.w5(32'h399253c6),
	.w6(32'hbb5259da),
	.w7(32'hbc20abe7),
	.w8(32'hbc44b062),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44543f),
	.w1(32'h3c06edc6),
	.w2(32'h3c3a09f8),
	.w3(32'hbb0d18bd),
	.w4(32'h3c3caa5a),
	.w5(32'h3c3dde1c),
	.w6(32'h3bd75ff1),
	.w7(32'h3c4d8c94),
	.w8(32'h3b0f6b9e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28bd0d),
	.w1(32'hbbda96d1),
	.w2(32'hbc1fca6e),
	.w3(32'h3c350686),
	.w4(32'hbb9665b6),
	.w5(32'hbc56d832),
	.w6(32'hbc07b898),
	.w7(32'hbc50baf7),
	.w8(32'hbc62283c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc884764),
	.w1(32'hbb606f39),
	.w2(32'hbb9b57e1),
	.w3(32'hbc79445c),
	.w4(32'hbbd7a018),
	.w5(32'hbb796c83),
	.w6(32'hbb68fafe),
	.w7(32'hbbb056ed),
	.w8(32'hbbfab8d4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe84dc5),
	.w1(32'h3bde9256),
	.w2(32'h3bb82650),
	.w3(32'hbac04aa6),
	.w4(32'h3c1c7341),
	.w5(32'h3c2ad853),
	.w6(32'h3a0aa030),
	.w7(32'h3a290f7b),
	.w8(32'hbb4ef934),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe53df6),
	.w1(32'hbc2bcce8),
	.w2(32'hbc8098c6),
	.w3(32'hbbca1456),
	.w4(32'hbbf9cf7e),
	.w5(32'hbc6f61f9),
	.w6(32'hb9a800c7),
	.w7(32'hbbf582cd),
	.w8(32'hbc2abdaf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2c7c4),
	.w1(32'h3baeaea6),
	.w2(32'h3b832d00),
	.w3(32'hbbfdc361),
	.w4(32'h3c03bbbd),
	.w5(32'h3bbe5b4f),
	.w6(32'h3b3fa91f),
	.w7(32'h3b4af144),
	.w8(32'hbb0c852a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1fff2),
	.w1(32'h3c099ac0),
	.w2(32'hba7c1889),
	.w3(32'h3bd39e05),
	.w4(32'h3c030be3),
	.w5(32'hbab33f1e),
	.w6(32'h3b8d6d68),
	.w7(32'hb9cd9d0f),
	.w8(32'h3b3bc1c9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb00f3),
	.w1(32'hbbac3eb2),
	.w2(32'hbb1ff434),
	.w3(32'h3b1b9813),
	.w4(32'hbc23c00d),
	.w5(32'hbb056818),
	.w6(32'hbb136df1),
	.w7(32'hbbcba01e),
	.w8(32'hbb88e682),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb703c0f),
	.w1(32'h3b82a3db),
	.w2(32'hbbb1380a),
	.w3(32'hb94e0910),
	.w4(32'hba94a8ee),
	.w5(32'hbb3c6440),
	.w6(32'hbb2b4a8c),
	.w7(32'hbb28deaf),
	.w8(32'hbb936588),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb381a46),
	.w1(32'h3bce13e9),
	.w2(32'h3b33194b),
	.w3(32'hbc225954),
	.w4(32'h3c20d851),
	.w5(32'h3c04fae7),
	.w6(32'h3c3ee07c),
	.w7(32'h3ca02951),
	.w8(32'h3c1ba084),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c240e12),
	.w1(32'hbc96fc92),
	.w2(32'hbbbe143d),
	.w3(32'h3c0eebf3),
	.w4(32'hbc5ac08e),
	.w5(32'hbb08971d),
	.w6(32'hbc1bdd6c),
	.w7(32'hbbbb3df1),
	.w8(32'h3a9e422f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9c1e8),
	.w1(32'h3b69efed),
	.w2(32'h3c08f284),
	.w3(32'h3bec483d),
	.w4(32'h3b79c33e),
	.w5(32'h3bde32fa),
	.w6(32'h3a087101),
	.w7(32'h3b97cca1),
	.w8(32'h3b31141d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7f9c7),
	.w1(32'hbb60aa17),
	.w2(32'hbc8c8f81),
	.w3(32'hbabf1b41),
	.w4(32'hbbc56183),
	.w5(32'hbc94722c),
	.w6(32'h38d8cbd6),
	.w7(32'hbc06b7b3),
	.w8(32'hbc15fba5),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd233f),
	.w1(32'hbb92b487),
	.w2(32'hbc559146),
	.w3(32'hbc11dcff),
	.w4(32'hbb8a2d6a),
	.w5(32'hbbee93d7),
	.w6(32'h3bd4ec65),
	.w7(32'hbb3ddb9f),
	.w8(32'hb9cae23c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d5e6a),
	.w1(32'hbc24352a),
	.w2(32'hbb33bf41),
	.w3(32'hbb2a3f02),
	.w4(32'hbbbc2009),
	.w5(32'h3ae5cb4e),
	.w6(32'hbbac606c),
	.w7(32'h39b8c4fe),
	.w8(32'h39180353),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9f6c),
	.w1(32'h3afabf4a),
	.w2(32'hbb97016e),
	.w3(32'h3b0bb0bc),
	.w4(32'hb95732fe),
	.w5(32'hbb960305),
	.w6(32'hb9aa4041),
	.w7(32'hbbdab609),
	.w8(32'hbc0e1470),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9cc01),
	.w1(32'hba3b0bed),
	.w2(32'hbc4a0ea6),
	.w3(32'hba96c165),
	.w4(32'hbc108e1d),
	.w5(32'hbc00144f),
	.w6(32'h3c3807bc),
	.w7(32'h3bd1aad3),
	.w8(32'h3acbf466),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b795268),
	.w1(32'h3b2a5f5f),
	.w2(32'hbb98e95e),
	.w3(32'hbbe08ac4),
	.w4(32'hbba9b9e4),
	.w5(32'hbb6ac674),
	.w6(32'hbb072995),
	.w7(32'hbb1d5f25),
	.w8(32'hbad226bd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e796a5),
	.w1(32'hbc1bb493),
	.w2(32'h3b91d63d),
	.w3(32'hbb303c98),
	.w4(32'hbc35c654),
	.w5(32'h3b68f5e3),
	.w6(32'hbb86fa8b),
	.w7(32'h3c7d8bb6),
	.w8(32'h3bc870bf),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb68fc7),
	.w1(32'h3cb8e2d0),
	.w2(32'h3c940335),
	.w3(32'h3c91cdb5),
	.w4(32'h3c831e23),
	.w5(32'h3c336230),
	.w6(32'h3c0d9ab4),
	.w7(32'h3c5d51f0),
	.w8(32'h3c3ffb01),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c88f3),
	.w1(32'hbcae903c),
	.w2(32'hbbe90f5f),
	.w3(32'hbbb457be),
	.w4(32'hbd171583),
	.w5(32'hbc8ea0a0),
	.w6(32'h3c1f36e0),
	.w7(32'h3b9db2ff),
	.w8(32'h3aca21fc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf263f3),
	.w1(32'hba6b2d02),
	.w2(32'hbb247364),
	.w3(32'h3bf20f7d),
	.w4(32'hbb7cea5c),
	.w5(32'hbb9e9ee1),
	.w6(32'h3bd256d0),
	.w7(32'hbabb2b38),
	.w8(32'h3a852375),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb542f64),
	.w1(32'hbb8f9814),
	.w2(32'hbc66a4c7),
	.w3(32'h3b361ef5),
	.w4(32'h3baf6556),
	.w5(32'hbaa0c616),
	.w6(32'hba35a617),
	.w7(32'hbc02fcf1),
	.w8(32'hbb9009ad),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9a2d6),
	.w1(32'h3bcdfd71),
	.w2(32'hbba3e266),
	.w3(32'hbbbcb7c2),
	.w4(32'hba1e3fc3),
	.w5(32'hbb8a301a),
	.w6(32'h39a97f81),
	.w7(32'hbb9ceb5d),
	.w8(32'hbc3942ff),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb481b6d),
	.w1(32'hbbded15a),
	.w2(32'hbcdbbe20),
	.w3(32'h3c29eaf0),
	.w4(32'h3b854173),
	.w5(32'hbc03d757),
	.w6(32'hbbafbafb),
	.w7(32'hbc2bbe3b),
	.w8(32'hbc0b0d17),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3887ed),
	.w1(32'hbc435868),
	.w2(32'hbbf7bd44),
	.w3(32'hbb85402a),
	.w4(32'hbb548286),
	.w5(32'hbbcf6114),
	.w6(32'hbbc892f2),
	.w7(32'hbc5aa3fc),
	.w8(32'hbc2708e4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99997b),
	.w1(32'hbbe24eb4),
	.w2(32'h3a833498),
	.w3(32'hbc99aced),
	.w4(32'hbc133f9a),
	.w5(32'hbb825cf3),
	.w6(32'hb9ec8073),
	.w7(32'hbb85d493),
	.w8(32'hbbf6fa8c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd82aa),
	.w1(32'hbb1feda2),
	.w2(32'hbbc8ee25),
	.w3(32'hbbbf4ebc),
	.w4(32'hbbc57352),
	.w5(32'hbbebb5c4),
	.w6(32'hbacfdbbb),
	.w7(32'hbbc9e7ad),
	.w8(32'hbbda0163),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ca1ea),
	.w1(32'h3a49a7cf),
	.w2(32'h3b6f5265),
	.w3(32'hbb648268),
	.w4(32'h3b68ccd1),
	.w5(32'h3bdc9ab1),
	.w6(32'hbab4e8e8),
	.w7(32'hb9e3dff1),
	.w8(32'h3ac8f09c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea1219),
	.w1(32'hbb90d4e6),
	.w2(32'hbbf28dfd),
	.w3(32'h3b7bc120),
	.w4(32'hbbd1657c),
	.w5(32'hbc34b0d3),
	.w6(32'h3b34ee05),
	.w7(32'h3a961ca3),
	.w8(32'h3bbd8b54),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73f5c5),
	.w1(32'h3b841783),
	.w2(32'hbb0f8acd),
	.w3(32'hbb6bdc00),
	.w4(32'h3bf0011e),
	.w5(32'hbb1b8238),
	.w6(32'hbacf6220),
	.w7(32'hbae5edb7),
	.w8(32'h3b1739f0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ebb6e),
	.w1(32'hbb3a7999),
	.w2(32'hbb1cacee),
	.w3(32'h3bb2102b),
	.w4(32'h3bd40f90),
	.w5(32'h3b9f49e4),
	.w6(32'h3c3ce575),
	.w7(32'h3c83eb71),
	.w8(32'h3bfff1b8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf5dfa),
	.w1(32'hbaa602e0),
	.w2(32'hba1255c0),
	.w3(32'h3bc63030),
	.w4(32'hbb8c43a4),
	.w5(32'hbaf5d9be),
	.w6(32'hbb0e92ee),
	.w7(32'hbb15cbbb),
	.w8(32'hbad7c599),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b330d19),
	.w1(32'h3b87e08b),
	.w2(32'h3aac79da),
	.w3(32'h3aa8c6da),
	.w4(32'h3b35c415),
	.w5(32'hb9ccb06b),
	.w6(32'h3adf8700),
	.w7(32'hbac6855d),
	.w8(32'hbb012934),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5e930),
	.w1(32'hbba76658),
	.w2(32'hbba82a90),
	.w3(32'h3aa66c55),
	.w4(32'hbbac6d69),
	.w5(32'hbc0ee437),
	.w6(32'h3b339b74),
	.w7(32'hbbe0f0bb),
	.w8(32'hbc2ad97e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c91ef9),
	.w1(32'h3c29391b),
	.w2(32'h3c06c87c),
	.w3(32'h3ae1a7c8),
	.w4(32'h3be5c912),
	.w5(32'hbac0d40a),
	.w6(32'h3c086bbe),
	.w7(32'h3c2aef17),
	.w8(32'h3ba37a53),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71b543),
	.w1(32'hbb802f33),
	.w2(32'hbbd10392),
	.w3(32'h3b681ae8),
	.w4(32'hbb47a488),
	.w5(32'hbb7ab110),
	.w6(32'hbc02ff19),
	.w7(32'hbb5e97ea),
	.w8(32'h3ab7e72a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6cc1f),
	.w1(32'h3bd71eb6),
	.w2(32'h39ee18ec),
	.w3(32'h3ae56c41),
	.w4(32'h3b92053b),
	.w5(32'h3b8f4a0a),
	.w6(32'hbaf671f4),
	.w7(32'h3aaf4cc6),
	.w8(32'h3c12152f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc120db),
	.w1(32'h3bc76d9b),
	.w2(32'hbc2e7590),
	.w3(32'h3c539eaa),
	.w4(32'hbc91af5a),
	.w5(32'hbc9ffdfc),
	.w6(32'hbbaaa82e),
	.w7(32'h3b5380fb),
	.w8(32'h3a12dfa5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58e212),
	.w1(32'h3be3e8e6),
	.w2(32'h3bd0c32f),
	.w3(32'h3b28624f),
	.w4(32'h3b6704fb),
	.w5(32'h3b6387ed),
	.w6(32'hba02fdf8),
	.w7(32'hba81be9e),
	.w8(32'h3b8d73a4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c379e78),
	.w1(32'hbc20a6cf),
	.w2(32'hbc589f70),
	.w3(32'h3c364e8c),
	.w4(32'hbade0507),
	.w5(32'hbbb1749a),
	.w6(32'hbb55d97e),
	.w7(32'hbc19ac2f),
	.w8(32'hbbf0947d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d0a3),
	.w1(32'h3b41de24),
	.w2(32'h3a7c465c),
	.w3(32'h3a4dc37a),
	.w4(32'h3b375421),
	.w5(32'h3a72f04d),
	.w6(32'h3bccca06),
	.w7(32'h3ad4e3b4),
	.w8(32'hbb094a20),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e54f09),
	.w1(32'h3b6c8e90),
	.w2(32'hbaa849b9),
	.w3(32'h3c1ca100),
	.w4(32'h3c068c0a),
	.w5(32'h3ba695b5),
	.w6(32'h3b2973fa),
	.w7(32'hbb019427),
	.w8(32'hbbaba6e6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a15b),
	.w1(32'hbc389804),
	.w2(32'hbb14ec7f),
	.w3(32'hbb53a4e7),
	.w4(32'hbb983f2f),
	.w5(32'hbadac76a),
	.w6(32'hbc1e9e4b),
	.w7(32'hbb680891),
	.w8(32'hbad4798b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc31a7),
	.w1(32'h3c3cdc33),
	.w2(32'h3c795161),
	.w3(32'h3bfb5ed9),
	.w4(32'h3c4a3214),
	.w5(32'h3c551ebb),
	.w6(32'h3c358811),
	.w7(32'h3c4992c7),
	.w8(32'h3c6dd84d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce69bda),
	.w1(32'h3a86ee66),
	.w2(32'h3b819cc4),
	.w3(32'h3caed022),
	.w4(32'hba64c22d),
	.w5(32'h3a1c0159),
	.w6(32'h3acb8abe),
	.w7(32'h3b4ba498),
	.w8(32'h3aaac654),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baeaafc),
	.w1(32'hbc051fee),
	.w2(32'hba3f39da),
	.w3(32'h3a49887b),
	.w4(32'hbc1254a1),
	.w5(32'hbb04723e),
	.w6(32'h3b14b777),
	.w7(32'h3c20c463),
	.w8(32'h3bfc1ffa),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25e124),
	.w1(32'hbc7c2325),
	.w2(32'hbc8fef90),
	.w3(32'hba6b83e4),
	.w4(32'hbc505a0f),
	.w5(32'hbbd7f516),
	.w6(32'hbbf363cc),
	.w7(32'hbc6e488b),
	.w8(32'hbbf57cea),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd368),
	.w1(32'hbade55e7),
	.w2(32'hbc209a09),
	.w3(32'h3920075b),
	.w4(32'hbab2f598),
	.w5(32'hbb881291),
	.w6(32'hbbc702b6),
	.w7(32'hbad0dd58),
	.w8(32'hbab1ac63),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ec8cb),
	.w1(32'hbb6b1944),
	.w2(32'hbc180991),
	.w3(32'hbbe6cccd),
	.w4(32'hbb7e6d1d),
	.w5(32'hbc1ac404),
	.w6(32'h3ba64341),
	.w7(32'hbb668f0a),
	.w8(32'h3bfd96b5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2ebba),
	.w1(32'hbad85087),
	.w2(32'h3badf31f),
	.w3(32'hbb8c0820),
	.w4(32'h3b5b9c84),
	.w5(32'h3b0ab81e),
	.w6(32'h398be679),
	.w7(32'hbbd1a01c),
	.w8(32'hbae4e3a2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e92e9),
	.w1(32'hbaf66a80),
	.w2(32'hbbb3ee60),
	.w3(32'h3c02844f),
	.w4(32'hbbc4b30a),
	.w5(32'hbb236635),
	.w6(32'h3bf217f7),
	.w7(32'h3c103318),
	.w8(32'h3c5a590a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ea3a4),
	.w1(32'hbc2af60b),
	.w2(32'hbc8e0733),
	.w3(32'h3b5a8627),
	.w4(32'h3a125b50),
	.w5(32'hbbebd9ca),
	.w6(32'h39d38e5e),
	.w7(32'h3ba90279),
	.w8(32'hbb1fb4fb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1809c),
	.w1(32'hbc69a2fe),
	.w2(32'hbcdd8815),
	.w3(32'hb996e7d1),
	.w4(32'hbc3b2883),
	.w5(32'hbc73a4ee),
	.w6(32'h3c4d6847),
	.w7(32'h3c316d6b),
	.w8(32'h3c0d40f1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8300a9),
	.w1(32'hbb0258e8),
	.w2(32'h3b7dcd51),
	.w3(32'h3c9ef700),
	.w4(32'h3bb8414d),
	.w5(32'hba3ccac4),
	.w6(32'h3c719150),
	.w7(32'h3b993859),
	.w8(32'hbb090a36),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb057298),
	.w1(32'hbaa03689),
	.w2(32'h3b6b7988),
	.w3(32'hbb0adfd3),
	.w4(32'hbb7e636d),
	.w5(32'h3b5619f8),
	.w6(32'hbb418b35),
	.w7(32'hbb46ac62),
	.w8(32'hbaca16c3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb02bc2),
	.w1(32'h3ab4637c),
	.w2(32'h391e9a0a),
	.w3(32'h3b92d103),
	.w4(32'h3c0faa2f),
	.w5(32'h3b853f6d),
	.w6(32'hbaa24b31),
	.w7(32'h3a8a26a4),
	.w8(32'hbaf83833),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62a8b2),
	.w1(32'hba7199e7),
	.w2(32'hbab3856a),
	.w3(32'h3b394dc3),
	.w4(32'h3a30432c),
	.w5(32'h3bde629f),
	.w6(32'hba3ea620),
	.w7(32'hbba4da0e),
	.w8(32'hbbac877f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f3db9),
	.w1(32'h3af9f698),
	.w2(32'hbb49a78f),
	.w3(32'h3bec84f7),
	.w4(32'hba82d4e0),
	.w5(32'h3ac8fdaa),
	.w6(32'h3bf73e5e),
	.w7(32'h3bc73058),
	.w8(32'h3b069cdf),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb237324),
	.w1(32'hbbc9b45e),
	.w2(32'hbbb8c483),
	.w3(32'h3b8936d0),
	.w4(32'h3a8ef5b9),
	.w5(32'h3aee47f5),
	.w6(32'hbb0a4ccf),
	.w7(32'h3ab84e5a),
	.w8(32'hbbf232f0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afee836),
	.w1(32'h39b3bfe7),
	.w2(32'hbb855794),
	.w3(32'h3af3823f),
	.w4(32'h3a22bf99),
	.w5(32'hbbeb130d),
	.w6(32'hbaab03b7),
	.w7(32'hbb55e9f9),
	.w8(32'hbc217521),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6611b9),
	.w1(32'h3b0e99cc),
	.w2(32'h3bb80f20),
	.w3(32'hbc38f13e),
	.w4(32'hba92e665),
	.w5(32'h3ba4aef5),
	.w6(32'hbb26c5a3),
	.w7(32'hbab49f81),
	.w8(32'hba87e9e3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6b919),
	.w1(32'h3ab95482),
	.w2(32'hbb0ef418),
	.w3(32'h3b97e85e),
	.w4(32'h3b2a7027),
	.w5(32'hbaa6cfe4),
	.w6(32'h3bb91978),
	.w7(32'h3b1048f5),
	.w8(32'hbb024172),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8472dc),
	.w1(32'h3cbbd091),
	.w2(32'h3d0bafd3),
	.w3(32'h3b196405),
	.w4(32'h3c92268e),
	.w5(32'h3cbdec75),
	.w6(32'h3c43ebb7),
	.w7(32'h3c943d7d),
	.w8(32'h3bcd3823),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc20fd9),
	.w1(32'h3ad02a24),
	.w2(32'hbb84781e),
	.w3(32'h3c7d08db),
	.w4(32'h3850508f),
	.w5(32'hbbace8f0),
	.w6(32'h3c19e9ca),
	.w7(32'h3babc713),
	.w8(32'hbbedbfc2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b484f7c),
	.w1(32'hbb6d8f2c),
	.w2(32'hbba2ba62),
	.w3(32'h3986025d),
	.w4(32'h3addb538),
	.w5(32'h3b8a39e2),
	.w6(32'h3c8d783d),
	.w7(32'h3b5dbb80),
	.w8(32'hbb8f2453),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb578dc6),
	.w1(32'h3a0c07c9),
	.w2(32'hbc56d8e1),
	.w3(32'hbc03b8d0),
	.w4(32'hbad0a9c2),
	.w5(32'hbc57fd76),
	.w6(32'hbbc1f2fa),
	.w7(32'hbc6ce7a5),
	.w8(32'hbc3b8f38),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c5e0d),
	.w1(32'hbbaafb2c),
	.w2(32'hbc2714ec),
	.w3(32'hbb83a62d),
	.w4(32'hbb89b398),
	.w5(32'hbbd039fe),
	.w6(32'hbb874c71),
	.w7(32'hbb9e3eed),
	.w8(32'hbbc1b6df),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63e9a4),
	.w1(32'hbb3abf54),
	.w2(32'h3a07a8cd),
	.w3(32'hbb8f6764),
	.w4(32'hbc0bb08d),
	.w5(32'hbc08b4e8),
	.w6(32'hbba33d0d),
	.w7(32'h3b7d9929),
	.w8(32'h3b7906fd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac37a3),
	.w1(32'hbb9ae4e3),
	.w2(32'hbc07f11c),
	.w3(32'hbbf8f6bd),
	.w4(32'hbbbb8d8f),
	.w5(32'hbbeb69da),
	.w6(32'hbc0103d4),
	.w7(32'hbc2b0fd3),
	.w8(32'h3b8bb038),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4ef6c),
	.w1(32'h3b06ce69),
	.w2(32'hb9bdf43c),
	.w3(32'h3bbc061b),
	.w4(32'h3bee9be5),
	.w5(32'h3b647d67),
	.w6(32'hbb5512f3),
	.w7(32'hbaa0d6cb),
	.w8(32'h399a3c9a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d65be),
	.w1(32'h3b9f1209),
	.w2(32'h3c0756cb),
	.w3(32'h3b1ebdc7),
	.w4(32'h3a3bff1f),
	.w5(32'hba69a4b7),
	.w6(32'h3b14d581),
	.w7(32'hbb3e9f93),
	.w8(32'h3ba27230),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa0e0c),
	.w1(32'hbbeb9f2b),
	.w2(32'h3b578de8),
	.w3(32'hbbd124ea),
	.w4(32'hbc0141d9),
	.w5(32'h3ba9aae4),
	.w6(32'hbc092c67),
	.w7(32'hbc16b203),
	.w8(32'hbbf08a47),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a044b),
	.w1(32'hbbd4b30a),
	.w2(32'hbb22a186),
	.w3(32'h3b51cb05),
	.w4(32'hbbd4494d),
	.w5(32'hbb6a2c2e),
	.w6(32'hbc2ad5a0),
	.w7(32'hbbd9a472),
	.w8(32'hbb0340fa),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22f5bf),
	.w1(32'hbbc0e570),
	.w2(32'hbc1422ca),
	.w3(32'hbbabfa18),
	.w4(32'hbc45ac91),
	.w5(32'hbc3d8630),
	.w6(32'hb92cad0d),
	.w7(32'h3a7c5bed),
	.w8(32'hbb384d1f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2ed6f),
	.w1(32'hbbc390cf),
	.w2(32'hbb919290),
	.w3(32'hba3af641),
	.w4(32'hbbc6be47),
	.w5(32'hb9f8586c),
	.w6(32'hbbcada2a),
	.w7(32'hbbee7ee4),
	.w8(32'hbc454681),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0517ab),
	.w1(32'h3a4bffa1),
	.w2(32'h3b9fb4bb),
	.w3(32'h3afcc0c6),
	.w4(32'h3b245833),
	.w5(32'h3a1ec15e),
	.w6(32'hbb2af47e),
	.w7(32'h3a99757b),
	.w8(32'h39d61164),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1791f),
	.w1(32'h3b8ace58),
	.w2(32'hba57e9bf),
	.w3(32'hbb29d4da),
	.w4(32'h3b4212d6),
	.w5(32'hbb477278),
	.w6(32'hbb9d6190),
	.w7(32'hbb87df6f),
	.w8(32'hbc232c7f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a670708),
	.w1(32'h3a9d60ad),
	.w2(32'h38950dfb),
	.w3(32'h3acf0fd9),
	.w4(32'h3b80ce91),
	.w5(32'hba020026),
	.w6(32'h3bc06cf3),
	.w7(32'hba694182),
	.w8(32'hbb1429e4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6af24),
	.w1(32'hbb2b4eff),
	.w2(32'hbba5ad7e),
	.w3(32'hb9cbdfcc),
	.w4(32'h3be3870f),
	.w5(32'hbb41785f),
	.w6(32'hbacb68f9),
	.w7(32'h3b94eb67),
	.w8(32'h3b31cb98),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6dd9),
	.w1(32'hbb742977),
	.w2(32'hbaee4789),
	.w3(32'hbba69b7a),
	.w4(32'hbaf78e39),
	.w5(32'hb956f198),
	.w6(32'h3a9cc8cc),
	.w7(32'h3b60f9f3),
	.w8(32'hbb5770d6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f1b68),
	.w1(32'h3b1743c9),
	.w2(32'h3b7f8823),
	.w3(32'hba19444b),
	.w4(32'h3a2c1759),
	.w5(32'h3aa16573),
	.w6(32'h3b40a7b2),
	.w7(32'hbc0de2d3),
	.w8(32'hbba41c68),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaec7c1),
	.w1(32'hbb81a13b),
	.w2(32'hbc20880d),
	.w3(32'hbb83081d),
	.w4(32'hbaf98ba5),
	.w5(32'hbb62731f),
	.w6(32'hba0f7497),
	.w7(32'hbbe9f255),
	.w8(32'hbbc5e93d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89b08d),
	.w1(32'hbbc1f652),
	.w2(32'hbb4fd2c5),
	.w3(32'h3ae9b98c),
	.w4(32'hbab53f75),
	.w5(32'h3b748cc5),
	.w6(32'hbb97c6d8),
	.w7(32'hbbd43e23),
	.w8(32'hbb918790),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5eca0),
	.w1(32'h3bb238a6),
	.w2(32'h3b733baa),
	.w3(32'h3c6f67a3),
	.w4(32'h3bbbfc89),
	.w5(32'h3b7be50c),
	.w6(32'h3bce9b5e),
	.w7(32'h3b8659ee),
	.w8(32'h3b1bb263),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae42641),
	.w1(32'hb82f1bb9),
	.w2(32'h3a18d72f),
	.w3(32'h3ab6298e),
	.w4(32'hbb20b01c),
	.w5(32'hbbe37308),
	.w6(32'hbb8b0154),
	.w7(32'hba787e4f),
	.w8(32'h3b9e8e3e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11f2ea),
	.w1(32'h3ae4e93d),
	.w2(32'hbb726016),
	.w3(32'h3ae0d84a),
	.w4(32'hbb84a1c5),
	.w5(32'hbc1d13c5),
	.w6(32'hbb0cef93),
	.w7(32'h3a93c169),
	.w8(32'hbb718734),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8caa30),
	.w1(32'hbb1869de),
	.w2(32'hbb103303),
	.w3(32'hbabf07b1),
	.w4(32'h3bbfe937),
	.w5(32'hbb35413a),
	.w6(32'hbab36e3a),
	.w7(32'hbbca2acc),
	.w8(32'hbbb22f98),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9776e),
	.w1(32'hbbdb0ca0),
	.w2(32'hbbbdd36e),
	.w3(32'h3a5151d4),
	.w4(32'hbb4f0d2f),
	.w5(32'hbb6f021f),
	.w6(32'hbb824eff),
	.w7(32'hbb814ec8),
	.w8(32'hb9bc706a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92b2a4),
	.w1(32'hbb3df1d5),
	.w2(32'hba1e6b52),
	.w3(32'h3bea1ee2),
	.w4(32'h3b866fd6),
	.w5(32'h3b059aad),
	.w6(32'hbbb9dde3),
	.w7(32'hbb92780c),
	.w8(32'h3a9f34bf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a2657),
	.w1(32'hba026cdc),
	.w2(32'h3b2e1ec8),
	.w3(32'hbb6b887a),
	.w4(32'h3b9277c7),
	.w5(32'h3c1241a4),
	.w6(32'h3bb4d1ce),
	.w7(32'h3bea8fb9),
	.w8(32'h3ab94549),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ea66c),
	.w1(32'hb9979f71),
	.w2(32'h3a43aa43),
	.w3(32'h3b4f25dd),
	.w4(32'h3aaa8195),
	.w5(32'h3ae3b729),
	.w6(32'hbaa7cdbe),
	.w7(32'hbafb444b),
	.w8(32'hbb92b1c2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9984b8),
	.w1(32'h3c0edaf0),
	.w2(32'h3b38ffd1),
	.w3(32'hba976a62),
	.w4(32'h3b8f87be),
	.w5(32'hba87eeca),
	.w6(32'hb9c05755),
	.w7(32'hb9b670c2),
	.w8(32'hbb8e069e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c482042),
	.w1(32'h3bb7cdd3),
	.w2(32'hba8b23b5),
	.w3(32'h3bfe1f45),
	.w4(32'h3b0ced37),
	.w5(32'hbb8a506a),
	.w6(32'h3bd46e8e),
	.w7(32'h3b5ae455),
	.w8(32'h3b2c66ab),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385ef42a),
	.w1(32'h3b7d8055),
	.w2(32'h3b1d4d84),
	.w3(32'hbb85109e),
	.w4(32'h3a6fa649),
	.w5(32'hb8e353d1),
	.w6(32'h3ac383bc),
	.w7(32'h3a07760e),
	.w8(32'hba807318),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72a602),
	.w1(32'hba9aa815),
	.w2(32'hbaee489b),
	.w3(32'h3bc6a764),
	.w4(32'h3b31d924),
	.w5(32'h39be85c1),
	.w6(32'hba773179),
	.w7(32'hba5a05f8),
	.w8(32'h3a281657),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fc05b),
	.w1(32'hbb96924d),
	.w2(32'h3c054e63),
	.w3(32'hbb2dc58c),
	.w4(32'hbc0714cd),
	.w5(32'h3b7f91b7),
	.w6(32'hbbae69bb),
	.w7(32'h3b9799fc),
	.w8(32'h3bc23a4f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule