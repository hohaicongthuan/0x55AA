module layer_10_featuremap_1(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d3500),
	.w1(32'hbb995ade),
	.w2(32'hbadb9dbe),
	.w3(32'h3c8215cf),
	.w4(32'hbc80f62c),
	.w5(32'hbb2ab9bd),
	.w6(32'h3aa2150c),
	.w7(32'hbc5089db),
	.w8(32'h3b1ee6df),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b3e8c),
	.w1(32'hbaaca337),
	.w2(32'h3a8fa037),
	.w3(32'h3c277e52),
	.w4(32'h3be66ccb),
	.w5(32'hba75b36f),
	.w6(32'h3bacfc7d),
	.w7(32'h3bb9756d),
	.w8(32'h3bce6903),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddbc10),
	.w1(32'h399512c4),
	.w2(32'h3a0f2579),
	.w3(32'hbbda4892),
	.w4(32'hbc03bb77),
	.w5(32'hbb873eda),
	.w6(32'hbc2a499b),
	.w7(32'hbbe687b1),
	.w8(32'h3b332f17),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0da27d),
	.w1(32'hbbb88686),
	.w2(32'hbafe2b10),
	.w3(32'h3b822bbd),
	.w4(32'hbb2a4ba2),
	.w5(32'hbb9279c5),
	.w6(32'hbb8c1911),
	.w7(32'hbbdeba7c),
	.w8(32'hbc1b49b7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aa909),
	.w1(32'hbc6e934d),
	.w2(32'hbc3499db),
	.w3(32'hbc8251bc),
	.w4(32'h3a94d43c),
	.w5(32'hbc42f226),
	.w6(32'hbbc77798),
	.w7(32'h3c330c36),
	.w8(32'hbbf8b3ed),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f1223),
	.w1(32'hbbfb99be),
	.w2(32'h3bb556c7),
	.w3(32'hbb0d5e64),
	.w4(32'h3bbb0299),
	.w5(32'h3bf63b87),
	.w6(32'hbb3950e8),
	.w7(32'hba82e57c),
	.w8(32'h3b871635),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09a03f),
	.w1(32'h3ad043a6),
	.w2(32'h3bd3df12),
	.w3(32'hba7c1309),
	.w4(32'hbb3265e1),
	.w5(32'h3b2355f4),
	.w6(32'hbb01aaa4),
	.w7(32'hbb77799a),
	.w8(32'hbb4c41cf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ac68d),
	.w1(32'hbc6a83c5),
	.w2(32'h3ba9a1db),
	.w3(32'hbaf3d90b),
	.w4(32'hbc91be75),
	.w5(32'h3bba9a78),
	.w6(32'hbc615b8a),
	.w7(32'hbc5ab122),
	.w8(32'h3912f4e5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b117194),
	.w1(32'h3a271f87),
	.w2(32'hba303708),
	.w3(32'hbb50ebb9),
	.w4(32'hbb5364e1),
	.w5(32'hbaaad1e3),
	.w6(32'hbc0db153),
	.w7(32'h3a9e8974),
	.w8(32'hbc29cc65),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e1f60),
	.w1(32'h3b1c6eac),
	.w2(32'hbbbd5e11),
	.w3(32'hbc05628e),
	.w4(32'h3b376c93),
	.w5(32'hbb9950be),
	.w6(32'hbc28106b),
	.w7(32'h3b9f95b9),
	.w8(32'hbb82c544),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af6e3f),
	.w1(32'hba1649df),
	.w2(32'hbba61e66),
	.w3(32'h3b8ba45f),
	.w4(32'hb9d40e6a),
	.w5(32'hbbb79349),
	.w6(32'h3aa4ca8b),
	.w7(32'hbb5a71d0),
	.w8(32'hbc17929c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8f719),
	.w1(32'h3bfff704),
	.w2(32'hbb1c3626),
	.w3(32'h3bdb4676),
	.w4(32'h3be725d7),
	.w5(32'hbb75b06a),
	.w6(32'hbb2d7ce7),
	.w7(32'h393de699),
	.w8(32'hbb397c09),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ec842),
	.w1(32'hbb2ecfe2),
	.w2(32'h3ba8822d),
	.w3(32'hbb0c53d8),
	.w4(32'hbba8f6e0),
	.w5(32'h3b0afe88),
	.w6(32'hbb2b98c9),
	.w7(32'hbb9f78a5),
	.w8(32'hbb07729f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc440884),
	.w1(32'h3a3734a1),
	.w2(32'hbb757e86),
	.w3(32'hbbe70198),
	.w4(32'hbba869b9),
	.w5(32'hbbf102eb),
	.w6(32'hbb806c11),
	.w7(32'h3b42ac65),
	.w8(32'hbca50f68),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb5c36),
	.w1(32'h3b8c0a45),
	.w2(32'hbc4f3ccb),
	.w3(32'h3b8d9056),
	.w4(32'hbacdd6d4),
	.w5(32'hbc7a538f),
	.w6(32'hba6c80f6),
	.w7(32'h3b17463b),
	.w8(32'hbb68e4d4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b2488),
	.w1(32'h3b17fe11),
	.w2(32'hb9167bda),
	.w3(32'hbbee1291),
	.w4(32'h3b476a1e),
	.w5(32'h3b0832b9),
	.w6(32'h3c01c97c),
	.w7(32'h3c6533e1),
	.w8(32'h3b49b1df),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb319b5),
	.w1(32'hbb49f76d),
	.w2(32'hbc58f204),
	.w3(32'h3c093d8e),
	.w4(32'hbb8cabfd),
	.w5(32'hbc312be6),
	.w6(32'h3b6b4b5c),
	.w7(32'hbbfe287e),
	.w8(32'hbc60ee81),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcbc06),
	.w1(32'h3c932901),
	.w2(32'hba3ae702),
	.w3(32'h3c310fdb),
	.w4(32'h3d101e26),
	.w5(32'hbb20435c),
	.w6(32'h3baea7fa),
	.w7(32'h3d1620c8),
	.w8(32'hbac30047),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf398a2),
	.w1(32'hbb044d34),
	.w2(32'h3a0b7449),
	.w3(32'hba55bc82),
	.w4(32'h3b03eaec),
	.w5(32'hbb2371f4),
	.w6(32'hbb284230),
	.w7(32'hbb25ad7a),
	.w8(32'hbb11c13a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cf853),
	.w1(32'hbc27d9b3),
	.w2(32'hbc9f23c4),
	.w3(32'hbba8d521),
	.w4(32'hbc10d13b),
	.w5(32'hbcb0bb7f),
	.w6(32'hbb2a46eb),
	.w7(32'hbc1de762),
	.w8(32'hbc208f4d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe59a96),
	.w1(32'h3b3882fa),
	.w2(32'hbb06c6f6),
	.w3(32'hb88cfa62),
	.w4(32'h3c46999b),
	.w5(32'h3b88fba5),
	.w6(32'h3bd8c772),
	.w7(32'h3c3562b4),
	.w8(32'hb9504260),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b604d86),
	.w1(32'h3bb0fd7e),
	.w2(32'hbb044c55),
	.w3(32'h3c18c671),
	.w4(32'h3c1a5e59),
	.w5(32'hba082140),
	.w6(32'h3bdd852d),
	.w7(32'h3b8b0bf0),
	.w8(32'hbaef9e54),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac03a6c),
	.w1(32'h39ca9fce),
	.w2(32'hbad3fe47),
	.w3(32'hba77c508),
	.w4(32'hbb8a9e88),
	.w5(32'hbaf44c35),
	.w6(32'hbc308678),
	.w7(32'hbc2dbd41),
	.w8(32'hbb7d631a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2c643),
	.w1(32'hbb4a0207),
	.w2(32'h3b581e58),
	.w3(32'h3ba171fb),
	.w4(32'hbbab6d4f),
	.w5(32'hbc12aa95),
	.w6(32'h39db3d8b),
	.w7(32'hbc02685c),
	.w8(32'hbb977460),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f4f50),
	.w1(32'hbaafa1d0),
	.w2(32'hbb02caea),
	.w3(32'hbae76cc4),
	.w4(32'hbba3f19f),
	.w5(32'hbbff61a3),
	.w6(32'hbc0dcc16),
	.w7(32'h3afd61ac),
	.w8(32'h3bb6f2c4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b3b55),
	.w1(32'hb9a49e04),
	.w2(32'hbb0cf966),
	.w3(32'h3c15c1cb),
	.w4(32'h3c158512),
	.w5(32'hbc34eac3),
	.w6(32'h3c514f5a),
	.w7(32'h3ba66559),
	.w8(32'hbc1bb339),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc254ba9),
	.w1(32'hbbac9617),
	.w2(32'h3bd94291),
	.w3(32'hbbfde463),
	.w4(32'h393841bf),
	.w5(32'h3b4cb213),
	.w6(32'hbca3c3dc),
	.w7(32'h3b98c0e9),
	.w8(32'h3b799473),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b538aaf),
	.w1(32'h3b216849),
	.w2(32'hbb85811e),
	.w3(32'hbbe7e6a6),
	.w4(32'hbb21f45b),
	.w5(32'hbbc41037),
	.w6(32'hbb3e0b93),
	.w7(32'hba4aa5eb),
	.w8(32'hbb35f793),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc57ee1),
	.w1(32'h3c40c1ff),
	.w2(32'hbb0d1ab7),
	.w3(32'hba7e057e),
	.w4(32'h3c5b9391),
	.w5(32'h3c073b86),
	.w6(32'h39e3ca42),
	.w7(32'h3c75a85d),
	.w8(32'h3bac3e2c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d452f),
	.w1(32'hbbb6941a),
	.w2(32'hbcbafef5),
	.w3(32'hb9537be6),
	.w4(32'hbb14bb82),
	.w5(32'hbc990049),
	.w6(32'h3b40073d),
	.w7(32'h3b04560b),
	.w8(32'hbcc8a56d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b2e7c),
	.w1(32'hbc6faa99),
	.w2(32'hbb952a37),
	.w3(32'hbb80ac9f),
	.w4(32'hbbe3e723),
	.w5(32'hb946fafe),
	.w6(32'hbc73bd4a),
	.w7(32'hbc93caa1),
	.w8(32'h3a20a4a5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3135bc),
	.w1(32'hb8313d40),
	.w2(32'hbafa933a),
	.w3(32'h3bd8ae15),
	.w4(32'h3bd9dbfc),
	.w5(32'hbab824db),
	.w6(32'h3c2e9f25),
	.w7(32'h3bb36f6d),
	.w8(32'hbbc8aa19),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004f0c),
	.w1(32'hbb553073),
	.w2(32'hbca6dedd),
	.w3(32'hbb6da5db),
	.w4(32'hbae5bfbb),
	.w5(32'hbae55063),
	.w6(32'hbafe8c66),
	.w7(32'h39ce2e0d),
	.w8(32'hbc220ed2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34ae51),
	.w1(32'h3ac9ac48),
	.w2(32'hba77434c),
	.w3(32'h3d228948),
	.w4(32'h3d0c02b9),
	.w5(32'h39a38374),
	.w6(32'h3cc241d1),
	.w7(32'h3c8ab94f),
	.w8(32'h3b5608f2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c015007),
	.w1(32'h3ba14d29),
	.w2(32'hba9a51c3),
	.w3(32'h3bdd6091),
	.w4(32'h3c097516),
	.w5(32'hb883426d),
	.w6(32'h3b2f8da7),
	.w7(32'h3bb8f988),
	.w8(32'h3b36e3db),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87345a7),
	.w1(32'h3b2b4739),
	.w2(32'hbaa24582),
	.w3(32'h3af6016a),
	.w4(32'h3b240ada),
	.w5(32'hb9c4e3c8),
	.w6(32'h3b932906),
	.w7(32'h3bcf34b9),
	.w8(32'hbb3520ca),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11a05b),
	.w1(32'hba47fa4a),
	.w2(32'h389ad2ec),
	.w3(32'h3bde16cd),
	.w4(32'hba66baf5),
	.w5(32'h3cd82045),
	.w6(32'h3bb6cb1d),
	.w7(32'h3c0c7f8f),
	.w8(32'h3c9c84d8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1f60be),
	.w1(32'h3d1b0bed),
	.w2(32'h3a7c74e2),
	.w3(32'h3daaa214),
	.w4(32'h3da44691),
	.w5(32'hbc080163),
	.w6(32'h3d8facb2),
	.w7(32'h3d7c6da5),
	.w8(32'hbc5e3f1c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a884fa9),
	.w1(32'h3a918b21),
	.w2(32'hbb96c99f),
	.w3(32'hbb0a09e3),
	.w4(32'hbbae7897),
	.w5(32'hb80d4839),
	.w6(32'hbc5149f9),
	.w7(32'hbc4b6f3f),
	.w8(32'h3bf549ed),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce32e1),
	.w1(32'h3b209b3b),
	.w2(32'h3acb1236),
	.w3(32'h3c0342df),
	.w4(32'h3bfda2bb),
	.w5(32'hbb2ff658),
	.w6(32'h3c42b64b),
	.w7(32'h3c157927),
	.w8(32'hbb2ea66d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5eb25),
	.w1(32'hbbbb3316),
	.w2(32'hba38fea3),
	.w3(32'hbb8b61f6),
	.w4(32'hbc450db8),
	.w5(32'hbb8f9edf),
	.w6(32'hbbfa72a8),
	.w7(32'hbc2f0ff7),
	.w8(32'hbc0698f2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a718bf3),
	.w1(32'h3b6c86a2),
	.w2(32'hbaa18b70),
	.w3(32'h3b14b3cc),
	.w4(32'h3b7b5af5),
	.w5(32'hba917a97),
	.w6(32'hbb05692e),
	.w7(32'hba86f8a2),
	.w8(32'hbb360bb8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb264638),
	.w1(32'h3ad7a6a8),
	.w2(32'h3cde3e98),
	.w3(32'hbb1664df),
	.w4(32'h3ae4c4ce),
	.w5(32'h3c6fe705),
	.w6(32'hba390a2f),
	.w7(32'h3b9caf77),
	.w8(32'h3cb00895),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59a543),
	.w1(32'h3c889331),
	.w2(32'h3b6c0cdb),
	.w3(32'hbc7a43d5),
	.w4(32'hbbc0d0ec),
	.w5(32'h3b482b9e),
	.w6(32'hbb30f9fe),
	.w7(32'h3bac5697),
	.w8(32'h3b2cb70a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00a0b1),
	.w1(32'h3b810ebd),
	.w2(32'hbac5ac63),
	.w3(32'hba632a85),
	.w4(32'h3b4af326),
	.w5(32'hb90d6d30),
	.w6(32'hbac6234c),
	.w7(32'h3abc3472),
	.w8(32'h39435080),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fdff17),
	.w1(32'hbab254df),
	.w2(32'hbb9a2696),
	.w3(32'h3b389718),
	.w4(32'hbb32e129),
	.w5(32'h3abae770),
	.w6(32'hbb6ba3e9),
	.w7(32'hbb33df41),
	.w8(32'h3a97eec4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a78d2),
	.w1(32'h3b26183e),
	.w2(32'hbb1c33f7),
	.w3(32'h3baee98f),
	.w4(32'h3b71ecd6),
	.w5(32'hba423cd9),
	.w6(32'h3ba7ff3b),
	.w7(32'h3b2e25a2),
	.w8(32'hbb19a682),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2f2ba),
	.w1(32'h3c60988e),
	.w2(32'h3c1d38d2),
	.w3(32'h3c003e59),
	.w4(32'h3c2bb876),
	.w5(32'h3be0b0a7),
	.w6(32'h3a8f6524),
	.w7(32'h3aad5bb4),
	.w8(32'h3c3b60ee),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c4dde),
	.w1(32'h3c22674f),
	.w2(32'h3ad15dde),
	.w3(32'h3afb6ae3),
	.w4(32'h3beae945),
	.w5(32'h3b5396ee),
	.w6(32'h3c6e781d),
	.w7(32'h3c9df091),
	.w8(32'h3aa18025),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54150a),
	.w1(32'h3b7425b6),
	.w2(32'h3b3ed4fc),
	.w3(32'h3c243ab8),
	.w4(32'h3c1e2ebc),
	.w5(32'hb9a200ae),
	.w6(32'h3ba73a70),
	.w7(32'h3c0fc2f6),
	.w8(32'h3a8ae198),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1afd32),
	.w1(32'hb9f7f0b7),
	.w2(32'hb982a68c),
	.w3(32'h39a98d32),
	.w4(32'h3b77ea70),
	.w5(32'hbb04fbe3),
	.w6(32'hbb2a9581),
	.w7(32'hbaa64c5c),
	.w8(32'h3a912be9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18c7c4),
	.w1(32'h3b0c0b2e),
	.w2(32'h3b7db6e0),
	.w3(32'hbb0b40b8),
	.w4(32'h3b629867),
	.w5(32'h3b38b9b5),
	.w6(32'hb9f73990),
	.w7(32'h3b7aaa9b),
	.w8(32'hba0b4a4c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1014e1),
	.w1(32'hbb175373),
	.w2(32'h3b77c710),
	.w3(32'h3c13d116),
	.w4(32'hb88aba8e),
	.w5(32'hba3d9410),
	.w6(32'h37432e8d),
	.w7(32'hbbb25886),
	.w8(32'hba838f82),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0121b6),
	.w1(32'h3bec0227),
	.w2(32'h3a59f39f),
	.w3(32'h3bbfb764),
	.w4(32'h3a651b87),
	.w5(32'h3afef9b6),
	.w6(32'hb94a76e4),
	.w7(32'hbbbe0cb4),
	.w8(32'h3b9c4897),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c19f),
	.w1(32'h3ba6f771),
	.w2(32'hbbce4dfe),
	.w3(32'h3c5916ef),
	.w4(32'h3c435911),
	.w5(32'hbb5aa6cb),
	.w6(32'h3c3214ad),
	.w7(32'h3c397cc4),
	.w8(32'hb97926fe),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b14a9),
	.w1(32'hbc1a6d62),
	.w2(32'hb97cd1d7),
	.w3(32'hbb0774d0),
	.w4(32'hbb542db6),
	.w5(32'h3a24120d),
	.w6(32'h3baa6946),
	.w7(32'h3bcdedd9),
	.w8(32'h3ad52dc8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ef1eb),
	.w1(32'h3b27c67c),
	.w2(32'hbc7e13e3),
	.w3(32'h3c14b94f),
	.w4(32'h3c487a3e),
	.w5(32'hbcabbd9c),
	.w6(32'h3c362724),
	.w7(32'h3c27875d),
	.w8(32'hbc9c2add),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9216ed),
	.w1(32'hbc1cd14c),
	.w2(32'h3bdedeab),
	.w3(32'hbcce9ff4),
	.w4(32'hbc3e0331),
	.w5(32'h3c363911),
	.w6(32'hbc9cedad),
	.w7(32'hbb87cc26),
	.w8(32'h3af26fa2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cd4b8),
	.w1(32'h3bb3cfde),
	.w2(32'hbadd9b60),
	.w3(32'h3c8c0067),
	.w4(32'h3c08f0e2),
	.w5(32'hbbbaa4d9),
	.w6(32'h3b92db1d),
	.w7(32'hbb095506),
	.w8(32'hbb8e58b3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8822a4),
	.w1(32'hbbf3a6f2),
	.w2(32'hbc4d723a),
	.w3(32'hbb673b1d),
	.w4(32'hbbb5bdbc),
	.w5(32'hbc0ad003),
	.w6(32'h3b33906c),
	.w7(32'h3ba5776f),
	.w8(32'hbbcd3b06),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83d831),
	.w1(32'h3c35c4c6),
	.w2(32'hbb8cbf16),
	.w3(32'h3bb71fca),
	.w4(32'h3bd980b1),
	.w5(32'hbbf293ff),
	.w6(32'h3b20d75b),
	.w7(32'h3bd59f1a),
	.w8(32'hbb52ac61),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b934),
	.w1(32'hbb968a5f),
	.w2(32'h3b00cc82),
	.w3(32'hba00c2d2),
	.w4(32'hbb4817c6),
	.w5(32'h38abd666),
	.w6(32'hbb01f409),
	.w7(32'hbb6bf67c),
	.w8(32'h3a7c2f64),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adecc78),
	.w1(32'h3b879140),
	.w2(32'h3a804691),
	.w3(32'h3b41df3b),
	.w4(32'h3bcda443),
	.w5(32'h3c110e47),
	.w6(32'h3af94b17),
	.w7(32'h3bd6d1aa),
	.w8(32'hba8f15fc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79eb5c),
	.w1(32'hbba800d5),
	.w2(32'hb9d14636),
	.w3(32'h3c5fd07f),
	.w4(32'h3bb79ee6),
	.w5(32'h3a1bac72),
	.w6(32'hb9c0e6c8),
	.w7(32'hbc01e3bb),
	.w8(32'h3a45a997),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9b30a),
	.w1(32'h3a34e3b4),
	.w2(32'hbb7bf293),
	.w3(32'h3b8bba43),
	.w4(32'h3ae46fd3),
	.w5(32'hbb679ff0),
	.w6(32'h3b1ecd3c),
	.w7(32'h3b3a94a7),
	.w8(32'hbbac5eea),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec9511),
	.w1(32'h3a88ee13),
	.w2(32'h3c77c608),
	.w3(32'hba9e4c00),
	.w4(32'h3ad1da15),
	.w5(32'h3bbc250f),
	.w6(32'hbb5490d1),
	.w7(32'h3a2c0d32),
	.w8(32'h3b110934),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e29a9),
	.w1(32'h368af613),
	.w2(32'h3b109f87),
	.w3(32'hbc96ce01),
	.w4(32'hbc696255),
	.w5(32'h3b5e4b86),
	.w6(32'hbc99b517),
	.w7(32'hbc77d6eb),
	.w8(32'h3afebd67),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3e4c4),
	.w1(32'hbb7e2b0f),
	.w2(32'h3ba700a7),
	.w3(32'h3bbe032c),
	.w4(32'h3a95ef2c),
	.w5(32'h3b04ecde),
	.w6(32'h3ba0aeed),
	.w7(32'hbb3caac5),
	.w8(32'hbb00c3b4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11d77e),
	.w1(32'h3b911f7a),
	.w2(32'hbc1b4ec7),
	.w3(32'h3bcebc43),
	.w4(32'h3ae2f037),
	.w5(32'hbc4d6737),
	.w6(32'h3b3804db),
	.w7(32'h3add0f59),
	.w8(32'hbc791a1f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87d40b),
	.w1(32'hbc8c6e0c),
	.w2(32'hbbf254b8),
	.w3(32'hbcad385e),
	.w4(32'hbcaa552e),
	.w5(32'hbbdc4807),
	.w6(32'hbcca9dd3),
	.w7(32'hbcb085fb),
	.w8(32'hbc06003e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c76d41),
	.w1(32'hbb9b94e6),
	.w2(32'h3b97610d),
	.w3(32'h3abcdc92),
	.w4(32'hbc38eb40),
	.w5(32'h3920d40e),
	.w6(32'hbb51efae),
	.w7(32'hbc4715c0),
	.w8(32'h3b8e2032),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad03189),
	.w1(32'h3aa15f35),
	.w2(32'hba589ede),
	.w3(32'hbbd9b5bc),
	.w4(32'h39ddb151),
	.w5(32'h3addfd82),
	.w6(32'hbabe6869),
	.w7(32'h3b3c5239),
	.w8(32'h3b0d2400),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc9f98),
	.w1(32'hb8ed7edd),
	.w2(32'h3b9ab42f),
	.w3(32'h3a28b384),
	.w4(32'hbb9edf33),
	.w5(32'h3afff78f),
	.w6(32'h3bd223f7),
	.w7(32'hbb90f36c),
	.w8(32'h3af36c88),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb068f),
	.w1(32'h3b8a304f),
	.w2(32'hbc17c5d9),
	.w3(32'h3c2f6c9c),
	.w4(32'h3c30d80f),
	.w5(32'hbc5a9673),
	.w6(32'h39106fd2),
	.w7(32'h3adb3469),
	.w8(32'hbc14117d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50c608),
	.w1(32'hbbbe081b),
	.w2(32'h3b4a97fa),
	.w3(32'hbca4ee66),
	.w4(32'hbc5d15e3),
	.w5(32'h3b62baa1),
	.w6(32'hbc69dc30),
	.w7(32'hbbb2c1f0),
	.w8(32'h3b45966b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7efb1a),
	.w1(32'h3be5177e),
	.w2(32'hbb876396),
	.w3(32'h3bef2034),
	.w4(32'h3c16a3d8),
	.w5(32'hbb038b61),
	.w6(32'h3af02069),
	.w7(32'h3b614cac),
	.w8(32'h39c2209b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adee8d5),
	.w1(32'hba9e6acc),
	.w2(32'h39807741),
	.w3(32'h3b34d55a),
	.w4(32'hbaf1bcd7),
	.w5(32'hbb585eb7),
	.w6(32'hb9bd4dbc),
	.w7(32'hba0d3d3e),
	.w8(32'hbb50fb08),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976d971),
	.w1(32'h3984b9a8),
	.w2(32'h3b3093a8),
	.w3(32'h3b44922f),
	.w4(32'h3ab0e469),
	.w5(32'h3bf379f2),
	.w6(32'h3b429f30),
	.w7(32'h3922b82b),
	.w8(32'hb98d69f9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba128f6),
	.w1(32'h3bfbb82c),
	.w2(32'h3c1eac2e),
	.w3(32'h3bfd4030),
	.w4(32'h3c383c36),
	.w5(32'h3b19e015),
	.w6(32'h3c709a38),
	.w7(32'h3c502b60),
	.w8(32'h3ba81253),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a46d8),
	.w1(32'h3b9bf509),
	.w2(32'h3b896056),
	.w3(32'hbc8837fc),
	.w4(32'hbbeec22d),
	.w5(32'h3b899159),
	.w6(32'hbc2f16ad),
	.w7(32'hbb00e315),
	.w8(32'h38e8fabb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6693f),
	.w1(32'h3a0dc3c2),
	.w2(32'h3ca443f7),
	.w3(32'h3bd3e2b3),
	.w4(32'hba86822a),
	.w5(32'h3c565b0d),
	.w6(32'hb97778e9),
	.w7(32'hbbe1158c),
	.w8(32'h3bb12f20),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bd313),
	.w1(32'h3bb2423a),
	.w2(32'h3b9cc378),
	.w3(32'hbc12b8ef),
	.w4(32'hbc4bfd8d),
	.w5(32'h3a867cbc),
	.w6(32'hbca24894),
	.w7(32'hbc9cc148),
	.w8(32'hbbbab2d7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdbdb5),
	.w1(32'h3ba35fc1),
	.w2(32'h38a1e322),
	.w3(32'h3b5956a8),
	.w4(32'h3bf53cce),
	.w5(32'hb883c076),
	.w6(32'h3a129bec),
	.w7(32'h3a6a69e0),
	.w8(32'hbb866383),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba513101),
	.w1(32'h3b00fd92),
	.w2(32'hbb08f289),
	.w3(32'h3ab901cb),
	.w4(32'h3bb9d1cd),
	.w5(32'hbbf9e394),
	.w6(32'h3b0ef7c5),
	.w7(32'hbb362826),
	.w8(32'hbaf299c4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aac56),
	.w1(32'hbb100483),
	.w2(32'h3c3f8f9c),
	.w3(32'hbba50706),
	.w4(32'hbb375352),
	.w5(32'h3b2f4d49),
	.w6(32'hba9c9567),
	.w7(32'hbb5463ac),
	.w8(32'h3b88400c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7dc1e9),
	.w1(32'h3b4f57ee),
	.w2(32'h3b0afc0f),
	.w3(32'hbafad2ab),
	.w4(32'h37636b8b),
	.w5(32'h3a2fdddc),
	.w6(32'hba8b4806),
	.w7(32'h3ad42351),
	.w8(32'h3b2e907a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9aa85),
	.w1(32'hbb1be433),
	.w2(32'hbb451fd6),
	.w3(32'h3bceb4d9),
	.w4(32'hba0d8361),
	.w5(32'hbc31b9e7),
	.w6(32'h3c00f32b),
	.w7(32'h3a2c8af3),
	.w8(32'hbc0174f0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc246c32),
	.w1(32'hbc16dcd3),
	.w2(32'h3b0ba61c),
	.w3(32'hbcad068b),
	.w4(32'hbca14e8b),
	.w5(32'hb8d1a926),
	.w6(32'hbc9f4ea1),
	.w7(32'hbc7d8a7b),
	.w8(32'h3a737ccb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88570c),
	.w1(32'h3b9a69f0),
	.w2(32'hbb920d12),
	.w3(32'h3acabcca),
	.w4(32'hb9e5b808),
	.w5(32'hbc3acd35),
	.w6(32'h3a4263db),
	.w7(32'h3a690d1a),
	.w8(32'hba85adcb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc183a63),
	.w1(32'hbb6dbb03),
	.w2(32'h3b21810b),
	.w3(32'hbc3f22ec),
	.w4(32'hbbacbafc),
	.w5(32'h3bb3909a),
	.w6(32'hbb57ad31),
	.w7(32'hbbb81095),
	.w8(32'hbb53eaa8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5408a9),
	.w1(32'h3c1c121e),
	.w2(32'hbba91d39),
	.w3(32'h3c83304b),
	.w4(32'h3c5865a7),
	.w5(32'hbb5bb90e),
	.w6(32'h3bb017dc),
	.w7(32'h3b661572),
	.w8(32'hbbaa88fb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a7c02),
	.w1(32'hb82ecaa1),
	.w2(32'hbb90afac),
	.w3(32'h3bae31c5),
	.w4(32'hbbcca6b5),
	.w5(32'hbbc86d71),
	.w6(32'hb9c15a65),
	.w7(32'hbbb20955),
	.w8(32'hbbe43993),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f20af),
	.w1(32'hbbb7704d),
	.w2(32'h3b87df78),
	.w3(32'hbbd2287a),
	.w4(32'hbbd11179),
	.w5(32'hbc4af3e9),
	.w6(32'hbbccb156),
	.w7(32'hbb9f3219),
	.w8(32'hbc19f342),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32f05e),
	.w1(32'hbc3fa47e),
	.w2(32'hbb087603),
	.w3(32'hbd33cb79),
	.w4(32'hbd1e6ef2),
	.w5(32'h39a76f3f),
	.w6(32'hbd1f1bcb),
	.w7(32'hbcfcaccd),
	.w8(32'hb72a41ed),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0df90d),
	.w1(32'h3a53f41e),
	.w2(32'h3b4acef9),
	.w3(32'h3b847ee8),
	.w4(32'h3b0940df),
	.w5(32'h3b4fb7c8),
	.w6(32'hbb17c689),
	.w7(32'hbb2db499),
	.w8(32'h3ad64cd3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93f4d7),
	.w1(32'h3a8edabb),
	.w2(32'h3925caf3),
	.w3(32'h3a400daa),
	.w4(32'h3a775652),
	.w5(32'h3b2a68fc),
	.w6(32'hbb1b4dc4),
	.w7(32'hbb91bfae),
	.w8(32'h3b094770),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbc5db),
	.w1(32'h3c180e0b),
	.w2(32'hbaf75f1b),
	.w3(32'h3c250611),
	.w4(32'h3c58176d),
	.w5(32'h3a847944),
	.w6(32'h3c1f2c62),
	.w7(32'h3c3fe12c),
	.w8(32'h3ab9abff),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e221a),
	.w1(32'h3b874c34),
	.w2(32'hb9f137a5),
	.w3(32'h3b7e6909),
	.w4(32'hbb05833c),
	.w5(32'h3b654504),
	.w6(32'h3abea475),
	.w7(32'h3b96da25),
	.w8(32'h3913cb0d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c145f43),
	.w1(32'h3bcd76a5),
	.w2(32'hb9aa2f2a),
	.w3(32'h3bb7dc92),
	.w4(32'h3c0f43f0),
	.w5(32'h3bc084e2),
	.w6(32'h3bd9e181),
	.w7(32'h3c116ed5),
	.w8(32'h3b6412f7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4be0bf),
	.w1(32'hb9b82c08),
	.w2(32'hbb3b7834),
	.w3(32'h3c7c94ee),
	.w4(32'hbb896aab),
	.w5(32'hbb8c4044),
	.w6(32'h3c222ca1),
	.w7(32'hbc2e4acc),
	.w8(32'hbabd94c0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980d2cc),
	.w1(32'hba31fd63),
	.w2(32'hbb7089e4),
	.w3(32'hba487a03),
	.w4(32'h3b63fb9a),
	.w5(32'hbb01c0ac),
	.w6(32'hbb140d49),
	.w7(32'hb99c7483),
	.w8(32'hbbc67df3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2f610),
	.w1(32'h3b8a1a73),
	.w2(32'hbb04eec0),
	.w3(32'hba73ff58),
	.w4(32'hba2eaee8),
	.w5(32'hbb820ae0),
	.w6(32'hbafb9f7c),
	.w7(32'hbb07d05d),
	.w8(32'hbbbfb884),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb60e6a),
	.w1(32'h39bcaa94),
	.w2(32'h3a9322a7),
	.w3(32'h3b9e3eb5),
	.w4(32'hbb5382d9),
	.w5(32'hbad17202),
	.w6(32'h3b471d63),
	.w7(32'hbbd52189),
	.w8(32'hbbaa83de),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be084f4),
	.w1(32'h3b0ebbdf),
	.w2(32'h3ba00f95),
	.w3(32'h3b57be82),
	.w4(32'hbb284467),
	.w5(32'h3c03584a),
	.w6(32'hbb35f766),
	.w7(32'hbbeb567a),
	.w8(32'h3b6a7d94),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01dd3b),
	.w1(32'h3be9e547),
	.w2(32'hbaa89cbc),
	.w3(32'h3c14ed00),
	.w4(32'h3c1f93f8),
	.w5(32'hba092bef),
	.w6(32'h3b768384),
	.w7(32'h3bb062c0),
	.w8(32'hbc1250eb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d19bfe),
	.w1(32'h3bc8cc4b),
	.w2(32'hbb8e3922),
	.w3(32'hb9e9bf45),
	.w4(32'h3c0285b6),
	.w5(32'hbbb91c64),
	.w6(32'hbbabb978),
	.w7(32'h3aeb0f6f),
	.w8(32'hbbf1316e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75908c),
	.w1(32'h3bbc670c),
	.w2(32'hbb0d6172),
	.w3(32'hbb889d79),
	.w4(32'h3c02fe9f),
	.w5(32'hbac7a6f7),
	.w6(32'hbb84ac3e),
	.w7(32'h3bf2b172),
	.w8(32'hbac386a5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e2cee),
	.w1(32'hbb2c825e),
	.w2(32'hbb4a6f30),
	.w3(32'h3adc1204),
	.w4(32'hbaf37fab),
	.w5(32'h3b194db6),
	.w6(32'h3bae5073),
	.w7(32'hb9e05b60),
	.w8(32'h3ba4f1a2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fc18b),
	.w1(32'hbaaade2f),
	.w2(32'h3aabf0a0),
	.w3(32'h3b4feed9),
	.w4(32'h3b98c147),
	.w5(32'hbb533b07),
	.w6(32'h39a09fb1),
	.w7(32'h3b4b365c),
	.w8(32'hbb8c2ede),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b376ef3),
	.w1(32'h3b549d82),
	.w2(32'hbbd161f5),
	.w3(32'h39ddb904),
	.w4(32'h3b8b14c9),
	.w5(32'hbb0b85a0),
	.w6(32'h3b9e930e),
	.w7(32'h3bd3b5fc),
	.w8(32'hbba8c4e3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91b01e),
	.w1(32'h3b0afe31),
	.w2(32'hbb373436),
	.w3(32'hba6cbb82),
	.w4(32'hbae99f0e),
	.w5(32'hbbac548b),
	.w6(32'hbb0da486),
	.w7(32'h38dc405c),
	.w8(32'hbb62b55f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32d0ee),
	.w1(32'h3bbf01a1),
	.w2(32'h3a015305),
	.w3(32'h3b855a4e),
	.w4(32'h3c1022e8),
	.w5(32'hbaec2578),
	.w6(32'h3bfa8c80),
	.w7(32'h3b3ea859),
	.w8(32'hbb803b43),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e4d87),
	.w1(32'hbb10a491),
	.w2(32'hb9ef4e62),
	.w3(32'h3a7c9101),
	.w4(32'h3b238c27),
	.w5(32'hba29e5c0),
	.w6(32'hba1aa491),
	.w7(32'h3b5caae4),
	.w8(32'hbb6a1084),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a4dbc),
	.w1(32'hba84f72c),
	.w2(32'hbb81d5ad),
	.w3(32'h3a0a2c56),
	.w4(32'h3be3f62e),
	.w5(32'hba94dbc7),
	.w6(32'h3b40617d),
	.w7(32'h3bcaf990),
	.w8(32'hbb1cb6d5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b324d5a),
	.w1(32'h3b2e5db8),
	.w2(32'hbc244ba8),
	.w3(32'h3b4b432a),
	.w4(32'h3b38d5eb),
	.w5(32'hbc0f4de7),
	.w6(32'h3b2702d2),
	.w7(32'h3bae4b3f),
	.w8(32'hbb6fc443),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9cf54),
	.w1(32'hbbeaacae),
	.w2(32'hbc0dcd42),
	.w3(32'hbb857605),
	.w4(32'hbb89b438),
	.w5(32'hbc7776af),
	.w6(32'h3a0e9687),
	.w7(32'h396befb8),
	.w8(32'hbc5b2b7d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8036a2),
	.w1(32'hb94d412d),
	.w2(32'hbb7889b6),
	.w3(32'hbbbb3720),
	.w4(32'hbc1ea18f),
	.w5(32'hbb187c1f),
	.w6(32'hbc5ff333),
	.w7(32'hbc7ab3ee),
	.w8(32'hbc0b909f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45c5fd),
	.w1(32'hba89eaab),
	.w2(32'h3ae0d767),
	.w3(32'h3a6bac50),
	.w4(32'h3b29905c),
	.w5(32'hb9e559fd),
	.w6(32'hbbad36d5),
	.w7(32'hbb4dd105),
	.w8(32'h3b459c37),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d50a8),
	.w1(32'h3a1f4883),
	.w2(32'hbb501ea2),
	.w3(32'hb936204e),
	.w4(32'h3ae73648),
	.w5(32'hbabe620f),
	.w6(32'h3b99fa2d),
	.w7(32'h3b05b200),
	.w8(32'hbb38c5a3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47b0bd),
	.w1(32'hbb37852e),
	.w2(32'hbb3a5f28),
	.w3(32'hbb449360),
	.w4(32'hbb802b6a),
	.w5(32'hb928948c),
	.w6(32'hb9fee76e),
	.w7(32'hbb3df5bb),
	.w8(32'h39142d0f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72ad88),
	.w1(32'h3b0a52b0),
	.w2(32'hbcd2586d),
	.w3(32'h3b70e6be),
	.w4(32'h39ab3706),
	.w5(32'hbcc49cfb),
	.w6(32'h3bb243e0),
	.w7(32'h3b7a98d5),
	.w8(32'hbcaf5ac0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0560f),
	.w1(32'hbc896fbc),
	.w2(32'hbc719772),
	.w3(32'hbc1b1acc),
	.w4(32'hbbd9e65e),
	.w5(32'hbc6929a0),
	.w6(32'hbc171ee7),
	.w7(32'hbbd95b9b),
	.w8(32'hbc8e48cd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc167467),
	.w1(32'hbc23a309),
	.w2(32'h3b35206f),
	.w3(32'hbb6c7eb9),
	.w4(32'hbbd57af6),
	.w5(32'h3bed12a5),
	.w6(32'hbc280830),
	.w7(32'hbc3d1497),
	.w8(32'h39c02b81),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babeefc),
	.w1(32'hb9687fe5),
	.w2(32'hbbbb3090),
	.w3(32'h3bc01a89),
	.w4(32'h3b6226d5),
	.w5(32'hbbc380cb),
	.w6(32'h3b142ab9),
	.w7(32'hbb189d07),
	.w8(32'hbb930b1b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb78ae7),
	.w1(32'h3ae5c2d4),
	.w2(32'h3b51d959),
	.w3(32'hbb1e184f),
	.w4(32'h3ba68b04),
	.w5(32'hbb37169b),
	.w6(32'hbb13a8b2),
	.w7(32'h3bd2af15),
	.w8(32'h39a9ba2d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03369e),
	.w1(32'h3bf860fe),
	.w2(32'hb8ee9a2b),
	.w3(32'h3b935b38),
	.w4(32'h3c3be13c),
	.w5(32'hba7c1829),
	.w6(32'h3be60592),
	.w7(32'h3c4e345e),
	.w8(32'h37e8dc13),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac33fc2),
	.w1(32'hbaff8f64),
	.w2(32'h3acc00fa),
	.w3(32'hbb505281),
	.w4(32'h3b2710e2),
	.w5(32'h399477fe),
	.w6(32'hba9cabd3),
	.w7(32'hbb2deb7f),
	.w8(32'hbb8d2026),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b955dbd),
	.w1(32'h3bb0af52),
	.w2(32'h39f2f7c5),
	.w3(32'h3b2eabe1),
	.w4(32'h3b4d54c2),
	.w5(32'h3b55ee4e),
	.w6(32'hba0442f5),
	.w7(32'hb90652ce),
	.w8(32'h3c0908c7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19aef9),
	.w1(32'hbbb5bc40),
	.w2(32'hba8380b0),
	.w3(32'hbad3b60f),
	.w4(32'hbb7af7e2),
	.w5(32'h3b70730e),
	.w6(32'h3bad9a24),
	.w7(32'h3b414551),
	.w8(32'h3af5bab7),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e79b8),
	.w1(32'h3c4a5336),
	.w2(32'h3bcb72c8),
	.w3(32'h3c86da4d),
	.w4(32'h3c8ca4a9),
	.w5(32'hba97ef91),
	.w6(32'h3c328484),
	.w7(32'h3c884168),
	.w8(32'hbaa8acdb),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a82f2),
	.w1(32'h3888fa4a),
	.w2(32'h3afee3cf),
	.w3(32'hb9ae6301),
	.w4(32'hbb5c74ed),
	.w5(32'hba752afc),
	.w6(32'hbb411319),
	.w7(32'hbb0a5a78),
	.w8(32'hbb5dca7c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b4054),
	.w1(32'h3a79325e),
	.w2(32'h3b204319),
	.w3(32'h3aa0f928),
	.w4(32'h3acd903b),
	.w5(32'hbbcaa5ef),
	.w6(32'hba4f873c),
	.w7(32'h3b868b50),
	.w8(32'hbad8e4e7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a1177),
	.w1(32'h3b812dd1),
	.w2(32'h39659c49),
	.w3(32'hba23b860),
	.w4(32'h3a45d021),
	.w5(32'hba1e4fb1),
	.w6(32'h39bcd440),
	.w7(32'hbb93f6c4),
	.w8(32'hb9ffea04),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a7bd8),
	.w1(32'hba60fca0),
	.w2(32'hbb29879a),
	.w3(32'h3b0c4026),
	.w4(32'h3baf4e5a),
	.w5(32'hbc80bac9),
	.w6(32'hba2c2fd0),
	.w7(32'h3abf5112),
	.w8(32'hbc4d6f14),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18cade),
	.w1(32'hbc41c1c5),
	.w2(32'hbb7c849a),
	.w3(32'hbd2c4077),
	.w4(32'hbd2c7e4a),
	.w5(32'hb9a8f0a9),
	.w6(32'hbd1ed674),
	.w7(32'hbd079abc),
	.w8(32'hbb92af0b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf690a4),
	.w1(32'h3ad3b823),
	.w2(32'hbb2b76d9),
	.w3(32'h3abf7a9f),
	.w4(32'h3b372875),
	.w5(32'hbbb868fb),
	.w6(32'hb96e7ddb),
	.w7(32'h3ae520df),
	.w8(32'hbb362994),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba463a77),
	.w1(32'hbb13de01),
	.w2(32'hbad5bd93),
	.w3(32'hb9a21d3a),
	.w4(32'hba490816),
	.w5(32'hba8e067a),
	.w6(32'h3b5f0f52),
	.w7(32'h3b1bc507),
	.w8(32'hbbc308e2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6e96f),
	.w1(32'h3ae34c79),
	.w2(32'hbb7d4fc8),
	.w3(32'h3afa9434),
	.w4(32'h3aa9ced7),
	.w5(32'hbbb36e69),
	.w6(32'hbbc89789),
	.w7(32'hbb6784ec),
	.w8(32'hbc6635d1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c0e42),
	.w1(32'hbbc8fb43),
	.w2(32'hbb734660),
	.w3(32'hbbe15545),
	.w4(32'hbc2dd3bb),
	.w5(32'hb9c52235),
	.w6(32'hbc7b6b67),
	.w7(32'hbc86ab59),
	.w8(32'hbba689b6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96f93b),
	.w1(32'hbb051e0c),
	.w2(32'hbc934fd4),
	.w3(32'h3b82dd8e),
	.w4(32'h3b558acd),
	.w5(32'hbca46645),
	.w6(32'h3b0f142e),
	.w7(32'hbabd7219),
	.w8(32'hbc962454),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ecebf),
	.w1(32'hbc56686e),
	.w2(32'hbbcebe70),
	.w3(32'hbc9e4b80),
	.w4(32'hbc77e457),
	.w5(32'hbb0e496b),
	.w6(32'hbc8a37ef),
	.w7(32'hbc247a23),
	.w8(32'hbb644e17),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb001e47),
	.w1(32'hbb19c067),
	.w2(32'h3b362d94),
	.w3(32'h3baa8583),
	.w4(32'hbb934ac8),
	.w5(32'h3ad7478b),
	.w6(32'h3a65d4f8),
	.w7(32'hbbfaed89),
	.w8(32'h3b849371),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b413925),
	.w1(32'h3bda35c2),
	.w2(32'h39d0839d),
	.w3(32'h3ba25164),
	.w4(32'h3adf8480),
	.w5(32'hbb1ef505),
	.w6(32'h3a95b316),
	.w7(32'h3b64e381),
	.w8(32'hbba4338e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93e4f8),
	.w1(32'h3ba15d51),
	.w2(32'h3c0e79d9),
	.w3(32'h3b3c78ba),
	.w4(32'h3ab9c4d6),
	.w5(32'h3ad6d251),
	.w6(32'h3a837dca),
	.w7(32'h390f0961),
	.w8(32'hbaef243b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b7687),
	.w1(32'hb7fdb1d2),
	.w2(32'hbb8cd1c8),
	.w3(32'hbc4c3673),
	.w4(32'hbc61a264),
	.w5(32'hba5f63ce),
	.w6(32'hbc84b0e5),
	.w7(32'hbc64f3d0),
	.w8(32'h3b1df41c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb017b3a),
	.w1(32'h3bcca9ba),
	.w2(32'hbb9a6770),
	.w3(32'h38bb256c),
	.w4(32'h3c24c30c),
	.w5(32'hbb94b0e6),
	.w6(32'h3b855324),
	.w7(32'h3c36ea5a),
	.w8(32'hbbc530bc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac86dec),
	.w1(32'hbb06ac17),
	.w2(32'h3a5fec55),
	.w3(32'h3b0bcee4),
	.w4(32'hbb8c0e27),
	.w5(32'h3bb9fa03),
	.w6(32'h3bc828ce),
	.w7(32'h3b83c511),
	.w8(32'h3b9a5ac8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7863f3),
	.w1(32'h3b49ca16),
	.w2(32'hbb929593),
	.w3(32'h3b2f4060),
	.w4(32'hbac5a5de),
	.w5(32'hbbb0022e),
	.w6(32'h3ba03a5f),
	.w7(32'h3b8cc6d6),
	.w8(32'hbb3ce3b8),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9823d37),
	.w1(32'h39534dd5),
	.w2(32'hba52ede6),
	.w3(32'h3b7213da),
	.w4(32'h3ad7dd6a),
	.w5(32'h3a63391a),
	.w6(32'h3af44a1d),
	.w7(32'hba36bf7e),
	.w8(32'hb861b22d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee05e3),
	.w1(32'h3af7bc22),
	.w2(32'hbbe8eff0),
	.w3(32'h3a960a03),
	.w4(32'hb8855088),
	.w5(32'hbb79fe5d),
	.w6(32'hba974b9d),
	.w7(32'h3b3f54e1),
	.w8(32'h3a0b441d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25d8e4),
	.w1(32'h3adf8c21),
	.w2(32'hbcb57ef6),
	.w3(32'hbbb4e806),
	.w4(32'hbb595923),
	.w5(32'hbc7deb51),
	.w6(32'hbbb42b40),
	.w7(32'hbadb7e6d),
	.w8(32'hbca11394),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5e4ec),
	.w1(32'hbc10b613),
	.w2(32'h39e05e55),
	.w3(32'h3c2d0d64),
	.w4(32'h3bca8cef),
	.w5(32'hbab8a746),
	.w6(32'hbb143916),
	.w7(32'hbb86ff16),
	.w8(32'hbc0ae5b6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b947493),
	.w1(32'hbb23d15d),
	.w2(32'hbb06442c),
	.w3(32'h3b9a5dd6),
	.w4(32'hbbac505f),
	.w5(32'hbbee0fa0),
	.w6(32'h3b569d1a),
	.w7(32'hbb16d55c),
	.w8(32'hb9afba50),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7bbe2),
	.w1(32'h3bc12735),
	.w2(32'hbb5bb442),
	.w3(32'hb9b625c6),
	.w4(32'h3b73e1f7),
	.w5(32'hbb012f62),
	.w6(32'h3a2be920),
	.w7(32'hba506aaf),
	.w8(32'hbb0c22ce),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbababe37),
	.w1(32'hbaebed30),
	.w2(32'h3a9ba310),
	.w3(32'hba108c7c),
	.w4(32'hbad38929),
	.w5(32'hba2b56b4),
	.w6(32'h393507ef),
	.w7(32'hbb3bedcf),
	.w8(32'h3ada7013),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987c0e),
	.w1(32'hba5f402b),
	.w2(32'hbb47f06c),
	.w3(32'h3b60c284),
	.w4(32'hbb80ebfd),
	.w5(32'hbc24e4ee),
	.w6(32'h3b95fcb6),
	.w7(32'hb9a18afb),
	.w8(32'hbbb19ae6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ed15a),
	.w1(32'h3be8356d),
	.w2(32'hbadf0d17),
	.w3(32'h3a85421e),
	.w4(32'h3c80eb06),
	.w5(32'hbbc957f9),
	.w6(32'h3c01c459),
	.w7(32'h3cbf44ac),
	.w8(32'h3b405a3f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab22fd),
	.w1(32'h3c3527b5),
	.w2(32'hbafb0f68),
	.w3(32'hbbf12e8b),
	.w4(32'hbc2fdb59),
	.w5(32'hbb18701c),
	.w6(32'hbbeec4ae),
	.w7(32'hbc16f34c),
	.w8(32'hbc0157f0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7468a9),
	.w1(32'hbc0c37f7),
	.w2(32'h3bf24e4d),
	.w3(32'hbc17a5a6),
	.w4(32'hbc8b3a79),
	.w5(32'h3c5a2b6d),
	.w6(32'hbc6e993a),
	.w7(32'hbca2cce9),
	.w8(32'h393a0794),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfed40b),
	.w1(32'h3b58911a),
	.w2(32'h3b24d6bc),
	.w3(32'h3b268409),
	.w4(32'hbba88a11),
	.w5(32'hbaedaff0),
	.w6(32'hbc65e18b),
	.w7(32'hbc1dcb43),
	.w8(32'h3b6543fa),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc61235),
	.w1(32'hbc1bd06a),
	.w2(32'hbbcb56d2),
	.w3(32'hbc394af0),
	.w4(32'hbc8574cf),
	.w5(32'hbae17d00),
	.w6(32'h3a8c6a6b),
	.w7(32'hbb5de07d),
	.w8(32'hbb151dd0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae8a6b),
	.w1(32'h3c1bc7dc),
	.w2(32'hbc67f49c),
	.w3(32'h3c900e0e),
	.w4(32'h3cb963e0),
	.w5(32'hbc8ad4a1),
	.w6(32'h3c861dfb),
	.w7(32'h3c9ebc78),
	.w8(32'hbc55f992),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34aba5),
	.w1(32'hbc314d81),
	.w2(32'hbc55b33f),
	.w3(32'hbc88609e),
	.w4(32'hbcb68a7b),
	.w5(32'hbc137b51),
	.w6(32'hbcba63d3),
	.w7(32'hbcacde66),
	.w8(32'hbb31663f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b983aea),
	.w1(32'h3c832277),
	.w2(32'h3c8075cb),
	.w3(32'h3c800ee4),
	.w4(32'h3d09119d),
	.w5(32'h3c8fbf03),
	.w6(32'h3cb6d8fb),
	.w7(32'h3d112517),
	.w8(32'h3c0a4e76),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3daa79),
	.w1(32'h3c3de104),
	.w2(32'hbb20f23c),
	.w3(32'h3c3d9a1a),
	.w4(32'h3b3823a6),
	.w5(32'hbbf9c137),
	.w6(32'h3bdd7a1a),
	.w7(32'h3ae45a8d),
	.w8(32'hbc3a5a20),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66a206),
	.w1(32'hbc036132),
	.w2(32'h3b8ee76c),
	.w3(32'hbc0e0703),
	.w4(32'hbc7181fa),
	.w5(32'hbb5a71a9),
	.w6(32'hbc25a82f),
	.w7(32'hbc9860ba),
	.w8(32'hbb0ebe7a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd82d44),
	.w1(32'h3bc29977),
	.w2(32'hbc227696),
	.w3(32'hbba61fae),
	.w4(32'h3a3df418),
	.w5(32'h393f7a31),
	.w6(32'hbb63a965),
	.w7(32'hbbf1e08d),
	.w8(32'h3b438b98),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7557462),
	.w1(32'h3afc3f60),
	.w2(32'hbc2878e3),
	.w3(32'h3c7cf01e),
	.w4(32'h3c0529d6),
	.w5(32'hbb8e7dea),
	.w6(32'h3ccc6d63),
	.w7(32'h3c70617c),
	.w8(32'hbbdda735),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba057d),
	.w1(32'hbb8b4e19),
	.w2(32'h391e9821),
	.w3(32'h3c7ad631),
	.w4(32'h3c3ad47b),
	.w5(32'hbbe20336),
	.w6(32'h3c0a86c2),
	.w7(32'h3c07e935),
	.w8(32'hbc07d016),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dc18b),
	.w1(32'h3b742b94),
	.w2(32'hbb8069d4),
	.w3(32'hba22d200),
	.w4(32'h3b79f743),
	.w5(32'h3a505463),
	.w6(32'hbb958598),
	.w7(32'hbc0b85b2),
	.w8(32'h3bfe107e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0af28),
	.w1(32'h3b6869a6),
	.w2(32'hbbb43df3),
	.w3(32'h3a4349ea),
	.w4(32'h3bb2921c),
	.w5(32'hbc0f0987),
	.w6(32'hbb23ca71),
	.w7(32'hbc140d13),
	.w8(32'hbb81851c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21a036),
	.w1(32'h3b990556),
	.w2(32'hbb9779bb),
	.w3(32'h3a344f5a),
	.w4(32'h3b75ae0a),
	.w5(32'hbcbf8029),
	.w6(32'h3b84b2db),
	.w7(32'h3bc14366),
	.w8(32'hbc704bba),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc807001),
	.w1(32'hbbb8f752),
	.w2(32'hbb627bcc),
	.w3(32'hbd39a941),
	.w4(32'hbce4e98e),
	.w5(32'hbc2d6cce),
	.w6(32'hbd23b30e),
	.w7(32'hbca42613),
	.w8(32'hbc1d88c5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843864),
	.w1(32'hbbb4dbfd),
	.w2(32'h3bbf1dc0),
	.w3(32'hbc3cb207),
	.w4(32'h3c07cf7b),
	.w5(32'h3c2259f7),
	.w6(32'h3c0f5876),
	.w7(32'h3c4c9b41),
	.w8(32'h3b962e5a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31faf7),
	.w1(32'hbaf5c648),
	.w2(32'hbc7b5c39),
	.w3(32'h3b7cfcee),
	.w4(32'hbc1c46ef),
	.w5(32'hbc7baa7d),
	.w6(32'hbbd9f8a6),
	.w7(32'hbcbf0b5c),
	.w8(32'hbc93679d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87ce10),
	.w1(32'hbb11e806),
	.w2(32'hbbc35e71),
	.w3(32'hbc924ad1),
	.w4(32'hbb404006),
	.w5(32'hbc2d8aea),
	.w6(32'hbc983703),
	.w7(32'hb9d093f9),
	.w8(32'hbb9ccb88),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a29eb),
	.w1(32'hbac02eeb),
	.w2(32'hbc1eeaea),
	.w3(32'hbc20d44c),
	.w4(32'hbba9e52d),
	.w5(32'hbc2fb2c9),
	.w6(32'hbbe42a01),
	.w7(32'hbb119484),
	.w8(32'hbbd74cb6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd08640),
	.w1(32'h39a41edf),
	.w2(32'hbbeacdf7),
	.w3(32'hbc62eaee),
	.w4(32'hbc49a174),
	.w5(32'hbaadda31),
	.w6(32'hbc1bb685),
	.w7(32'h395a97fd),
	.w8(32'hbc08c1f4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d7864),
	.w1(32'h3c33f2ab),
	.w2(32'h3c6a4bdd),
	.w3(32'h3b1a9838),
	.w4(32'hbab3af54),
	.w5(32'h3c5a8af6),
	.w6(32'hbb962d62),
	.w7(32'hbafa1751),
	.w8(32'h3ad0d9bf),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7879d),
	.w1(32'h3c55c383),
	.w2(32'hbbd69df5),
	.w3(32'h3ca61198),
	.w4(32'h3cc25643),
	.w5(32'hbb670966),
	.w6(32'h3c640a47),
	.w7(32'h3cbd9b7d),
	.w8(32'hbc41f1ef),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81c102),
	.w1(32'h39a1a40c),
	.w2(32'hba095647),
	.w3(32'h3bf175f0),
	.w4(32'h3c0bd467),
	.w5(32'hbac909b9),
	.w6(32'hbb5740bc),
	.w7(32'h3ba8d1d7),
	.w8(32'h3c44c3d8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba34b88),
	.w1(32'hbbcd3784),
	.w2(32'hbb9ad9f2),
	.w3(32'hbadce1b9),
	.w4(32'hba6d7f45),
	.w5(32'h389d97d1),
	.w6(32'h3bcff800),
	.w7(32'hb88303b3),
	.w8(32'hb79f2d82),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebe9b6),
	.w1(32'h3bdc8fa6),
	.w2(32'hbc1fc146),
	.w3(32'h3b05e7f2),
	.w4(32'h3bb21ddd),
	.w5(32'hbc587c78),
	.w6(32'h3b69a070),
	.w7(32'h3a35d14f),
	.w8(32'hbc25e996),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02ed4a),
	.w1(32'hbc362c46),
	.w2(32'hbb29b8bf),
	.w3(32'hbc81e694),
	.w4(32'hbcacad2e),
	.w5(32'h3b93c3f9),
	.w6(32'hbc42d222),
	.w7(32'hbaf2db7c),
	.w8(32'h3c02f8ec),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64c130),
	.w1(32'h3c55250d),
	.w2(32'hbc506ece),
	.w3(32'h3bafcb34),
	.w4(32'h3a3595e3),
	.w5(32'hbc82b800),
	.w6(32'h3ba2fabe),
	.w7(32'h3ba76041),
	.w8(32'hbc6bf483),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9d8d3),
	.w1(32'h3b16b10a),
	.w2(32'hbaedc332),
	.w3(32'h3b353218),
	.w4(32'hbc324be7),
	.w5(32'h3b280476),
	.w6(32'hbba60468),
	.w7(32'hbc6e1134),
	.w8(32'h3be6d796),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb079a8),
	.w1(32'h3c75354d),
	.w2(32'h3c15f608),
	.w3(32'h3c7c03fa),
	.w4(32'h3cdfdc6f),
	.w5(32'h3bc1356e),
	.w6(32'h3ca2e75d),
	.w7(32'h3ce1a1a9),
	.w8(32'h3a6eb971),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d9f67),
	.w1(32'h3c0f3897),
	.w2(32'hbc7cba66),
	.w3(32'h3c4d863b),
	.w4(32'h3c370097),
	.w5(32'hbcd82937),
	.w6(32'hbb736df3),
	.w7(32'hbc1d5b33),
	.w8(32'hbcbca337),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc248b4c),
	.w1(32'h3a13e465),
	.w2(32'h3b7090b5),
	.w3(32'hbc665067),
	.w4(32'hba985f98),
	.w5(32'h3ae414d9),
	.w6(32'hbc519502),
	.w7(32'hbb7fb632),
	.w8(32'h3b875187),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb93c0d),
	.w1(32'hbc22da1c),
	.w2(32'hbbf8acbb),
	.w3(32'hbcb919df),
	.w4(32'hbd07ad70),
	.w5(32'hbbc4e8cf),
	.w6(32'hbc19fce5),
	.w7(32'hbcf350bc),
	.w8(32'hbbbb47e3),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c873f),
	.w1(32'hba7d322f),
	.w2(32'h3c41e092),
	.w3(32'h3bfe9ad4),
	.w4(32'h3cb346c4),
	.w5(32'h3c2bfb06),
	.w6(32'h3c40c7ce),
	.w7(32'h3c8aead9),
	.w8(32'h3bd3d269),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07a668),
	.w1(32'hbbf1c486),
	.w2(32'hbc33e8a9),
	.w3(32'hbbe6a3ce),
	.w4(32'hbc771801),
	.w5(32'hbc3225cb),
	.w6(32'hbc40c678),
	.w7(32'hbc9f9ff7),
	.w8(32'hbc0ae7a7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e3465),
	.w1(32'hbbfd0024),
	.w2(32'h3b77ff69),
	.w3(32'h3b23a0e5),
	.w4(32'h3c650250),
	.w5(32'h3a734aa7),
	.w6(32'h3c645588),
	.w7(32'h3cb31b3b),
	.w8(32'hbb36c03e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39265da9),
	.w1(32'hbb9179b8),
	.w2(32'h3c56aa1f),
	.w3(32'hbb823741),
	.w4(32'hbc11d4ea),
	.w5(32'h3be670d1),
	.w6(32'hbc02a66b),
	.w7(32'hbc2959f9),
	.w8(32'h3b71b509),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98b275),
	.w1(32'hbc22d20b),
	.w2(32'hbbdd7e4b),
	.w3(32'hbb959151),
	.w4(32'hbcb3ffab),
	.w5(32'hbbfce057),
	.w6(32'hbc006551),
	.w7(32'hbcb97177),
	.w8(32'hbb3e0bea),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83bdfb),
	.w1(32'h3b740288),
	.w2(32'hbccf2bcf),
	.w3(32'h3c407caf),
	.w4(32'h3c369d96),
	.w5(32'hbc9e64c4),
	.w6(32'h3bbfb0c9),
	.w7(32'h3c094135),
	.w8(32'hbc02789e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2debdd),
	.w1(32'h3af7b213),
	.w2(32'h3b873a76),
	.w3(32'h3ad426b8),
	.w4(32'h3ca54b87),
	.w5(32'hbaad2668),
	.w6(32'h3c182a7f),
	.w7(32'h3c6f272a),
	.w8(32'hbbbb51b6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc584be8),
	.w1(32'hbca31646),
	.w2(32'h3b98fe73),
	.w3(32'hbcace315),
	.w4(32'hbd038456),
	.w5(32'hbc0fa836),
	.w6(32'hbce8235c),
	.w7(32'hbd1a8692),
	.w8(32'hbc70c2e6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95e7c7),
	.w1(32'h3c737aaf),
	.w2(32'h3848099e),
	.w3(32'hbb876ec9),
	.w4(32'h3c6917bd),
	.w5(32'h3a980b97),
	.w6(32'hbc26691c),
	.w7(32'h3bf9d9fd),
	.w8(32'hbb2e0a49),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50b959),
	.w1(32'h3be4062e),
	.w2(32'hbc051c09),
	.w3(32'h3b69ae3b),
	.w4(32'h3c041e40),
	.w5(32'hbc0c2434),
	.w6(32'h3a9cbfec),
	.w7(32'h3b856580),
	.w8(32'hbc33d3b6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab11712),
	.w1(32'h3a39b23c),
	.w2(32'hbb312243),
	.w3(32'h3ba1b4b0),
	.w4(32'h3c2859ba),
	.w5(32'h3bb74e92),
	.w6(32'h3a765090),
	.w7(32'hb9e3d16b),
	.w8(32'h3c3b626b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33e941),
	.w1(32'hbcb12b2a),
	.w2(32'hbc43edf0),
	.w3(32'hbc550a8f),
	.w4(32'hbcecc054),
	.w5(32'hbc67e250),
	.w6(32'h3a4a70af),
	.w7(32'hbc0fdf5a),
	.w8(32'hbc1b7474),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2e2a4),
	.w1(32'h3bd04485),
	.w2(32'hbd26ca02),
	.w3(32'hbaca3ccd),
	.w4(32'h3b220ed6),
	.w5(32'hbcf535a7),
	.w6(32'hba40fa86),
	.w7(32'h3baafde4),
	.w8(32'hbc9e29a0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98add1),
	.w1(32'h3d18dd15),
	.w2(32'hbc23f6e7),
	.w3(32'h3d281103),
	.w4(32'h3da9f73e),
	.w5(32'hbbf56fb4),
	.w6(32'h3d45628c),
	.w7(32'h3daf8ed8),
	.w8(32'hbc34b0f5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc290edf),
	.w1(32'hbb03c463),
	.w2(32'h3bb0e373),
	.w3(32'hbb883252),
	.w4(32'h3a5c5775),
	.w5(32'h3b5a46d1),
	.w6(32'hbb4ae98d),
	.w7(32'h3c39dcbd),
	.w8(32'hba6d212a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d4db6),
	.w1(32'h3c30ee33),
	.w2(32'hbbc1b785),
	.w3(32'hb965ebaf),
	.w4(32'h3bf5a3b5),
	.w5(32'hbbfd666f),
	.w6(32'hbbecbdbc),
	.w7(32'hbaf86be9),
	.w8(32'hbc0d5900),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abea80c),
	.w1(32'h3b2eecd1),
	.w2(32'h3a275a23),
	.w3(32'hbbb96c57),
	.w4(32'hbb3a6088),
	.w5(32'h3635815a),
	.w6(32'hbc70280a),
	.w7(32'hbc817198),
	.w8(32'h3b1dc43f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2757f4),
	.w1(32'hbb4fc079),
	.w2(32'h3a90593d),
	.w3(32'h3bf955ab),
	.w4(32'hbb9f7f1e),
	.w5(32'h3a16572a),
	.w6(32'h3b962774),
	.w7(32'hbb389bcd),
	.w8(32'hbba6d095),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d6c88),
	.w1(32'hbb13034b),
	.w2(32'hbb3c96f4),
	.w3(32'hbb3e2a24),
	.w4(32'h3ae6924d),
	.w5(32'h3a35470b),
	.w6(32'hbafb4595),
	.w7(32'h3a77153a),
	.w8(32'h3928c6fb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0f774),
	.w1(32'hba412a35),
	.w2(32'h3ae519ab),
	.w3(32'h3bf4ce6f),
	.w4(32'h3b0fc397),
	.w5(32'h3c6f4214),
	.w6(32'h3c073655),
	.w7(32'h3b64f9c4),
	.w8(32'h3c2383fb),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa30edd),
	.w1(32'h3ac84ed2),
	.w2(32'h3b05ca32),
	.w3(32'h3bf9c0f9),
	.w4(32'hbb904ed4),
	.w5(32'hba494555),
	.w6(32'h3b2b4591),
	.w7(32'hbc3de188),
	.w8(32'hbb233b28),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5e9e8),
	.w1(32'h39554aa8),
	.w2(32'hbb758f86),
	.w3(32'hbb8f02cc),
	.w4(32'hbc2291e4),
	.w5(32'hbbe9467e),
	.w6(32'hbc90aa43),
	.w7(32'hbc981a71),
	.w8(32'hbb7a4197),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a7dad),
	.w1(32'h3bd1983c),
	.w2(32'h3c11200d),
	.w3(32'h3c0b848d),
	.w4(32'h3c293366),
	.w5(32'h3c43aa0f),
	.w6(32'h3abafc2b),
	.w7(32'hbbaf6756),
	.w8(32'hbbbf2038),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48417e),
	.w1(32'h3c5ca129),
	.w2(32'hbb945428),
	.w3(32'h3c72ef78),
	.w4(32'h3c98fe96),
	.w5(32'hbaf1b11e),
	.w6(32'h3bab4959),
	.w7(32'h3c80e93b),
	.w8(32'hbab5f5bb),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c744e),
	.w1(32'hbb1027cd),
	.w2(32'hbb234b8c),
	.w3(32'h3bcaa9b4),
	.w4(32'hbadc3bf8),
	.w5(32'hba22f219),
	.w6(32'h3b28af3a),
	.w7(32'h3aa77ec2),
	.w8(32'hbabe9eae),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e196e),
	.w1(32'h3ba966c1),
	.w2(32'hb814a78b),
	.w3(32'h3b8fcce7),
	.w4(32'h3bee8687),
	.w5(32'hb87c67df),
	.w6(32'h3bbe08ab),
	.w7(32'h3bb3275b),
	.w8(32'hbb7cc880),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52dfa),
	.w1(32'h3bfbd55c),
	.w2(32'h3b1b214d),
	.w3(32'h3b2114d6),
	.w4(32'h3b8c90a7),
	.w5(32'hbc5604f7),
	.w6(32'h3adf6a30),
	.w7(32'h3bb0db0a),
	.w8(32'hbbf2ec45),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb67d12),
	.w1(32'hbb29e969),
	.w2(32'hbc17ed50),
	.w3(32'hbb9f7aa1),
	.w4(32'hbb67efb1),
	.w5(32'hbc492dd7),
	.w6(32'hbc798af9),
	.w7(32'hbc5af061),
	.w8(32'hbc52d57f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae94a0e),
	.w1(32'h3c1ea9e6),
	.w2(32'hba63c47b),
	.w3(32'h3b9be9fd),
	.w4(32'h3c5e5770),
	.w5(32'hbc55ff4b),
	.w6(32'hbba3e9fc),
	.w7(32'hbb65f66c),
	.w8(32'hbc86cf4a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14aee2),
	.w1(32'hbc83b16d),
	.w2(32'h3b268d08),
	.w3(32'hbc9a208b),
	.w4(32'hbcc1cb27),
	.w5(32'h3b425908),
	.w6(32'hbcb7ae84),
	.w7(32'hbcd4d508),
	.w8(32'hbb1e09e6),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02cab0),
	.w1(32'h3b8951fc),
	.w2(32'h3aecd717),
	.w3(32'h3bf2a7fb),
	.w4(32'h3ba3af74),
	.w5(32'hbb30e66a),
	.w6(32'h3b6bdd6d),
	.w7(32'h3a8095b2),
	.w8(32'hba9e87a7),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae77d56),
	.w1(32'h392d1cc9),
	.w2(32'hbca6788b),
	.w3(32'hbba5bf6f),
	.w4(32'hbc131b32),
	.w5(32'hbc9f9259),
	.w6(32'hbbe249d4),
	.w7(32'hbc274d18),
	.w8(32'hbcaa957a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02dbd1),
	.w1(32'h394b86b9),
	.w2(32'hbc5a4287),
	.w3(32'h3b00976d),
	.w4(32'h3c43240e),
	.w5(32'hbb97e1ed),
	.w6(32'h3bdcdac0),
	.w7(32'h3c3b5f57),
	.w8(32'hbbbb4f05),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58200e),
	.w1(32'hbbd8762c),
	.w2(32'hbcbaf5ed),
	.w3(32'hbc42663a),
	.w4(32'hbc8cc1e1),
	.w5(32'hbc8d0e0c),
	.w6(32'hb9fe634f),
	.w7(32'hbb55ef36),
	.w8(32'hbbe56941),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e3bd6),
	.w1(32'h3c3c697e),
	.w2(32'hbb9e52e3),
	.w3(32'h3c878b84),
	.w4(32'h3d138645),
	.w5(32'hbb645b6d),
	.w6(32'h3ca79bd2),
	.w7(32'h3cf89798),
	.w8(32'hb9135f9b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c35b6),
	.w1(32'h3c445a3a),
	.w2(32'h3c79611b),
	.w3(32'hba1f1265),
	.w4(32'h3c37c6eb),
	.w5(32'h3c95de0d),
	.w6(32'h3bc02662),
	.w7(32'h3bfbf46d),
	.w8(32'h3afdb7f2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c643930),
	.w1(32'hbb1a9831),
	.w2(32'hbbbb3215),
	.w3(32'hbc03fef7),
	.w4(32'hbcad363b),
	.w5(32'hbc17becb),
	.w6(32'hbc2a0c18),
	.w7(32'hbc4067c9),
	.w8(32'hbc20b397),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a56c3),
	.w1(32'hbc0e8407),
	.w2(32'hbc2876ba),
	.w3(32'hba8117de),
	.w4(32'hbbb93858),
	.w5(32'hbc11a181),
	.w6(32'h3b030f73),
	.w7(32'hbb9a1c35),
	.w8(32'hbb04b223),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89a818),
	.w1(32'h3bbaf7b2),
	.w2(32'hbb893010),
	.w3(32'h3c1b9b08),
	.w4(32'h3c7d2712),
	.w5(32'hbc2811d7),
	.w6(32'h3bfbe579),
	.w7(32'h3c98dcec),
	.w8(32'hbc60b175),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f4d29),
	.w1(32'hbb003376),
	.w2(32'h3bcf8328),
	.w3(32'hbabe4017),
	.w4(32'h3c1bf7c3),
	.w5(32'h3b55243e),
	.w6(32'h3a9780f2),
	.w7(32'h3befa034),
	.w8(32'h3b9e6fe3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77733e),
	.w1(32'hbbc3fd24),
	.w2(32'h3b79dc13),
	.w3(32'h3ba7ca07),
	.w4(32'hbb9b91a2),
	.w5(32'h39c486c9),
	.w6(32'h3b9a14fe),
	.w7(32'h3a4eb47a),
	.w8(32'hbbb32557),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88837af),
	.w1(32'hbbcdb830),
	.w2(32'h3c8758f9),
	.w3(32'hbb65caf2),
	.w4(32'hbc26fffd),
	.w5(32'h3c8d1f80),
	.w6(32'hbba34075),
	.w7(32'hbc15f72b),
	.w8(32'h3c16996f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e1895),
	.w1(32'h3aa17eae),
	.w2(32'h3be11eeb),
	.w3(32'h3c83b45d),
	.w4(32'hbbc20bd3),
	.w5(32'h3ba1f018),
	.w6(32'h3b41038e),
	.w7(32'hbc4d3f3e),
	.w8(32'h3b97388e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba09a53),
	.w1(32'h3b4c8abb),
	.w2(32'h3b93b697),
	.w3(32'h3c04fd09),
	.w4(32'h3bedbdd0),
	.w5(32'h3a65dd18),
	.w6(32'h3bec0fcb),
	.w7(32'h3c08a336),
	.w8(32'hbb62bbde),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14a2fa),
	.w1(32'h3c552c36),
	.w2(32'h3b93cea4),
	.w3(32'hb99d7d56),
	.w4(32'h3c597377),
	.w5(32'h3b872e1c),
	.w6(32'hbb39b911),
	.w7(32'h3c404901),
	.w8(32'h3c3da787),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1351a0),
	.w1(32'hbba441bd),
	.w2(32'hbb043166),
	.w3(32'h3b409e57),
	.w4(32'hbc1202cf),
	.w5(32'h3b0301a4),
	.w6(32'h3b875988),
	.w7(32'hbb2062fe),
	.w8(32'h3a94ba11),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c075186),
	.w1(32'h3c65f1d7),
	.w2(32'h3b6f0064),
	.w3(32'h3c21d87c),
	.w4(32'h3c39c46d),
	.w5(32'hb8bb7636),
	.w6(32'h3c33b115),
	.w7(32'h3bbc011c),
	.w8(32'h3ba9d130),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec868a),
	.w1(32'h3b557c19),
	.w2(32'h3853bbe2),
	.w3(32'hbc152194),
	.w4(32'hbc3c5f3c),
	.w5(32'hbbc4da8e),
	.w6(32'hbc0739de),
	.w7(32'hbc01db8b),
	.w8(32'h3be8f431),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39771ec4),
	.w1(32'h3c123bb8),
	.w2(32'h3c66a716),
	.w3(32'h3bbaf966),
	.w4(32'h3c27e27c),
	.w5(32'h3c9e12a5),
	.w6(32'h3c4d6106),
	.w7(32'h3c240614),
	.w8(32'h3c46d6f3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a228f),
	.w1(32'hbc28353a),
	.w2(32'hbc3c5f88),
	.w3(32'hbb9d3d65),
	.w4(32'hbd025312),
	.w5(32'hbc5a90df),
	.w6(32'hbc878b64),
	.w7(32'hbcd2cd2f),
	.w8(32'hbc59b69b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf90acd),
	.w1(32'hbbc3931e),
	.w2(32'h3c07794f),
	.w3(32'hbba7b0ac),
	.w4(32'hbc0bff29),
	.w5(32'h3c138891),
	.w6(32'hbc5b0be3),
	.w7(32'hbca9e31d),
	.w8(32'h3c4bb149),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8e1d4),
	.w1(32'h3ad2da3a),
	.w2(32'hbc95a920),
	.w3(32'hba94e7b5),
	.w4(32'hbbd511d5),
	.w5(32'hbcafac1b),
	.w6(32'hbb9d72de),
	.w7(32'hbc01ff49),
	.w8(32'hbc89c1b2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b0cd7),
	.w1(32'hbc7c6049),
	.w2(32'h3a14be67),
	.w3(32'hbcc52963),
	.w4(32'hbcb67db9),
	.w5(32'hbaaca995),
	.w6(32'hbca0591d),
	.w7(32'hbc3c0cd9),
	.w8(32'h3acead88),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28d862),
	.w1(32'h3a37a78c),
	.w2(32'h3b169b51),
	.w3(32'hbb101f93),
	.w4(32'hbadf12a5),
	.w5(32'hbb2c12e7),
	.w6(32'hbb147b15),
	.w7(32'hbaf776a5),
	.w8(32'hbb99e0a4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad11b56),
	.w1(32'hbbac756b),
	.w2(32'hbb580eb7),
	.w3(32'h3b2ceabb),
	.w4(32'hbbb042c2),
	.w5(32'hba6eba94),
	.w6(32'h3bf83246),
	.w7(32'h3b99ad5c),
	.w8(32'h3bc708bd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67d25d),
	.w1(32'hbb8171af),
	.w2(32'h3c9eb682),
	.w3(32'h3b795d3d),
	.w4(32'h3b86ad5d),
	.w5(32'h3c52927a),
	.w6(32'h3ba9cd65),
	.w7(32'h3b1f65ec),
	.w8(32'h3c0c17e2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97d2d0),
	.w1(32'h3bed7602),
	.w2(32'hbc82da5b),
	.w3(32'h3c5911f5),
	.w4(32'hbb8e5875),
	.w5(32'hbc559764),
	.w6(32'h3b92f29d),
	.w7(32'h3a9310e9),
	.w8(32'hbc5c1f58),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb897dd9),
	.w1(32'h3af44fd6),
	.w2(32'hbc891789),
	.w3(32'h3bf5652f),
	.w4(32'h3c894f77),
	.w5(32'hbc4ae18f),
	.w6(32'h3c1588a0),
	.w7(32'h3c9ab843),
	.w8(32'hbc1057bc),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bb90a),
	.w1(32'h3b8cb02c),
	.w2(32'hbab90b8c),
	.w3(32'h3c708845),
	.w4(32'h3cda50bf),
	.w5(32'hbb5e76ce),
	.w6(32'h3c84c3a6),
	.w7(32'h3cec1cc5),
	.w8(32'hbba95b39),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ac637),
	.w1(32'hbb449537),
	.w2(32'hbc260a46),
	.w3(32'hbbc8d90e),
	.w4(32'hbbb7c1db),
	.w5(32'hbc151d43),
	.w6(32'hbc13bc6e),
	.w7(32'hbbb47953),
	.w8(32'hbc125078),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bd165),
	.w1(32'h3bffc0ac),
	.w2(32'hbc80aeab),
	.w3(32'h3b6c68ef),
	.w4(32'h3c5c7e5e),
	.w5(32'hbcb8f595),
	.w6(32'h3b1ef8a3),
	.w7(32'h3c480fdb),
	.w8(32'hbcb751bc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb541aa),
	.w1(32'hbc93b023),
	.w2(32'hb6e47181),
	.w3(32'hbcbd8d9f),
	.w4(32'hbcc21207),
	.w5(32'h3a55d2d8),
	.w6(32'hbcc058f5),
	.w7(32'hbca9e1d6),
	.w8(32'h3b8e436f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba6abe),
	.w1(32'hbab0ff38),
	.w2(32'h3bfcd22a),
	.w3(32'h3acd1693),
	.w4(32'h3a8c217b),
	.w5(32'h3bf9122c),
	.w6(32'h3bb1c623),
	.w7(32'h3b29d161),
	.w8(32'h3be4d880),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f8537),
	.w1(32'hb947bc21),
	.w2(32'hbb88d74a),
	.w3(32'h3aa749de),
	.w4(32'hbc34033c),
	.w5(32'hbb9f7b75),
	.w6(32'hbbfd4de5),
	.w7(32'hbc5205d7),
	.w8(32'h3ba8ea15),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81c2ec),
	.w1(32'h3b38bbe9),
	.w2(32'hbae7143f),
	.w3(32'h3b1685ac),
	.w4(32'hbc2b7f1d),
	.w5(32'hbb0885f7),
	.w6(32'hbb985d2a),
	.w7(32'hbc8a16fa),
	.w8(32'hbbbd3fba),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33e93d),
	.w1(32'h3bc14ed2),
	.w2(32'h3bad51d8),
	.w3(32'h3c5eb5ca),
	.w4(32'h3c82aeab),
	.w5(32'h3c638da3),
	.w6(32'h3b9ab31c),
	.w7(32'h3b4c6044),
	.w8(32'h3c1a93cd),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule