module layer_8_featuremap_248(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba61f7),
	.w1(32'hbbada56b),
	.w2(32'h3b40a40d),
	.w3(32'h3c5ce49f),
	.w4(32'hbb44e8c4),
	.w5(32'h3b386ed0),
	.w6(32'hbbda2f4a),
	.w7(32'hb9b78080),
	.w8(32'h3c3e4c7b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b942e47),
	.w1(32'hbb7c6406),
	.w2(32'hbb009d26),
	.w3(32'h3b39445c),
	.w4(32'hbad8909b),
	.w5(32'hba874ddf),
	.w6(32'hbb75d95b),
	.w7(32'hbb12e8c8),
	.w8(32'hba9d62c3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a3524),
	.w1(32'hbaac90be),
	.w2(32'hbbe58223),
	.w3(32'h3a5ff298),
	.w4(32'hbbb8d424),
	.w5(32'hbbd738e6),
	.w6(32'hbbd8cce9),
	.w7(32'hbbc34f5b),
	.w8(32'hbb45aeed),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a98b6),
	.w1(32'h3b2f44ea),
	.w2(32'h3b902d69),
	.w3(32'h3a904eb2),
	.w4(32'h3b2261e3),
	.w5(32'hbbdafbd4),
	.w6(32'hbbcc8aa9),
	.w7(32'hbac1bdf1),
	.w8(32'h3b210519),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68a351),
	.w1(32'h3abe68e4),
	.w2(32'h3b76ced0),
	.w3(32'hbc47d8a1),
	.w4(32'h3b2642ac),
	.w5(32'h3b365474),
	.w6(32'hba581818),
	.w7(32'h3a8fc8cb),
	.w8(32'hba106cfb),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9aaa7),
	.w1(32'h3c042cc4),
	.w2(32'hbcbbe654),
	.w3(32'hbb471425),
	.w4(32'h3bb739ee),
	.w5(32'hbcf94217),
	.w6(32'h3c484295),
	.w7(32'hbc491ce7),
	.w8(32'hbd05989f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3146a8),
	.w1(32'hba96ce88),
	.w2(32'hbaf0324f),
	.w3(32'hbcd794b6),
	.w4(32'hbb80ae82),
	.w5(32'hbb7748b6),
	.w6(32'hbb22c991),
	.w7(32'hbb06da56),
	.w8(32'hbb8f3cf8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b91c4),
	.w1(32'hbc029f5b),
	.w2(32'hbb42a4c5),
	.w3(32'hbc05a21e),
	.w4(32'hbbb3c348),
	.w5(32'hbb19dc98),
	.w6(32'hbb74106d),
	.w7(32'hbc044f39),
	.w8(32'hb9d28bc4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4118f8),
	.w1(32'h3b262ea0),
	.w2(32'h3b6e64cd),
	.w3(32'hb8c269d5),
	.w4(32'h3b80ee34),
	.w5(32'h3b1f8227),
	.w6(32'hbb697758),
	.w7(32'hbacfd531),
	.w8(32'hbbcb48be),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5856f),
	.w1(32'hbb5cd830),
	.w2(32'hbc0b1be6),
	.w3(32'hbc1bb605),
	.w4(32'hbafda9b1),
	.w5(32'hbb1fdd65),
	.w6(32'hbc21a211),
	.w7(32'hbbe8ccd8),
	.w8(32'h3b858028),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6badb),
	.w1(32'hbaa8c543),
	.w2(32'h3b7f47fa),
	.w3(32'h3c89b275),
	.w4(32'hbbebf285),
	.w5(32'hbb180bc6),
	.w6(32'hbb7e3fa5),
	.w7(32'h3b4493e6),
	.w8(32'h3c308d6c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96aa4b),
	.w1(32'h3b1f6328),
	.w2(32'h39d3681c),
	.w3(32'h3c4057a7),
	.w4(32'hbb972771),
	.w5(32'hbb9daef6),
	.w6(32'h3aca2bbf),
	.w7(32'h3b89cec5),
	.w8(32'h3bf6d600),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e9e1d),
	.w1(32'h3b6cdbec),
	.w2(32'hbb3e2752),
	.w3(32'h3ba37d1c),
	.w4(32'hbb6b73dc),
	.w5(32'hbae6741e),
	.w6(32'hba0f5686),
	.w7(32'hb94c532a),
	.w8(32'h39fc7f48),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be22d96),
	.w1(32'hbaa90e65),
	.w2(32'h3b839288),
	.w3(32'h39ea8c34),
	.w4(32'hb89b8041),
	.w5(32'hbbf23f35),
	.w6(32'hbb94886c),
	.w7(32'hba3fd22b),
	.w8(32'h3a831221),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba735fc),
	.w1(32'h3bae44fa),
	.w2(32'h3b26d9e7),
	.w3(32'hbb836d92),
	.w4(32'h3b664a57),
	.w5(32'h3aa365d1),
	.w6(32'h3b144d8b),
	.w7(32'h3b0443e9),
	.w8(32'hbac6d34d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86c7a6),
	.w1(32'hbbcd767f),
	.w2(32'h3bae09fc),
	.w3(32'hbb6523af),
	.w4(32'hbbb144eb),
	.w5(32'h3b0325ed),
	.w6(32'h39dabeb7),
	.w7(32'h3a513966),
	.w8(32'h3a39fdd2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1ce36),
	.w1(32'h3b625de9),
	.w2(32'hbb6a7a63),
	.w3(32'hbbb908f0),
	.w4(32'h39893a81),
	.w5(32'h3c28e2e4),
	.w6(32'h3c239903),
	.w7(32'h38ac189d),
	.w8(32'h3b9dff84),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2e565),
	.w1(32'hbb6218c1),
	.w2(32'hbb5c871f),
	.w3(32'hba6b1b66),
	.w4(32'hbb823025),
	.w5(32'hbbf448eb),
	.w6(32'hbc7b41c2),
	.w7(32'hbb89585d),
	.w8(32'hba9b5ec9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe543e2),
	.w1(32'hbb88bf05),
	.w2(32'hbcd30f9f),
	.w3(32'hbbbd136d),
	.w4(32'hbbe63ab3),
	.w5(32'hbcd0701e),
	.w6(32'hbaf76f1d),
	.w7(32'hbc718834),
	.w8(32'hbc7fdf7e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd15a6),
	.w1(32'hbbb96c6e),
	.w2(32'hbb6531f9),
	.w3(32'hbc694544),
	.w4(32'hba9c39fc),
	.w5(32'hb9b2c203),
	.w6(32'hbb6c3b07),
	.w7(32'hbad05e7c),
	.w8(32'hbb81d8ef),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa841c),
	.w1(32'h3be3acb6),
	.w2(32'h3c1c08e8),
	.w3(32'hbaf08cb1),
	.w4(32'h3b651eae),
	.w5(32'h3c17914e),
	.w6(32'h3b41f92d),
	.w7(32'h3b4c93ba),
	.w8(32'hbb3058a9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae44ba),
	.w1(32'hbbfd13c0),
	.w2(32'hbc08a7c4),
	.w3(32'hbb539454),
	.w4(32'hbb0fea5e),
	.w5(32'hbb8cd90d),
	.w6(32'hbbec8664),
	.w7(32'hba5b4082),
	.w8(32'hbc4527a0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc652b76),
	.w1(32'hbc728b7f),
	.w2(32'hbc362a9a),
	.w3(32'hbb0ca37d),
	.w4(32'hbbdfdbb2),
	.w5(32'h3b38ebd4),
	.w6(32'hbc9be486),
	.w7(32'hbc207c0e),
	.w8(32'h3b5c3002),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc84931),
	.w1(32'h3b1e0f85),
	.w2(32'h38c52266),
	.w3(32'h3cbb72fe),
	.w4(32'hbb748182),
	.w5(32'hba7f4822),
	.w6(32'h3b925771),
	.w7(32'h3b389ffc),
	.w8(32'hbc4533ca),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e0ef5),
	.w1(32'hbb2da191),
	.w2(32'hbc01d00b),
	.w3(32'h3b517837),
	.w4(32'hba756086),
	.w5(32'hb9d8c7a3),
	.w6(32'hbb9ecbdc),
	.w7(32'hbc1e69cd),
	.w8(32'hbc0fc426),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47553d),
	.w1(32'h3b631b77),
	.w2(32'h3c21f402),
	.w3(32'hbadafad0),
	.w4(32'h3c575ff3),
	.w5(32'h3c58c900),
	.w6(32'h3b658546),
	.w7(32'h3bd6932e),
	.w8(32'h3ba06fdd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897bd3),
	.w1(32'h3bdbf15f),
	.w2(32'h3c66ce38),
	.w3(32'h3ab6aaf5),
	.w4(32'h3c0187a3),
	.w5(32'h3c371578),
	.w6(32'h3bc9a328),
	.w7(32'h3bffc9f2),
	.w8(32'h3c2af5cf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cb8a5),
	.w1(32'hbbcd3443),
	.w2(32'hbd146e06),
	.w3(32'h3c8988ad),
	.w4(32'h3a7f04eb),
	.w5(32'hbcb666c8),
	.w6(32'h3b0e3faf),
	.w7(32'hbcb4a174),
	.w8(32'hbd055a22),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2aec9f),
	.w1(32'h3a1cac8f),
	.w2(32'h3c58f036),
	.w3(32'hbce10746),
	.w4(32'h3bdcfc8b),
	.w5(32'h3c765694),
	.w6(32'hbbee6477),
	.w7(32'h3ba8d1c4),
	.w8(32'h3bcce146),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c932d6f),
	.w1(32'hbb12fc80),
	.w2(32'h38eb02f7),
	.w3(32'h3c73882c),
	.w4(32'h3afd74c9),
	.w5(32'h3bf9d0c5),
	.w6(32'hbbaee697),
	.w7(32'hbb867319),
	.w8(32'h3b993d37),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd96e0c),
	.w1(32'hbaa3661b),
	.w2(32'h3b8b4f12),
	.w3(32'h3c708e4f),
	.w4(32'h3b25aa4c),
	.w5(32'h3b99fe04),
	.w6(32'hbbbc1045),
	.w7(32'h39b6e574),
	.w8(32'hbba2a784),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae88ed),
	.w1(32'hbcea03bc),
	.w2(32'hbd035798),
	.w3(32'hbb268f12),
	.w4(32'hbcb3658f),
	.w5(32'hbcd9473f),
	.w6(32'hbc45c9f5),
	.w7(32'hbc9bf1d5),
	.w8(32'h3b36de2f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb1d82),
	.w1(32'hbbb0877f),
	.w2(32'h3ca89f5a),
	.w3(32'h3bf83dfd),
	.w4(32'hba438f1c),
	.w5(32'h3caa8361),
	.w6(32'hbb788ac1),
	.w7(32'h3bdb9da9),
	.w8(32'h3c90dac1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf7debe),
	.w1(32'h3c00fef4),
	.w2(32'h3c2acd46),
	.w3(32'h3c6a340e),
	.w4(32'h3bca0487),
	.w5(32'h3bfd37ee),
	.w6(32'h3bddb4d9),
	.w7(32'h3b6b0036),
	.w8(32'h3be21e1f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf9dad),
	.w1(32'hb9f0d805),
	.w2(32'h3bfa398a),
	.w3(32'hbb5348bf),
	.w4(32'hbbbf2796),
	.w5(32'h3b95fea0),
	.w6(32'hbbce3992),
	.w7(32'h3af99af6),
	.w8(32'hbb4c267f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e0548),
	.w1(32'h39fd9685),
	.w2(32'hbbc920a8),
	.w3(32'h3b5a3bf0),
	.w4(32'hba9baa37),
	.w5(32'hbb7f8a89),
	.w6(32'hba20ba13),
	.w7(32'h3b8d28e6),
	.w8(32'hb9414809),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc545e25),
	.w1(32'h388a16ac),
	.w2(32'h3bcd1fce),
	.w3(32'hbb9fc348),
	.w4(32'hbb0df445),
	.w5(32'h3bbdab3b),
	.w6(32'hbb844db5),
	.w7(32'h3ada016f),
	.w8(32'h3b62929a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be35a69),
	.w1(32'h3bbfe3f9),
	.w2(32'h3b48cdbb),
	.w3(32'h3bb085b8),
	.w4(32'h3b84d65f),
	.w5(32'h3a348a1f),
	.w6(32'hbacfa423),
	.w7(32'hbab22f0b),
	.w8(32'hbbe1330e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84136f),
	.w1(32'h3bd4aa14),
	.w2(32'h3c0c852c),
	.w3(32'hbbc4ad25),
	.w4(32'h3b9fe7c0),
	.w5(32'h3b99e02d),
	.w6(32'hbb02554b),
	.w7(32'h3a7fdf75),
	.w8(32'h395f8f5d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa444b),
	.w1(32'h3c070327),
	.w2(32'h3c27aee7),
	.w3(32'h3ba9d980),
	.w4(32'h3b9aec56),
	.w5(32'h3afeda5c),
	.w6(32'h3b34eb6b),
	.w7(32'h3b3f64cd),
	.w8(32'h3b137d7c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3c891),
	.w1(32'h3a407212),
	.w2(32'h3a74f3cb),
	.w3(32'h3a064c08),
	.w4(32'hba45c58b),
	.w5(32'h3a273908),
	.w6(32'hbb0133cc),
	.w7(32'hbb65f036),
	.w8(32'hbb78cf92),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76c810),
	.w1(32'h3c655706),
	.w2(32'hbcb557fb),
	.w3(32'h3b4c9248),
	.w4(32'h3c43be9d),
	.w5(32'hbcab3b4b),
	.w6(32'h3c6e80ec),
	.w7(32'hbc8baf3f),
	.w8(32'hbc5e353f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf42ab),
	.w1(32'h3aa067ef),
	.w2(32'h3c2a4183),
	.w3(32'hbc6fa137),
	.w4(32'h3bc0583b),
	.w5(32'h3c75c83d),
	.w6(32'hbbd74590),
	.w7(32'h39d84b46),
	.w8(32'h3c5578aa),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0c8cd),
	.w1(32'hbbf3e667),
	.w2(32'hbc32b31a),
	.w3(32'h3c9aa641),
	.w4(32'hbb4a7a5b),
	.w5(32'hbbe32d7b),
	.w6(32'hbac7fa17),
	.w7(32'hbc0cb771),
	.w8(32'hb9e4e5c8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b759359),
	.w1(32'hbb001047),
	.w2(32'h399c6244),
	.w3(32'h3a6f6af7),
	.w4(32'h3ac3cc51),
	.w5(32'h3b82284e),
	.w6(32'hbbce96b4),
	.w7(32'h3bcde0a5),
	.w8(32'hbba0213f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7e93d),
	.w1(32'h3b3aa9a2),
	.w2(32'hb9d8c977),
	.w3(32'hbb9a4c90),
	.w4(32'h3ba14a6c),
	.w5(32'h3a9aa3dc),
	.w6(32'h3b464111),
	.w7(32'h3b1a636b),
	.w8(32'h399d59d9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa239f),
	.w1(32'h38dd825f),
	.w2(32'h3aad916e),
	.w3(32'hbb34e7f8),
	.w4(32'hbb447f10),
	.w5(32'hbb8c60c8),
	.w6(32'hbb1c308b),
	.w7(32'hba638df7),
	.w8(32'hbb0e0636),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf75b2),
	.w1(32'h3c086d63),
	.w2(32'h3b4bccdf),
	.w3(32'hbbe91e9b),
	.w4(32'h3bab22ac),
	.w5(32'h3a56fa96),
	.w6(32'h3b817733),
	.w7(32'h3c26219d),
	.w8(32'hbb87ddf6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc304b0),
	.w1(32'h3be43212),
	.w2(32'hbb242fad),
	.w3(32'h3b9aef6d),
	.w4(32'hbbb5336d),
	.w5(32'hbc339d77),
	.w6(32'h3bb9429a),
	.w7(32'hbabfcb15),
	.w8(32'hbb0b3711),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc493ddd),
	.w1(32'h3c5b3160),
	.w2(32'hbc3da847),
	.w3(32'hbacbb900),
	.w4(32'h3bb88ec9),
	.w5(32'hbc10e2af),
	.w6(32'h3bf554ec),
	.w7(32'hbc140367),
	.w8(32'hbcad5a9b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1f2f54),
	.w1(32'h3bd84fec),
	.w2(32'h3bbef4cc),
	.w3(32'hbcfd8925),
	.w4(32'hbaa58a28),
	.w5(32'hbabce476),
	.w6(32'hbb4408ff),
	.w7(32'hba0df63c),
	.w8(32'h39847478),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7fb9e),
	.w1(32'hbc80e03e),
	.w2(32'hbc6d5e6d),
	.w3(32'hba1ab54c),
	.w4(32'hbc3c57e9),
	.w5(32'hbc4403bf),
	.w6(32'hbc068d4e),
	.w7(32'hbc11746e),
	.w8(32'hbc7ae4e3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94b140),
	.w1(32'hbb1d6728),
	.w2(32'hbb8f5b52),
	.w3(32'hbc6b1b80),
	.w4(32'hbb4082d6),
	.w5(32'hbb89943e),
	.w6(32'hbb693315),
	.w7(32'hbb154c7e),
	.w8(32'hbb973339),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f0b18),
	.w1(32'hba0020ee),
	.w2(32'hbba95ae8),
	.w3(32'hbb00edd7),
	.w4(32'hbbde6960),
	.w5(32'hbacd6067),
	.w6(32'h3ab09fbd),
	.w7(32'h3b194559),
	.w8(32'hbc0ff752),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3607c),
	.w1(32'hbb8f30c4),
	.w2(32'h3d0ebe8d),
	.w3(32'h3b2d5e79),
	.w4(32'h3b38c375),
	.w5(32'h3d0bb3b6),
	.w6(32'hbc404dc6),
	.w7(32'h3c2cf8e2),
	.w8(32'h3cc27b55),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d27b0ba),
	.w1(32'h387c4bbc),
	.w2(32'h3b390de5),
	.w3(32'h3d01936b),
	.w4(32'hbaad2b76),
	.w5(32'h3821ee7d),
	.w6(32'hbaff0dc7),
	.w7(32'h3b1161b3),
	.w8(32'h3b43e42a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb631aab),
	.w1(32'h3bf271a4),
	.w2(32'hbbff2694),
	.w3(32'hbb16c414),
	.w4(32'hbb8a0752),
	.w5(32'hbb6ab997),
	.w6(32'h3c0ba250),
	.w7(32'hba9c90a6),
	.w8(32'hbc2fbacb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d56f9),
	.w1(32'h3b4828d1),
	.w2(32'h3b8bf5f0),
	.w3(32'h3b1018eb),
	.w4(32'h3bbadb12),
	.w5(32'h3c2dbd04),
	.w6(32'hbb05f1d9),
	.w7(32'h3ac0124a),
	.w8(32'h3c2734d8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c602480),
	.w1(32'h3b2d7b28),
	.w2(32'hbb37f7bb),
	.w3(32'h3c941cc6),
	.w4(32'h3a63081d),
	.w5(32'hbaf24045),
	.w6(32'h3aa760bd),
	.w7(32'hbb481cd3),
	.w8(32'hbbb0bd18),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc460),
	.w1(32'hbbdd8f35),
	.w2(32'h3bdcde38),
	.w3(32'hbba2229f),
	.w4(32'hbac23f16),
	.w5(32'h3c2003bc),
	.w6(32'hbbc9c6a6),
	.w7(32'hbafe7a8a),
	.w8(32'h3ad98e35),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb3065),
	.w1(32'hb932d560),
	.w2(32'hbc1ba428),
	.w3(32'hb9acdcba),
	.w4(32'hbbb29002),
	.w5(32'hbc4e4241),
	.w6(32'h3adbb38f),
	.w7(32'hbb8b2b2e),
	.w8(32'hbb9946f6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc222e42),
	.w1(32'h3b5602c6),
	.w2(32'hba9f2df8),
	.w3(32'hbb9a90be),
	.w4(32'hbb469f94),
	.w5(32'hb98883c7),
	.w6(32'hbb54c48a),
	.w7(32'h3ad974de),
	.w8(32'hba6a85eb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc364a9b),
	.w1(32'hbbc8f50b),
	.w2(32'hbbced9ab),
	.w3(32'hbb1a2caf),
	.w4(32'hb9cf3446),
	.w5(32'h3b809ea2),
	.w6(32'hbb964c2f),
	.w7(32'h388cc1c7),
	.w8(32'hbb256c7d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12392b),
	.w1(32'h3c028561),
	.w2(32'h3c0309e3),
	.w3(32'h3ac30404),
	.w4(32'h3bfe9c9b),
	.w5(32'h3c1136fe),
	.w6(32'h3b14d6a3),
	.w7(32'h3b5d3400),
	.w8(32'h3ad8ed69),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7de04),
	.w1(32'hbba70579),
	.w2(32'hbbcdd675),
	.w3(32'h3bbffc5a),
	.w4(32'hbb9c56f9),
	.w5(32'hbb9122c0),
	.w6(32'hbbb7200c),
	.w7(32'hbbdf0b35),
	.w8(32'hbba1261c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba633d06),
	.w1(32'h3b7dd297),
	.w2(32'h3c43f669),
	.w3(32'hbb037a67),
	.w4(32'h3bbb1cca),
	.w5(32'h3bde2ca5),
	.w6(32'h3b327eee),
	.w7(32'h3c19df0d),
	.w8(32'h3b608c19),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2275e2),
	.w1(32'hbb999e62),
	.w2(32'h3c80f8ec),
	.w3(32'hbadaeb5e),
	.w4(32'hbb90881b),
	.w5(32'h3c099df4),
	.w6(32'hbb30e6e1),
	.w7(32'h3c376c6a),
	.w8(32'h3c11ecd4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdc7b1),
	.w1(32'h3bcf1669),
	.w2(32'h3c3fe239),
	.w3(32'h3c666cf3),
	.w4(32'h3bc43ed6),
	.w5(32'h3a094968),
	.w6(32'hb9f2be5f),
	.w7(32'h3b9311d4),
	.w8(32'h3af6d142),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb771670),
	.w1(32'hbbab2bfb),
	.w2(32'hbc193bc1),
	.w3(32'h3a7c7def),
	.w4(32'hbbfe9401),
	.w5(32'hbbb8866a),
	.w6(32'hbc04af1f),
	.w7(32'hbaae2e61),
	.w8(32'h3bf7f2e9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904a36e),
	.w1(32'hbc17ad03),
	.w2(32'hbb5e38bd),
	.w3(32'hbb82afbb),
	.w4(32'hbc55f3e0),
	.w5(32'hbc3c7662),
	.w6(32'hbc4cb643),
	.w7(32'hbc145b3c),
	.w8(32'hbc7053bd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e67b6),
	.w1(32'h3bf030f2),
	.w2(32'hbc17a4e9),
	.w3(32'hbc6f0d6f),
	.w4(32'h3b902f3d),
	.w5(32'hbc576cb6),
	.w6(32'h3be44b8e),
	.w7(32'hbbe86c04),
	.w8(32'hbc63b5ba),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0f9f4),
	.w1(32'h3b2d97bd),
	.w2(32'hbb15aa28),
	.w3(32'hbcb37671),
	.w4(32'h3b3470e5),
	.w5(32'h3aa06343),
	.w6(32'h3b967062),
	.w7(32'h3c1c5e13),
	.w8(32'h3bcecc8f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3737),
	.w1(32'hbb6a5dbe),
	.w2(32'h3a861bf7),
	.w3(32'h3b94ea48),
	.w4(32'h3bc41557),
	.w5(32'hbb7e9ad8),
	.w6(32'h3b1d7134),
	.w7(32'h3bd0732e),
	.w8(32'h3c031437),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5cad),
	.w1(32'hbb74c1c0),
	.w2(32'hbb853512),
	.w3(32'hbb93864e),
	.w4(32'hbaf7703d),
	.w5(32'hbbf8db66),
	.w6(32'hbc075287),
	.w7(32'hbb9868df),
	.w8(32'hbb53e20c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb620b7c),
	.w1(32'hba939308),
	.w2(32'hbcd7b057),
	.w3(32'hbb4e137a),
	.w4(32'hbb3ae22f),
	.w5(32'hbcb63542),
	.w6(32'h3ba83d02),
	.w7(32'hbc82ee23),
	.w8(32'hbc7acb2f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb5d50),
	.w1(32'h3b2b848f),
	.w2(32'hbb38e942),
	.w3(32'hbc955fd5),
	.w4(32'h3b1f4be2),
	.w5(32'h3beba95d),
	.w6(32'hbab7c911),
	.w7(32'h39845f98),
	.w8(32'h3b80a25f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60e073),
	.w1(32'h3b7dde55),
	.w2(32'h3b6ec3a8),
	.w3(32'h3c847b2b),
	.w4(32'h3bc0d1e7),
	.w5(32'h3ba43fd6),
	.w6(32'hbacc50d7),
	.w7(32'h3b0e1e58),
	.w8(32'h3bd6da7e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c29b5),
	.w1(32'hbb212dfd),
	.w2(32'h3bc33202),
	.w3(32'h3c8c14e9),
	.w4(32'hb789536f),
	.w5(32'h3bf15ed8),
	.w6(32'hbbd93bff),
	.w7(32'h3b29c5a1),
	.w8(32'h3be322e3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f2a22),
	.w1(32'hbbade1c7),
	.w2(32'hbbf2ca1b),
	.w3(32'h3c5da9e3),
	.w4(32'hbc460ad9),
	.w5(32'hbc6b41f5),
	.w6(32'hbb8be8fd),
	.w7(32'hbc6788fa),
	.w8(32'hbca4e182),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5a07e),
	.w1(32'hbbbaffbf),
	.w2(32'h3b8e0f68),
	.w3(32'hbc161f69),
	.w4(32'hbb036231),
	.w5(32'h3c070e33),
	.w6(32'hbb80e664),
	.w7(32'hba4ea626),
	.w8(32'hba6a43fa),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c281b),
	.w1(32'hbb59dae4),
	.w2(32'h3c180bec),
	.w3(32'h3b68d356),
	.w4(32'h3bbf2206),
	.w5(32'h3a52c5ea),
	.w6(32'h3b2227c7),
	.w7(32'h3bb053f0),
	.w8(32'h3a2e7ddd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa0f6b),
	.w1(32'h3b84664b),
	.w2(32'h3c5892dc),
	.w3(32'hbc1bcf84),
	.w4(32'h3acf7145),
	.w5(32'h3c0af1b7),
	.w6(32'h3b0a3aff),
	.w7(32'h3ba83a74),
	.w8(32'h3b0697a7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31271e),
	.w1(32'hbc170b2f),
	.w2(32'hbcc87408),
	.w3(32'h3be74e61),
	.w4(32'hbc2fe09a),
	.w5(32'hbc69ee19),
	.w6(32'hbbf21837),
	.w7(32'hbc422b62),
	.w8(32'hbc871707),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98cbc9),
	.w1(32'h3b23f21a),
	.w2(32'h3c959316),
	.w3(32'hbc11beb0),
	.w4(32'h3b93aa3c),
	.w5(32'h3c78ba5b),
	.w6(32'hb9e18927),
	.w7(32'h3c41886e),
	.w8(32'h3c676ad5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb26766),
	.w1(32'hbc30657c),
	.w2(32'hbbfad5f7),
	.w3(32'h3c6a48b7),
	.w4(32'hbc6583ed),
	.w5(32'hbc6bdf68),
	.w6(32'hbc3c0b2a),
	.w7(32'hbc4ead74),
	.w8(32'hbc115522),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a0e5f),
	.w1(32'hbbcc9127),
	.w2(32'hbbe0746f),
	.w3(32'hbbcdd5fb),
	.w4(32'hbabb4fe0),
	.w5(32'hbabd8712),
	.w6(32'hbb081bfb),
	.w7(32'h3c05ae93),
	.w8(32'hbbeb87d0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7ea60),
	.w1(32'hbafc03ae),
	.w2(32'hbb2cb32b),
	.w3(32'hbc2e407e),
	.w4(32'hbb8b3a55),
	.w5(32'hbb6f51ec),
	.w6(32'hba85e7ab),
	.w7(32'hbb291f1a),
	.w8(32'h39f863b7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25ef1f),
	.w1(32'h3b387855),
	.w2(32'hbb2e98a2),
	.w3(32'hba1176fe),
	.w4(32'hbb94f7bd),
	.w5(32'hbb90a38e),
	.w6(32'h3b70586b),
	.w7(32'h3aabd43f),
	.w8(32'hba93a246),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6d3da),
	.w1(32'h3b8f2b75),
	.w2(32'h3bd0ad80),
	.w3(32'h3ada49bf),
	.w4(32'hbabeed8b),
	.w5(32'h3b022591),
	.w6(32'h3b99426b),
	.w7(32'h3c02b618),
	.w8(32'h3ba7d693),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47d7fc),
	.w1(32'hbc255eb6),
	.w2(32'hbc1c7829),
	.w3(32'h3b79a805),
	.w4(32'hbc4c3a9d),
	.w5(32'hbbf0c021),
	.w6(32'hbc34e0b3),
	.w7(32'hbc1eca0d),
	.w8(32'hbc30caef),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb698e4e),
	.w1(32'h3b929893),
	.w2(32'hba0c7558),
	.w3(32'hba0319bc),
	.w4(32'h3ad6337e),
	.w5(32'h398bb10a),
	.w6(32'h3a3e113e),
	.w7(32'hbb046083),
	.w8(32'hbb83b01d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cd8d8),
	.w1(32'h3bd101ff),
	.w2(32'h3b5f8077),
	.w3(32'hbb955a96),
	.w4(32'h3bf236d5),
	.w5(32'h3bbb0b8d),
	.w6(32'h3b3f8f31),
	.w7(32'h3c341b32),
	.w8(32'h3b8768d6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeac69f),
	.w1(32'hbb3ba8da),
	.w2(32'hbb12f824),
	.w3(32'hbaca2a8d),
	.w4(32'h3a0890e0),
	.w5(32'h3ac8a88f),
	.w6(32'hba00a0f2),
	.w7(32'h3948a8ad),
	.w8(32'hb8c6ce7a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40ebcd),
	.w1(32'hbbdb6340),
	.w2(32'hbbceb75a),
	.w3(32'h3a355c8c),
	.w4(32'hbbe6fab9),
	.w5(32'hbbce2c58),
	.w6(32'hbbe71c01),
	.w7(32'hbba091c5),
	.w8(32'hbb4fd705),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e4603),
	.w1(32'hbcd42603),
	.w2(32'h3c5ce5a3),
	.w3(32'hbb0f6459),
	.w4(32'hbcb53d2d),
	.w5(32'h3cafd9b7),
	.w6(32'hbcdd1d00),
	.w7(32'hb8b5f5af),
	.w8(32'h3c6b4298),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c376b9d),
	.w1(32'hba104c71),
	.w2(32'h3c287c9f),
	.w3(32'h3c734cca),
	.w4(32'h3b3e9ecf),
	.w5(32'h3c03116c),
	.w6(32'hbb8745b6),
	.w7(32'h3baa2b9a),
	.w8(32'h3b99e2b4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccc55c),
	.w1(32'hbbc3a26c),
	.w2(32'h3d0bb7a5),
	.w3(32'h3b960c58),
	.w4(32'hbb402b2b),
	.w5(32'h3d15884f),
	.w6(32'hbc4a0f8f),
	.w7(32'h3c9895cd),
	.w8(32'h3caa3c56),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf4e37),
	.w1(32'h3b3936b8),
	.w2(32'h3c8ce580),
	.w3(32'h3c445886),
	.w4(32'h3b014df3),
	.w5(32'h3c52dc25),
	.w6(32'h3bac61b6),
	.w7(32'h3bafe93c),
	.w8(32'h3c905029),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1bccd),
	.w1(32'h3b9c89d9),
	.w2(32'hbbffd957),
	.w3(32'h3c725921),
	.w4(32'h3ba28bca),
	.w5(32'hbbe5ac14),
	.w6(32'h3b607822),
	.w7(32'hbb5606d0),
	.w8(32'hb98640c0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22700e),
	.w1(32'hbc342f6c),
	.w2(32'hbc56dc74),
	.w3(32'hbbebd188),
	.w4(32'hbc0e3198),
	.w5(32'hbb03ac84),
	.w6(32'hbc897ba4),
	.w7(32'hbc00ef15),
	.w8(32'h3c468018),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4b9c2),
	.w1(32'h3b9aba3c),
	.w2(32'hbb7e3d47),
	.w3(32'h3caaa4c6),
	.w4(32'h3adeeee5),
	.w5(32'hbb20e8aa),
	.w6(32'h3b7a635e),
	.w7(32'hbb081836),
	.w8(32'hbafd98c3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cedaa),
	.w1(32'h3a2a1d1d),
	.w2(32'hbb8644ca),
	.w3(32'hbb118ee3),
	.w4(32'hbaa8cd33),
	.w5(32'h3aab7938),
	.w6(32'h3bd491c6),
	.w7(32'hbba48e27),
	.w8(32'h3a1c777e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff576f),
	.w1(32'hba880920),
	.w2(32'h3b496e0f),
	.w3(32'h3a637328),
	.w4(32'hbb982f03),
	.w5(32'h3abb4ca5),
	.w6(32'hbb7bcd41),
	.w7(32'h3b85aa01),
	.w8(32'h3bbcd152),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad59613),
	.w1(32'h3b066451),
	.w2(32'hbcef38ed),
	.w3(32'h3b50ca2b),
	.w4(32'hbc71c8e5),
	.w5(32'hbcc83464),
	.w6(32'hbb9d512c),
	.w7(32'hbc59415b),
	.w8(32'hbc76aaa8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadbea8),
	.w1(32'h3b184f45),
	.w2(32'h3b37414e),
	.w3(32'hbbbad571),
	.w4(32'h3b17bb2d),
	.w5(32'h3b0a3d61),
	.w6(32'hba39c0ef),
	.w7(32'h3aee0f83),
	.w8(32'hbb5586ce),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d6fe2),
	.w1(32'hbb38f1e4),
	.w2(32'hbc356a25),
	.w3(32'hbb3f8f09),
	.w4(32'hba0a0ca2),
	.w5(32'hbc3d3aa2),
	.w6(32'hba165f53),
	.w7(32'hbbcecf3e),
	.w8(32'hbbec0fb0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d6d18),
	.w1(32'h3b5ad8a3),
	.w2(32'h3c09124c),
	.w3(32'hbbfcb213),
	.w4(32'hbb899ef5),
	.w5(32'hba0ab734),
	.w6(32'hbb6af350),
	.w7(32'h3bfff0c4),
	.w8(32'h3bb47a16),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b674489),
	.w1(32'hbb2dc845),
	.w2(32'h3b97c8d8),
	.w3(32'hbb0fe245),
	.w4(32'hbbb65db5),
	.w5(32'h3bdcc100),
	.w6(32'hbc221d0c),
	.w7(32'hbb9075a7),
	.w8(32'h3b09f2fc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07b72c),
	.w1(32'h3b95d5c1),
	.w2(32'hbacf8693),
	.w3(32'h3af13614),
	.w4(32'h3b391e8c),
	.w5(32'hbab85143),
	.w6(32'h3a26fb64),
	.w7(32'h3b8e2f7c),
	.w8(32'hbbcaf688),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eee37),
	.w1(32'hbac0922b),
	.w2(32'hbb64cd88),
	.w3(32'hbc385535),
	.w4(32'hba72a5c8),
	.w5(32'hbb32d55d),
	.w6(32'hbb50a728),
	.w7(32'hbb3da824),
	.w8(32'hbab05057),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19a87a),
	.w1(32'h3bdc6f64),
	.w2(32'h3b8b0070),
	.w3(32'h3b27d34b),
	.w4(32'h3bdcaf72),
	.w5(32'h3acfa402),
	.w6(32'hb9cfaefa),
	.w7(32'h3968878b),
	.w8(32'h3aebe8de),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe11ca9),
	.w1(32'hbbea0c49),
	.w2(32'hbbaa0595),
	.w3(32'hbc029250),
	.w4(32'hbb9a9b2b),
	.w5(32'hbb40374e),
	.w6(32'hbc044d89),
	.w7(32'hbb83330e),
	.w8(32'hbb73c1af),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba354519),
	.w1(32'hbb8a17f5),
	.w2(32'h3bca798f),
	.w3(32'h3a5d9334),
	.w4(32'hbbd1ae94),
	.w5(32'hbaf5895d),
	.w6(32'hbb688c23),
	.w7(32'h3b16429f),
	.w8(32'h3c097fb0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b264eff),
	.w1(32'h3c89b507),
	.w2(32'h3ca1ac0e),
	.w3(32'h3b6fc710),
	.w4(32'h3c2690f8),
	.w5(32'h3c8a0190),
	.w6(32'h3c688cae),
	.w7(32'h3cc693da),
	.w8(32'h3bf96e79),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ad057),
	.w1(32'hb833df9f),
	.w2(32'hbc6386ee),
	.w3(32'h3af956d8),
	.w4(32'h3ac58431),
	.w5(32'hbc0b3879),
	.w6(32'h3b6442bb),
	.w7(32'hbbf16f7d),
	.w8(32'hbc1618a5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6edfd6),
	.w1(32'hbaab6627),
	.w2(32'h388ead8d),
	.w3(32'hbbfa0dbd),
	.w4(32'hbacd70d5),
	.w5(32'h3b06a6ac),
	.w6(32'hbb26508f),
	.w7(32'hbab75817),
	.w8(32'h3abcd51d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be03e8d),
	.w1(32'hbbcbb4f5),
	.w2(32'hbbc691b8),
	.w3(32'h3be8d5fa),
	.w4(32'h3b67bfea),
	.w5(32'hb9935711),
	.w6(32'hbb98af93),
	.w7(32'hbbecc4ad),
	.w8(32'hbbeacf64),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28c5a3),
	.w1(32'hbafad3f2),
	.w2(32'h3b043076),
	.w3(32'hbc6eee5b),
	.w4(32'h39c49480),
	.w5(32'hbb87369b),
	.w6(32'hbb1b3241),
	.w7(32'hbb12e9fb),
	.w8(32'h3a3e3e75),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb4951),
	.w1(32'hbaa29bff),
	.w2(32'hbc2ebd4b),
	.w3(32'hbb8031fb),
	.w4(32'h3b693669),
	.w5(32'hbc02c172),
	.w6(32'h3b84afd9),
	.w7(32'hbbced3b4),
	.w8(32'hbbd1a142),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d1407),
	.w1(32'hbb4e9784),
	.w2(32'hbc2c7233),
	.w3(32'hbc0c3eeb),
	.w4(32'hbaa8b505),
	.w5(32'hbc1284c4),
	.w6(32'hbb0d0027),
	.w7(32'hbbe8ba03),
	.w8(32'hbb8f654e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66cbad),
	.w1(32'h39f87789),
	.w2(32'hb8830bd5),
	.w3(32'hbc49710d),
	.w4(32'h3bb1fa8c),
	.w5(32'hba94c61c),
	.w6(32'hbb0d4d6a),
	.w7(32'hbb866429),
	.w8(32'h3b4e7c10),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43672e),
	.w1(32'hbbb7d92f),
	.w2(32'hbac547e1),
	.w3(32'hbc101253),
	.w4(32'hbbded4a1),
	.w5(32'hbb313735),
	.w6(32'hbbc69dc5),
	.w7(32'hb9213fec),
	.w8(32'h3b8e256e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1df8b9),
	.w1(32'hbc22f207),
	.w2(32'hbbcb8eb0),
	.w3(32'h3bd9be1f),
	.w4(32'hbbe8f51d),
	.w5(32'hbbbdc951),
	.w6(32'hbc0a13e3),
	.w7(32'hbb9f1e19),
	.w8(32'hbb6244ed),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc011843),
	.w1(32'hbacae907),
	.w2(32'hb99735fc),
	.w3(32'hbbc54af1),
	.w4(32'h39154032),
	.w5(32'hbbae7f8e),
	.w6(32'hbb9e04b2),
	.w7(32'h3967fefd),
	.w8(32'hbc1028a2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb039b33),
	.w1(32'hbb852d66),
	.w2(32'hbbd578cd),
	.w3(32'hbc499001),
	.w4(32'hbb068db5),
	.w5(32'h3bb6efdb),
	.w6(32'hbaab1fab),
	.w7(32'hbbbd8a3a),
	.w8(32'hbc0d4f27),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09dd2b),
	.w1(32'h3b6c6e72),
	.w2(32'h3bb82b76),
	.w3(32'hbc5351ab),
	.w4(32'hbab34578),
	.w5(32'h3c240865),
	.w6(32'hbb978081),
	.w7(32'h3bc586d2),
	.w8(32'h3b6247c6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07a18d),
	.w1(32'hbaa9624a),
	.w2(32'hbbe1de5a),
	.w3(32'h3bcc4ec6),
	.w4(32'h3b37a461),
	.w5(32'hbb162c47),
	.w6(32'hbac8f5f7),
	.w7(32'hbbf0d5f0),
	.w8(32'h3b344a88),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cc7bb),
	.w1(32'h3c836ec4),
	.w2(32'hbb41d013),
	.w3(32'h3bd42bde),
	.w4(32'h3c3cc3db),
	.w5(32'hba75d1b9),
	.w6(32'h3c8e69e4),
	.w7(32'h3c567bdd),
	.w8(32'h3aee84d8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule