module layer_8_featuremap_104(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea2b2c),
	.w1(32'h3b971510),
	.w2(32'h3cdd4c78),
	.w3(32'hbc12cff6),
	.w4(32'h3c489d28),
	.w5(32'h3ca8f8ad),
	.w6(32'h3c72f04f),
	.w7(32'h3c7c00a1),
	.w8(32'hbae1b4e6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48d5dd),
	.w1(32'h3b470aab),
	.w2(32'h3a51fa59),
	.w3(32'hbb5639bc),
	.w4(32'hbb3af06e),
	.w5(32'hbb941ed1),
	.w6(32'hbb99c1c2),
	.w7(32'hbbb16a90),
	.w8(32'hbb9fb709),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cb504),
	.w1(32'h3b896d2c),
	.w2(32'h3b8e3b2c),
	.w3(32'hba733e27),
	.w4(32'h3842675e),
	.w5(32'hbb429f5f),
	.w6(32'hbb1f9720),
	.w7(32'hbaa623ae),
	.w8(32'hbacadf34),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb9d8f3),
	.w1(32'hbb6ca914),
	.w2(32'hbbcc5932),
	.w3(32'hbacf2f16),
	.w4(32'hbaaa38b0),
	.w5(32'hbb90e56b),
	.w6(32'hbc5e1040),
	.w7(32'hbc47cca6),
	.w8(32'hbbdfe57e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab947b2),
	.w1(32'h396aced9),
	.w2(32'h3af9718f),
	.w3(32'h3a3fe37b),
	.w4(32'hba909f4f),
	.w5(32'h3abfebbd),
	.w6(32'hbb08df2a),
	.w7(32'h3a5dfb8b),
	.w8(32'h3b05b426),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53e9ce),
	.w1(32'h3b8909af),
	.w2(32'hbc985708),
	.w3(32'h3c9ea0ee),
	.w4(32'hbc39780c),
	.w5(32'hbbbfc6d7),
	.w6(32'hbc9903a8),
	.w7(32'hbc2bc112),
	.w8(32'h3c1fcdef),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f8f4f),
	.w1(32'h38d295eb),
	.w2(32'h397e506d),
	.w3(32'h383b7627),
	.w4(32'h38222162),
	.w5(32'h39235376),
	.w6(32'h37fdecf4),
	.w7(32'hb70709bf),
	.w8(32'h393dccd1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc1765),
	.w1(32'h3bfd313e),
	.w2(32'h3c4edbd7),
	.w3(32'hbb9c5905),
	.w4(32'h3c1e3edf),
	.w5(32'h3c6f568b),
	.w6(32'h3b96cf6f),
	.w7(32'h3bcad7db),
	.w8(32'h3b735177),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10e43a),
	.w1(32'h3b7c3515),
	.w2(32'h3be8c3be),
	.w3(32'hbb31c2ec),
	.w4(32'hbac4ad4e),
	.w5(32'h3b45d953),
	.w6(32'hb94e2b4a),
	.w7(32'hbaf90c48),
	.w8(32'h3ae76b2d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefa173),
	.w1(32'h3ac62862),
	.w2(32'h3c3963db),
	.w3(32'hbc3a1d73),
	.w4(32'h3b3475f6),
	.w5(32'h3bd174dd),
	.w6(32'h3a482146),
	.w7(32'hbb2d2350),
	.w8(32'hbc22adb9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb606b6a),
	.w1(32'h3be10c05),
	.w2(32'h3cb5dd9e),
	.w3(32'hbbf90e96),
	.w4(32'h3c840683),
	.w5(32'h3ca2b131),
	.w6(32'h3c260b33),
	.w7(32'h3c7d6d5f),
	.w8(32'h3a8d4bae),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69a3c6),
	.w1(32'hbbc3234a),
	.w2(32'hbac48c13),
	.w3(32'hbbf3625f),
	.w4(32'hbc2d58ab),
	.w5(32'hbbba2254),
	.w6(32'h39d0729c),
	.w7(32'hbc1e1535),
	.w8(32'hbc49dd6d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e32fe),
	.w1(32'h3afffc1a),
	.w2(32'h3b0f6f49),
	.w3(32'h3a19fe8f),
	.w4(32'hbb96ac99),
	.w5(32'hbc5d9aa0),
	.w6(32'hbaa99878),
	.w7(32'hbb0ace2d),
	.w8(32'hbb325671),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40c7c4),
	.w1(32'h39f66f40),
	.w2(32'hbbae19f6),
	.w3(32'h3855f065),
	.w4(32'hbb94bb1f),
	.w5(32'hbc21249b),
	.w6(32'h3ac5a817),
	.w7(32'h3a687d09),
	.w8(32'h3c9067fc),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f35c0),
	.w1(32'hbae5b5f3),
	.w2(32'hbb426b98),
	.w3(32'h3b55ef5e),
	.w4(32'hba144bde),
	.w5(32'hbb992f5f),
	.w6(32'h3c4bee25),
	.w7(32'h3b4b0ad9),
	.w8(32'h3aa10f1e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba302e8),
	.w1(32'hbb22b9d3),
	.w2(32'hba6bd1bb),
	.w3(32'h39928f31),
	.w4(32'hbb3914cf),
	.w5(32'h399f6a15),
	.w6(32'h39b89ecf),
	.w7(32'hba9e724b),
	.w8(32'hbc127908),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41274b),
	.w1(32'h3b820342),
	.w2(32'hbbc9d66d),
	.w3(32'h3a54965e),
	.w4(32'hbc36692a),
	.w5(32'h3c1fc296),
	.w6(32'hbc35b8a1),
	.w7(32'h3cc93418),
	.w8(32'h3c5599cd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced13c8),
	.w1(32'h3ba6eb19),
	.w2(32'h3c7d017c),
	.w3(32'hbc634ef2),
	.w4(32'h3c3ba8cb),
	.w5(32'h3b7457de),
	.w6(32'h3c9a76a8),
	.w7(32'hbc30bb31),
	.w8(32'hbd7b2bc7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda17412),
	.w1(32'hbc2605f1),
	.w2(32'h3d806a82),
	.w3(32'hbd8d6df4),
	.w4(32'h3d067e76),
	.w5(32'h3cf7056f),
	.w6(32'h3d0ffa1e),
	.w7(32'h3c7cb5cf),
	.w8(32'hbd56c708),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1272e9),
	.w1(32'hbcba259a),
	.w2(32'hbad22823),
	.w3(32'hbb369d50),
	.w4(32'h3c15438a),
	.w5(32'hbba9278f),
	.w6(32'h3c3192fb),
	.w7(32'hbbebc946),
	.w8(32'hbcc70597),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0b24f),
	.w1(32'h3c49c431),
	.w2(32'h3c21c5e2),
	.w3(32'hb9c1a37c),
	.w4(32'hbbc17cf4),
	.w5(32'h3c1fe65d),
	.w6(32'h3beddedf),
	.w7(32'h3ca51d53),
	.w8(32'h3ca0129c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c799aac),
	.w1(32'hbb5f899c),
	.w2(32'h3c03d57d),
	.w3(32'h3b8a4d42),
	.w4(32'hbc506d9e),
	.w5(32'hbb52f822),
	.w6(32'hbbb7a856),
	.w7(32'hbc6b2b67),
	.w8(32'hbd3c2cdf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b408150),
	.w1(32'hbc563f9e),
	.w2(32'h3d842e01),
	.w3(32'hbcd99c9f),
	.w4(32'h3d222ab2),
	.w5(32'h3da2a3db),
	.w6(32'hbb90a916),
	.w7(32'h3d093a2c),
	.w8(32'h3bfbe48e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0df9b),
	.w1(32'h3c26f29b),
	.w2(32'hbc61ad5a),
	.w3(32'h3c9159fb),
	.w4(32'hbb58fc56),
	.w5(32'hbbf45922),
	.w6(32'h3bfba9d0),
	.w7(32'hba649b9f),
	.w8(32'hbaf40c25),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaf73a),
	.w1(32'h3accfbab),
	.w2(32'hbac4594f),
	.w3(32'h3ad35b14),
	.w4(32'hbb820a25),
	.w5(32'hbc18f86c),
	.w6(32'h3bc5d08b),
	.w7(32'hbb0aa176),
	.w8(32'hbbf1b2de),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24ad38),
	.w1(32'hba967c86),
	.w2(32'h3c747b9d),
	.w3(32'hbc9bd065),
	.w4(32'hbc032e3c),
	.w5(32'h3c36a496),
	.w6(32'h3b04d6d4),
	.w7(32'h3c5cb65a),
	.w8(32'hbc2ab887),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca42ac),
	.w1(32'h3b5b87c3),
	.w2(32'hbc250731),
	.w3(32'h3b2e178e),
	.w4(32'hbc69b99d),
	.w5(32'hbc8d346a),
	.w6(32'h39d1e347),
	.w7(32'hbcacc85e),
	.w8(32'h3dd51c11),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd89e41),
	.w1(32'hbe52b8b2),
	.w2(32'h3d92f309),
	.w3(32'hbeb31bf9),
	.w4(32'h3dae2857),
	.w5(32'h3e52a598),
	.w6(32'hbd9ff9c6),
	.w7(32'h3d94d70f),
	.w8(32'hbd04476e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85beb3),
	.w1(32'h3c303f17),
	.w2(32'h3c955d2d),
	.w3(32'hbb05cffc),
	.w4(32'h3a76ed17),
	.w5(32'h3b28ca95),
	.w6(32'hbc4020c8),
	.w7(32'hbb7a9375),
	.w8(32'hbcdd0d2c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6f1e7),
	.w1(32'hbc70a4d8),
	.w2(32'hbc62d483),
	.w3(32'h3c2a8d8c),
	.w4(32'hbc1dafb2),
	.w5(32'hbbb5a809),
	.w6(32'h3bf54a1a),
	.w7(32'h3b06f66e),
	.w8(32'h3cdf5bde),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a0ecc),
	.w1(32'h3bccd145),
	.w2(32'h392898d6),
	.w3(32'hbc2e9d51),
	.w4(32'hb9ff9fa8),
	.w5(32'hba4d0606),
	.w6(32'hbc3b5023),
	.w7(32'h3af1ea0a),
	.w8(32'h3ac87c89),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93b58b),
	.w1(32'hba85d44e),
	.w2(32'hbd07fdde),
	.w3(32'h3b862731),
	.w4(32'hbc378fa3),
	.w5(32'hbc461d88),
	.w6(32'h3c097cd4),
	.w7(32'hbbafa939),
	.w8(32'h3cd38064),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9241f7),
	.w1(32'hbcb2af7a),
	.w2(32'h3cab3f74),
	.w3(32'hbc556d20),
	.w4(32'hba98cfd5),
	.w5(32'hb98fbcf1),
	.w6(32'hbcd7ea78),
	.w7(32'hb96f9e7e),
	.w8(32'hbc8e1d6e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d008b40),
	.w1(32'hbb46ca00),
	.w2(32'hbc24b13d),
	.w3(32'hbc30a4a4),
	.w4(32'hba948411),
	.w5(32'hbbf504ad),
	.w6(32'h3a44a83b),
	.w7(32'h3bc0e781),
	.w8(32'hbbab9a2e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ee7f3),
	.w1(32'h3bb3dcae),
	.w2(32'h3b2f580f),
	.w3(32'h3b6f4edf),
	.w4(32'hbb6e70d1),
	.w5(32'hbc995b14),
	.w6(32'h3ca0438a),
	.w7(32'hbbd2d451),
	.w8(32'hbd050bf7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeb67b),
	.w1(32'hbaa2bed4),
	.w2(32'h3bb2d208),
	.w3(32'hbcd4f21a),
	.w4(32'h3c0f023d),
	.w5(32'h3c2bdff9),
	.w6(32'hba2699aa),
	.w7(32'hbc62c271),
	.w8(32'hbd8565ba),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cde8404),
	.w1(32'hba858e40),
	.w2(32'hbc2002f9),
	.w3(32'h3c18846e),
	.w4(32'hba949ec8),
	.w5(32'h3c00e6c4),
	.w6(32'hbc40df60),
	.w7(32'hbbd64e6e),
	.w8(32'h3cb9f4c6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57f46b),
	.w1(32'hbc4b5a46),
	.w2(32'h3c2d0237),
	.w3(32'hbc1eaacd),
	.w4(32'h3b5f2e64),
	.w5(32'h3ba81dbb),
	.w6(32'h3cba682c),
	.w7(32'h3ca1cfe8),
	.w8(32'h3c435c38),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43965a),
	.w1(32'hbc1dfc70),
	.w2(32'h3b4607bc),
	.w3(32'hbc2efad3),
	.w4(32'hbbf319d4),
	.w5(32'hbbf248af),
	.w6(32'h3afac35f),
	.w7(32'h3b007157),
	.w8(32'h3c3f3fd9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba32090),
	.w1(32'hbce87c1f),
	.w2(32'h3afedee8),
	.w3(32'h3bc8fc3e),
	.w4(32'h3b987518),
	.w5(32'h3c915b60),
	.w6(32'hbb6f0f94),
	.w7(32'hbc1ff4b0),
	.w8(32'hbb6a147a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc222af9),
	.w1(32'hbc222c2d),
	.w2(32'hbc67bcca),
	.w3(32'hbc0f78ef),
	.w4(32'h3bbe6de3),
	.w5(32'hbca8d2a0),
	.w6(32'hbb7c6c8c),
	.w7(32'hbb94b469),
	.w8(32'hbd858688),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf861c0),
	.w1(32'h3bd5bb4b),
	.w2(32'h3c12c8a0),
	.w3(32'hba60c964),
	.w4(32'h3b32dea1),
	.w5(32'h3c940bb2),
	.w6(32'hba00775e),
	.w7(32'hbc837d7c),
	.w8(32'hbce52291),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf52268),
	.w1(32'h3c414238),
	.w2(32'h3c0f654d),
	.w3(32'hbb9d45b4),
	.w4(32'hbc631a57),
	.w5(32'hbba430ba),
	.w6(32'hbb1239c4),
	.w7(32'hbc68d844),
	.w8(32'hbca905bb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c373a42),
	.w1(32'hbb8bcdbe),
	.w2(32'h3b806146),
	.w3(32'hbc8477c9),
	.w4(32'hbad26924),
	.w5(32'h3ac802b8),
	.w6(32'h3a8cf617),
	.w7(32'h3c26c87d),
	.w8(32'h3b31e83e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd2488),
	.w1(32'hbc35d75a),
	.w2(32'h3cf1c23d),
	.w3(32'hbcb06ef3),
	.w4(32'h3b7dbf22),
	.w5(32'h3d197a0e),
	.w6(32'h3b768201),
	.w7(32'h3ce3cb82),
	.w8(32'h3bdb0edd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccf8372),
	.w1(32'hb93966ee),
	.w2(32'h39c0aca5),
	.w3(32'hba54463c),
	.w4(32'h3c45280c),
	.w5(32'hbbe80bd0),
	.w6(32'h3b30d029),
	.w7(32'hbb12453f),
	.w8(32'hbd11a5f0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c1763),
	.w1(32'h3b937a60),
	.w2(32'h3c6d8b04),
	.w3(32'h3beeae9b),
	.w4(32'h3893cbcb),
	.w5(32'h3b4050d7),
	.w6(32'hbc2ad897),
	.w7(32'h3b05160e),
	.w8(32'hbc52d338),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05e958),
	.w1(32'hbc7306c2),
	.w2(32'h3cee385e),
	.w3(32'hbca27fcc),
	.w4(32'h3ca25569),
	.w5(32'h3ce752ca),
	.w6(32'hbc48c2c6),
	.w7(32'h3cd8e6cf),
	.w8(32'hbb05b5ca),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb227e1),
	.w1(32'hbbf44842),
	.w2(32'hbccc370e),
	.w3(32'h3b89daf3),
	.w4(32'h3b625eb3),
	.w5(32'hbbcd5bff),
	.w6(32'h3c548374),
	.w7(32'hbc21d01f),
	.w8(32'h3b1eb6dc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62d475),
	.w1(32'h3c5105f1),
	.w2(32'hbd113117),
	.w3(32'hbc8a2370),
	.w4(32'hbcd396dd),
	.w5(32'hbbf8bd7e),
	.w6(32'hbcafdeeb),
	.w7(32'hbc984c5e),
	.w8(32'h3d1e597b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce008d4),
	.w1(32'hbd4e2baa),
	.w2(32'hbceca166),
	.w3(32'hbc0d6acf),
	.w4(32'hbca8b1b7),
	.w5(32'hbce5ae9b),
	.w6(32'h3b94a9ea),
	.w7(32'hbcc52c16),
	.w8(32'hbd227455),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc859322),
	.w1(32'hba5def69),
	.w2(32'h3c21621b),
	.w3(32'hbcf6281e),
	.w4(32'h3d0b1555),
	.w5(32'h3d2af798),
	.w6(32'h3d0c7f1b),
	.w7(32'h3cfd6393),
	.w8(32'hbda942e7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba727b8),
	.w1(32'h3b82b84c),
	.w2(32'hbbe157c9),
	.w3(32'h3c0b194b),
	.w4(32'hba1ffa4b),
	.w5(32'h3979a0ec),
	.w6(32'hbca0aff7),
	.w7(32'h3b5c85d3),
	.w8(32'h3d691c0e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6cbda),
	.w1(32'hbc09b84d),
	.w2(32'h3cdab4ab),
	.w3(32'hbd01a6a8),
	.w4(32'h3c7f30a8),
	.w5(32'h3c2ffc71),
	.w6(32'h3ce84ad7),
	.w7(32'h3c8627a8),
	.w8(32'h3c503b71),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e868b),
	.w1(32'h3ad4a492),
	.w2(32'hbc14fa79),
	.w3(32'h3a23fbc4),
	.w4(32'hbc71f7d9),
	.w5(32'hbbe72e8b),
	.w6(32'h3bdb9272),
	.w7(32'hbba0065f),
	.w8(32'h3ce17b9b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65a1b3),
	.w1(32'hbccdfedd),
	.w2(32'h3ca11333),
	.w3(32'hbd64ff41),
	.w4(32'hb9b8adf1),
	.w5(32'h3ca33bd0),
	.w6(32'h3beb42be),
	.w7(32'hb962836f),
	.w8(32'h3c786667),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb68e83),
	.w1(32'hbbcff3ec),
	.w2(32'h3c751fbe),
	.w3(32'hbc1302db),
	.w4(32'hbaf452d6),
	.w5(32'h3c6b912f),
	.w6(32'hbb824539),
	.w7(32'h3c0d89b2),
	.w8(32'h3c4d7a5b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ef4fb),
	.w1(32'h3c30d81e),
	.w2(32'h3c0dfc2f),
	.w3(32'hbcb8502b),
	.w4(32'h3cae321d),
	.w5(32'h3cef6b39),
	.w6(32'hbc8631a3),
	.w7(32'h3c38d7f5),
	.w8(32'hbd32f529),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd722ba9),
	.w1(32'hbba36760),
	.w2(32'h3c372421),
	.w3(32'hb97e1223),
	.w4(32'h3bafd2e1),
	.w5(32'h3c8fed7d),
	.w6(32'h3ca954d2),
	.w7(32'h3c8b1021),
	.w8(32'h3c82d152),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8bd19),
	.w1(32'hbbc0173f),
	.w2(32'hbb38668e),
	.w3(32'hb9cddd31),
	.w4(32'h3bea081e),
	.w5(32'h3c89dd7f),
	.w6(32'h3c6182ff),
	.w7(32'h3b77d670),
	.w8(32'hbcd61aa2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29b709),
	.w1(32'h3be64dc5),
	.w2(32'hba94fe34),
	.w3(32'hbae12d3d),
	.w4(32'h393ba843),
	.w5(32'h3b84e75b),
	.w6(32'h3b6633a4),
	.w7(32'hbbbe1d75),
	.w8(32'hbc81ba53),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37cb26),
	.w1(32'h3c49bb0f),
	.w2(32'hbb110bd5),
	.w3(32'hbc301fc4),
	.w4(32'hbb480cd4),
	.w5(32'h3bdd9b1d),
	.w6(32'h3bbc5846),
	.w7(32'hbc2f312b),
	.w8(32'hbbb40b4a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86a477),
	.w1(32'hbc289a5d),
	.w2(32'hb829b562),
	.w3(32'hbc1c50ba),
	.w4(32'hbc267c03),
	.w5(32'hbc2e4ed9),
	.w6(32'h3cede269),
	.w7(32'hbc2670e9),
	.w8(32'hbd6a1d42),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f5ddf),
	.w1(32'hbba7021e),
	.w2(32'h3c4ced04),
	.w3(32'h3c7f6c48),
	.w4(32'h3b8216ae),
	.w5(32'h3b50baa3),
	.w6(32'hbc16193e),
	.w7(32'h3c36f0d4),
	.w8(32'h3d2a4d70),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc765a4),
	.w1(32'hbb3ef860),
	.w2(32'h3ca67648),
	.w3(32'h3c202181),
	.w4(32'h3c5b7e87),
	.w5(32'h3ca7c60e),
	.w6(32'hbbb6b288),
	.w7(32'hbc10754d),
	.w8(32'hbc80b722),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb15e54),
	.w1(32'h3b7abcda),
	.w2(32'h3c97e26e),
	.w3(32'h3bff2afd),
	.w4(32'h3c7ed3ff),
	.w5(32'h3cc7ad38),
	.w6(32'hbc7670e2),
	.w7(32'h3ca2955d),
	.w8(32'hbc46f3a1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11da11),
	.w1(32'h3c1894c1),
	.w2(32'hbc5975a7),
	.w3(32'h3c0d16c8),
	.w4(32'h3c4955cd),
	.w5(32'hbb8aec36),
	.w6(32'h3c12ff7e),
	.w7(32'h3914245e),
	.w8(32'hbaa29db6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51da34),
	.w1(32'hbca21554),
	.w2(32'h3c3dc12d),
	.w3(32'h3a6c4a6c),
	.w4(32'hbbcd90e9),
	.w5(32'hbc88c9ca),
	.w6(32'h3cf0a2d4),
	.w7(32'h3c0caa28),
	.w8(32'hbc73f191),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d33f65e),
	.w1(32'h3c4f10b9),
	.w2(32'hbbf0ac5c),
	.w3(32'hbb856945),
	.w4(32'h3bf7ce07),
	.w5(32'h3ba9e35d),
	.w6(32'hbc919541),
	.w7(32'hbb5dd6ea),
	.w8(32'h3c0fa582),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5d855),
	.w1(32'hbd27ff88),
	.w2(32'h3d235f7c),
	.w3(32'hbd70f65b),
	.w4(32'h3d04609d),
	.w5(32'h3d9db5f4),
	.w6(32'h3c0e1252),
	.w7(32'h3d8b5db6),
	.w8(32'h3d120286),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad50098),
	.w1(32'h3c053990),
	.w2(32'hbc485ce1),
	.w3(32'hbb165a69),
	.w4(32'h3c83be00),
	.w5(32'h3c803cf2),
	.w6(32'hbb67f8ef),
	.w7(32'hbba53882),
	.w8(32'hbc7d790f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad544cf),
	.w1(32'h3cbdee2f),
	.w2(32'hbd14277a),
	.w3(32'h3bf3ca1a),
	.w4(32'hbc7cf134),
	.w5(32'hbc99fef4),
	.w6(32'h3bf5752f),
	.w7(32'h3d092aad),
	.w8(32'h3db5b8a5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd050b2c),
	.w1(32'hbb15353a),
	.w2(32'hbcd56dbb),
	.w3(32'h3aff4e38),
	.w4(32'h3bed11aa),
	.w5(32'h3c5b21c8),
	.w6(32'hbc63f62d),
	.w7(32'hbc5ed712),
	.w8(32'hbcae4ef4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09d7f7),
	.w1(32'hbc61eb73),
	.w2(32'h3c811053),
	.w3(32'hbbdf2602),
	.w4(32'h3c1c24af),
	.w5(32'h3ca02dd4),
	.w6(32'hbccaeda2),
	.w7(32'hbb8f9370),
	.w8(32'hbd7d91b9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31fa2a),
	.w1(32'h3c7ba59c),
	.w2(32'h3b9fdea4),
	.w3(32'h3a5ab18a),
	.w4(32'hbcb0d0fa),
	.w5(32'hbcc15e35),
	.w6(32'hbc73cd09),
	.w7(32'hbc653b46),
	.w8(32'h3d7b6264),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51d835),
	.w1(32'hbd09b87a),
	.w2(32'h39dfc72f),
	.w3(32'hbcdd2100),
	.w4(32'h3c7d3c95),
	.w5(32'h3c10e5bf),
	.w6(32'hbbf79624),
	.w7(32'h3cd65baf),
	.w8(32'h3c0bad3a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb829e4c),
	.w1(32'h3bdf62a5),
	.w2(32'h3b7ee2a8),
	.w3(32'h3c1a4caa),
	.w4(32'hbaa3af64),
	.w5(32'h3c025728),
	.w6(32'hbc0b5b9d),
	.w7(32'h3bd727c1),
	.w8(32'h3a16a638),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ee537),
	.w1(32'hbc160b35),
	.w2(32'h3c96d7c8),
	.w3(32'hbcef2dd3),
	.w4(32'h3c28ab23),
	.w5(32'h3cbd5522),
	.w6(32'h3c6dc6a4),
	.w7(32'h3c340c14),
	.w8(32'hbbfdfaf4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc6edd),
	.w1(32'h3accc216),
	.w2(32'h3b68dcfb),
	.w3(32'hbc664bb0),
	.w4(32'hbc00cee2),
	.w5(32'h3bc6c42f),
	.w6(32'h3b4a2c4f),
	.w7(32'hba9bfe64),
	.w8(32'hbb95d7dd),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9215c),
	.w1(32'h3b8421ef),
	.w2(32'hbca6141c),
	.w3(32'h3ba1b9a3),
	.w4(32'h3b3eb476),
	.w5(32'hbc7a6fed),
	.w6(32'h3b1e2f65),
	.w7(32'hbbe6016e),
	.w8(32'hbc6bc488),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3bb34),
	.w1(32'hbc5d8939),
	.w2(32'hbc62d643),
	.w3(32'hb9216ea4),
	.w4(32'h3c36f8c7),
	.w5(32'hbc844207),
	.w6(32'h3b6f07c2),
	.w7(32'h3be81732),
	.w8(32'hbc011e24),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d11e7a4),
	.w1(32'h3c280c39),
	.w2(32'h3bdffb39),
	.w3(32'h3b35b131),
	.w4(32'hbc7374eb),
	.w5(32'h3c1686c5),
	.w6(32'hbc90cf16),
	.w7(32'hbb0ce322),
	.w8(32'h3d2d3cd2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdbb177),
	.w1(32'hbac9696a),
	.w2(32'hbc21f299),
	.w3(32'hbcc569d4),
	.w4(32'h3caecd34),
	.w5(32'hbc8a4764),
	.w6(32'hbcb6b179),
	.w7(32'h3ca56a49),
	.w8(32'hbd047117),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a2aa1),
	.w1(32'hbd3e975d),
	.w2(32'hbd7dadd2),
	.w3(32'hbd2620d2),
	.w4(32'hbc702e77),
	.w5(32'hbd878a05),
	.w6(32'h3cf1f7ae),
	.w7(32'hbcb5dbf6),
	.w8(32'hbd5070a1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee082a),
	.w1(32'h3a613d82),
	.w2(32'h3cb2fbc3),
	.w3(32'hbc65de40),
	.w4(32'h3cb2cd0a),
	.w5(32'h3c528b30),
	.w6(32'hba9dcd6e),
	.w7(32'h3ca389bb),
	.w8(32'hbcbdca4c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccf3b3d),
	.w1(32'h3bd98167),
	.w2(32'h3c8eaca9),
	.w3(32'hbc48706e),
	.w4(32'hbc7f72d3),
	.w5(32'h3c36324f),
	.w6(32'hbbbdddf2),
	.w7(32'hbbf06bcd),
	.w8(32'h3c651ff0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb217a73),
	.w1(32'h3abb1bb1),
	.w2(32'h3b8232a7),
	.w3(32'hbc0ac719),
	.w4(32'h39fab3ea),
	.w5(32'h3c828ea9),
	.w6(32'h3c1d0bf6),
	.w7(32'h3c7ced2e),
	.w8(32'hbb60df67),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94f038),
	.w1(32'h3a9d59b3),
	.w2(32'h3c16fd43),
	.w3(32'h3aca58c5),
	.w4(32'hbb0a48f4),
	.w5(32'h3cb30ce6),
	.w6(32'h3b24cf1b),
	.w7(32'h3bcd5ba1),
	.w8(32'h3c15ab34),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb984862),
	.w1(32'h38a3e849),
	.w2(32'hbc26f630),
	.w3(32'hbb49f537),
	.w4(32'hbb673eb7),
	.w5(32'hbb2f798f),
	.w6(32'h38d09450),
	.w7(32'h3b054c0f),
	.w8(32'hbbe8593b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accdfa4),
	.w1(32'h3bb21fbf),
	.w2(32'hbcb3e31a),
	.w3(32'hbb82acd8),
	.w4(32'h3cb325af),
	.w5(32'hbcf3500a),
	.w6(32'h3c02cc14),
	.w7(32'h3b865bef),
	.w8(32'hbca0e468),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d784320),
	.w1(32'hbc5db4be),
	.w2(32'h3bfb5ddb),
	.w3(32'h3c50327d),
	.w4(32'hbc132d4b),
	.w5(32'h3bb54274),
	.w6(32'h3ca1c804),
	.w7(32'hbbd340fc),
	.w8(32'h3c872e84),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a5c4d),
	.w1(32'hbbe5026d),
	.w2(32'hbbee07d7),
	.w3(32'h3bcd9956),
	.w4(32'hbaf1152e),
	.w5(32'hbb22de00),
	.w6(32'hbcc39b65),
	.w7(32'hbbc1df35),
	.w8(32'hbae93385),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce880d6),
	.w1(32'h3c49cc19),
	.w2(32'hbc6c5c1c),
	.w3(32'h3c5e226d),
	.w4(32'h394a007f),
	.w5(32'h3c892017),
	.w6(32'hbb160936),
	.w7(32'h3cb66f53),
	.w8(32'hbc8e240a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12ef7f),
	.w1(32'h3ba17a88),
	.w2(32'hbc0e09d6),
	.w3(32'hbc3b9497),
	.w4(32'h3be8b25c),
	.w5(32'h3cb60a8f),
	.w6(32'h3ce3a79f),
	.w7(32'h3d49ef09),
	.w8(32'hbdc27626),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0053b0),
	.w1(32'hbc809a0e),
	.w2(32'h3ad77bdc),
	.w3(32'hbcf870c9),
	.w4(32'hbb24fc4b),
	.w5(32'hbc15dd57),
	.w6(32'h3cde0e1d),
	.w7(32'hbc1cc7c6),
	.w8(32'hbc2b7f6c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd1a17),
	.w1(32'hbc211d57),
	.w2(32'h3c0e6eb8),
	.w3(32'hbc96ef60),
	.w4(32'hbc2a8aaf),
	.w5(32'hbc6738a1),
	.w6(32'hbbbc896d),
	.w7(32'hba7a8166),
	.w8(32'hbad3e25e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3e4b0),
	.w1(32'h39e7db04),
	.w2(32'h3bc7f523),
	.w3(32'hbbc03c44),
	.w4(32'h3b9ce2be),
	.w5(32'h3cb4b6f1),
	.w6(32'hbc27d640),
	.w7(32'h3d0ff4f2),
	.w8(32'hbce5f561),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cb1b0),
	.w1(32'h3c4d94a9),
	.w2(32'hbc9133a4),
	.w3(32'hbcbd08ce),
	.w4(32'hbb463b4d),
	.w5(32'hbc858179),
	.w6(32'hbc34e450),
	.w7(32'hbc0d1e6d),
	.w8(32'hbc4c8bf6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d168c29),
	.w1(32'hbc4ed219),
	.w2(32'h3c02d34a),
	.w3(32'h3bc485da),
	.w4(32'h3c166c74),
	.w5(32'hbb9d2f2c),
	.w6(32'hbbeae680),
	.w7(32'h3c041b3a),
	.w8(32'hbc42e632),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeea414),
	.w1(32'hbb447580),
	.w2(32'h3ad63a01),
	.w3(32'h3b862d44),
	.w4(32'hbc89b76e),
	.w5(32'h3cf20a14),
	.w6(32'h3b0c9c4e),
	.w7(32'h3d10fc03),
	.w8(32'hbcc57e6d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf4494b),
	.w1(32'h3ca354d1),
	.w2(32'hbc43941a),
	.w3(32'hbca36689),
	.w4(32'hbb58cf4e),
	.w5(32'hbbb5e733),
	.w6(32'hbc8c5c3b),
	.w7(32'h3bb2a8c3),
	.w8(32'hbd0c9fc3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10da1b),
	.w1(32'h3bef0877),
	.w2(32'h3c21a397),
	.w3(32'h39ed42e6),
	.w4(32'h3b791ab8),
	.w5(32'hbaa2b307),
	.w6(32'h3c841eac),
	.w7(32'hbae3f43f),
	.w8(32'h3c95245e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b728c58),
	.w1(32'h3ba0c861),
	.w2(32'h3c03b85b),
	.w3(32'h3c26f7e3),
	.w4(32'hbbda9ef7),
	.w5(32'hbb2a19d3),
	.w6(32'h3bebd390),
	.w7(32'h3bba84cb),
	.w8(32'hbbeb2873),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c260fe3),
	.w1(32'h3b513a6e),
	.w2(32'h3884fc70),
	.w3(32'h3b9d7256),
	.w4(32'h3c37abea),
	.w5(32'h3bd9959a),
	.w6(32'hba49e745),
	.w7(32'h3c730c14),
	.w8(32'h3b394c68),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb5d4),
	.w1(32'hbb940476),
	.w2(32'hbc9cb3a3),
	.w3(32'hbbe3fc08),
	.w4(32'h3a63f5ce),
	.w5(32'hbcf2e568),
	.w6(32'hbc7089ae),
	.w7(32'hbd2d5657),
	.w8(32'h3d06a5b0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c872722),
	.w1(32'hbcb677eb),
	.w2(32'h3cf08eac),
	.w3(32'hbcc1c45a),
	.w4(32'h3caf6072),
	.w5(32'h3d5627a2),
	.w6(32'hbc846364),
	.w7(32'h3cdb8ec0),
	.w8(32'h3be82fb4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb523ea9),
	.w1(32'hbbadf42d),
	.w2(32'h3cca0788),
	.w3(32'h3b4ae2cb),
	.w4(32'hbc227ca4),
	.w5(32'h3d050998),
	.w6(32'h3c00e909),
	.w7(32'h39e872c1),
	.w8(32'h3c8c4b71),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5a0951),
	.w1(32'h3ce513bd),
	.w2(32'h3b5ec491),
	.w3(32'hbc60d2fd),
	.w4(32'h3b525e3d),
	.w5(32'h3c1e4556),
	.w6(32'hbc2532a9),
	.w7(32'h3c3f26a1),
	.w8(32'hb98f4d5f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1953b3),
	.w1(32'h3ac61c11),
	.w2(32'hbb48e24a),
	.w3(32'hbab9d441),
	.w4(32'hbbe51829),
	.w5(32'hbb50e867),
	.w6(32'hbc00e21e),
	.w7(32'h3bf6306b),
	.w8(32'hbcb5252f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc318f70),
	.w1(32'h3b8e2584),
	.w2(32'h3d190bde),
	.w3(32'hbc019d5a),
	.w4(32'hbc866e63),
	.w5(32'h3d3d68c0),
	.w6(32'hbab71b4e),
	.w7(32'h3c2421b0),
	.w8(32'h3c4f312b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd654889),
	.w1(32'h3c55ccd2),
	.w2(32'hb888a39c),
	.w3(32'hbca3168f),
	.w4(32'h3bc97f2b),
	.w5(32'hbc8efbfd),
	.w6(32'hbc0a2869),
	.w7(32'h3baf5040),
	.w8(32'hbc6033f7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a5caf),
	.w1(32'h39a7b754),
	.w2(32'hbbddbdf9),
	.w3(32'hbbd54484),
	.w4(32'h3b1bbb2c),
	.w5(32'hba906dee),
	.w6(32'h3b9df97e),
	.w7(32'hbb96dbd3),
	.w8(32'hbd54d6ed),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956d074),
	.w1(32'h3cb1d43b),
	.w2(32'hbc0f763f),
	.w3(32'hbc8db2d0),
	.w4(32'hbc8ad994),
	.w5(32'hbb449f9d),
	.w6(32'h3c24cdfb),
	.w7(32'hbb29c028),
	.w8(32'hbb8a89fc),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5ec21),
	.w1(32'hbc8286cb),
	.w2(32'hbc6ad23f),
	.w3(32'hbc07c86c),
	.w4(32'hbccb6c41),
	.w5(32'hbcb57600),
	.w6(32'hbc4d6260),
	.w7(32'hbcf22351),
	.w8(32'hbaa275be),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe9298),
	.w1(32'hbd0f1dc5),
	.w2(32'hbcfc073e),
	.w3(32'hbcb6dd83),
	.w4(32'hb91a9598),
	.w5(32'hbc87055a),
	.w6(32'hbcf382d5),
	.w7(32'hbb1957fb),
	.w8(32'h3c6fcf4a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba714c0),
	.w1(32'h3aaf9add),
	.w2(32'hbc01a7b9),
	.w3(32'hbbab6e22),
	.w4(32'h3c13f735),
	.w5(32'hbbaa1b0c),
	.w6(32'h3c9fb84f),
	.w7(32'hbc883502),
	.w8(32'hbb24ea79),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c173de5),
	.w1(32'h3c0d0218),
	.w2(32'hbc102b2a),
	.w3(32'hbc3b2a6b),
	.w4(32'h3cb0da85),
	.w5(32'hbc55e4b1),
	.w6(32'h3d15f9a5),
	.w7(32'hbb9a7fce),
	.w8(32'h3d15ce55),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcccd51b),
	.w1(32'hbcb3812b),
	.w2(32'hba577ba2),
	.w3(32'hbd07aaf8),
	.w4(32'h3add8078),
	.w5(32'h3c4b2ab8),
	.w6(32'hbca7a00a),
	.w7(32'h3b822380),
	.w8(32'hbbcdc767),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7250a),
	.w1(32'h3b147a91),
	.w2(32'hbc38b9fe),
	.w3(32'h38931380),
	.w4(32'h3b9931dc),
	.w5(32'h3c7f8cf5),
	.w6(32'hbb1f147f),
	.w7(32'h3cb90f56),
	.w8(32'hbd5531a8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40f8f0),
	.w1(32'hbba23bcf),
	.w2(32'hbbc482e9),
	.w3(32'hbc2a3e58),
	.w4(32'hbbccd144),
	.w5(32'h3be74be8),
	.w6(32'h3c92c7fc),
	.w7(32'hbbeccd09),
	.w8(32'h3cd23801),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac25d8d),
	.w1(32'h3b67abd5),
	.w2(32'h3c010f93),
	.w3(32'hbba9630d),
	.w4(32'h3b7797c6),
	.w5(32'h3cbb6996),
	.w6(32'hbc14a303),
	.w7(32'h3c8cf92a),
	.w8(32'h3c8bdfcd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75ef31),
	.w1(32'h3b8b4abb),
	.w2(32'hbc23622e),
	.w3(32'hbbbcc6c3),
	.w4(32'hbb0cd465),
	.w5(32'hbc0e6549),
	.w6(32'hbacc2ef5),
	.w7(32'hbc0778cf),
	.w8(32'h3bce9e21),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f2e4a),
	.w1(32'h3b80375b),
	.w2(32'h3b8456d3),
	.w3(32'hbb949210),
	.w4(32'hbaa52eeb),
	.w5(32'h3c054ed8),
	.w6(32'h3ad70c48),
	.w7(32'h3bb133f4),
	.w8(32'hbb8bd131),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c519c),
	.w1(32'h3bdb10ad),
	.w2(32'hbbd21ebf),
	.w3(32'h3b0b626e),
	.w4(32'hbb98a6c9),
	.w5(32'hbcb917de),
	.w6(32'hbb18c4d8),
	.w7(32'hbd2ab45b),
	.w8(32'h3d74ac2e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09b676),
	.w1(32'h3af2a082),
	.w2(32'h3befb7e3),
	.w3(32'h3c3b06ba),
	.w4(32'h3a925835),
	.w5(32'h3c425e86),
	.w6(32'hbcbde81d),
	.w7(32'hbcf1c387),
	.w8(32'h3d5baeb7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4cdcb1),
	.w1(32'hba5598f7),
	.w2(32'hbb311da8),
	.w3(32'hbc81133d),
	.w4(32'h394da282),
	.w5(32'h3aa008b4),
	.w6(32'hbd04a28f),
	.w7(32'h3c4da5ba),
	.w8(32'hbb8d32b2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc033998),
	.w1(32'h3bab13d2),
	.w2(32'hbc18e8bf),
	.w3(32'hbae54f99),
	.w4(32'h3bb0a8b5),
	.w5(32'hbc7571c7),
	.w6(32'h3b11fb79),
	.w7(32'hbcbabb6a),
	.w8(32'hbc8d83f5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adacb81),
	.w1(32'h3c091dba),
	.w2(32'h3cb783a2),
	.w3(32'hbce9ffa0),
	.w4(32'h3c00d61c),
	.w5(32'h3beb9077),
	.w6(32'h3c0f91af),
	.w7(32'h3c92e5ab),
	.w8(32'h3c30766a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule