module layer_6_featuremap_86(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b762c3c),
	.w1(32'h3b6d6d32),
	.w2(32'hbc0732c2),
	.w3(32'hb8a902e4),
	.w4(32'hb9aaee9b),
	.w5(32'hbb740609),
	.w6(32'h3a345890),
	.w7(32'hbb2d5cdb),
	.w8(32'hbb8cd082),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb84521),
	.w1(32'h3a9fb269),
	.w2(32'hbb29afb3),
	.w3(32'hbbd495ee),
	.w4(32'hbb657531),
	.w5(32'hbb9ce52e),
	.w6(32'h3b01f337),
	.w7(32'hbb24f400),
	.w8(32'hbb568b06),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3ba4e),
	.w1(32'h3bf525f4),
	.w2(32'hbbcbf613),
	.w3(32'hbb8aaed4),
	.w4(32'h3bbcb8e4),
	.w5(32'hbc0010cc),
	.w6(32'h3b7eedf5),
	.w7(32'hbba4b403),
	.w8(32'hbc093f04),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc207bb8),
	.w1(32'hbb135b95),
	.w2(32'h3b88714f),
	.w3(32'hbae78dff),
	.w4(32'hba633d9d),
	.w5(32'h39266fb5),
	.w6(32'hbb2dccb2),
	.w7(32'h3b6dd3ac),
	.w8(32'hbb1945e8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fa8b7),
	.w1(32'h3d041a86),
	.w2(32'hbd810044),
	.w3(32'hbd236070),
	.w4(32'h3c35ee73),
	.w5(32'h3a5e30fc),
	.w6(32'h3a8c7ddf),
	.w7(32'hbd397727),
	.w8(32'h3d29632a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d326605),
	.w1(32'h3a793d4b),
	.w2(32'hbb83e241),
	.w3(32'hb885f257),
	.w4(32'hba498668),
	.w5(32'hba28cf25),
	.w6(32'hb9b20765),
	.w7(32'hbac6ea30),
	.w8(32'hbb117abb),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbce9b7),
	.w1(32'hbbbcc85e),
	.w2(32'h3c2e5559),
	.w3(32'hbb797e89),
	.w4(32'hba7b8a83),
	.w5(32'h3bcf059d),
	.w6(32'hbba2312d),
	.w7(32'h3a3d9eb3),
	.w8(32'h3a4de156),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4871f9),
	.w1(32'hbd2e18e6),
	.w2(32'h3d19f7ed),
	.w3(32'h3acf5f65),
	.w4(32'h3c7f8cca),
	.w5(32'hbc524eb5),
	.w6(32'hbca8cc4a),
	.w7(32'h3d31faf1),
	.w8(32'hbd301641),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5b663),
	.w1(32'h3ca0130a),
	.w2(32'hbd1c46b2),
	.w3(32'hbb12897a),
	.w4(32'hbc219b06),
	.w5(32'h3c0c79d1),
	.w6(32'h3cf063aa),
	.w7(32'hbd80bf69),
	.w8(32'h3cc1cae9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38a838),
	.w1(32'hbaa895c8),
	.w2(32'hbb8c7bba),
	.w3(32'h398d629c),
	.w4(32'h3960ac6e),
	.w5(32'hbb30ba7d),
	.w6(32'hbaba4176),
	.w7(32'hbb504e07),
	.w8(32'hbb76438e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cd18a),
	.w1(32'hbb1f2f32),
	.w2(32'hbcdbf037),
	.w3(32'hbc230f35),
	.w4(32'hbcdc5e29),
	.w5(32'hbb88f4d0),
	.w6(32'hbc04e19d),
	.w7(32'hbd4f5611),
	.w8(32'hbd19cb29),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd060e13),
	.w1(32'h3c02f302),
	.w2(32'hbc2ea772),
	.w3(32'h3b0a83a1),
	.w4(32'h3b06600a),
	.w5(32'hba599597),
	.w6(32'h3a906510),
	.w7(32'hbbe7ea53),
	.w8(32'hbac5c716),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6697cd),
	.w1(32'hbb3e0dcc),
	.w2(32'h3c17947d),
	.w3(32'hbb8cf8df),
	.w4(32'h3c42134a),
	.w5(32'h39ca537e),
	.w6(32'h3a2f1b6d),
	.w7(32'h3c0764c0),
	.w8(32'hbb94a33a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb2d07),
	.w1(32'h3c72ecac),
	.w2(32'hbbd1eacc),
	.w3(32'hbbedd7a9),
	.w4(32'hbb50dafa),
	.w5(32'hbc198ef7),
	.w6(32'hbba8bca0),
	.w7(32'hbc89bee7),
	.w8(32'hbc7ff7c5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c6a5d),
	.w1(32'hbbfc0e17),
	.w2(32'hba9aa253),
	.w3(32'hbc02f228),
	.w4(32'hbbcf8521),
	.w5(32'h3c51afb8),
	.w6(32'hbc2467f9),
	.w7(32'hbb0e5628),
	.w8(32'h3ba98fec),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba075ef0),
	.w1(32'hba980114),
	.w2(32'h3b106dc7),
	.w3(32'h3b60f90c),
	.w4(32'h3a8327a5),
	.w5(32'h3a1a1baa),
	.w6(32'hb8f60a57),
	.w7(32'h3b3bf1e4),
	.w8(32'hbbafaf7a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc85d09),
	.w1(32'h3b4e90ab),
	.w2(32'h3c67ff16),
	.w3(32'h3a632d58),
	.w4(32'h3c66208d),
	.w5(32'hbc11d8ef),
	.w6(32'h3cab7669),
	.w7(32'h3cb8b08b),
	.w8(32'h3c462276),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897de5),
	.w1(32'hb9269452),
	.w2(32'hba1c93e2),
	.w3(32'h3b629d7d),
	.w4(32'hbbcbbe56),
	.w5(32'hba951c94),
	.w6(32'hb9713a01),
	.w7(32'hbb489f72),
	.w8(32'hbc01d430),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95faf0),
	.w1(32'hb9ac7f6d),
	.w2(32'hba383761),
	.w3(32'h3b7c4666),
	.w4(32'h3af951fd),
	.w5(32'h3a5529ce),
	.w6(32'h3ad6944c),
	.w7(32'h39b94577),
	.w8(32'h3adfc79c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31f9b8),
	.w1(32'h3bb66c8a),
	.w2(32'hbcb71a7c),
	.w3(32'h3bd6c120),
	.w4(32'h3c34b5e8),
	.w5(32'hbc322c6e),
	.w6(32'h3d1824e9),
	.w7(32'hbc7077f2),
	.w8(32'h3c4dd931),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e6af3),
	.w1(32'hbae72f45),
	.w2(32'hbb0fe064),
	.w3(32'hbba07458),
	.w4(32'hbb46a743),
	.w5(32'hb909362b),
	.w6(32'hbbbc46a3),
	.w7(32'hbaeb965d),
	.w8(32'hbb7fa4cc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff9791),
	.w1(32'h3ad6e388),
	.w2(32'hbba877b4),
	.w3(32'hbbac3f40),
	.w4(32'h3bbfe6ec),
	.w5(32'h3bc68375),
	.w6(32'h3afdca5a),
	.w7(32'h3b4422e0),
	.w8(32'hbaf50c6e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999f190),
	.w1(32'h3b82dbc3),
	.w2(32'h3b250b53),
	.w3(32'hbc8da24a),
	.w4(32'h3cb7b3b3),
	.w5(32'hbc8290a6),
	.w6(32'hbca37b0b),
	.w7(32'h3d110606),
	.w8(32'hbcc85714),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9f2ad),
	.w1(32'hbb528fab),
	.w2(32'h3c47719b),
	.w3(32'h3d18c6af),
	.w4(32'hbcbc71e3),
	.w5(32'h3c6dd484),
	.w6(32'h3c226e82),
	.w7(32'hb93c3d28),
	.w8(32'h3bd104c3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca66a3a),
	.w1(32'h3b85de97),
	.w2(32'hbc09ef75),
	.w3(32'h3ba60f43),
	.w4(32'hbc3851a4),
	.w5(32'h3a758eb2),
	.w6(32'h3bfabfbc),
	.w7(32'hbc140d49),
	.w8(32'hbb24913a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce5fcc7),
	.w1(32'h3c00d335),
	.w2(32'h3aa2c035),
	.w3(32'hbbcfaeee),
	.w4(32'h3b29b8e3),
	.w5(32'h3a773426),
	.w6(32'hba598167),
	.w7(32'h3c1ee4bc),
	.w8(32'h3c100085),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b04b9),
	.w1(32'hb9a2d6f1),
	.w2(32'h3b545ce7),
	.w3(32'h3b4a0061),
	.w4(32'hba2607c5),
	.w5(32'hbb17b38b),
	.w6(32'hbbed76aa),
	.w7(32'h3ba8f07a),
	.w8(32'hbac414fd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82f34f),
	.w1(32'hbb9ff612),
	.w2(32'h3b0e41ef),
	.w3(32'h39fbe5c9),
	.w4(32'hbb29bc5f),
	.w5(32'h3b0ab4e1),
	.w6(32'hbab2e7c0),
	.w7(32'hbb005d0a),
	.w8(32'h3b89c024),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af21149),
	.w1(32'hbb45cd71),
	.w2(32'hba851b97),
	.w3(32'h3ab0bd07),
	.w4(32'h39423379),
	.w5(32'h3a8277ec),
	.w6(32'hba859072),
	.w7(32'hb7eb53aa),
	.w8(32'h3a20e76b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51c494),
	.w1(32'hbc669182),
	.w2(32'h3c842e7e),
	.w3(32'h3bfda514),
	.w4(32'hbcda6775),
	.w5(32'h3aeaa45d),
	.w6(32'h3c273514),
	.w7(32'hbbb04c14),
	.w8(32'h3a871c73),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9853107),
	.w1(32'h3c69d8d8),
	.w2(32'hbcc2f816),
	.w3(32'hbd2bec55),
	.w4(32'h3c9943f7),
	.w5(32'h3c427506),
	.w6(32'hbc87dd61),
	.w7(32'hbc59a9a6),
	.w8(32'h3cb5bf28),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdd811b),
	.w1(32'h3c47fe63),
	.w2(32'hbc47b9ec),
	.w3(32'hbbfeed51),
	.w4(32'hbc3bdb2e),
	.w5(32'h3b2750e7),
	.w6(32'h3b55e862),
	.w7(32'hbc2ba7a1),
	.w8(32'h3b55ad78),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11df50),
	.w1(32'hbd00073b),
	.w2(32'h3c9b471b),
	.w3(32'h3c292a28),
	.w4(32'hbcafaf70),
	.w5(32'h395dfe8e),
	.w6(32'hbb67daaf),
	.w7(32'h3c97129c),
	.w8(32'hbce1dbc0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd207293),
	.w1(32'h3cac29ac),
	.w2(32'h3d0a0234),
	.w3(32'hbb01c0f7),
	.w4(32'h3d2e12ca),
	.w5(32'hbc3305d1),
	.w6(32'h3c8bcc72),
	.w7(32'h3d90158d),
	.w8(32'h3cdf97b5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb886ac),
	.w1(32'h3b986f10),
	.w2(32'hba2c498d),
	.w3(32'h3ad8732a),
	.w4(32'h3c093055),
	.w5(32'hbab411ca),
	.w6(32'h3b069dfb),
	.w7(32'h3b92eafc),
	.w8(32'hbb542fd8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac77f53),
	.w1(32'hbb9fec47),
	.w2(32'h3b31a0a9),
	.w3(32'h3b0ffb91),
	.w4(32'h3c497197),
	.w5(32'hbab67c94),
	.w6(32'hbc2f42d0),
	.w7(32'h3c0d3cc7),
	.w8(32'hbbb31e41),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98bd87),
	.w1(32'h3bd67198),
	.w2(32'hbc2b4c4c),
	.w3(32'hbb2da1f9),
	.w4(32'h3aeef961),
	.w5(32'hbb6e94ff),
	.w6(32'h39e1e831),
	.w7(32'hbaf5a502),
	.w8(32'h3b1e4608),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecb47d),
	.w1(32'h3a69b23f),
	.w2(32'hbb9e007d),
	.w3(32'hba6077a6),
	.w4(32'h393383a4),
	.w5(32'h38bbdfb7),
	.w6(32'hbad03aef),
	.w7(32'hbb20ddaf),
	.w8(32'h3adcec73),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8378c3),
	.w1(32'h3b906a68),
	.w2(32'hbc6e635e),
	.w3(32'h3b881a1e),
	.w4(32'hbc31814e),
	.w5(32'hbbc1dec7),
	.w6(32'h3b8133bf),
	.w7(32'hbcb8b625),
	.w8(32'hbba63d24),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ce3b6),
	.w1(32'h3c86ecd9),
	.w2(32'hbae460dd),
	.w3(32'h3d0849d8),
	.w4(32'hbd876ddc),
	.w5(32'h3cd9f381),
	.w6(32'h3d885219),
	.w7(32'hbdb2fc97),
	.w8(32'h3cfa0314),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca623e6),
	.w1(32'h3a847476),
	.w2(32'hbcca4aed),
	.w3(32'hbcb7123b),
	.w4(32'h3c741053),
	.w5(32'hbb0a1202),
	.w6(32'hbc7f2df5),
	.w7(32'hbbcc6b9a),
	.w8(32'hbb0d339d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9181c3),
	.w1(32'hbb7d347e),
	.w2(32'h3b9d82be),
	.w3(32'hbb208ac1),
	.w4(32'h3a86348d),
	.w5(32'h3b07af08),
	.w6(32'hbb2d6556),
	.w7(32'h3b352544),
	.w8(32'hba9f9263),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cb053),
	.w1(32'h3bc8137d),
	.w2(32'hbbcb4868),
	.w3(32'h3ac192ca),
	.w4(32'h3b63fbe3),
	.w5(32'hbc280d0d),
	.w6(32'h3a0beef2),
	.w7(32'hba588369),
	.w8(32'hbba72f4f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeeadc4),
	.w1(32'hbb0ceb7c),
	.w2(32'hba9fa464),
	.w3(32'hbaf7e980),
	.w4(32'hbb86c59e),
	.w5(32'hbbf126a5),
	.w6(32'hbb7f3767),
	.w7(32'hbc2a72a9),
	.w8(32'hbad6c6c7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e9b5e),
	.w1(32'hba1280eb),
	.w2(32'hbba30be5),
	.w3(32'h3b0fd8e6),
	.w4(32'hbb2eae66),
	.w5(32'h3b4651ea),
	.w6(32'hbb143089),
	.w7(32'hbbb20a05),
	.w8(32'hbaf8af35),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c8686),
	.w1(32'hbc20c6c2),
	.w2(32'hbc2ad6c6),
	.w3(32'hbccdc118),
	.w4(32'hbc539297),
	.w5(32'h3af8cd2b),
	.w6(32'hbcb95cf4),
	.w7(32'hbcd68825),
	.w8(32'hbc7e0230),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba60ba),
	.w1(32'hbbf6a8d0),
	.w2(32'h3c8ace1a),
	.w3(32'hbc1042ae),
	.w4(32'h3b0716ed),
	.w5(32'h3c9eb05a),
	.w6(32'hba41c6c9),
	.w7(32'h3bd88f84),
	.w8(32'h3c11a7d8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cbac9),
	.w1(32'h3cc621c5),
	.w2(32'hbbab9c95),
	.w3(32'h3c392359),
	.w4(32'hba23c5aa),
	.w5(32'hbbe1f6df),
	.w6(32'h3c99eb61),
	.w7(32'hbb78c280),
	.w8(32'h3b28b930),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f8248),
	.w1(32'h3a6ba134),
	.w2(32'hbb596a8e),
	.w3(32'hba0ebfdb),
	.w4(32'h3ac990ce),
	.w5(32'h3bc68a35),
	.w6(32'hba85b1ee),
	.w7(32'hba110e39),
	.w8(32'h3b2eeb2b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0214b7),
	.w1(32'hbcdd4443),
	.w2(32'h3d288e62),
	.w3(32'hbc1fd780),
	.w4(32'h3d0c2b83),
	.w5(32'hbc5b21a9),
	.w6(32'hbd2e43a1),
	.w7(32'h3d86e79c),
	.w8(32'hbcab7d0c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3e562),
	.w1(32'hbb91c62d),
	.w2(32'h3c4ce174),
	.w3(32'hbba7a642),
	.w4(32'h3b5bfa51),
	.w5(32'h3b4c7094),
	.w6(32'hbb94c95b),
	.w7(32'h3c02f85d),
	.w8(32'hbb747fe2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b25d1),
	.w1(32'hbb9e5713),
	.w2(32'h3ad4f132),
	.w3(32'hbaf284d2),
	.w4(32'h3af0d154),
	.w5(32'h3b14f05a),
	.w6(32'hbb479f68),
	.w7(32'h3b22f08c),
	.w8(32'h3a30df34),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac92d41),
	.w1(32'hbbf234f3),
	.w2(32'h3b3bcaa0),
	.w3(32'h39bf4de3),
	.w4(32'hbb826fc9),
	.w5(32'h3a790965),
	.w6(32'hbb877c6b),
	.w7(32'h39bed3af),
	.w8(32'hbb88ad28),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb849bfd),
	.w1(32'hba992c99),
	.w2(32'hb7e80d91),
	.w3(32'h3a919286),
	.w4(32'hbaa5afc1),
	.w5(32'h3bcc98c3),
	.w6(32'h3abda1c2),
	.w7(32'h3a03f150),
	.w8(32'h3b04a571),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e17bd),
	.w1(32'h3b124ea3),
	.w2(32'h3c15b697),
	.w3(32'h3b8a26a9),
	.w4(32'h3b2d9e79),
	.w5(32'h3c0c6185),
	.w6(32'h3b80410b),
	.w7(32'h3b838f6f),
	.w8(32'h3a0590be),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad670ca),
	.w1(32'h3b917a67),
	.w2(32'hbb189db1),
	.w3(32'hbca0ff48),
	.w4(32'hbcafc0b3),
	.w5(32'h3c2e5d61),
	.w6(32'hbcbbdf21),
	.w7(32'h3c38b2b3),
	.w8(32'h3b4d3b3a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc9c292),
	.w1(32'h3aad52d3),
	.w2(32'hbacef1d5),
	.w3(32'h3a07324c),
	.w4(32'hbc0601d5),
	.w5(32'hbb0f7ec1),
	.w6(32'hbad4374e),
	.w7(32'hbb94c7f8),
	.w8(32'h3b383e38),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d8553),
	.w1(32'hba0a4701),
	.w2(32'h3b34a43f),
	.w3(32'hbc43cdc2),
	.w4(32'hbce2ec8c),
	.w5(32'hbc260b6e),
	.w6(32'hbc23fbcd),
	.w7(32'hbcf33641),
	.w8(32'h3947a11c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6420e4),
	.w1(32'h3a501560),
	.w2(32'hbab2949d),
	.w3(32'h3af260cb),
	.w4(32'h3afa37cb),
	.w5(32'hbb0c001e),
	.w6(32'h3b0ad332),
	.w7(32'h39348a03),
	.w8(32'hbbee4a69),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9dc9c),
	.w1(32'h3b4c65f6),
	.w2(32'h3b0347ef),
	.w3(32'hbd09021e),
	.w4(32'h3c9be3a4),
	.w5(32'hbc1ef646),
	.w6(32'hbc3ff9a7),
	.w7(32'h3d1fd151),
	.w8(32'hbcc38214),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7891d),
	.w1(32'hbc248bb0),
	.w2(32'hbbb74735),
	.w3(32'hbc393332),
	.w4(32'hbc4350a6),
	.w5(32'hbc3284d8),
	.w6(32'hbc3275d3),
	.w7(32'hbc128cd2),
	.w8(32'hbbecaf46),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6a16a),
	.w1(32'hbd02b9e6),
	.w2(32'hbc7c470e),
	.w3(32'hbcabec5b),
	.w4(32'hbccc4f9e),
	.w5(32'h3c97ff1b),
	.w6(32'hbce54350),
	.w7(32'hbcf3cf4e),
	.w8(32'h3c9e88eb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63c037),
	.w1(32'hbb1b824b),
	.w2(32'hbc270880),
	.w3(32'hbc24a8f2),
	.w4(32'h3c780c90),
	.w5(32'hbaa38869),
	.w6(32'hbc3cc0ec),
	.w7(32'h3c5cdef6),
	.w8(32'h3ab72aab),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75f778),
	.w1(32'h3bc1cd2c),
	.w2(32'hba146c0c),
	.w3(32'h376dcfdb),
	.w4(32'h3c148718),
	.w5(32'hbab04d97),
	.w6(32'h3bc6db4e),
	.w7(32'h3bcbccff),
	.w8(32'hbc4bae82),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule