module layer_10_featuremap_421(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae484c7),
	.w1(32'hbb89534e),
	.w2(32'h39cc2e31),
	.w3(32'hbb924f0e),
	.w4(32'h3a652ed0),
	.w5(32'h398ee14e),
	.w6(32'hbba5a167),
	.w7(32'hbb6861c6),
	.w8(32'hb5e4f8a9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa16556),
	.w1(32'h3af70f05),
	.w2(32'h3b1eb7b5),
	.w3(32'hbac14ebf),
	.w4(32'h3b4ef0d8),
	.w5(32'h3a34aea7),
	.w6(32'h39e1d6da),
	.w7(32'h3a48d261),
	.w8(32'hba2a2159),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b8320),
	.w1(32'h3b7d9cc1),
	.w2(32'h3c577018),
	.w3(32'hbbc25160),
	.w4(32'h3b104d72),
	.w5(32'h3c850003),
	.w6(32'hbb00fa00),
	.w7(32'h39cb4e26),
	.w8(32'h3bc70751),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3be3d6),
	.w1(32'hbbb8ee5a),
	.w2(32'hba9d7026),
	.w3(32'h3afcf2cb),
	.w4(32'hbb5866ca),
	.w5(32'hbc295f13),
	.w6(32'h3b047577),
	.w7(32'hbba67164),
	.w8(32'hbaaaad6e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67958d),
	.w1(32'hbb178c0f),
	.w2(32'h3b595b99),
	.w3(32'hbb4ea280),
	.w4(32'hbafa1af0),
	.w5(32'h3b89cc5e),
	.w6(32'hbb813cd2),
	.w7(32'hb9e8f9e2),
	.w8(32'h397172dc),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b638045),
	.w1(32'hbbd2df88),
	.w2(32'hbc35e632),
	.w3(32'h3b831ecc),
	.w4(32'h3c090487),
	.w5(32'h3c8e688f),
	.w6(32'hbac4a2af),
	.w7(32'hba15c36a),
	.w8(32'h3a103b10),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393fda7a),
	.w1(32'hbbcbf3ce),
	.w2(32'hbc0149eb),
	.w3(32'hbbdc150d),
	.w4(32'hbb160d7d),
	.w5(32'hbb5bced0),
	.w6(32'h3a877648),
	.w7(32'hbb779bcf),
	.w8(32'hbb981af3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb499bc6),
	.w1(32'hbaffa6e2),
	.w2(32'h399f59ca),
	.w3(32'h3a0d8100),
	.w4(32'hba6bb309),
	.w5(32'h3c1c9e9f),
	.w6(32'hba966a75),
	.w7(32'h3abe8442),
	.w8(32'hbaa57b50),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf08b13),
	.w1(32'h3a3a6014),
	.w2(32'h3bc5964b),
	.w3(32'hbbe7328f),
	.w4(32'h38a1e26a),
	.w5(32'h3be2f59c),
	.w6(32'hbb665412),
	.w7(32'h3b03d6e2),
	.w8(32'h3b918de2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73deb0),
	.w1(32'hbad6ccc4),
	.w2(32'hba8428c0),
	.w3(32'hbad34184),
	.w4(32'h3bc4321d),
	.w5(32'h3ba409a3),
	.w6(32'hba375d2e),
	.w7(32'h3b7ed84d),
	.w8(32'hbacc9add),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988c627),
	.w1(32'hbb3d8392),
	.w2(32'hba9ea343),
	.w3(32'hbae5f9b7),
	.w4(32'hb9a0ee84),
	.w5(32'h3a8dd0b9),
	.w6(32'hbb77e3f3),
	.w7(32'hbb1c82bc),
	.w8(32'hb69371c6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb23a63),
	.w1(32'hbb350172),
	.w2(32'h3b168227),
	.w3(32'hbb103d80),
	.w4(32'h3b81dcba),
	.w5(32'h3c29a03b),
	.w6(32'hb9a98570),
	.w7(32'hbb3ee8f3),
	.w8(32'h37f59907),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8661dd),
	.w1(32'h3a7f4d6b),
	.w2(32'hba958975),
	.w3(32'h3c092a10),
	.w4(32'hba45c66c),
	.w5(32'hbb44c152),
	.w6(32'hbafbf3ee),
	.w7(32'h38f677b0),
	.w8(32'hbb4d7e92),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33ad37),
	.w1(32'h39971634),
	.w2(32'hba8fb37b),
	.w3(32'hbc4d7392),
	.w4(32'h389416b5),
	.w5(32'h3b2c10fd),
	.w6(32'hbc3661b9),
	.w7(32'hbb895c9c),
	.w8(32'hbb8c2024),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc302ea7),
	.w1(32'hbc3961c3),
	.w2(32'hbc139877),
	.w3(32'hbb802edd),
	.w4(32'hbb8eb052),
	.w5(32'hbc7c92dc),
	.w6(32'hbbacc002),
	.w7(32'hbb9728e8),
	.w8(32'hbbc69aef),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30910a),
	.w1(32'hbb644a98),
	.w2(32'hbc18ca8a),
	.w3(32'hbbf6be5d),
	.w4(32'hba2f59e2),
	.w5(32'hbb9b61d5),
	.w6(32'hbc41afdc),
	.w7(32'hbb11e105),
	.w8(32'hbbe3d5b4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30c23c),
	.w1(32'h3ba191a0),
	.w2(32'h3b4d15fa),
	.w3(32'hbb041c4e),
	.w4(32'h3b9149d3),
	.w5(32'hbb077d0b),
	.w6(32'hbc089b56),
	.w7(32'h39ebdb6e),
	.w8(32'h3a96203a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73b5a9),
	.w1(32'h3bc132ff),
	.w2(32'h3bd94087),
	.w3(32'h39ca75f0),
	.w4(32'h3c2a0038),
	.w5(32'h3ca9d8e2),
	.w6(32'hba59dde2),
	.w7(32'h3b38a3ac),
	.w8(32'h3b929328),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbb332),
	.w1(32'hbb5933d9),
	.w2(32'h39259e1d),
	.w3(32'h3c628900),
	.w4(32'h391a7f20),
	.w5(32'hbbab8f4f),
	.w6(32'h3c2d368e),
	.w7(32'hb8b716f7),
	.w8(32'hbb40c813),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3fe0b),
	.w1(32'hbb84e6c5),
	.w2(32'hbbc29b59),
	.w3(32'hbc010670),
	.w4(32'hb98ae740),
	.w5(32'h3c028147),
	.w6(32'hbb13bb23),
	.w7(32'hbc091615),
	.w8(32'h3b0314ce),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90a1a7),
	.w1(32'hbb83643a),
	.w2(32'h3b0eef08),
	.w3(32'hbbd88c74),
	.w4(32'h3a7b57c9),
	.w5(32'h3c33a613),
	.w6(32'hbb95c328),
	.w7(32'h3a82c095),
	.w8(32'h3b9c0fb6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70f330),
	.w1(32'hbbefbd98),
	.w2(32'h3b8cf50e),
	.w3(32'h3b63a623),
	.w4(32'hbbaee7b6),
	.w5(32'h3b66dc88),
	.w6(32'h384c68b6),
	.w7(32'hbb2df786),
	.w8(32'h3c0167a3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00d065),
	.w1(32'h39f922c2),
	.w2(32'hbb2bd9ba),
	.w3(32'hbbe6dd39),
	.w4(32'h395442af),
	.w5(32'hbb5e61df),
	.w6(32'hbbea51ef),
	.w7(32'hbbc3c274),
	.w8(32'hbc1826dd),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cacb0),
	.w1(32'h3b3072b4),
	.w2(32'h3b6f0490),
	.w3(32'hbb3d591f),
	.w4(32'h3b71b983),
	.w5(32'h3bab4d4c),
	.w6(32'hbbf252fe),
	.w7(32'hb84126c5),
	.w8(32'h3bce6cd7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fb460),
	.w1(32'h3b98d1c2),
	.w2(32'h3b97183e),
	.w3(32'h3bf87521),
	.w4(32'h3a88db63),
	.w5(32'h3ac91198),
	.w6(32'h3b336db4),
	.w7(32'h3ade82b5),
	.w8(32'h3af9042a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fffc4),
	.w1(32'hbbbc94bf),
	.w2(32'hbbb8d00e),
	.w3(32'h3c055c25),
	.w4(32'hbbe856e8),
	.w5(32'hbb51da0e),
	.w6(32'hbbae5c9d),
	.w7(32'hbc387ec1),
	.w8(32'hbbec35b9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb974ef8),
	.w1(32'hbb9d430c),
	.w2(32'hbb8e8e39),
	.w3(32'hbbb7fb82),
	.w4(32'hbbb6d679),
	.w5(32'h3b8a9a44),
	.w6(32'hbc3c6fde),
	.w7(32'h3a94cbe9),
	.w8(32'hba2a142c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb850af5),
	.w1(32'h3b9e0117),
	.w2(32'h3b2c358f),
	.w3(32'h393dba16),
	.w4(32'h3ba83177),
	.w5(32'hbb28f698),
	.w6(32'hb9f7cdce),
	.w7(32'h3ac40577),
	.w8(32'hba8983f0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68fd262),
	.w1(32'h3b023084),
	.w2(32'hbbc5ed9f),
	.w3(32'hba6621e2),
	.w4(32'hbb6211b1),
	.w5(32'h3a8ec6e0),
	.w6(32'hbb38b363),
	.w7(32'hbbd00035),
	.w8(32'hbb414200),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf293a6),
	.w1(32'h3bcafbfc),
	.w2(32'h3bd068d3),
	.w3(32'h3b4b2deb),
	.w4(32'h3b65c113),
	.w5(32'h3c6972ba),
	.w6(32'hbb03efef),
	.w7(32'h3b8467bf),
	.w8(32'h3b88c8ea),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbe244),
	.w1(32'h3b159abb),
	.w2(32'hba9ea397),
	.w3(32'h3bde845a),
	.w4(32'h3c10eeec),
	.w5(32'h3c51c98e),
	.w6(32'hbadc9a8f),
	.w7(32'hb9b01fde),
	.w8(32'hba997854),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ef4bc),
	.w1(32'hbb667b72),
	.w2(32'hbb605254),
	.w3(32'h3b6c6571),
	.w4(32'hbbe84c48),
	.w5(32'hbbb0dee2),
	.w6(32'h3884cd57),
	.w7(32'h398b8ea9),
	.w8(32'hb98f019d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc00f59),
	.w1(32'hbbf17948),
	.w2(32'hbb91bdcb),
	.w3(32'hbae0a83e),
	.w4(32'h38bca4f3),
	.w5(32'hba6de9b2),
	.w6(32'hbb59ec13),
	.w7(32'hbb46ede8),
	.w8(32'hbbe2848d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb534237),
	.w1(32'hbb18acfd),
	.w2(32'h3a2cd137),
	.w3(32'h3b4627ab),
	.w4(32'h3b35ece4),
	.w5(32'h3b9f7f49),
	.w6(32'hbb80aac9),
	.w7(32'hbba20953),
	.w8(32'hbc1e51f0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2841fa),
	.w1(32'hba83ded9),
	.w2(32'h3b6a85c7),
	.w3(32'hbb8f862a),
	.w4(32'h3c249eea),
	.w5(32'h3c95f0c4),
	.w6(32'hbc41f73c),
	.w7(32'h3bed12b0),
	.w8(32'h3baa0afb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b1649),
	.w1(32'h3ad1c37d),
	.w2(32'h3a78d351),
	.w3(32'h3b76c1cf),
	.w4(32'h3c0406ca),
	.w5(32'h3a1e3e35),
	.w6(32'h39cbfcd6),
	.w7(32'h3b09952c),
	.w8(32'h3b1cf722),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3ece9),
	.w1(32'h3b267c76),
	.w2(32'hbb50d363),
	.w3(32'hba6fa0c2),
	.w4(32'hbbf93eef),
	.w5(32'hbc21ae38),
	.w6(32'h3b89b0d0),
	.w7(32'hbb527a57),
	.w8(32'hbbfdd080),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc921b3),
	.w1(32'hbbe4fa2e),
	.w2(32'hbbe454f9),
	.w3(32'hbbc9d094),
	.w4(32'hbbdc103a),
	.w5(32'hbb4eee79),
	.w6(32'hbb95fe98),
	.w7(32'hbb6754b1),
	.w8(32'h3b0ace38),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09ee97),
	.w1(32'h3b1bcf63),
	.w2(32'h3a76429e),
	.w3(32'hbc0b8dfe),
	.w4(32'h3bcf8fe6),
	.w5(32'h3bc60374),
	.w6(32'hbc021b75),
	.w7(32'hbb62902b),
	.w8(32'h3b0d646b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f545a),
	.w1(32'h3b017606),
	.w2(32'hba5e8dcc),
	.w3(32'hbc095d27),
	.w4(32'h3ad12aaf),
	.w5(32'h39be43f3),
	.w6(32'hbbdc7f98),
	.w7(32'hbb56b874),
	.w8(32'hbb3e1aa7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e4f79),
	.w1(32'h3b236b4a),
	.w2(32'h3b5d4584),
	.w3(32'hbc2817e8),
	.w4(32'h3c184309),
	.w5(32'h3c4b896e),
	.w6(32'hbc2e1973),
	.w7(32'h3bcc4741),
	.w8(32'h3c0ff082),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b994ec8),
	.w1(32'hbbf67f09),
	.w2(32'hbb443d04),
	.w3(32'h3c1707ab),
	.w4(32'hbbd0b5d7),
	.w5(32'h3a9c905c),
	.w6(32'h3bc1b450),
	.w7(32'hbbb755de),
	.w8(32'hbbaf5ae7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5802e8),
	.w1(32'hbc029277),
	.w2(32'hbb79043d),
	.w3(32'hbc0743d4),
	.w4(32'hbc1367f2),
	.w5(32'h36e28ffa),
	.w6(32'hbc1ae30c),
	.w7(32'hbbe5f3a7),
	.w8(32'hbb872043),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c08c28),
	.w1(32'h380af243),
	.w2(32'h3ba59620),
	.w3(32'hb9c4a6d3),
	.w4(32'h3b871b76),
	.w5(32'h3c2fe5be),
	.w6(32'hbabae5ea),
	.w7(32'hba837c3f),
	.w8(32'h3ad44c13),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb186849),
	.w1(32'hbc27e566),
	.w2(32'hbac71fa3),
	.w3(32'hba8b658a),
	.w4(32'hbbbde4ab),
	.w5(32'h3aa7d098),
	.w6(32'hbb9ed4cc),
	.w7(32'hbaefe512),
	.w8(32'h3a20d2bd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f651c),
	.w1(32'hbb9d9cab),
	.w2(32'hbb9bb568),
	.w3(32'hba5cc5f8),
	.w4(32'hb9c06535),
	.w5(32'h3a8d96ae),
	.w6(32'hbb057401),
	.w7(32'hbb8e9ad0),
	.w8(32'hbae4e081),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc3b28),
	.w1(32'hbb7eda3a),
	.w2(32'hbba1dc20),
	.w3(32'h3b199b11),
	.w4(32'h39f5d4eb),
	.w5(32'hbbf952bb),
	.w6(32'hbb82104c),
	.w7(32'h393b358d),
	.w8(32'hbb90ec39),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc533578),
	.w1(32'hba71255e),
	.w2(32'h3aeff0aa),
	.w3(32'hba9a8c0b),
	.w4(32'h3b70d772),
	.w5(32'hb859e557),
	.w6(32'hbadcac62),
	.w7(32'hbb498448),
	.w8(32'h3abb108a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb740b2),
	.w1(32'hbac5067a),
	.w2(32'hbc06457b),
	.w3(32'hbc165212),
	.w4(32'h3a307dd7),
	.w5(32'hba2dd814),
	.w6(32'hbc067613),
	.w7(32'h3b54efa3),
	.w8(32'hb9b51f89),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3ad71),
	.w1(32'hbb0a320d),
	.w2(32'hbc15f07d),
	.w3(32'h3ba0bc07),
	.w4(32'h3b5fb5ba),
	.w5(32'h3a5994ba),
	.w6(32'h3ace819c),
	.w7(32'h3be434f5),
	.w8(32'h398e1772),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52fdd),
	.w1(32'hbb65f07a),
	.w2(32'hbae55323),
	.w3(32'hb77bfdd9),
	.w4(32'hbbd68d38),
	.w5(32'hbba9d477),
	.w6(32'h3afc2dc6),
	.w7(32'hbbce8211),
	.w8(32'hbbb6d283),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf68ef8),
	.w1(32'hba8ad8b0),
	.w2(32'hbbe2a2db),
	.w3(32'hbc17609b),
	.w4(32'hbaed3a30),
	.w5(32'hbc304fb0),
	.w6(32'hbbc95f04),
	.w7(32'hbabf73a2),
	.w8(32'hbb95f052),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba605f41),
	.w1(32'h3be3660b),
	.w2(32'h3bb1afda),
	.w3(32'hbb2e9dd6),
	.w4(32'h3c417520),
	.w5(32'h3c756dcc),
	.w6(32'h3aee33a9),
	.w7(32'h3c063da2),
	.w8(32'hba54f6b0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4762),
	.w1(32'hbae2b554),
	.w2(32'h3935a930),
	.w3(32'h3c0c26a2),
	.w4(32'hb9ea6077),
	.w5(32'h3c1c6e94),
	.w6(32'h3ab97a3d),
	.w7(32'hb9fddf59),
	.w8(32'h3b12e5f5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33030c),
	.w1(32'h38824f2e),
	.w2(32'h3afa308a),
	.w3(32'h3b94a54a),
	.w4(32'hbb562370),
	.w5(32'h3b9c7378),
	.w6(32'h3a9c14aa),
	.w7(32'hba86ef21),
	.w8(32'h3b16a636),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bfd91),
	.w1(32'hbc31b6c2),
	.w2(32'hbbdae6c7),
	.w3(32'hbacec838),
	.w4(32'hbc1a44b1),
	.w5(32'h3b0afbf0),
	.w6(32'hbb361e50),
	.w7(32'hbc1dce7a),
	.w8(32'hba834568),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e6228),
	.w1(32'hbb694721),
	.w2(32'hbb8d7f72),
	.w3(32'hbbb68014),
	.w4(32'hbb1cfbed),
	.w5(32'hbba4c2f8),
	.w6(32'hbb3731cd),
	.w7(32'hbb953fa8),
	.w8(32'hbbba853b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26d95f),
	.w1(32'hba0dbdd5),
	.w2(32'hbb765c09),
	.w3(32'hbb2f7ed4),
	.w4(32'h3b8ea979),
	.w5(32'h3a56e61e),
	.w6(32'hbb6184ba),
	.w7(32'h3b743478),
	.w8(32'h3a970f3a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb769ffb),
	.w1(32'hbbc2fe4a),
	.w2(32'hbb57bdb1),
	.w3(32'hbb9432fc),
	.w4(32'hbc087834),
	.w5(32'h3a8c05d9),
	.w6(32'hbbec296b),
	.w7(32'hbba604ce),
	.w8(32'hbb6c99df),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc605e4),
	.w1(32'h3b900d92),
	.w2(32'h3a9993d1),
	.w3(32'h3bea5123),
	.w4(32'h3b26f4fd),
	.w5(32'hbbf15d48),
	.w6(32'h3ad68548),
	.w7(32'hbbb32529),
	.w8(32'h3a41853c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd84b81),
	.w1(32'hb9e35dce),
	.w2(32'h3b24e63a),
	.w3(32'hba846fb4),
	.w4(32'hbbd3f8f7),
	.w5(32'hbb0e2e86),
	.w6(32'hbbbe2480),
	.w7(32'hbc185b4f),
	.w8(32'hbb4ab37d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2a16c),
	.w1(32'hbb5851f8),
	.w2(32'h3b98cf40),
	.w3(32'hbb03612f),
	.w4(32'hbbe99a68),
	.w5(32'h3ba598ea),
	.w6(32'hbbcc587b),
	.w7(32'hbb8da307),
	.w8(32'h3a1d9477),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993276f),
	.w1(32'hbb8f09fe),
	.w2(32'h39e9abd4),
	.w3(32'hb996b94f),
	.w4(32'hbad5c70c),
	.w5(32'h3a0624c1),
	.w6(32'h3b65f5e0),
	.w7(32'h3a639296),
	.w8(32'h3bf4b512),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c367763),
	.w1(32'hbc2f3a3c),
	.w2(32'hbc20894b),
	.w3(32'h3c9e17e5),
	.w4(32'hbc12c04e),
	.w5(32'hbbb0d5b6),
	.w6(32'h3c4378ee),
	.w7(32'hbc2b10ff),
	.w8(32'hbbdbe778),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbded5cc),
	.w1(32'hbc9e4ae0),
	.w2(32'hbca77f46),
	.w3(32'hb8ad4f6e),
	.w4(32'hbba22f05),
	.w5(32'hbb5432f9),
	.w6(32'hbb8c95fa),
	.w7(32'hbb9150ab),
	.w8(32'hbaeda18a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e0938),
	.w1(32'hbb043738),
	.w2(32'h3b7e4896),
	.w3(32'hbb9921f6),
	.w4(32'h3a92a543),
	.w5(32'h3c070dfa),
	.w6(32'hbb0f1b2a),
	.w7(32'hbb2485e1),
	.w8(32'hbb08b947),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ae22e),
	.w1(32'h3bdbbb5f),
	.w2(32'h3b8dad49),
	.w3(32'h3b0291af),
	.w4(32'hbaec8b0d),
	.w5(32'h3b1d3b14),
	.w6(32'h3b8716e7),
	.w7(32'hbc147fc3),
	.w8(32'hbc6c7ef5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9b405),
	.w1(32'h3ad8bea0),
	.w2(32'h3b1acbb0),
	.w3(32'hbc2e4de5),
	.w4(32'hbb07958f),
	.w5(32'h3ba86b1f),
	.w6(32'hbc508c39),
	.w7(32'hbc0c14c9),
	.w8(32'hbbe50ebc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03450f),
	.w1(32'hbbfed450),
	.w2(32'h3afd3272),
	.w3(32'h3bca6aaf),
	.w4(32'hbbbb4d2f),
	.w5(32'hbb6f76af),
	.w6(32'h3a908a5f),
	.w7(32'h39554989),
	.w8(32'h3b581be4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb0da8),
	.w1(32'hbc35154f),
	.w2(32'hbb28b206),
	.w3(32'h3a32eb8c),
	.w4(32'hbc0ffbbe),
	.w5(32'hbb14aace),
	.w6(32'h3a8377f1),
	.w7(32'hbc268ca5),
	.w8(32'hbb3d4bc5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5b9fa),
	.w1(32'h3c26aa2f),
	.w2(32'h3babe86d),
	.w3(32'h3aa4b0b1),
	.w4(32'h3b8212ce),
	.w5(32'hbae3d087),
	.w6(32'hbaa6baa9),
	.w7(32'h3b9a8748),
	.w8(32'h3bb110ba),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b930965),
	.w1(32'h3ac25687),
	.w2(32'hbc072d7c),
	.w3(32'h3b231515),
	.w4(32'h3b168c72),
	.w5(32'h3b982761),
	.w6(32'h3c5e1606),
	.w7(32'h3bc158ec),
	.w8(32'h3c3768d4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1615b8),
	.w1(32'h3bb7b772),
	.w2(32'h3bb56b60),
	.w3(32'h3c1e6030),
	.w4(32'h3b361fbb),
	.w5(32'h3b2ffdbd),
	.w6(32'h3b71aa0b),
	.w7(32'hb93e4688),
	.w8(32'h3bdd9144),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af13ee0),
	.w1(32'hbb3bcb21),
	.w2(32'hbb83b111),
	.w3(32'hbb33da9c),
	.w4(32'hbb9417c6),
	.w5(32'hbb218161),
	.w6(32'h3b43c71d),
	.w7(32'hbbd7e312),
	.w8(32'hba44a95c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc045bc7),
	.w1(32'hbb5a3e33),
	.w2(32'hbaf3a8a0),
	.w3(32'hbbb26753),
	.w4(32'hbb1bde25),
	.w5(32'h3b84b067),
	.w6(32'h3a27a4b2),
	.w7(32'h37144609),
	.w8(32'hbbc6b248),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6149ca),
	.w1(32'hbb4cb71c),
	.w2(32'hbb6a6bc3),
	.w3(32'h3b8c8e85),
	.w4(32'hbc0cd91a),
	.w5(32'hbb445a3b),
	.w6(32'hbb39ff08),
	.w7(32'hbbbd9a88),
	.w8(32'hba1a8b29),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89bedd),
	.w1(32'hbc09b192),
	.w2(32'hbbdabb34),
	.w3(32'hbb98e617),
	.w4(32'hbc412074),
	.w5(32'hbc96b4b6),
	.w6(32'hbb319f09),
	.w7(32'hbb427556),
	.w8(32'hbba8ea53),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4e59a),
	.w1(32'hbc19078b),
	.w2(32'hbc5dc4d7),
	.w3(32'h39ee8e51),
	.w4(32'h3bff5b32),
	.w5(32'h3beacec0),
	.w6(32'h3aceb306),
	.w7(32'h3c031ff7),
	.w8(32'h3c0b3db4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92adbd),
	.w1(32'h397fb27a),
	.w2(32'h3beddd13),
	.w3(32'h3a8a37aa),
	.w4(32'hbb66f3ce),
	.w5(32'hbb3b5445),
	.w6(32'hbb646e7a),
	.w7(32'h3b254c02),
	.w8(32'h3aa5faeb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ec253),
	.w1(32'hbba3cd4f),
	.w2(32'h3abf1c5c),
	.w3(32'h3bcb19c4),
	.w4(32'hbbb7ab8f),
	.w5(32'hbab50e2b),
	.w6(32'h3b84efc6),
	.w7(32'h39c4247e),
	.w8(32'hbb3b4be7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b1f72),
	.w1(32'h3a86c77f),
	.w2(32'h3b89da0c),
	.w3(32'h3c1b350d),
	.w4(32'hbb11ede7),
	.w5(32'hbb5f61f6),
	.w6(32'h3aec484a),
	.w7(32'h3b4c6be6),
	.w8(32'h3bb5dff2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be92f0f),
	.w1(32'h3ba6be24),
	.w2(32'hbbb86585),
	.w3(32'h3bb6be3a),
	.w4(32'h3c65bf38),
	.w5(32'hb9cad88d),
	.w6(32'h3b766405),
	.w7(32'h3c64aebb),
	.w8(32'h3c1ab51c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8f73e),
	.w1(32'h3bd94269),
	.w2(32'h3bdaa472),
	.w3(32'hbb9d638f),
	.w4(32'h3a10246c),
	.w5(32'hbb04fc8a),
	.w6(32'h3b3a5949),
	.w7(32'hbc30d614),
	.w8(32'hbc304873),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e742a),
	.w1(32'h3c562390),
	.w2(32'h3c678a4a),
	.w3(32'hbbbe6e22),
	.w4(32'h3c3a027d),
	.w5(32'h3c44b43a),
	.w6(32'hbc003af2),
	.w7(32'h3b6b7e28),
	.w8(32'h3b98b235),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cbe74),
	.w1(32'hba83ed35),
	.w2(32'hbc11410a),
	.w3(32'h3bb2bd03),
	.w4(32'h3ad0bdea),
	.w5(32'hbaf82c29),
	.w6(32'h3c2eb889),
	.w7(32'h3bfd55e3),
	.w8(32'h3b90f3be),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab705bd),
	.w1(32'h3b167d45),
	.w2(32'h3c6a2d6c),
	.w3(32'h3b5dc3a2),
	.w4(32'h3bbdc1eb),
	.w5(32'h3bbb93d1),
	.w6(32'h3c117325),
	.w7(32'hbc2d7c75),
	.w8(32'hbc03a961),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68f5c5),
	.w1(32'hba9798e2),
	.w2(32'h3b999e46),
	.w3(32'hbc335cbd),
	.w4(32'hbbc31a43),
	.w5(32'hbab1e453),
	.w6(32'hbbe65f6f),
	.w7(32'hb9a68ab0),
	.w8(32'hbbf1b67a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba082076),
	.w1(32'h3b69a155),
	.w2(32'h3c279666),
	.w3(32'h39ff792b),
	.w4(32'hbc0fa240),
	.w5(32'h3969d9aa),
	.w6(32'hbbe9edff),
	.w7(32'hbc57b30a),
	.w8(32'hbc9c1a62),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da02a7),
	.w1(32'hba0a2811),
	.w2(32'hbbe26178),
	.w3(32'hbbbcb19f),
	.w4(32'hbbb700bc),
	.w5(32'hbc2dae1b),
	.w6(32'hbbd28d05),
	.w7(32'hb94fe63b),
	.w8(32'hbbcff4c9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b5a8a),
	.w1(32'hbabd1e1e),
	.w2(32'hbb793b57),
	.w3(32'h3a1b84f0),
	.w4(32'h3b5cb375),
	.w5(32'hbb4f5f3b),
	.w6(32'hb9c85c8e),
	.w7(32'h3b0daa0b),
	.w8(32'h3a930972),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb022e0),
	.w1(32'h3b550d23),
	.w2(32'h3b2f1337),
	.w3(32'hbb0b11b3),
	.w4(32'h3bff8bea),
	.w5(32'h3bd7cca8),
	.w6(32'h3ae0def8),
	.w7(32'h3b81dda6),
	.w8(32'hbabd0842),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89674d),
	.w1(32'hbbab27b5),
	.w2(32'hbbc56c86),
	.w3(32'hbb8096a8),
	.w4(32'hbbd8d574),
	.w5(32'hbb18dff2),
	.w6(32'hbb3fb5d5),
	.w7(32'h3abe11de),
	.w8(32'h3b71e104),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad972be),
	.w1(32'h3bc488dd),
	.w2(32'h3ab63769),
	.w3(32'hbb2e0a0f),
	.w4(32'hbad72a83),
	.w5(32'h3a1f5f06),
	.w6(32'h3b9cf48c),
	.w7(32'h3aefa4ea),
	.w8(32'h3c05f8e1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb89839),
	.w1(32'h3a64e8fe),
	.w2(32'h3a32795a),
	.w3(32'h38810c67),
	.w4(32'hbac02095),
	.w5(32'hbbc37414),
	.w6(32'h3bb691c3),
	.w7(32'hbb8fac20),
	.w8(32'hbb976a06),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b4eec),
	.w1(32'h3b845e41),
	.w2(32'h3b0b50b6),
	.w3(32'hb9789c95),
	.w4(32'hbb947845),
	.w5(32'h3adf4868),
	.w6(32'h397341b2),
	.w7(32'h3bd2826a),
	.w8(32'hb96a482e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d3d47),
	.w1(32'hbbeab187),
	.w2(32'hba50d52d),
	.w3(32'h3c515da3),
	.w4(32'hbbba8263),
	.w5(32'h3c1a8774),
	.w6(32'h3c7bc083),
	.w7(32'hbc63d70b),
	.w8(32'hbb83ca77),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32bf7b),
	.w1(32'h3b6d5be5),
	.w2(32'h384a562b),
	.w3(32'h3b874e91),
	.w4(32'hba5d5b00),
	.w5(32'hbc25fdfc),
	.w6(32'hbadd0a25),
	.w7(32'hbbe01094),
	.w8(32'hbc5cff38),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cd480),
	.w1(32'hbb0b3ebd),
	.w2(32'h3b865340),
	.w3(32'hbb65264d),
	.w4(32'hbc1dd261),
	.w5(32'h3ba72447),
	.w6(32'hbb2c7ca7),
	.w7(32'hbbe3d7c5),
	.w8(32'h39bb2b6c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb712e9b1),
	.w1(32'h3c12f3ee),
	.w2(32'h3c0b30e0),
	.w3(32'hbb200f59),
	.w4(32'h3bfb36e0),
	.w5(32'h3b781ed9),
	.w6(32'h3b18c45f),
	.w7(32'h3c0c99e3),
	.w8(32'h3a1af861),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c682b69),
	.w1(32'h3bcd9c8b),
	.w2(32'h3bf8d917),
	.w3(32'h3c36d4b2),
	.w4(32'h3b97f968),
	.w5(32'h3c903d4e),
	.w6(32'h3c432962),
	.w7(32'h3be07325),
	.w8(32'h3a2cf194),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7febf),
	.w1(32'h3bd71afe),
	.w2(32'h3bf76d68),
	.w3(32'h3c13639f),
	.w4(32'hbb8da280),
	.w5(32'hbba29842),
	.w6(32'hbb9b5796),
	.w7(32'hbb6d2413),
	.w8(32'hbbb76d13),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c8133),
	.w1(32'hb99af2a9),
	.w2(32'hb8ac7c0c),
	.w3(32'hbabea696),
	.w4(32'hb976792c),
	.w5(32'h3b54fe2d),
	.w6(32'h3b2ed6a9),
	.w7(32'h3b1c2a7b),
	.w8(32'hba081431),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e5f06),
	.w1(32'hbabc461d),
	.w2(32'h3a30cc5a),
	.w3(32'hbb3e6094),
	.w4(32'hbb464516),
	.w5(32'h3977b3f5),
	.w6(32'h3b0aed30),
	.w7(32'hbadc63f6),
	.w8(32'hbbbbfbd2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaad595),
	.w1(32'h3ace9e74),
	.w2(32'hbc0b1824),
	.w3(32'hbae3c0f3),
	.w4(32'h3ba24270),
	.w5(32'hbba0024a),
	.w6(32'h3b47929d),
	.w7(32'h3c0b53cb),
	.w8(32'hba97659f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd25800),
	.w1(32'h38c751d5),
	.w2(32'h3b2c5e6e),
	.w3(32'hb91e1a32),
	.w4(32'hbb27d002),
	.w5(32'h3ad7da8b),
	.w6(32'hbac2aa64),
	.w7(32'hbc1e8d74),
	.w8(32'hbbec895e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91b96e),
	.w1(32'h3c4182b1),
	.w2(32'h3c071eb6),
	.w3(32'hbbc091ee),
	.w4(32'h3c0b06b0),
	.w5(32'h3af9f138),
	.w6(32'hbba2771e),
	.w7(32'hbab43e03),
	.w8(32'hbba61eb7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97d9f0),
	.w1(32'hbb3b0df1),
	.w2(32'hbb2a2d63),
	.w3(32'hbb08ee1e),
	.w4(32'h3b011c62),
	.w5(32'hbb91a85a),
	.w6(32'hbbdb2f30),
	.w7(32'hba037a47),
	.w8(32'h3b08ed00),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d0ea2),
	.w1(32'h3b42d635),
	.w2(32'h3c2f9c0e),
	.w3(32'hbb4b48d9),
	.w4(32'hbb6e6be6),
	.w5(32'h3bf3eef3),
	.w6(32'hba2add4c),
	.w7(32'hbba2463b),
	.w8(32'hbaacac94),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d52d),
	.w1(32'h3b02db1d),
	.w2(32'hbb101304),
	.w3(32'h3b369471),
	.w4(32'hbb5b3cd3),
	.w5(32'h3b39cd2d),
	.w6(32'hbb48a18d),
	.w7(32'hbc06c322),
	.w8(32'hbbb9bb3f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b767e39),
	.w1(32'h3b6de432),
	.w2(32'h38598162),
	.w3(32'h3a9f1d95),
	.w4(32'hbb88a02f),
	.w5(32'h3bcda875),
	.w6(32'hbb93dd59),
	.w7(32'hbc054c14),
	.w8(32'hbc305976),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a64f9),
	.w1(32'hb88be174),
	.w2(32'hb9e706e2),
	.w3(32'hbb045de3),
	.w4(32'hbb319434),
	.w5(32'hbbfc814c),
	.w6(32'hbc2eba6b),
	.w7(32'hbb78169b),
	.w8(32'h3a8fc185),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba16be1),
	.w1(32'hbb1797f4),
	.w2(32'hbc530c79),
	.w3(32'hbb9ba048),
	.w4(32'h3c3cc570),
	.w5(32'hbb96c16c),
	.w6(32'h3bc8f459),
	.w7(32'h3b03ff6d),
	.w8(32'hbb0b228a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a620a),
	.w1(32'h3b427551),
	.w2(32'h3b95aa26),
	.w3(32'hbc8244e6),
	.w4(32'h3b951c9e),
	.w5(32'h3b546b7c),
	.w6(32'hbc044f3b),
	.w7(32'hbb5ddef4),
	.w8(32'hbafab347),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cf37c),
	.w1(32'hbaed5e87),
	.w2(32'hbb5fe9cc),
	.w3(32'hbbf1f52a),
	.w4(32'h3ab709d4),
	.w5(32'hbb2ffe9d),
	.w6(32'hba31560c),
	.w7(32'h3b1a9ac3),
	.w8(32'h3ac47f49),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b089c25),
	.w1(32'h3b985c8d),
	.w2(32'h3b865e40),
	.w3(32'h3b2c748e),
	.w4(32'h3b4ae41b),
	.w5(32'hba631a0f),
	.w6(32'h3bc0b545),
	.w7(32'hbbff6e3c),
	.w8(32'hbbaffb87),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407574),
	.w1(32'h3bead4b7),
	.w2(32'hbb8484ad),
	.w3(32'h39b3e05f),
	.w4(32'h3ba19e6d),
	.w5(32'hbc81994f),
	.w6(32'h3b384c99),
	.w7(32'hba7834d0),
	.w8(32'hbbbf8f82),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83af79),
	.w1(32'h3b3007e7),
	.w2(32'hbb2f9b70),
	.w3(32'hbbd28ef3),
	.w4(32'h3c053e33),
	.w5(32'h3c3daac4),
	.w6(32'hbadb2d9f),
	.w7(32'h39b12ed9),
	.w8(32'h3bf16017),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f3152),
	.w1(32'hbbb898ef),
	.w2(32'hbc23ab92),
	.w3(32'hbb36dc6e),
	.w4(32'hba03ecd7),
	.w5(32'hbae736de),
	.w6(32'hbad8a45c),
	.w7(32'h3b86feee),
	.w8(32'h3bfd7811),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bec1b),
	.w1(32'hbba734cd),
	.w2(32'hbb94e003),
	.w3(32'hb87a07da),
	.w4(32'hbb85338b),
	.w5(32'h39f668d9),
	.w6(32'h3b8ce5f3),
	.w7(32'h3aec4637),
	.w8(32'h3bf36906),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936c37),
	.w1(32'h3ab5e522),
	.w2(32'h3a2a43dd),
	.w3(32'hbae33e15),
	.w4(32'h3aa6a6ba),
	.w5(32'h3b36c416),
	.w6(32'h3ba57a39),
	.w7(32'h3b3c15b5),
	.w8(32'hbb194ef9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31f62f),
	.w1(32'hbb82402c),
	.w2(32'hbb8f5091),
	.w3(32'hbadeeda8),
	.w4(32'hbb9917d3),
	.w5(32'hbc339bbc),
	.w6(32'hb9cfbd26),
	.w7(32'hbb6d3424),
	.w8(32'h3b0a1148),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9cfb0),
	.w1(32'hbbf057e8),
	.w2(32'hbaaf77db),
	.w3(32'hba817a1a),
	.w4(32'hbb30b3f3),
	.w5(32'h3be1e6ce),
	.w6(32'h3bcfed56),
	.w7(32'hbb6bdf1a),
	.w8(32'h39156cec),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7761a),
	.w1(32'hbad6e393),
	.w2(32'h3a2920e6),
	.w3(32'h3ae663cd),
	.w4(32'h3a2f7439),
	.w5(32'hbc35aea7),
	.w6(32'hbb5870f2),
	.w7(32'hbb9d96d7),
	.w8(32'hbc1c4a25),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc138a4),
	.w1(32'h3a604955),
	.w2(32'hbb88d689),
	.w3(32'hbc346853),
	.w4(32'h3c3f1474),
	.w5(32'h3ba8d1dc),
	.w6(32'h39911622),
	.w7(32'h3bab7cb6),
	.w8(32'h3b8e092e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb0143),
	.w1(32'hbc2a50ce),
	.w2(32'hbc8e2310),
	.w3(32'hbbc6b848),
	.w4(32'hbb10c48a),
	.w5(32'h3b9c9ed3),
	.w6(32'h3a8176b0),
	.w7(32'h3c24c397),
	.w8(32'h3c8c44c0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9ef95),
	.w1(32'h3b70d98d),
	.w2(32'hb92755f2),
	.w3(32'hbaef1e74),
	.w4(32'hb97a1509),
	.w5(32'h3b11336c),
	.w6(32'h3bc052c1),
	.w7(32'hbb1cd8e3),
	.w8(32'h3b3645a8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a6bd1),
	.w1(32'hbc077dae),
	.w2(32'hbc35e28b),
	.w3(32'h3becab6d),
	.w4(32'hbbae98aa),
	.w5(32'hbbbeb2a1),
	.w6(32'h3c0fac33),
	.w7(32'hbc2b4b9a),
	.w8(32'hbc6a4d12),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa8d9e),
	.w1(32'hbab2537d),
	.w2(32'h3b02d01e),
	.w3(32'hbc6e76b8),
	.w4(32'h37b7d56c),
	.w5(32'hbadba13c),
	.w6(32'hbc8ced65),
	.w7(32'hbb9b48ac),
	.w8(32'hbb371844),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a138aa3),
	.w1(32'hbbc364fb),
	.w2(32'h3bba4b08),
	.w3(32'hbbcc8430),
	.w4(32'hbc677b8c),
	.w5(32'hbb1c1d81),
	.w6(32'hb9312f67),
	.w7(32'hbc2224e1),
	.w8(32'hbbe37f90),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf3ac3),
	.w1(32'hbb00d743),
	.w2(32'h38f68811),
	.w3(32'h3ca5905c),
	.w4(32'h3a10ed53),
	.w5(32'h3b0ded53),
	.w6(32'h3b944b97),
	.w7(32'h3b5f1f62),
	.w8(32'hba72fd81),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7142f8),
	.w1(32'h3ace8be9),
	.w2(32'h3aed1de7),
	.w3(32'hba8f47e6),
	.w4(32'h3b36c4dc),
	.w5(32'h3b4a27f5),
	.w6(32'hbab0979d),
	.w7(32'hbb43ef81),
	.w8(32'h3b417a3c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f2554),
	.w1(32'h39daed93),
	.w2(32'hbb3ce97c),
	.w3(32'hba598bd7),
	.w4(32'hbb6c9d47),
	.w5(32'hbaea7deb),
	.w6(32'hb8e74214),
	.w7(32'hbbb7c5c7),
	.w8(32'hbbff897a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67ba1e),
	.w1(32'h3aeb3c1d),
	.w2(32'hba3399b3),
	.w3(32'hbafd04db),
	.w4(32'h3b1c4198),
	.w5(32'h3b14eb22),
	.w6(32'hbbb6d6e0),
	.w7(32'hbb9055b0),
	.w8(32'hbb0e9d8d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4332e),
	.w1(32'h3c258996),
	.w2(32'h3b05319f),
	.w3(32'h3a397312),
	.w4(32'h3c3c89c0),
	.w5(32'h3c317789),
	.w6(32'h3b76b0b0),
	.w7(32'h3be4b3d4),
	.w8(32'hba69746b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0268fa),
	.w1(32'hbaaed1d5),
	.w2(32'hbb843eed),
	.w3(32'hbba4d81e),
	.w4(32'hbbb344b7),
	.w5(32'h39c1467b),
	.w6(32'hbbb53a88),
	.w7(32'hbc1f7439),
	.w8(32'h3b581e79),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4fe86),
	.w1(32'h3b00f60f),
	.w2(32'hbaf96494),
	.w3(32'hbb4175ec),
	.w4(32'h3bbf2fcd),
	.w5(32'hbbd5b253),
	.w6(32'hbb1c2b98),
	.w7(32'h3bc0ac9d),
	.w8(32'h3b4a68c5),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca172e),
	.w1(32'hbb9c71c6),
	.w2(32'h3b143872),
	.w3(32'hbc015fae),
	.w4(32'hbb810086),
	.w5(32'h3a8c7859),
	.w6(32'h3b1decac),
	.w7(32'hbb6e90db),
	.w8(32'hbb7cb1cc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44f232),
	.w1(32'h3c0790e6),
	.w2(32'h3c1b56cf),
	.w3(32'h3a9ee737),
	.w4(32'h3b5dbb3f),
	.w5(32'h3c191f56),
	.w6(32'hbb85a74d),
	.w7(32'hb9a55890),
	.w8(32'hbbb6f89e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44fba1),
	.w1(32'hba9029cb),
	.w2(32'h3b987d95),
	.w3(32'hba8d14e6),
	.w4(32'hbb06d55a),
	.w5(32'h3b3e3637),
	.w6(32'hbba10ebf),
	.w7(32'hbaf9d146),
	.w8(32'hbb4a4b96),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b184dac),
	.w1(32'h3a09a7ae),
	.w2(32'hbc42abb1),
	.w3(32'hba88d689),
	.w4(32'h3b84957c),
	.w5(32'hbc9a4346),
	.w6(32'h3aab4c6a),
	.w7(32'h3c4aa189),
	.w8(32'h3bf3785b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf268d5),
	.w1(32'hba6d7992),
	.w2(32'hbb8db049),
	.w3(32'hbc163952),
	.w4(32'h3c114417),
	.w5(32'hbc00ec52),
	.w6(32'h3bb61438),
	.w7(32'hbbabe882),
	.w8(32'hbb93c085),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3cc9),
	.w1(32'hba803de0),
	.w2(32'h3bced7ed),
	.w3(32'hbba59a93),
	.w4(32'hbc1d96a0),
	.w5(32'h3afb77b6),
	.w6(32'h3a900b2e),
	.w7(32'hbc875b2a),
	.w8(32'hbc588902),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4b37b),
	.w1(32'hbbe51a53),
	.w2(32'hbc5f7288),
	.w3(32'hbb48dad6),
	.w4(32'h3b805088),
	.w5(32'hba2ac9ba),
	.w6(32'hbc2dec53),
	.w7(32'h3ba9e246),
	.w8(32'h3b90a27a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f7fb5),
	.w1(32'hbb14bca9),
	.w2(32'hbbfb00d2),
	.w3(32'hbb5c7bd9),
	.w4(32'h3a403775),
	.w5(32'hbc6cfe72),
	.w6(32'h3b4acecf),
	.w7(32'h3ba946e7),
	.w8(32'h3c063241),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50cbdf),
	.w1(32'hbc419c41),
	.w2(32'hbc7026da),
	.w3(32'h3bd4d69e),
	.w4(32'hbb382a4a),
	.w5(32'hbbfa8f49),
	.w6(32'h3c551323),
	.w7(32'h3c4ca08e),
	.w8(32'h3c0dc5be),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafae6b5),
	.w1(32'hbc603a9e),
	.w2(32'hb9ebd0ad),
	.w3(32'hbb443961),
	.w4(32'hbc789c3e),
	.w5(32'h399e1499),
	.w6(32'h3b994383),
	.w7(32'hbbae94ed),
	.w8(32'h3b1f0fdc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95f324),
	.w1(32'hba4a80b9),
	.w2(32'hbba631b5),
	.w3(32'h3ca49893),
	.w4(32'h3a28fd2d),
	.w5(32'hbc12609c),
	.w6(32'h3c8b2e68),
	.w7(32'h3b9af451),
	.w8(32'h3af7ea89),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb430b0d),
	.w1(32'h3c042448),
	.w2(32'hbb19ffa3),
	.w3(32'hbb8d2832),
	.w4(32'h3c3eb291),
	.w5(32'h3be7aade),
	.w6(32'h3be643a0),
	.w7(32'h3c4df168),
	.w8(32'h3c1ab8f6),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b7d0a),
	.w1(32'h3b8336bc),
	.w2(32'hbb302ee8),
	.w3(32'h3c067944),
	.w4(32'h3b74bd3a),
	.w5(32'hbbeb6f05),
	.w6(32'h3c1b7a76),
	.w7(32'h3b07dbaa),
	.w8(32'hbb646298),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe99f2d),
	.w1(32'h3a168994),
	.w2(32'h39eaae9c),
	.w3(32'hbc6ff844),
	.w4(32'h3b8819e3),
	.w5(32'h3baa97fc),
	.w6(32'hbbe68a65),
	.w7(32'hbbc58130),
	.w8(32'hbb8f7056),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4495f6),
	.w1(32'hbbefa6f4),
	.w2(32'h360d0f25),
	.w3(32'hbbb3b6c2),
	.w4(32'h3a549cbd),
	.w5(32'h3bcae360),
	.w6(32'h3b1eed84),
	.w7(32'h3b9ee7af),
	.w8(32'h3b885c22),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973c56),
	.w1(32'h3b16c08b),
	.w2(32'h3bed8a4d),
	.w3(32'hbb7b5d45),
	.w4(32'h3c2787a4),
	.w5(32'h3c639860),
	.w6(32'hb9dd6f26),
	.w7(32'h3baf7b6e),
	.w8(32'h3c07cbc3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb089e7d),
	.w1(32'hbb144364),
	.w2(32'hbb6941a5),
	.w3(32'h3b2f2985),
	.w4(32'h3b71b0e9),
	.w5(32'h3bcb7d61),
	.w6(32'hbb9969a3),
	.w7(32'hbc675271),
	.w8(32'hbc8e7047),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc801948),
	.w1(32'h3b899a10),
	.w2(32'hba064ba0),
	.w3(32'hbc9d6e0e),
	.w4(32'hbafcadab),
	.w5(32'hbbe6ba3a),
	.w6(32'hbca94b7c),
	.w7(32'hbae6b40e),
	.w8(32'hbb8cb8ab),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fa40c),
	.w1(32'hba6368e3),
	.w2(32'hbaa7106b),
	.w3(32'hbc095575),
	.w4(32'hbc445f65),
	.w5(32'hbb94ef2e),
	.w6(32'hbab6c204),
	.w7(32'h3b1f469f),
	.w8(32'h3b92b579),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba576d37),
	.w1(32'hbb8968a5),
	.w2(32'h3b3c849d),
	.w3(32'hbab00aa7),
	.w4(32'hbb0872fb),
	.w5(32'h3c182a7e),
	.w6(32'h3be095c6),
	.w7(32'hbb1f13fb),
	.w8(32'hb903f905),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b5696),
	.w1(32'hbba89286),
	.w2(32'h3aa3ff20),
	.w3(32'hbb8b1a12),
	.w4(32'h3ac5f765),
	.w5(32'h3beb112e),
	.w6(32'hbbd6e805),
	.w7(32'h3b86335b),
	.w8(32'h3c137ed9),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55a431),
	.w1(32'hb94c77f1),
	.w2(32'hbc30596a),
	.w3(32'h3c461681),
	.w4(32'h3bb35c1e),
	.w5(32'hbb872589),
	.w6(32'h3c15ca0e),
	.w7(32'h3c8b83af),
	.w8(32'h3c178427),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e43e1),
	.w1(32'h399f976d),
	.w2(32'hbb14d310),
	.w3(32'hbbe4edff),
	.w4(32'hbbbac6d1),
	.w5(32'hbc58126b),
	.w6(32'h3b0a5762),
	.w7(32'hbb3a9d80),
	.w8(32'hbb5ae744),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63747b),
	.w1(32'hba3d58b7),
	.w2(32'hbba9fcb4),
	.w3(32'h3ba05c0a),
	.w4(32'h3bd0b204),
	.w5(32'hba6897fd),
	.w6(32'hbb1a0300),
	.w7(32'h3bdf53da),
	.w8(32'hbaa9fe7e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3e79c),
	.w1(32'h3b47e428),
	.w2(32'h3b57cda8),
	.w3(32'hbb301b1b),
	.w4(32'hbbb5ee95),
	.w5(32'hbb9c4794),
	.w6(32'hbb8cf071),
	.w7(32'hba11d31a),
	.w8(32'hbba2b912),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95af9f2),
	.w1(32'hba99962b),
	.w2(32'h3b157062),
	.w3(32'hbb581d6f),
	.w4(32'h3bace911),
	.w5(32'h3c3c8a41),
	.w6(32'hbbda6303),
	.w7(32'h3b5b07b6),
	.w8(32'h3bbf65d4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6908ae),
	.w1(32'h3bddd2af),
	.w2(32'h3b453ee0),
	.w3(32'h3bda9d14),
	.w4(32'hba49ab6c),
	.w5(32'hbbfea38e),
	.w6(32'h3bff7402),
	.w7(32'hba8a74e6),
	.w8(32'hbb734fee),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ed55b),
	.w1(32'hbc36d55c),
	.w2(32'hbb38c786),
	.w3(32'hbadd3178),
	.w4(32'hbbce4c52),
	.w5(32'hb9e95ddc),
	.w6(32'hbb4b7184),
	.w7(32'h3a089704),
	.w8(32'h3b81ba6a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ba708),
	.w1(32'h390bbc5a),
	.w2(32'h3c05e944),
	.w3(32'h3c214ded),
	.w4(32'hbb54dd6b),
	.w5(32'h3b90b01b),
	.w6(32'h3b4bc605),
	.w7(32'hbaab9dea),
	.w8(32'hbb3c4f46),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab1e86),
	.w1(32'hbc0cfe72),
	.w2(32'hbbea85bc),
	.w3(32'hbb1acbcf),
	.w4(32'hba5d5694),
	.w5(32'hbb3a1fa4),
	.w6(32'hbb035959),
	.w7(32'hbb8655ad),
	.w8(32'hbb7bbfa1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe76225),
	.w1(32'hb9851546),
	.w2(32'h3b3088a1),
	.w3(32'hbb9ce559),
	.w4(32'hbbbc6039),
	.w5(32'h3ba67fef),
	.w6(32'hbbb138a4),
	.w7(32'hbc26935a),
	.w8(32'hbbf8a3b7),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c1f09),
	.w1(32'hb9b8a52a),
	.w2(32'h3ba3ca1d),
	.w3(32'h3c0cc6b0),
	.w4(32'hbb9c23d7),
	.w5(32'h3b7beccf),
	.w6(32'hbb3e07e1),
	.w7(32'hbbbe4ad2),
	.w8(32'hbb9f38c3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cbab3),
	.w1(32'hbbf9aa5d),
	.w2(32'hb9c1b7da),
	.w3(32'hbb17a1f1),
	.w4(32'hbbe37f00),
	.w5(32'h3a918e9b),
	.w6(32'hbb37e246),
	.w7(32'hbc2fce6f),
	.w8(32'hbb4f4e3f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba65934),
	.w1(32'hbbe1bfd7),
	.w2(32'hbbc8f8cc),
	.w3(32'hbb648a9a),
	.w4(32'hbb97b512),
	.w5(32'hbba6e626),
	.w6(32'hbb9a7062),
	.w7(32'hb8950b79),
	.w8(32'hbb5b5466),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf32a7b),
	.w1(32'h3be86ff2),
	.w2(32'h3bc2746c),
	.w3(32'hbaeb1e34),
	.w4(32'h3b18b18f),
	.w5(32'hb8ce98fb),
	.w6(32'h3b73542d),
	.w7(32'hbae2b042),
	.w8(32'hbb8ad531),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb27807),
	.w1(32'h3a6a98b1),
	.w2(32'h3b7ab7c6),
	.w3(32'h3bf6560d),
	.w4(32'hbc151c61),
	.w5(32'h3b481a56),
	.w6(32'h3ba76f93),
	.w7(32'hbc12419b),
	.w8(32'hbba04d72),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6033da),
	.w1(32'h3b188b21),
	.w2(32'h3b8891a9),
	.w3(32'h3ac8e6c6),
	.w4(32'h3a1bc498),
	.w5(32'hbb20d430),
	.w6(32'hbbb4d60b),
	.w7(32'h3a52435e),
	.w8(32'h3afd8e03),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f12a7),
	.w1(32'h3b9e1cb8),
	.w2(32'h3abc5df2),
	.w3(32'h3adf8a05),
	.w4(32'h3bbc0c2e),
	.w5(32'hbc14071c),
	.w6(32'h3c076aa9),
	.w7(32'h3ca9048c),
	.w8(32'h3c9348ab),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c238bfa),
	.w1(32'h3bdea183),
	.w2(32'h3bd0b50d),
	.w3(32'h3c7d6dad),
	.w4(32'h3b5fb0d9),
	.w5(32'h3b864d98),
	.w6(32'h3c96c9a2),
	.w7(32'hbc422a79),
	.w8(32'hbc22d572),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02c78b),
	.w1(32'hbbec27b9),
	.w2(32'h3bbe79a2),
	.w3(32'hbacd97f9),
	.w4(32'hbc0dca00),
	.w5(32'h3bea666d),
	.w6(32'hbbe49df5),
	.w7(32'hba2461d3),
	.w8(32'h3c00ce0a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba333ac),
	.w1(32'hbb609dfd),
	.w2(32'hba35f836),
	.w3(32'h3c64f9ae),
	.w4(32'hbb921c16),
	.w5(32'h3aada2e7),
	.w6(32'h3b9f0fe1),
	.w7(32'hbb87bca9),
	.w8(32'h3ba1de85),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2a15e),
	.w1(32'h3a838244),
	.w2(32'hbbbf6696),
	.w3(32'h3b5137e9),
	.w4(32'h3ae5ff68),
	.w5(32'hbbf84052),
	.w6(32'h3bdbdb72),
	.w7(32'h3bea2ebc),
	.w8(32'h3a3496e7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d516f),
	.w1(32'hbb99bb89),
	.w2(32'hbc241b31),
	.w3(32'hbb2cba1f),
	.w4(32'h3a8961dc),
	.w5(32'hbc739052),
	.w6(32'h3b3f9e60),
	.w7(32'hbbecd7ba),
	.w8(32'hbbe0981c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e7a7e),
	.w1(32'h3b6d4545),
	.w2(32'h3c5b3ee0),
	.w3(32'hbc558f89),
	.w4(32'hbbaba4b7),
	.w5(32'h3bd0fd68),
	.w6(32'hbc31fdae),
	.w7(32'h3bed71c4),
	.w8(32'h3ba8b486),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c34e1),
	.w1(32'h39f53232),
	.w2(32'h3ab0cbbe),
	.w3(32'h3c64fd67),
	.w4(32'h39f0c91c),
	.w5(32'h3b1e4467),
	.w6(32'h3b8ea5c9),
	.w7(32'h3b004f41),
	.w8(32'h3bcb6240),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92503b),
	.w1(32'h3c2a3b18),
	.w2(32'h3c9d2127),
	.w3(32'hbafacb62),
	.w4(32'hbbd2e857),
	.w5(32'hbb82321f),
	.w6(32'h3ab5c994),
	.w7(32'hbbef4cda),
	.w8(32'hbc5b2c09),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17a68d),
	.w1(32'h3bab7b37),
	.w2(32'hbad5a76c),
	.w3(32'hbb8bb54f),
	.w4(32'h3bee80c1),
	.w5(32'hbb6230e9),
	.w6(32'hbc15c933),
	.w7(32'h3b83466a),
	.w8(32'hbb227f67),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2ab54),
	.w1(32'hbadd91e7),
	.w2(32'h3bbdaec8),
	.w3(32'hbc1b58a6),
	.w4(32'hbb5f9c83),
	.w5(32'h3bae283a),
	.w6(32'hbba1f719),
	.w7(32'hba1e90d3),
	.w8(32'hbb371052),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be91cc4),
	.w1(32'hb92ab583),
	.w2(32'hbbd365b1),
	.w3(32'h3c64522d),
	.w4(32'h3b081aa9),
	.w5(32'hbb60665c),
	.w6(32'h3a7415d7),
	.w7(32'hbb6932f9),
	.w8(32'hbba596a5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaea8cb),
	.w1(32'h3a198b93),
	.w2(32'hbb66830a),
	.w3(32'hbb80b77c),
	.w4(32'hba896c72),
	.w5(32'h39db0820),
	.w6(32'hbbac1987),
	.w7(32'hbb775ee8),
	.w8(32'hbb909d3d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989871),
	.w1(32'hb8da87c1),
	.w2(32'hba8fd8aa),
	.w3(32'hbb6355fc),
	.w4(32'h39f197d2),
	.w5(32'hbb871ba9),
	.w6(32'h3b37ed1a),
	.w7(32'hba5f3cac),
	.w8(32'h3b143836),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b16c9),
	.w1(32'h3b6bd338),
	.w2(32'h3b8f77e7),
	.w3(32'hbb030f4f),
	.w4(32'h3a619938),
	.w5(32'h3be853cc),
	.w6(32'h3b48d82d),
	.w7(32'h3adc3432),
	.w8(32'hbb05ae49),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0f179),
	.w1(32'hba05c5d1),
	.w2(32'h3ab3c146),
	.w3(32'h3b0bc605),
	.w4(32'h3b4a6532),
	.w5(32'hba6c303b),
	.w6(32'hbbaac8b2),
	.w7(32'h3b95f3a4),
	.w8(32'h3b0c1ee5),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2b1d6),
	.w1(32'h3b8005cf),
	.w2(32'hbaa3e344),
	.w3(32'h3aa3b9dd),
	.w4(32'h3ba6b754),
	.w5(32'h3b78f883),
	.w6(32'h3bf9f915),
	.w7(32'h3bac3a93),
	.w8(32'h3b08fd64),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac36d2),
	.w1(32'hbabf177a),
	.w2(32'h3a88cbe3),
	.w3(32'hbc0c0533),
	.w4(32'hbb592352),
	.w5(32'h3ba60960),
	.w6(32'hbb347f81),
	.w7(32'hbbbe8f18),
	.w8(32'hbad3400b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eb5d7),
	.w1(32'h3bcf962c),
	.w2(32'hbb8a2d9e),
	.w3(32'h3b26508a),
	.w4(32'hba1652f8),
	.w5(32'hbc924668),
	.w6(32'hbb31fb43),
	.w7(32'h3bb1c5cf),
	.w8(32'hbb1dc07a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a4b17),
	.w1(32'hbb1caab6),
	.w2(32'h3a832389),
	.w3(32'hbb953772),
	.w4(32'hbaeb65fa),
	.w5(32'h3b21c95c),
	.w6(32'h3b4e69ad),
	.w7(32'hbae30835),
	.w8(32'h3aa768a0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b826e3e),
	.w1(32'hbbedb125),
	.w2(32'hbbf63f53),
	.w3(32'h3bc3c660),
	.w4(32'hbc2b4e72),
	.w5(32'hbbc78827),
	.w6(32'h3ad6791b),
	.w7(32'hbbed4fce),
	.w8(32'hba82c80b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdfddc),
	.w1(32'hbb922762),
	.w2(32'hba33063e),
	.w3(32'h3b840e0d),
	.w4(32'h3a1fabd0),
	.w5(32'h3ae17421),
	.w6(32'h3c047629),
	.w7(32'hbbad9f22),
	.w8(32'hbbe78798),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb85723),
	.w1(32'hbb79c800),
	.w2(32'hba4b2cb8),
	.w3(32'hbbe4f141),
	.w4(32'hb9d75441),
	.w5(32'h3b8a856a),
	.w6(32'hbc1185dd),
	.w7(32'h3b9c670b),
	.w8(32'h3b0bef32),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37416a),
	.w1(32'h3b9c5e3f),
	.w2(32'h3bed11ae),
	.w3(32'h3c31bbc2),
	.w4(32'h3a86f635),
	.w5(32'h3bd5e1c0),
	.w6(32'h3bc7e908),
	.w7(32'h39cae6c0),
	.w8(32'h3b878be0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe0225),
	.w1(32'hb7e200c6),
	.w2(32'h36ff7295),
	.w3(32'h3a08a769),
	.w4(32'h3765fdcc),
	.w5(32'h386d6bdf),
	.w6(32'hbc101a12),
	.w7(32'h38144d8e),
	.w8(32'h38931992),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7719e55),
	.w1(32'hb7204347),
	.w2(32'hb7e3f206),
	.w3(32'hb73d955f),
	.w4(32'h371ab1a5),
	.w5(32'hb6cf8256),
	.w6(32'hb5996d08),
	.w7(32'h367b08e4),
	.w8(32'hb78137d2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb51051bf),
	.w1(32'hb592879e),
	.w2(32'hb5664820),
	.w3(32'h33a54ea6),
	.w4(32'hb544f56e),
	.w5(32'hb4b66631),
	.w6(32'h35067f52),
	.w7(32'hb4a756fd),
	.w8(32'hb554d82f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3811d335),
	.w1(32'h3830801c),
	.w2(32'h375c5d74),
	.w3(32'h381adf38),
	.w4(32'h380c617b),
	.w5(32'h36b30169),
	.w6(32'h378ef7e2),
	.w7(32'h37b10c07),
	.w8(32'hb724df74),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb54e5199),
	.w1(32'h34af6ea4),
	.w2(32'hb574f315),
	.w3(32'hb5045f8d),
	.w4(32'h33d0702a),
	.w5(32'hb5a366d1),
	.w6(32'hb40c3994),
	.w7(32'hb5136a56),
	.w8(32'hb61c31e0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f7bbd3),
	.w1(32'h37419d9c),
	.w2(32'hb7a46b58),
	.w3(32'h378351f1),
	.w4(32'h38045401),
	.w5(32'hb73224fc),
	.w6(32'h3693e0c2),
	.w7(32'hb67ab5ce),
	.w8(32'hb813c1a8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a43417),
	.w1(32'hb7a75e8d),
	.w2(32'hb8028ea7),
	.w3(32'hb7aa3c87),
	.w4(32'hb81f711a),
	.w5(32'hb8328db1),
	.w6(32'hb78338c3),
	.w7(32'hb76d1c80),
	.w8(32'hb7a1e431),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80b5e92),
	.w1(32'hb8013467),
	.w2(32'hb7d2626f),
	.w3(32'hb76dbefa),
	.w4(32'hb6b305c7),
	.w5(32'hb663cf8a),
	.w6(32'h361d2ad7),
	.w7(32'h3786ec6a),
	.w8(32'h3756e304),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb687b3bb),
	.w1(32'hb697ad43),
	.w2(32'hb6917a44),
	.w3(32'hb6c1440b),
	.w4(32'hb6b93390),
	.w5(32'hb6f69b6c),
	.w6(32'hb746344f),
	.w7(32'hb7207b65),
	.w8(32'hb733a1c6),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb823d072),
	.w1(32'hb8377bc0),
	.w2(32'hb86d83d6),
	.w3(32'hb7c3bea8),
	.w4(32'hb788e77f),
	.w5(32'hb7db830c),
	.w6(32'hb5bf800d),
	.w7(32'h3788fea3),
	.w8(32'hb6ba2b3e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d002f2),
	.w1(32'h3707bbf3),
	.w2(32'h3774649b),
	.w3(32'h383dc365),
	.w4(32'h37f72603),
	.w5(32'h37f0b0b4),
	.w6(32'h3820ff0e),
	.w7(32'h38177c4a),
	.w8(32'h38280a03),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb96be),
	.w1(32'hb8cdc300),
	.w2(32'hb8c7c46b),
	.w3(32'hb7d304e7),
	.w4(32'hb755acc9),
	.w5(32'hb80b4a9a),
	.w6(32'hb4a86f9a),
	.w7(32'h3772fbf2),
	.w8(32'h3731f6c9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb51b8181),
	.w1(32'h3500e5d8),
	.w2(32'h3514d647),
	.w3(32'hb5852763),
	.w4(32'hb526fb85),
	.w5(32'h34097959),
	.w6(32'hb5cb2e13),
	.w7(32'hb4fc67fc),
	.w8(32'h33171b3b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb49abc67),
	.w1(32'hb5bf287b),
	.w2(32'hb631540d),
	.w3(32'hb4b0bc2e),
	.w4(32'h35700990),
	.w5(32'hb4825cbe),
	.w6(32'h34ff42be),
	.w7(32'hb5538d23),
	.w8(32'hb5c1b384),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb862246d),
	.w1(32'hb7595f83),
	.w2(32'h37cdc439),
	.w3(32'hb88128f2),
	.w4(32'h36308a21),
	.w5(32'h384f3a46),
	.w6(32'hb75aafec),
	.w7(32'h376ed6b8),
	.w8(32'h37d97589),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6db3b25),
	.w1(32'h37a0ef1d),
	.w2(32'h380f36df),
	.w3(32'h38145fb5),
	.w4(32'h38354ed8),
	.w5(32'h389fc6e1),
	.w6(32'h38710722),
	.w7(32'h38683e89),
	.w8(32'h383ea409),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82943f2),
	.w1(32'hb82d10e0),
	.w2(32'hb86059fd),
	.w3(32'hb70f09f0),
	.w4(32'hb73637ca),
	.w5(32'hb7b97719),
	.w6(32'h37de4dec),
	.w7(32'h37f204fd),
	.w8(32'h37502d60),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375af00e),
	.w1(32'hb71fb977),
	.w2(32'h37049b1b),
	.w3(32'h3793ce74),
	.w4(32'h386a887c),
	.w5(32'h3737ec87),
	.w6(32'h374c93b2),
	.w7(32'h381dcc72),
	.w8(32'h38817384),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361fc70d),
	.w1(32'h370dc4fe),
	.w2(32'h36c2e84f),
	.w3(32'h3690cda8),
	.w4(32'h36f1ebca),
	.w5(32'h3621a948),
	.w6(32'h35b50ab3),
	.w7(32'h36b5520b),
	.w8(32'h369032b7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372e42d1),
	.w1(32'h37a81a04),
	.w2(32'h37990f4c),
	.w3(32'h36cb5dd5),
	.w4(32'h37a1bc42),
	.w5(32'h37667ec8),
	.w6(32'h3702fe5b),
	.w7(32'h373f7901),
	.w8(32'h35eaa0e3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71ed85b),
	.w1(32'h37e8017d),
	.w2(32'h386efb3d),
	.w3(32'hb8186d9f),
	.w4(32'h38768454),
	.w5(32'h3881d7a7),
	.w6(32'hb72f148c),
	.w7(32'hb64d72af),
	.w8(32'h38215643),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb823b2b7),
	.w1(32'hb815d547),
	.w2(32'hb63957ef),
	.w3(32'h37b898b4),
	.w4(32'h37a63cc8),
	.w5(32'h38777385),
	.w6(32'h38060aa6),
	.w7(32'h3825c3bc),
	.w8(32'h389bcdde),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372f5d2b),
	.w1(32'h3824c14e),
	.w2(32'h384e7aa3),
	.w3(32'h35c82415),
	.w4(32'h385ebc93),
	.w5(32'h388fa899),
	.w6(32'h37877005),
	.w7(32'h37bdece3),
	.w8(32'h385fcefe),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5501792),
	.w1(32'hb78fc05d),
	.w2(32'hb7bb066b),
	.w3(32'h3720cc1c),
	.w4(32'hb7757bd0),
	.w5(32'hb75978c5),
	.w6(32'h35bf7424),
	.w7(32'h3691c78a),
	.w8(32'hb74b738e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a89f4d),
	.w1(32'hb81002c2),
	.w2(32'hb8288bc1),
	.w3(32'hb29b2048),
	.w4(32'hb7a01fd9),
	.w5(32'hb8208c32),
	.w6(32'h3787f19f),
	.w7(32'h36cb9658),
	.w8(32'hb7a50dbd),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb533bcb7),
	.w1(32'hb4d710e4),
	.w2(32'hb5869a73),
	.w3(32'hb4f79e01),
	.w4(32'hb4a4c71a),
	.w5(32'hb5a2fbce),
	.w6(32'hb52c9fc2),
	.w7(32'hb5373c55),
	.w8(32'hb5a9c086),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c5bb20),
	.w1(32'hb50ce99c),
	.w2(32'h34a302f6),
	.w3(32'hb4a3a37d),
	.w4(32'hb588fdfc),
	.w5(32'hb46c02e1),
	.w6(32'hb56532e0),
	.w7(32'hb549faf2),
	.w8(32'hb4b0fd44),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75c5319),
	.w1(32'hb75bdcea),
	.w2(32'hb7225788),
	.w3(32'hb6f75a1e),
	.w4(32'h35ca73ac),
	.w5(32'h36bc0a85),
	.w6(32'hb6a0c5ea),
	.w7(32'h363c2e13),
	.w8(32'h373f2f2e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3479ca0),
	.w1(32'hb427caef),
	.w2(32'hb5143271),
	.w3(32'hb4868a24),
	.w4(32'hb5364a18),
	.w5(32'hb4e83dd1),
	.w6(32'h344868d6),
	.w7(32'hb4dabc32),
	.w8(32'hb586bf52),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bc5243),
	.w1(32'h37b65253),
	.w2(32'h37f9e58c),
	.w3(32'hb7063277),
	.w4(32'h37af086f),
	.w5(32'h37f48f57),
	.w6(32'hb70281a0),
	.w7(32'h370541dc),
	.w8(32'h379dc53c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3635e192),
	.w1(32'h372daa22),
	.w2(32'h379d8113),
	.w3(32'h37c8aaab),
	.w4(32'h37f9991d),
	.w5(32'h381d2698),
	.w6(32'h383c3cf5),
	.w7(32'h383f940d),
	.w8(32'h37f56115),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76de71b),
	.w1(32'hb652c0c1),
	.w2(32'hb6900e9e),
	.w3(32'hb627b80d),
	.w4(32'h373f5334),
	.w5(32'h37833bb3),
	.w6(32'h36626b82),
	.w7(32'h37bf47f6),
	.w8(32'h37b94547),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4f3140a),
	.w1(32'hb4d0ca49),
	.w2(32'hb51cbd9f),
	.w3(32'hb398e063),
	.w4(32'hb606a4e7),
	.w5(32'hb63fb157),
	.w6(32'h34299f29),
	.w7(32'hb5e44ed1),
	.w8(32'hb6004c26),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378639a0),
	.w1(32'h381e88ac),
	.w2(32'h38839375),
	.w3(32'h3483c627),
	.w4(32'h38732431),
	.w5(32'h3890d5f4),
	.w6(32'h37a64358),
	.w7(32'h379169df),
	.w8(32'h3895e625),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36df1c74),
	.w1(32'h369bac2c),
	.w2(32'h373f6514),
	.w3(32'h37600721),
	.w4(32'h37a6be8d),
	.w5(32'h37912985),
	.w6(32'h3730455f),
	.w7(32'h3788d290),
	.w8(32'h37ce3486),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34233dad),
	.w1(32'hb33c18ff),
	.w2(32'hb56fb905),
	.w3(32'hb3239c70),
	.w4(32'hb5c88004),
	.w5(32'hb67ed73c),
	.w6(32'hb5f83de3),
	.w7(32'hb5884609),
	.w8(32'hb6642508),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37017cad),
	.w1(32'h37a4c99c),
	.w2(32'h3832d484),
	.w3(32'h37af5013),
	.w4(32'h37d70244),
	.w5(32'h3815a0e4),
	.w6(32'h3798fc29),
	.w7(32'h3775bad9),
	.w8(32'h381376a4),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69471fa),
	.w1(32'hb6b35841),
	.w2(32'hb6607d72),
	.w3(32'hb6ca095a),
	.w4(32'hb6d71eb0),
	.w5(32'hb68b515a),
	.w6(32'hb65477a7),
	.w7(32'hb6430c92),
	.w8(32'hb5251945),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h363bb590),
	.w1(32'h368c4c89),
	.w2(32'hb3b71f17),
	.w3(32'h36692eb8),
	.w4(32'h363b0203),
	.w5(32'h35c1e199),
	.w6(32'h360eb197),
	.w7(32'h355f738c),
	.w8(32'h35a4174d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h343a05a0),
	.w1(32'hb555b407),
	.w2(32'hb5025591),
	.w3(32'h330e8d43),
	.w4(32'hb57f8e00),
	.w5(32'hb44566ec),
	.w6(32'hb3b9e392),
	.w7(32'hb47a9ebc),
	.w8(32'h350286c2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb51e9a03),
	.w1(32'hb584b1ba),
	.w2(32'hb562036f),
	.w3(32'hb4f92e9a),
	.w4(32'hb58e54d5),
	.w5(32'hb41d5237),
	.w6(32'hb4854819),
	.w7(32'h33394e98),
	.w8(32'h34b294a2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cefe47),
	.w1(32'hb7be8ee3),
	.w2(32'hb7bdadde),
	.w3(32'hb7795c74),
	.w4(32'hb78f4ea2),
	.w5(32'hb792a973),
	.w6(32'hb7a7eb74),
	.w7(32'hb7320fd3),
	.w8(32'hb7589145),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367da689),
	.w1(32'hb743f9cf),
	.w2(32'h38052cbe),
	.w3(32'h386a0d80),
	.w4(32'h38300758),
	.w5(32'h37fc4820),
	.w6(32'h3825d982),
	.w7(32'h3850d79d),
	.w8(32'h38904f7f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d6cf6b),
	.w1(32'h37bd2867),
	.w2(32'h3839fa10),
	.w3(32'h382c38df),
	.w4(32'h382f561d),
	.w5(32'h384f0902),
	.w6(32'h37fbf8ab),
	.w7(32'h37f56182),
	.w8(32'h3841e3b1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7633b46),
	.w1(32'hb7734968),
	.w2(32'h38152558),
	.w3(32'h381ab27c),
	.w4(32'h3804767c),
	.w5(32'h3807329a),
	.w6(32'h3802b521),
	.w7(32'h383b43d5),
	.w8(32'h3895ed14),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35edb716),
	.w1(32'h35143ff0),
	.w2(32'h35260c96),
	.w3(32'h35d001d5),
	.w4(32'h35a98e66),
	.w5(32'h33de5cc5),
	.w6(32'h3532d316),
	.w7(32'h3543d8cd),
	.w8(32'h34a0b78d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36704531),
	.w1(32'h36af045e),
	.w2(32'h36ba0964),
	.w3(32'h3626201f),
	.w4(32'h3691cb8f),
	.w5(32'h364d2ef1),
	.w6(32'h35929821),
	.w7(32'h36925edc),
	.w8(32'h35f164ff),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h355e7da2),
	.w1(32'h351c6a80),
	.w2(32'h33d2f816),
	.w3(32'h34fb9531),
	.w4(32'h350a6c52),
	.w5(32'h355b3c6b),
	.w6(32'h35dc546d),
	.w7(32'h35884a82),
	.w8(32'h354158ac),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3512a11d),
	.w1(32'h3338d312),
	.w2(32'hb526196c),
	.w3(32'h33cdecea),
	.w4(32'hb42ec7ee),
	.w5(32'h345d0345),
	.w6(32'hb4a865ea),
	.w7(32'hb4ed4121),
	.w8(32'hb503bb1a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812234e),
	.w1(32'h37d8fe7d),
	.w2(32'h37f3641c),
	.w3(32'h37ff9b48),
	.w4(32'h380b6b1a),
	.w5(32'h37c6d776),
	.w6(32'h37e1ec34),
	.w7(32'h381fd2f5),
	.w8(32'h37f147be),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37636cc1),
	.w1(32'h37126def),
	.w2(32'h370e1777),
	.w3(32'h37157581),
	.w4(32'h36a55384),
	.w5(32'h36f46ee0),
	.w6(32'h36ff35e6),
	.w7(32'h369ccf2d),
	.w8(32'h36f5c8e3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d9248c),
	.w1(32'hb7218499),
	.w2(32'hb6d98bc5),
	.w3(32'hb755032f),
	.w4(32'hb7387894),
	.w5(32'hb7303adf),
	.w6(32'hb7b3b008),
	.w7(32'hb789befa),
	.w8(32'hb74b3ea6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3754eb2c),
	.w1(32'h37a7f7b7),
	.w2(32'h35d31600),
	.w3(32'h3795a022),
	.w4(32'h377d559c),
	.w5(32'h358e3fa2),
	.w6(32'h36d696a6),
	.w7(32'h3707817b),
	.w8(32'hb7436ec0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34121290),
	.w1(32'hb5039c8c),
	.w2(32'h36046c30),
	.w3(32'hb621dabf),
	.w4(32'hb609ce23),
	.w5(32'h35d3735a),
	.w6(32'hb5fe56d0),
	.w7(32'hb5b0e94c),
	.w8(32'h35aff0b0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a28f1e),
	.w1(32'hb76bf70f),
	.w2(32'hb703e135),
	.w3(32'hb6e2de9e),
	.w4(32'hb53c8562),
	.w5(32'h361c9d00),
	.w6(32'hb69d8eb3),
	.w7(32'h35fc7a69),
	.w8(32'h373d87db),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c8dd5b),
	.w1(32'h36c38053),
	.w2(32'h3656c8e3),
	.w3(32'h36886a08),
	.w4(32'h36ce4bee),
	.w5(32'h365f9c92),
	.w6(32'h3613a7e0),
	.w7(32'h36b4e8dc),
	.w8(32'h365e0647),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38926b37),
	.w1(32'h3846f01f),
	.w2(32'h388a52f2),
	.w3(32'h38d5b6f3),
	.w4(32'h388a5b3a),
	.w5(32'h37ff82d6),
	.w6(32'h38863a59),
	.w7(32'h38941646),
	.w8(32'h383e1af2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6069e38),
	.w1(32'hb60310a1),
	.w2(32'h35afaa5b),
	.w3(32'hb5dd0c87),
	.w4(32'hb5caa486),
	.w5(32'h361c611c),
	.w6(32'hb5a8e52a),
	.w7(32'h3570d925),
	.w8(32'h366ffb7c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375c1187),
	.w1(32'h3777e80b),
	.w2(32'h381bef33),
	.w3(32'h37cfd253),
	.w4(32'h37c8c0af),
	.w5(32'h37a16a93),
	.w6(32'h37225851),
	.w7(32'hb70b3b8d),
	.w8(32'hb81af36f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule