module layer_10_featuremap_253(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c863d),
	.w1(32'hbb11a36e),
	.w2(32'hbb370131),
	.w3(32'hbb4918ee),
	.w4(32'hbaf0b317),
	.w5(32'h3a4c8bfa),
	.w6(32'hbb1640fd),
	.w7(32'hbaa92a49),
	.w8(32'hb9d4ae86),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a955a7c),
	.w1(32'h3a6bc3bf),
	.w2(32'hb99b4936),
	.w3(32'hba271513),
	.w4(32'hba406f17),
	.w5(32'hba6a7382),
	.w6(32'hba2a11a3),
	.w7(32'h39a23090),
	.w8(32'hba391188),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27a752),
	.w1(32'h3a3ef1d6),
	.w2(32'h3b26d36c),
	.w3(32'h38f23819),
	.w4(32'h3a924111),
	.w5(32'hbaa6746d),
	.w6(32'h3b655580),
	.w7(32'h3b806c71),
	.w8(32'hba806cd5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c00087),
	.w1(32'hbaa9b846),
	.w2(32'hba825154),
	.w3(32'hba914699),
	.w4(32'h394b35bd),
	.w5(32'hba45c7c4),
	.w6(32'h3730b866),
	.w7(32'hb7d81ad1),
	.w8(32'hbb02d6ee),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4604c9),
	.w1(32'hbba2c854),
	.w2(32'hbb5a74df),
	.w3(32'hbaa0f9f6),
	.w4(32'h3aafc975),
	.w5(32'h39cf5a3a),
	.w6(32'hba963312),
	.w7(32'hbb283584),
	.w8(32'h3a570d22),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5df0f0),
	.w1(32'hb8920d20),
	.w2(32'h36ec25a8),
	.w3(32'h3a3cf64e),
	.w4(32'h3a8428df),
	.w5(32'hba19ab4d),
	.w6(32'h3a445860),
	.w7(32'h3ac4fddc),
	.w8(32'h36790cf8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de93b7),
	.w1(32'hb9c4219d),
	.w2(32'hb9904b02),
	.w3(32'h3a1c4d32),
	.w4(32'h39a6964d),
	.w5(32'hbad3a769),
	.w6(32'h39641fe3),
	.w7(32'h36d41d6e),
	.w8(32'hbb062e70),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c84c0),
	.w1(32'hbb77286a),
	.w2(32'hbb4f9b5c),
	.w3(32'hbabf7673),
	.w4(32'hbac05ff9),
	.w5(32'hba99c58a),
	.w6(32'hbb0d8ce6),
	.w7(32'hbb46506b),
	.w8(32'hba4db644),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf5296),
	.w1(32'hbab5e871),
	.w2(32'hba97ba45),
	.w3(32'hbaf58894),
	.w4(32'hbac90fa7),
	.w5(32'h3a8b9bee),
	.w6(32'hba77b820),
	.w7(32'hba3e763c),
	.w8(32'h3a89b502),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b004ac4),
	.w1(32'h39cd3916),
	.w2(32'h3a34984a),
	.w3(32'h3aebf005),
	.w4(32'h3a89d12a),
	.w5(32'hba38e762),
	.w6(32'h3aba78fb),
	.w7(32'h3ac4ff18),
	.w8(32'hba86d7e2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aaa773),
	.w1(32'hb9214870),
	.w2(32'hb99dd1fd),
	.w3(32'h3986519a),
	.w4(32'h3a97c186),
	.w5(32'hb8aa62d5),
	.w6(32'h398466e6),
	.w7(32'h3a85fe20),
	.w8(32'h39cc4509),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bfbef),
	.w1(32'h3a283d9a),
	.w2(32'hb7024fb4),
	.w3(32'hb9035a1b),
	.w4(32'hbace8932),
	.w5(32'h3a93a0c4),
	.w6(32'hba40ac16),
	.w7(32'h3a753497),
	.w8(32'h3b0302e3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eb9c7),
	.w1(32'h3b4b3fa3),
	.w2(32'h3adaa456),
	.w3(32'h3ac57bab),
	.w4(32'h3a8ffe50),
	.w5(32'h3b08dd56),
	.w6(32'h3b4fc7e7),
	.w7(32'h3a3b5758),
	.w8(32'hb9489b8c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f43de1),
	.w1(32'hbadbb720),
	.w2(32'hba61b639),
	.w3(32'h3a7fb9ae),
	.w4(32'h3a994307),
	.w5(32'h3947efcb),
	.w6(32'hba033173),
	.w7(32'h399592d4),
	.w8(32'h3a0a81b0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a856b8d),
	.w1(32'h399204c0),
	.w2(32'h3a34a114),
	.w3(32'h3a8c2299),
	.w4(32'h3a4212ec),
	.w5(32'h3adcbdbc),
	.w6(32'h3a556577),
	.w7(32'h3a1e793f),
	.w8(32'h3a2fa958),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac076d5),
	.w1(32'hbb01c4f9),
	.w2(32'hba835bdc),
	.w3(32'hb9bfb719),
	.w4(32'h3ab168bc),
	.w5(32'h3908b1a5),
	.w6(32'hb9959f59),
	.w7(32'hbb0404e7),
	.w8(32'h386838cc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd1dac),
	.w1(32'hba9e247b),
	.w2(32'hbb0c5735),
	.w3(32'h392e4dc3),
	.w4(32'h393b3324),
	.w5(32'h3a00c5aa),
	.w6(32'hbab0d3fb),
	.w7(32'hba9897ef),
	.w8(32'h3a9e8026),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e8282),
	.w1(32'h3aca199f),
	.w2(32'h3b080ca5),
	.w3(32'h3a2ebcfd),
	.w4(32'h3a88c384),
	.w5(32'hba32af9c),
	.w6(32'h3abc3817),
	.w7(32'h3a7aaa8f),
	.w8(32'hba7f4427),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c38677),
	.w1(32'hb9432326),
	.w2(32'h3a83399b),
	.w3(32'hb93c1387),
	.w4(32'hb98b8308),
	.w5(32'h38f51997),
	.w6(32'hbb03cbd3),
	.w7(32'hba8fadb7),
	.w8(32'h393b8292),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff9b66),
	.w1(32'h3b152d3f),
	.w2(32'hba1d9984),
	.w3(32'h3a92cfb0),
	.w4(32'h3b18d64e),
	.w5(32'h3b55b43f),
	.w6(32'h3a0807c1),
	.w7(32'h39d33bd2),
	.w8(32'h3a614be4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b089db9),
	.w1(32'hba3fecb3),
	.w2(32'hbaea4748),
	.w3(32'h38eec341),
	.w4(32'h3a344026),
	.w5(32'hb81c45d9),
	.w6(32'h39f9d20a),
	.w7(32'hbae8786e),
	.w8(32'hba0260c7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7715a9),
	.w1(32'hba613d64),
	.w2(32'hba689abd),
	.w3(32'h388b25c8),
	.w4(32'hba54a685),
	.w5(32'hb911702f),
	.w6(32'hba3c8855),
	.w7(32'hba4312b5),
	.w8(32'h39d988fd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a58da),
	.w1(32'h3b5aa12f),
	.w2(32'h3ae28a13),
	.w3(32'h3b25bf94),
	.w4(32'h3a3a0724),
	.w5(32'h3b23ec7c),
	.w6(32'h3b0949eb),
	.w7(32'h3a9b0afd),
	.w8(32'h3b31c57d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ac6fa),
	.w1(32'hba84add6),
	.w2(32'hba534f4c),
	.w3(32'h39b87057),
	.w4(32'h3b048cd5),
	.w5(32'hbaf51a63),
	.w6(32'hb91174ee),
	.w7(32'hb7c5e6b9),
	.w8(32'hbae2894b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0af7a),
	.w1(32'hbab24a3d),
	.w2(32'h3aaec1ad),
	.w3(32'hba335fb4),
	.w4(32'h3a3cf7b4),
	.w5(32'hba071ada),
	.w6(32'h3b2ff3e4),
	.w7(32'hb98606a4),
	.w8(32'h3adc50c8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03161a),
	.w1(32'hb810df94),
	.w2(32'h38840082),
	.w3(32'h3aeebdca),
	.w4(32'h3b1b49a3),
	.w5(32'hb930d0ea),
	.w6(32'h3a3710e0),
	.w7(32'h3ab81823),
	.w8(32'h37cc3de8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70edef),
	.w1(32'hb8f99ea6),
	.w2(32'h3a6eb80d),
	.w3(32'hb768f8bf),
	.w4(32'h39080de0),
	.w5(32'hb8c44c66),
	.w6(32'h38a9f9fb),
	.w7(32'h393c9bf1),
	.w8(32'h39709542),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2343ea),
	.w1(32'hbae0b614),
	.w2(32'hba906167),
	.w3(32'hbadaec0a),
	.w4(32'hbaea0574),
	.w5(32'h3aef4e80),
	.w6(32'hba114d79),
	.w7(32'hba998ec1),
	.w8(32'hba0f869c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46697c),
	.w1(32'hbabbaa57),
	.w2(32'h3a87809a),
	.w3(32'hb8761cc0),
	.w4(32'h3a8b0216),
	.w5(32'hbb09f543),
	.w6(32'h3b34e1a3),
	.w7(32'h3aa6e802),
	.w8(32'hbb0ae88c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5bf85d6),
	.w1(32'h3b03ba99),
	.w2(32'h3af55185),
	.w3(32'hba225979),
	.w4(32'h39effda0),
	.w5(32'hbaea6553),
	.w6(32'hb9a2a879),
	.w7(32'h39c75f54),
	.w8(32'hbb0f8b64),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb475843),
	.w1(32'hbb4f43c7),
	.w2(32'hba3b8eec),
	.w3(32'hba635a72),
	.w4(32'hbb36b434),
	.w5(32'hb8da03de),
	.w6(32'h3a203ce0),
	.w7(32'hba98040f),
	.w8(32'h3a133144),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a97c0),
	.w1(32'h39f0ff9f),
	.w2(32'h3a069bee),
	.w3(32'h3b58ce91),
	.w4(32'hb9cbfc0d),
	.w5(32'hbaf82782),
	.w6(32'h3b054454),
	.w7(32'h3b29593a),
	.w8(32'hbaaa45d3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e3735),
	.w1(32'hb6d2ef94),
	.w2(32'h3b0c194f),
	.w3(32'hbaea484a),
	.w4(32'h39eef229),
	.w5(32'h3ada987d),
	.w6(32'hba397f29),
	.w7(32'h3aa52b84),
	.w8(32'h3a202014),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9eb65),
	.w1(32'h3b04d345),
	.w2(32'h389cbcd5),
	.w3(32'h392b6930),
	.w4(32'h3aa3238a),
	.w5(32'hb94977f4),
	.w6(32'h3b64b91b),
	.w7(32'h39a4002d),
	.w8(32'h3a170625),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782f1e1),
	.w1(32'hba21cd0e),
	.w2(32'hba94b27c),
	.w3(32'hba282834),
	.w4(32'h3ac4dc3b),
	.w5(32'hbaaeb7be),
	.w6(32'h3ab3b674),
	.w7(32'hba7d1317),
	.w8(32'hba299577),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93e146),
	.w1(32'h3a297260),
	.w2(32'h3a903daf),
	.w3(32'hba02ceec),
	.w4(32'h3b29c762),
	.w5(32'hbb01a8d2),
	.w6(32'hb9ee739a),
	.w7(32'h39e4583e),
	.w8(32'hb9dc5f75),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b383517),
	.w1(32'h3b449e0b),
	.w2(32'h3ac6628b),
	.w3(32'hba2d8351),
	.w4(32'h3b64748e),
	.w5(32'h3a8a076a),
	.w6(32'h3b70506c),
	.w7(32'h3a42197f),
	.w8(32'h3aa7820d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af341c),
	.w1(32'hba74c2cb),
	.w2(32'hba352efb),
	.w3(32'hb8a5fa9c),
	.w4(32'h3afecfef),
	.w5(32'hb8d06a97),
	.w6(32'h3a426b61),
	.w7(32'h3ac1651d),
	.w8(32'h398825fe),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1567ab),
	.w1(32'h3a65eaa3),
	.w2(32'hbaa94bed),
	.w3(32'h3a1c20f6),
	.w4(32'h3a15eec5),
	.w5(32'hba3f0b01),
	.w6(32'h3a8c4609),
	.w7(32'hba38deb6),
	.w8(32'hb8e07a84),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e2099),
	.w1(32'hbb48b549),
	.w2(32'hbb872291),
	.w3(32'hba8adeb7),
	.w4(32'hba07a195),
	.w5(32'h39e8ed0f),
	.w6(32'hbab1b504),
	.w7(32'hba528f18),
	.w8(32'hba716522),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f5157),
	.w1(32'hb90b2292),
	.w2(32'h39502676),
	.w3(32'h3a2adf66),
	.w4(32'h3a44cb15),
	.w5(32'h3a51f1d2),
	.w6(32'h3ab518b5),
	.w7(32'hb98a3106),
	.w8(32'h3ae90f38),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cee23),
	.w1(32'hba538d7f),
	.w2(32'hba22173d),
	.w3(32'h3b0b78d1),
	.w4(32'h3ac6456f),
	.w5(32'hba2f5956),
	.w6(32'h3a8e21ee),
	.w7(32'h3a913fcf),
	.w8(32'h3ab3aa63),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a505b8b),
	.w1(32'h3a6789e5),
	.w2(32'h3b2f2371),
	.w3(32'hbad7a19b),
	.w4(32'h39a28f2b),
	.w5(32'h3a37e0b6),
	.w6(32'h39b642ef),
	.w7(32'h3a93e4d3),
	.w8(32'h3a81ca70),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae93537),
	.w1(32'h3b13067b),
	.w2(32'h3b1a3291),
	.w3(32'h3a19513e),
	.w4(32'h3af6404c),
	.w5(32'hbb1511a1),
	.w6(32'hba260a3b),
	.w7(32'hbabc380f),
	.w8(32'hbacf260d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba857ef2),
	.w1(32'hbb4f9062),
	.w2(32'hbb5289c1),
	.w3(32'hbb5d1498),
	.w4(32'hbb4dd2db),
	.w5(32'hba6bb443),
	.w6(32'hbadf8d9b),
	.w7(32'hbb4f8916),
	.w8(32'hba93d171),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3815cd19),
	.w1(32'h388ceeb4),
	.w2(32'h3a2dc4cc),
	.w3(32'h39378789),
	.w4(32'hb9f74387),
	.w5(32'hbac44b13),
	.w6(32'h3a61bb24),
	.w7(32'hba3cbcdd),
	.w8(32'hbb5431c4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2dd50),
	.w1(32'hbae78c57),
	.w2(32'hba6f5027),
	.w3(32'hbb02ed73),
	.w4(32'hbae835d8),
	.w5(32'hba26344f),
	.w6(32'hbaefa1ed),
	.w7(32'hbb02d94c),
	.w8(32'h3a400e9d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23fb52),
	.w1(32'h3a4ed8f3),
	.w2(32'h3a999663),
	.w3(32'h3b11170b),
	.w4(32'hb8a95f9c),
	.w5(32'hba8a5886),
	.w6(32'h3a598726),
	.w7(32'h38652152),
	.w8(32'h3aedd73c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dcf85),
	.w1(32'h3af49157),
	.w2(32'h3a7ee106),
	.w3(32'hbaaa681d),
	.w4(32'hbace8366),
	.w5(32'h38d36a65),
	.w6(32'h3a9064c3),
	.w7(32'h39c1220b),
	.w8(32'hb8db64e7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72a510),
	.w1(32'hbad3d9aa),
	.w2(32'hbaacdda7),
	.w3(32'h37478e67),
	.w4(32'h3a02da27),
	.w5(32'h3a9b29e1),
	.w6(32'h381065cb),
	.w7(32'hba2251f1),
	.w8(32'h3af0e412),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3e508),
	.w1(32'h3a934e0b),
	.w2(32'hb9aeeb92),
	.w3(32'h3ac3dad2),
	.w4(32'h39761faa),
	.w5(32'h3acbb527),
	.w6(32'h3a9afb31),
	.w7(32'h3a3b8002),
	.w8(32'h3a89fd49),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ef569),
	.w1(32'h3af23481),
	.w2(32'h399e1d97),
	.w3(32'h3afc6edd),
	.w4(32'h3b0a4d5e),
	.w5(32'h3a71e6e0),
	.w6(32'hba8e5691),
	.w7(32'h3a80a41a),
	.w8(32'h3a102ce9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a023ae1),
	.w1(32'hba7838ae),
	.w2(32'hb805f0cd),
	.w3(32'h384eefe7),
	.w4(32'h3895c079),
	.w5(32'hb989bb96),
	.w6(32'h38dfa088),
	.w7(32'h3a3d358f),
	.w8(32'hbab70f22),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae1646),
	.w1(32'hba8c2453),
	.w2(32'h3a90d88e),
	.w3(32'h3a8b70e3),
	.w4(32'hba2028de),
	.w5(32'h39d73d14),
	.w6(32'h398254c3),
	.w7(32'hb80f75c4),
	.w8(32'h3a0509ce),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af27f05),
	.w1(32'h3ad4a436),
	.w2(32'h39fd5f96),
	.w3(32'h39e17929),
	.w4(32'h3b0fe58c),
	.w5(32'h3a32cd61),
	.w6(32'hbac3d11e),
	.w7(32'hb99b80b0),
	.w8(32'hb9e1a175),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d25fa2),
	.w1(32'hbac5fbdb),
	.w2(32'hba2bbd55),
	.w3(32'hba9b38ba),
	.w4(32'hba159f3b),
	.w5(32'h3a0216ae),
	.w6(32'h3996e132),
	.w7(32'hbb02d5df),
	.w8(32'hb8d2b79e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d65314),
	.w1(32'hba53f7f5),
	.w2(32'hba5ce518),
	.w3(32'hb9aee596),
	.w4(32'hba0b6d34),
	.w5(32'h3ad2a465),
	.w6(32'h3a506104),
	.w7(32'hba83d5d9),
	.w8(32'hba0df136),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49fbe9),
	.w1(32'hba8c922d),
	.w2(32'hbae3ba3e),
	.w3(32'hbaa96b20),
	.w4(32'hba1b1575),
	.w5(32'h3a158f34),
	.w6(32'hbaeaee9c),
	.w7(32'hb9f2469b),
	.w8(32'h39dbb07f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b615ab),
	.w1(32'hbabb2c14),
	.w2(32'hba919409),
	.w3(32'h3a46ee7c),
	.w4(32'h3a41cb09),
	.w5(32'hbb8d2b87),
	.w6(32'h3a16fe43),
	.w7(32'h39b0d541),
	.w8(32'hbb52d604),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c4050),
	.w1(32'hbb33a783),
	.w2(32'hba994e02),
	.w3(32'hbb2f816d),
	.w4(32'hbb555725),
	.w5(32'hba753ee4),
	.w6(32'hb9f7a13a),
	.w7(32'hba94bd51),
	.w8(32'h3a8e2f4f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b9258),
	.w1(32'h3aeb3d56),
	.w2(32'h3a64cc47),
	.w3(32'hba59360c),
	.w4(32'h39b77c75),
	.w5(32'h3a7e4e7a),
	.w6(32'h3a67d991),
	.w7(32'hbaae0b93),
	.w8(32'h38fa8abc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe1c59),
	.w1(32'hbb09db0e),
	.w2(32'hba92d991),
	.w3(32'h3ab2c9c5),
	.w4(32'h3ad986b2),
	.w5(32'h3b030200),
	.w6(32'hb991bf31),
	.w7(32'hb91b4132),
	.w8(32'hba221b3b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd232f),
	.w1(32'hbb1b9564),
	.w2(32'hbaa2378d),
	.w3(32'h3a1bfdb2),
	.w4(32'h3aaab3f9),
	.w5(32'h3ac23f46),
	.w6(32'hbb1783ec),
	.w7(32'hbb62b916),
	.w8(32'h3a2294ae),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02aed7),
	.w1(32'h3a756203),
	.w2(32'h3a0668c9),
	.w3(32'h3a49b5a7),
	.w4(32'h3af6dff5),
	.w5(32'h3a97c4a9),
	.w6(32'h3b206993),
	.w7(32'hb8b63c6e),
	.w8(32'hbaf2a494),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94b4d8),
	.w1(32'h3a087c80),
	.w2(32'h3a41434b),
	.w3(32'h3a0467a2),
	.w4(32'h3b7bcbd7),
	.w5(32'hbab9a702),
	.w6(32'hbab45e58),
	.w7(32'h3a2129f8),
	.w8(32'hba30d299),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00996b),
	.w1(32'h39e1694c),
	.w2(32'h3a770cdb),
	.w3(32'hba931f6b),
	.w4(32'hb91e7ee5),
	.w5(32'hbac7fc9e),
	.w6(32'hba65bfee),
	.w7(32'h3858c95d),
	.w8(32'h367a8c64),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae177c2),
	.w1(32'hbac164f8),
	.w2(32'hbac5264d),
	.w3(32'h3a6794b8),
	.w4(32'h3a1cf3b6),
	.w5(32'hba7dc1f5),
	.w6(32'h3a4520ba),
	.w7(32'hb8e8ace3),
	.w8(32'h3a6f4d0f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b153f8c),
	.w1(32'h3a936d14),
	.w2(32'h3b12f5e7),
	.w3(32'hb75b8b9e),
	.w4(32'hba5e5648),
	.w5(32'h3aa4b24e),
	.w6(32'h3a0d25a8),
	.w7(32'hba97be21),
	.w8(32'hb9714c9a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8dfad),
	.w1(32'h3aa72535),
	.w2(32'hba087079),
	.w3(32'h3a999dbb),
	.w4(32'h3b32b80a),
	.w5(32'hb94ab278),
	.w6(32'h3a17c0a8),
	.w7(32'h3a3d4f2f),
	.w8(32'h388e3528),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d41385),
	.w1(32'h3b072b46),
	.w2(32'h3a191428),
	.w3(32'hbb0f59e9),
	.w4(32'hba7fdec5),
	.w5(32'hbadf9855),
	.w6(32'hbaa68b75),
	.w7(32'hbac486c0),
	.w8(32'hba9a5273),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5acd07),
	.w1(32'h3a50b2ec),
	.w2(32'h3a99a710),
	.w3(32'hb9be7776),
	.w4(32'h399e979d),
	.w5(32'h38f6a6aa),
	.w6(32'h38a4fdb3),
	.w7(32'hb84e0a84),
	.w8(32'hba5c93e2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdceed),
	.w1(32'hba13839d),
	.w2(32'hba1fe1b7),
	.w3(32'hba82cf36),
	.w4(32'hbabad85a),
	.w5(32'hb97370fe),
	.w6(32'hbb1b5ac4),
	.w7(32'hbac281af),
	.w8(32'h3abae069),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a80c4),
	.w1(32'hbaf7e8db),
	.w2(32'hba097c38),
	.w3(32'hbb213d18),
	.w4(32'hbb154de0),
	.w5(32'h3aeaa2da),
	.w6(32'h3b02ab5a),
	.w7(32'h3ab57a6a),
	.w8(32'hbaac7bd6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28ecb1),
	.w1(32'h3a705f4d),
	.w2(32'h3aa20ecc),
	.w3(32'hb9b25c4f),
	.w4(32'h39028302),
	.w5(32'hbaa0d1d7),
	.w6(32'h3ae89490),
	.w7(32'h3aca80bc),
	.w8(32'h3a24a4d3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9703cdf),
	.w1(32'hba8e8768),
	.w2(32'hba2fc0dd),
	.w3(32'hba634241),
	.w4(32'h3a1d5afb),
	.w5(32'h39bb4395),
	.w6(32'h38faa578),
	.w7(32'h39c8997b),
	.w8(32'h3ac6eb96),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb63c4),
	.w1(32'h3b15e4e2),
	.w2(32'h3b368e3d),
	.w3(32'h39116abf),
	.w4(32'hb9fea67a),
	.w5(32'hb9908f09),
	.w6(32'h3b4025ad),
	.w7(32'h3aa2e037),
	.w8(32'h386401f6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d0e1d),
	.w1(32'hba4f72ea),
	.w2(32'hb8cdb12b),
	.w3(32'h39a78d73),
	.w4(32'h391b3960),
	.w5(32'h3850d765),
	.w6(32'h39c0bbb5),
	.w7(32'hba36a132),
	.w8(32'hba1ae5bc),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a943650),
	.w1(32'hb918c13c),
	.w2(32'hbb5cfa6d),
	.w3(32'hb987d7d1),
	.w4(32'h3a12c9f3),
	.w5(32'hb7361a89),
	.w6(32'hbb018032),
	.w7(32'hbaa8f5e4),
	.w8(32'h3866b96d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02e569),
	.w1(32'hbb03bc7a),
	.w2(32'hba16e9bb),
	.w3(32'h3ad80c1f),
	.w4(32'h387c0e23),
	.w5(32'hbaba0413),
	.w6(32'h3a4a4879),
	.w7(32'hb9564af8),
	.w8(32'hb94057cc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a18da),
	.w1(32'hbaae5b0b),
	.w2(32'hbae83b9e),
	.w3(32'h39bc6b72),
	.w4(32'hba8b8d5c),
	.w5(32'hb9de9619),
	.w6(32'h39eac091),
	.w7(32'h3861f132),
	.w8(32'hb8f61366),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f59fd),
	.w1(32'hbada4b23),
	.w2(32'h3ab8ba27),
	.w3(32'hbb1a7143),
	.w4(32'hbb3886bd),
	.w5(32'hba706718),
	.w6(32'hbb108dfd),
	.w7(32'hba2094f0),
	.w8(32'h3a88c67a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba903cff),
	.w1(32'hb8a1c0ef),
	.w2(32'h3a788454),
	.w3(32'hbaebfa39),
	.w4(32'hba9d0dae),
	.w5(32'h39b67308),
	.w6(32'h3b262e21),
	.w7(32'h3ac577c4),
	.w8(32'h3ac2936d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99dcb2),
	.w1(32'h3aa20046),
	.w2(32'hba06e1f1),
	.w3(32'h3a762157),
	.w4(32'h3a8b9945),
	.w5(32'h3ad75e54),
	.w6(32'h3b662968),
	.w7(32'h3b107fdf),
	.w8(32'h3b5d9c0c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92d95d),
	.w1(32'h3b57a3a5),
	.w2(32'h3ba6069a),
	.w3(32'h3b07ca8d),
	.w4(32'h3b818d60),
	.w5(32'hba7ea71c),
	.w6(32'h3b4e0873),
	.w7(32'h3ba6187c),
	.w8(32'h38b30c69),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17eec0),
	.w1(32'h3b00a714),
	.w2(32'h3aec2ffc),
	.w3(32'h3a5f286e),
	.w4(32'h3a8839a9),
	.w5(32'hbb189f77),
	.w6(32'h3b69f019),
	.w7(32'h3b3092d2),
	.w8(32'hba356f43),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e157bc),
	.w1(32'hba800e52),
	.w2(32'hbb0a80c3),
	.w3(32'h3a032110),
	.w4(32'hba376365),
	.w5(32'h3b1127a4),
	.w6(32'h3b11eba2),
	.w7(32'hba3c5661),
	.w8(32'h3a0fcba8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc662e),
	.w1(32'hb8e20665),
	.w2(32'h3a21cc13),
	.w3(32'h394faf08),
	.w4(32'h3a963922),
	.w5(32'hba9b735a),
	.w6(32'h3a8fa8a7),
	.w7(32'h3a0b0906),
	.w8(32'hb9c0eae4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08045c),
	.w1(32'hb9f39706),
	.w2(32'h3945e753),
	.w3(32'hba4dfea9),
	.w4(32'h39c0c0f2),
	.w5(32'h393fa8b1),
	.w6(32'h3a6372a3),
	.w7(32'hb9af8249),
	.w8(32'h3a3ee03a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa15cf5),
	.w1(32'hbacae3e8),
	.w2(32'hbac965aa),
	.w3(32'hb881ce0a),
	.w4(32'hb9d240bc),
	.w5(32'hbaebcc19),
	.w6(32'hba029344),
	.w7(32'hba3660be),
	.w8(32'hbabe9004),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac540f1),
	.w1(32'h3b935387),
	.w2(32'h396738ba),
	.w3(32'h3b5794b3),
	.w4(32'h3ad22e0a),
	.w5(32'hbade557d),
	.w6(32'h3b0f8ca9),
	.w7(32'h3a81baa9),
	.w8(32'h3ab31293),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10763e),
	.w1(32'hb9a4dd6b),
	.w2(32'h38961e8f),
	.w3(32'hbab2009d),
	.w4(32'h3a30210c),
	.w5(32'hbaa4b64b),
	.w6(32'hbb45e599),
	.w7(32'h398e4815),
	.w8(32'hba77a8e5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5aa75),
	.w1(32'h3b6df70f),
	.w2(32'hb9221a46),
	.w3(32'h3987638f),
	.w4(32'h3b93101d),
	.w5(32'hba0bf28e),
	.w6(32'h39a2a785),
	.w7(32'h39efb8fd),
	.w8(32'hbb4861ff),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b154bee),
	.w1(32'h39e8c2ac),
	.w2(32'hb9ddb9a1),
	.w3(32'hba41a47c),
	.w4(32'hba35f741),
	.w5(32'h3a872db2),
	.w6(32'hbad905bc),
	.w7(32'hbb2592b9),
	.w8(32'h3a727a75),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1adb24),
	.w1(32'h3a9dab26),
	.w2(32'h3b0d2ca5),
	.w3(32'h3b3dd27d),
	.w4(32'h3b61aa10),
	.w5(32'h3a2b6d82),
	.w6(32'h3b02fee0),
	.w7(32'h3b227aee),
	.w8(32'h393e07d8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e91584),
	.w1(32'hb93d5c3f),
	.w2(32'hba8f402c),
	.w3(32'h3a9d3ec6),
	.w4(32'h3ade9cc7),
	.w5(32'hbaba9376),
	.w6(32'h3931a3cd),
	.w7(32'h3a479627),
	.w8(32'hb6c09c57),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad15050),
	.w1(32'hba6a07f4),
	.w2(32'hba90da13),
	.w3(32'hb9802413),
	.w4(32'h3abada81),
	.w5(32'h3a9f66da),
	.w6(32'h3aa2184a),
	.w7(32'h3b19dbdd),
	.w8(32'h3a8c2de1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba686d),
	.w1(32'hba0c2507),
	.w2(32'h3a80984a),
	.w3(32'h3b3c23c2),
	.w4(32'h3a4cb359),
	.w5(32'h3b2618a7),
	.w6(32'h3ac924e1),
	.w7(32'h3aed3563),
	.w8(32'h3ac45351),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4f462),
	.w1(32'hba86e501),
	.w2(32'h3a0103a8),
	.w3(32'h3b651b97),
	.w4(32'h3b2b1a98),
	.w5(32'hbaee9cbf),
	.w6(32'h3ab687cc),
	.w7(32'h3a4c01d9),
	.w8(32'h3ba6c662),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f32dd),
	.w1(32'hbc5806ae),
	.w2(32'hbc813582),
	.w3(32'h3c8520ba),
	.w4(32'hbb42a157),
	.w5(32'h3c8c4dcd),
	.w6(32'h3b0f949d),
	.w7(32'hbbcc9bab),
	.w8(32'h3c37647e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2278fd),
	.w1(32'hbcc87000),
	.w2(32'hbc363496),
	.w3(32'h3d140b78),
	.w4(32'h3b98a55d),
	.w5(32'h3c7fdae0),
	.w6(32'hbbab69ca),
	.w7(32'hba20d4a2),
	.w8(32'h3c47359a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16d186),
	.w1(32'hbcfe8553),
	.w2(32'hbc9d7d51),
	.w3(32'h3cd2d751),
	.w4(32'h3c28ae9a),
	.w5(32'h3bb0fe5d),
	.w6(32'hb9cb428c),
	.w7(32'hbc437257),
	.w8(32'hbc54df83),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd88ab2),
	.w1(32'hbae48034),
	.w2(32'hbbd8e222),
	.w3(32'hbc166dd2),
	.w4(32'hbb339577),
	.w5(32'h3944d6a4),
	.w6(32'hbbaa1050),
	.w7(32'hba82d567),
	.w8(32'hbaf57b1b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39362bb0),
	.w1(32'h3a66451b),
	.w2(32'h3b391a84),
	.w3(32'h39eea044),
	.w4(32'hbb951b19),
	.w5(32'h3d452c3b),
	.w6(32'h3bfc1132),
	.w7(32'h3b3c56bc),
	.w8(32'h3cb1c515),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c45cd),
	.w1(32'hbd91abe2),
	.w2(32'hbd3d240a),
	.w3(32'h3d8bc032),
	.w4(32'h3ce75326),
	.w5(32'hbb941d08),
	.w6(32'hbc295b95),
	.w7(32'hbccb5339),
	.w8(32'h3ab052e4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9e482),
	.w1(32'h3b04189b),
	.w2(32'h3a8ad51f),
	.w3(32'hbc07d6b4),
	.w4(32'hbbe9b703),
	.w5(32'h3c21368f),
	.w6(32'hbb4b7fa5),
	.w7(32'hbc27736d),
	.w8(32'h3c016925),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa19723),
	.w1(32'hbc4f071a),
	.w2(32'hbc8889bc),
	.w3(32'h3c5dcca7),
	.w4(32'h3b1712f9),
	.w5(32'hbc191ada),
	.w6(32'h3b43beed),
	.w7(32'hbb9c8df4),
	.w8(32'hbada7ae1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9385f0),
	.w1(32'h3ac0ba5e),
	.w2(32'hbbb756ae),
	.w3(32'h3c087061),
	.w4(32'h39f1ca3f),
	.w5(32'h3bc7ee90),
	.w6(32'h3c9f7b74),
	.w7(32'h3bcc5ad8),
	.w8(32'h3c515a3b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c218f2c),
	.w1(32'h3c21e1d7),
	.w2(32'hbb462a9d),
	.w3(32'hb9ae2671),
	.w4(32'hbb8a869e),
	.w5(32'h3c441188),
	.w6(32'h3bcf304e),
	.w7(32'h358f49f1),
	.w8(32'h3c55ea6f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf149e7),
	.w1(32'hbbf8a01e),
	.w2(32'hbc3b4376),
	.w3(32'h3cb60d14),
	.w4(32'h3c06db11),
	.w5(32'hbc6a4996),
	.w6(32'h3bfaea65),
	.w7(32'h3b3f5350),
	.w8(32'hbb9e8a89),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b049f),
	.w1(32'h3c0737c0),
	.w2(32'h3bfbb920),
	.w3(32'hbca156e8),
	.w4(32'hbc875cca),
	.w5(32'hbbec63dc),
	.w6(32'hbb42837f),
	.w7(32'h3a5a5272),
	.w8(32'h3b222636),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fe6d6),
	.w1(32'h3c339ac4),
	.w2(32'hbbf49b86),
	.w3(32'h3c38d5ba),
	.w4(32'hba75a340),
	.w5(32'hbba7d277),
	.w6(32'h3c04b128),
	.w7(32'h3b4dcc34),
	.w8(32'h3b1d4651),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb424a3b),
	.w1(32'h37b4432c),
	.w2(32'h3b32cedf),
	.w3(32'h3a18dfdf),
	.w4(32'h3b4d5df8),
	.w5(32'hbd14c02b),
	.w6(32'h3c693cb6),
	.w7(32'h3be1a2ab),
	.w8(32'hbc5efdb7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cf75c),
	.w1(32'h3d2b0336),
	.w2(32'h3cce9318),
	.w3(32'hbd210507),
	.w4(32'hbc7b5166),
	.w5(32'h384f7da8),
	.w6(32'h3bb7ad6f),
	.w7(32'h3bdb9b0d),
	.w8(32'hbb958e11),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37dbc7),
	.w1(32'hbbb08ab8),
	.w2(32'hbb9fb2cc),
	.w3(32'hbb4163d0),
	.w4(32'hbb28c135),
	.w5(32'h3c69e18b),
	.w6(32'h3c09fb66),
	.w7(32'hbb5c19c6),
	.w8(32'h3c1d4712),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5814d),
	.w1(32'hbc26c56d),
	.w2(32'hbc871b48),
	.w3(32'h3cdc035a),
	.w4(32'hba6da100),
	.w5(32'hbbfdef87),
	.w6(32'h39e8df42),
	.w7(32'hbc036bcb),
	.w8(32'hbbc6f78b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab62f6),
	.w1(32'hbb9140fe),
	.w2(32'hbb5be39e),
	.w3(32'hbafeaa4f),
	.w4(32'hbc355743),
	.w5(32'h3a986d4a),
	.w6(32'h3c87e936),
	.w7(32'hbb2eee3f),
	.w8(32'h3ae15ac6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf9cc9),
	.w1(32'hb9806c21),
	.w2(32'hbba8e5d2),
	.w3(32'hbb0718a9),
	.w4(32'hbbc67dea),
	.w5(32'h3c48d513),
	.w6(32'hb90034fb),
	.w7(32'h3a8bef6a),
	.w8(32'h3b04ed10),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0d11d),
	.w1(32'hbc356a93),
	.w2(32'hbbd91a5a),
	.w3(32'h3c3368a5),
	.w4(32'h3acd49f9),
	.w5(32'hbb0f54ac),
	.w6(32'hb9334af6),
	.w7(32'hbbf2bbfc),
	.w8(32'hbac8acb0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e766b),
	.w1(32'hbce12478),
	.w2(32'hbc8230c6),
	.w3(32'h3c96bd2d),
	.w4(32'hbb88fa6c),
	.w5(32'h3c8c7e85),
	.w6(32'hbbf23604),
	.w7(32'hbc395212),
	.w8(32'h3ca33c64),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1b053),
	.w1(32'hbd640c31),
	.w2(32'hbd0d4a92),
	.w3(32'h3d380b65),
	.w4(32'h3c898e59),
	.w5(32'h3b2b3e55),
	.w6(32'hbbed7cc5),
	.w7(32'hbc541b88),
	.w8(32'hbaffe77f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39291d9e),
	.w1(32'h3b5d0e39),
	.w2(32'hbbdf94c4),
	.w3(32'hbb8cd8a9),
	.w4(32'hba9ada95),
	.w5(32'hbbc08b5b),
	.w6(32'h3ca666dd),
	.w7(32'hb9bbbc64),
	.w8(32'hbb879586),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9949b1),
	.w1(32'h3c5a2ce0),
	.w2(32'h3cb90765),
	.w3(32'hbc621ec4),
	.w4(32'hbc2b92a1),
	.w5(32'hbc116fe2),
	.w6(32'hbbeaaec6),
	.w7(32'h3c8fd854),
	.w8(32'hbc28a84a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d1c02),
	.w1(32'h3ca5c0d8),
	.w2(32'h3c64d434),
	.w3(32'hbca68707),
	.w4(32'hbb4f09f3),
	.w5(32'hbc8f6d1c),
	.w6(32'h3c00cb35),
	.w7(32'h3c894220),
	.w8(32'hbc19e146),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17868a),
	.w1(32'h3d0279a5),
	.w2(32'h3c9fefcb),
	.w3(32'hbcb7e5fa),
	.w4(32'hbb7590b9),
	.w5(32'hbb783241),
	.w6(32'h3bf20ec9),
	.w7(32'h3c46f2c9),
	.w8(32'hbc6d4686),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd0a78),
	.w1(32'h3ca84fa0),
	.w2(32'h3c7876dc),
	.w3(32'hbc506a37),
	.w4(32'h39ea960b),
	.w5(32'hbb0c0453),
	.w6(32'hbc18c1be),
	.w7(32'h3aa3a3d6),
	.w8(32'hbbaf45cb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e150),
	.w1(32'hbb363e28),
	.w2(32'h3aecec89),
	.w3(32'hbb7001f1),
	.w4(32'hbae8cd84),
	.w5(32'hb917fc3e),
	.w6(32'hbb521881),
	.w7(32'hbb0f54fc),
	.w8(32'hbbb44030),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb671770),
	.w1(32'h3c09b5c4),
	.w2(32'h3bedef77),
	.w3(32'hba32a654),
	.w4(32'h3a16b6c7),
	.w5(32'hba1a1bab),
	.w6(32'h3a87c0a7),
	.w7(32'h39c91e23),
	.w8(32'h3a9e3757),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4eed9c),
	.w1(32'h39865d2b),
	.w2(32'hbb498977),
	.w3(32'h3ba071b9),
	.w4(32'h3c3855a6),
	.w5(32'hbc27ed3c),
	.w6(32'hbc031e94),
	.w7(32'hbb0964de),
	.w8(32'hb7741874),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2634a),
	.w1(32'h3c236295),
	.w2(32'h3b462399),
	.w3(32'hbc38814a),
	.w4(32'hbc5e4ce8),
	.w5(32'hbc95676e),
	.w6(32'h3b3cb070),
	.w7(32'hba144e48),
	.w8(32'hbb3eed4b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc5360),
	.w1(32'h3ca302d6),
	.w2(32'h3c7496a8),
	.w3(32'hbc95c1a3),
	.w4(32'h398fc82e),
	.w5(32'h3bc318b3),
	.w6(32'h3bbf065b),
	.w7(32'h3a87b205),
	.w8(32'hbb31e210),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e184e),
	.w1(32'hbbf113d6),
	.w2(32'h3c3fdcd5),
	.w3(32'h3c13098b),
	.w4(32'h3b882e75),
	.w5(32'h3c04caf7),
	.w6(32'hbb764dbe),
	.w7(32'h3b0d12aa),
	.w8(32'h3b4e9dc9),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98983c),
	.w1(32'hbbadc0c5),
	.w2(32'hbc4e4342),
	.w3(32'h3beaafbc),
	.w4(32'h3b963d1d),
	.w5(32'h3b04510e),
	.w6(32'h3b40babf),
	.w7(32'hba9fd441),
	.w8(32'hbd3a0a3e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5aef6c),
	.w1(32'hb944d9f2),
	.w2(32'h3c5fe387),
	.w3(32'h39bc9927),
	.w4(32'h3b25a235),
	.w5(32'hbc008bb8),
	.w6(32'hbcaad6f7),
	.w7(32'hbcb8d797),
	.w8(32'hbba7b6c9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42f6c8),
	.w1(32'hb994ebb1),
	.w2(32'hbbd27878),
	.w3(32'hbc807693),
	.w4(32'hbc649ddb),
	.w5(32'hbb35946d),
	.w6(32'hbb9f92b9),
	.w7(32'hbac9cba0),
	.w8(32'hbb147ffc),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d1f71),
	.w1(32'h3ba5c7d4),
	.w2(32'h3af0638e),
	.w3(32'hbc1097d6),
	.w4(32'hbc0b3bf9),
	.w5(32'hbb17bb10),
	.w6(32'hbb459e2c),
	.w7(32'h3a7b3633),
	.w8(32'h3bf6ad4f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd71f32),
	.w1(32'h3b54825a),
	.w2(32'hbb43f7ec),
	.w3(32'h3a24169d),
	.w4(32'hbb146823),
	.w5(32'hbca0351c),
	.w6(32'h3adb921a),
	.w7(32'h3b0e6b80),
	.w8(32'hbbc2ed8e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b483fc5),
	.w1(32'h3cb0f080),
	.w2(32'h3c85a983),
	.w3(32'hbcb61337),
	.w4(32'hbc80956d),
	.w5(32'hbbc19611),
	.w6(32'h3b5b2620),
	.w7(32'h3beb830e),
	.w8(32'hbb642773),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e0203),
	.w1(32'hb9a6d595),
	.w2(32'hbbbb49d2),
	.w3(32'hbc218242),
	.w4(32'hbc3c8a8d),
	.w5(32'h3c1c1e62),
	.w6(32'hbb81e934),
	.w7(32'hbb649190),
	.w8(32'hb9e0411d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89ef57),
	.w1(32'hbb89b36b),
	.w2(32'hbc78026b),
	.w3(32'hbad578d3),
	.w4(32'hbbcc6d32),
	.w5(32'h3bb612d5),
	.w6(32'hbbf39c92),
	.w7(32'h3af64c01),
	.w8(32'hba8dc1a1),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabee785),
	.w1(32'hbc072c3c),
	.w2(32'h3b80d2f5),
	.w3(32'h3ba4442f),
	.w4(32'h3b55febd),
	.w5(32'hbcaa019d),
	.w6(32'h399b168c),
	.w7(32'hbc84a1de),
	.w8(32'hbc91608c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5371ad),
	.w1(32'h3cb95a0d),
	.w2(32'h3ccd6fd0),
	.w3(32'hbd0e8b42),
	.w4(32'hbc2ec8aa),
	.w5(32'h3b5517a5),
	.w6(32'hba2a0783),
	.w7(32'h3c04ae89),
	.w8(32'h3aca6b5d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c6361),
	.w1(32'h3a53e949),
	.w2(32'hbaf37785),
	.w3(32'h396d6113),
	.w4(32'h39d16310),
	.w5(32'hbb396f4a),
	.w6(32'hba391ad5),
	.w7(32'hbc170938),
	.w8(32'hbbfa953f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d6ac8),
	.w1(32'h3c071f6e),
	.w2(32'hbc16885f),
	.w3(32'hbbfc52eb),
	.w4(32'hbbbbfd94),
	.w5(32'hbc491e45),
	.w6(32'hbbbd96a1),
	.w7(32'hbb91aaf9),
	.w8(32'hbbf604ec),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398530be),
	.w1(32'h3c8640ed),
	.w2(32'h3c4e1e7a),
	.w3(32'hbc5e5e20),
	.w4(32'hbc1761a5),
	.w5(32'hbc4d00cb),
	.w6(32'hb9c8fc72),
	.w7(32'h3c0de5e2),
	.w8(32'h3acaade8),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8539ea),
	.w1(32'h3c97c08f),
	.w2(32'h3b568de3),
	.w3(32'hbcc1c5b7),
	.w4(32'hbbc87e1b),
	.w5(32'h3c148c9b),
	.w6(32'h3c030213),
	.w7(32'h3c3fa905),
	.w8(32'h3bf2db6f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bd2eb),
	.w1(32'hbc039fef),
	.w2(32'hbbaa3526),
	.w3(32'h3c8fb22e),
	.w4(32'h3bf7d7be),
	.w5(32'h3c0997c4),
	.w6(32'h3ba23b16),
	.w7(32'h3bdf945c),
	.w8(32'hbad827cd),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc103f77),
	.w1(32'hbcc4b325),
	.w2(32'hbcc3d136),
	.w3(32'h3c9762eb),
	.w4(32'h3c1176cb),
	.w5(32'hbb4feff3),
	.w6(32'h3b2375f5),
	.w7(32'hbb859617),
	.w8(32'hbb02c24d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5307e),
	.w1(32'hbbe1a400),
	.w2(32'hbb9c502a),
	.w3(32'hb9c7f68f),
	.w4(32'h3babcada),
	.w5(32'hbaba8361),
	.w6(32'hbba5c51b),
	.w7(32'h39588ef7),
	.w8(32'hbc1991b5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8feb829),
	.w1(32'h3c946b74),
	.w2(32'h3c80fe49),
	.w3(32'hbc3cef1f),
	.w4(32'hbbe66991),
	.w5(32'h3bfa901e),
	.w6(32'hbbfed1cc),
	.w7(32'h3c05ce5c),
	.w8(32'h3bd8909e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb756d59),
	.w1(32'hbc2b07b1),
	.w2(32'hbc5df34a),
	.w3(32'h3c4168f8),
	.w4(32'h3a84f83a),
	.w5(32'h3ae0acf2),
	.w6(32'h3a8bb26c),
	.w7(32'hbb8dbe58),
	.w8(32'hbb76cd6e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf1216),
	.w1(32'hbb34ec64),
	.w2(32'h3b90e605),
	.w3(32'h39ba9a6b),
	.w4(32'hb793489c),
	.w5(32'hbc2551f3),
	.w6(32'h3bffc883),
	.w7(32'h3b4983a8),
	.w8(32'hbc15863e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab850b),
	.w1(32'h3ce7d73e),
	.w2(32'h3b143cdc),
	.w3(32'hbcae60b9),
	.w4(32'hbc05b68c),
	.w5(32'hbb32c7ed),
	.w6(32'h3b3e362a),
	.w7(32'h39a7158e),
	.w8(32'hb91c1749),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde3647),
	.w1(32'hbbb53d39),
	.w2(32'hbb11d073),
	.w3(32'hbbcc68a5),
	.w4(32'hbbe9f293),
	.w5(32'hb99e2dbc),
	.w6(32'h3cbaf70d),
	.w7(32'h3b7f2622),
	.w8(32'h3b59dbf3),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb0b4a),
	.w1(32'h3b8d108d),
	.w2(32'hbc446ce7),
	.w3(32'hbbb76b76),
	.w4(32'h3ac30a06),
	.w5(32'h3c134b9b),
	.w6(32'hbafe56b0),
	.w7(32'hbaefcd17),
	.w8(32'h3b8cd8f7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7baa84),
	.w1(32'hbbc9bdfd),
	.w2(32'hbaf36b72),
	.w3(32'h3c2092d3),
	.w4(32'h3bfd50bd),
	.w5(32'hbca19021),
	.w6(32'h3b9b24ae),
	.w7(32'h3b2a1c91),
	.w8(32'hbc05d811),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bcba8),
	.w1(32'h3c62bb0f),
	.w2(32'h3c5323d6),
	.w3(32'hbcc28c31),
	.w4(32'hbc9a1599),
	.w5(32'h3a74f584),
	.w6(32'hba2ffb33),
	.w7(32'h3b06b33c),
	.w8(32'hbbc580a6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092e65),
	.w1(32'hbb81ccc4),
	.w2(32'hbb620c47),
	.w3(32'h3b4869cd),
	.w4(32'hbb84dbe0),
	.w5(32'hbc1af017),
	.w6(32'h3b384c67),
	.w7(32'h3bdadcb1),
	.w8(32'hbb8e0621),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984a53d),
	.w1(32'h3c79bb75),
	.w2(32'h3c04dba4),
	.w3(32'hbc861948),
	.w4(32'hbb7ebe88),
	.w5(32'h3bfb4c14),
	.w6(32'hb82ca4ee),
	.w7(32'h3bbfc909),
	.w8(32'hbbc01f87),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1b1f3),
	.w1(32'h3b831c0f),
	.w2(32'h3c4db0bc),
	.w3(32'h3ba4af9c),
	.w4(32'h3ad7cefe),
	.w5(32'hbb0dd7ff),
	.w6(32'hb9f6e1f6),
	.w7(32'hbba84a52),
	.w8(32'hbb0cfa51),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa1e61),
	.w1(32'h3ae93482),
	.w2(32'h3bff8c3a),
	.w3(32'h3bc1f2f9),
	.w4(32'hbb67a2c6),
	.w5(32'h3bf2b48a),
	.w6(32'hbc3a21ec),
	.w7(32'hbc5e44e4),
	.w8(32'h3ad31d9e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36e8ce),
	.w1(32'hbc3635ae),
	.w2(32'h3bc67052),
	.w3(32'h3c000da9),
	.w4(32'h3b6d8129),
	.w5(32'h3c1b54d0),
	.w6(32'h3aabc155),
	.w7(32'hbb8ab6a8),
	.w8(32'h3bd826a0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd189d),
	.w1(32'hbc08fda8),
	.w2(32'hbc874f31),
	.w3(32'h3c6c9576),
	.w4(32'h3be60a53),
	.w5(32'h3be688e1),
	.w6(32'h3b3c7fa8),
	.w7(32'h3911a904),
	.w8(32'h3abe9385),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e89ea),
	.w1(32'hbc351dc9),
	.w2(32'hbbdf3de7),
	.w3(32'hbb8073a6),
	.w4(32'hbb4b4ed8),
	.w5(32'hbbcda6d4),
	.w6(32'h39f77b5f),
	.w7(32'hbb680533),
	.w8(32'hbbe498cc),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb03af3),
	.w1(32'h3bd3aa43),
	.w2(32'h39fedfc6),
	.w3(32'h39442b26),
	.w4(32'h39d0bd3b),
	.w5(32'h3ae6dddb),
	.w6(32'h3a177329),
	.w7(32'hbad54864),
	.w8(32'hbb20ec2e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a8d91),
	.w1(32'hb98c27c8),
	.w2(32'hbb63d0ca),
	.w3(32'h3ab1afdf),
	.w4(32'h3b866d09),
	.w5(32'h3ba02b10),
	.w6(32'hbb00173d),
	.w7(32'hbc25012a),
	.w8(32'h3b88c187),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a3e3a),
	.w1(32'hbb3bf554),
	.w2(32'hbbc37786),
	.w3(32'h3c1fae8f),
	.w4(32'h3bbfdb28),
	.w5(32'hbc3996f8),
	.w6(32'h3c216608),
	.w7(32'h3b036a99),
	.w8(32'hbc5791dd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda52b6),
	.w1(32'h3cb69c2b),
	.w2(32'h3be75207),
	.w3(32'hbc85de7c),
	.w4(32'hbb967c7f),
	.w5(32'h3cb37cd3),
	.w6(32'h3bff3be1),
	.w7(32'h3be661df),
	.w8(32'h3c9db56a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8582b5),
	.w1(32'hbd507d79),
	.w2(32'hbcd2b6e6),
	.w3(32'h3d25b761),
	.w4(32'h3c78c974),
	.w5(32'hbc0bb027),
	.w6(32'hbc0fa859),
	.w7(32'hbab55dab),
	.w8(32'hbabbba5c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83861f),
	.w1(32'hbaaa2c5d),
	.w2(32'h3b216109),
	.w3(32'hbbc0fc89),
	.w4(32'hbb8eaa4f),
	.w5(32'h3bbcba05),
	.w6(32'h3ba63da5),
	.w7(32'h3a035f9a),
	.w8(32'h3b463141),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8dbe9),
	.w1(32'hbb777002),
	.w2(32'hbc62fb8b),
	.w3(32'h3b3e76b2),
	.w4(32'h3b71b267),
	.w5(32'h3a498297),
	.w6(32'hbba15d65),
	.w7(32'hbc12c3d2),
	.w8(32'h3c360d56),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0f627),
	.w1(32'hbbf80c0a),
	.w2(32'h3b1e3610),
	.w3(32'h3c6c69a0),
	.w4(32'h3b65b16b),
	.w5(32'hbb93a8da),
	.w6(32'h3a842011),
	.w7(32'hbb68d174),
	.w8(32'hbb1e6718),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70558b),
	.w1(32'h3bc28015),
	.w2(32'h3b471d85),
	.w3(32'hbbb7032a),
	.w4(32'hbb8498a9),
	.w5(32'h3c917111),
	.w6(32'h3b9181cb),
	.w7(32'h3c30b74d),
	.w8(32'h3c95607f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c3c2a),
	.w1(32'hbd4dc8d8),
	.w2(32'hbd26bb5f),
	.w3(32'h3d2cd5a6),
	.w4(32'h3c49283c),
	.w5(32'h3beec4e3),
	.w6(32'hbc1f4aa6),
	.w7(32'hbc9685f6),
	.w8(32'h3aef9f61),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9328f),
	.w1(32'hba45b18a),
	.w2(32'h383d85b6),
	.w3(32'h3ba2e0da),
	.w4(32'h38b62a78),
	.w5(32'h3cb111ce),
	.w6(32'h3add0f02),
	.w7(32'hbc01a8d9),
	.w8(32'h3b928dc5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50ecd4),
	.w1(32'hbd0c68b7),
	.w2(32'hbca0a24b),
	.w3(32'h3ce66907),
	.w4(32'h3c80af2c),
	.w5(32'hbc9a7bb1),
	.w6(32'hbba380cb),
	.w7(32'hbc62df74),
	.w8(32'hbc7f1c25),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b2e63),
	.w1(32'h3d1dde12),
	.w2(32'h3d040e8c),
	.w3(32'hbce6afea),
	.w4(32'hbc24f989),
	.w5(32'hbc78b503),
	.w6(32'h3b794a9e),
	.w7(32'h3c2cf9d1),
	.w8(32'hbc3f4a98),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5393a8),
	.w1(32'h3ce08e91),
	.w2(32'h3ce8ef2b),
	.w3(32'hbca199bd),
	.w4(32'hbc1c9afc),
	.w5(32'h3c0f6f8a),
	.w6(32'hbb9834dd),
	.w7(32'h3c1ca188),
	.w8(32'h3bbc16e3),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb656a1f),
	.w1(32'hbbf3e53b),
	.w2(32'hbc2b4315),
	.w3(32'h3c36cc66),
	.w4(32'h3b963bc9),
	.w5(32'h3c3ef809),
	.w6(32'h3bb54e81),
	.w7(32'hb98948a3),
	.w8(32'hbb3b252d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1bdec),
	.w1(32'h3bca53f0),
	.w2(32'hba951455),
	.w3(32'h3b65190a),
	.w4(32'hbc840ae1),
	.w5(32'h3c9ef7e1),
	.w6(32'hbbded7c9),
	.w7(32'hbb66aa0f),
	.w8(32'hba9111ec),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9004d2),
	.w1(32'hbc77a55c),
	.w2(32'hbc637f94),
	.w3(32'h3ca85afb),
	.w4(32'hb9ac9daa),
	.w5(32'h3c190ca1),
	.w6(32'h398cd2aa),
	.w7(32'hbc89e6ac),
	.w8(32'hbb150914),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74309a),
	.w1(32'hba491c2d),
	.w2(32'hbbd46076),
	.w3(32'h3b1931ed),
	.w4(32'hbb1c6dd3),
	.w5(32'h3b9436c2),
	.w6(32'h3be74d07),
	.w7(32'hb9bf1c86),
	.w8(32'hbb0b0eb3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba568dc),
	.w1(32'hbc56094a),
	.w2(32'h3a7df876),
	.w3(32'hbb42e693),
	.w4(32'h3bf946ad),
	.w5(32'h39cf45cf),
	.w6(32'hbc2555a9),
	.w7(32'hbb90a7f0),
	.w8(32'h3a2b703b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22845a),
	.w1(32'hbbe6df44),
	.w2(32'hbc08790d),
	.w3(32'hb78eb09d),
	.w4(32'h3b587d96),
	.w5(32'h3b8e47f5),
	.w6(32'h3aa09175),
	.w7(32'h3b19ca43),
	.w8(32'h3b60d1a5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cb8b8),
	.w1(32'h37e5478e),
	.w2(32'h392c90a0),
	.w3(32'h3b110367),
	.w4(32'hbba60857),
	.w5(32'hbbb5dd28),
	.w6(32'h3c1d89f0),
	.w7(32'h3a40ed99),
	.w8(32'hbbefa5f4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89cb4a),
	.w1(32'h3b1bd18f),
	.w2(32'h3baee1c6),
	.w3(32'hbc09e4c4),
	.w4(32'hbb7899e8),
	.w5(32'h3b841c6f),
	.w6(32'hbba10bbc),
	.w7(32'hb910939f),
	.w8(32'h3b2fcc58),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395759f2),
	.w1(32'hba86edce),
	.w2(32'h3aca4fa0),
	.w3(32'h3c13b216),
	.w4(32'h3bd488aa),
	.w5(32'h3b68e43e),
	.w6(32'hbb5c8094),
	.w7(32'h3b4df7d9),
	.w8(32'h3b91e269),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48fde6),
	.w1(32'hbb468f1d),
	.w2(32'hbbf0298c),
	.w3(32'h3b369f12),
	.w4(32'h3a081957),
	.w5(32'h3c453e5c),
	.w6(32'h3bcb7c41),
	.w7(32'h3b8648e5),
	.w8(32'h3b4bc925),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8583a),
	.w1(32'hbcead19a),
	.w2(32'hbbe9f978),
	.w3(32'h3cd923a6),
	.w4(32'h3cc13e93),
	.w5(32'hbc07d0d9),
	.w6(32'h3bb2c640),
	.w7(32'h3868b9e6),
	.w8(32'hbb91a198),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6a7e2),
	.w1(32'h3c3ffe37),
	.w2(32'h3ade1c04),
	.w3(32'hbc0bd2ef),
	.w4(32'hba468516),
	.w5(32'hbb1b9e79),
	.w6(32'h3c33b023),
	.w7(32'h3c376978),
	.w8(32'hbc0f7f2d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8db7a),
	.w1(32'h3c6c140b),
	.w2(32'h3ab3fda8),
	.w3(32'h38b33c29),
	.w4(32'h3b16c0cb),
	.w5(32'hbb964586),
	.w6(32'hba226245),
	.w7(32'h3a3fb7da),
	.w8(32'hbcb88529),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4729b0),
	.w1(32'hbc09af61),
	.w2(32'hbb516418),
	.w3(32'hbc4decf7),
	.w4(32'hbbe3ebdb),
	.w5(32'h3b07102f),
	.w6(32'h3c14d73a),
	.w7(32'hbb835d07),
	.w8(32'hbc04f3a7),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d928cb),
	.w1(32'hbc10d954),
	.w2(32'hbad24be2),
	.w3(32'hbbf4965c),
	.w4(32'hba4d0681),
	.w5(32'h3b8b17d5),
	.w6(32'hbc47ffde),
	.w7(32'hbb7fb7a4),
	.w8(32'hbb30d76e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d1088),
	.w1(32'hba743281),
	.w2(32'hbbcde407),
	.w3(32'h3b8bd203),
	.w4(32'h3c05cdac),
	.w5(32'h3ad42452),
	.w6(32'hbbe7057d),
	.w7(32'hbb7b4b56),
	.w8(32'h3a98ab61),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8fe2a),
	.w1(32'hba5ef944),
	.w2(32'hbb9f896c),
	.w3(32'hbb331b52),
	.w4(32'hbbb896ec),
	.w5(32'hba696cf4),
	.w6(32'h3c9ae52b),
	.w7(32'hbb4bc0ed),
	.w8(32'hbc07dbd8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2acbb),
	.w1(32'h3c71e1d2),
	.w2(32'hba478a4e),
	.w3(32'hbc103e9d),
	.w4(32'hbb88f308),
	.w5(32'hbcd5aec4),
	.w6(32'hbb0bec90),
	.w7(32'hbc0886ab),
	.w8(32'hbca3cdf7),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90cbe86),
	.w1(32'h3d0a2e2d),
	.w2(32'h3cc3360d),
	.w3(32'hbd3f7f1c),
	.w4(32'hbc1ae73b),
	.w5(32'h3b0d82aa),
	.w6(32'hbc7f9f57),
	.w7(32'h3baddc54),
	.w8(32'h3b16762c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb806ba),
	.w1(32'h3b902ccf),
	.w2(32'hbbb58898),
	.w3(32'hbafa34df),
	.w4(32'hbb06c83a),
	.w5(32'hbae9978b),
	.w6(32'h3b121b89),
	.w7(32'h3b082639),
	.w8(32'h3b90fec5),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5f85a),
	.w1(32'hbc5ab95a),
	.w2(32'hbc03ac4f),
	.w3(32'h3c8396ca),
	.w4(32'h392d7a3c),
	.w5(32'h3becfba2),
	.w6(32'hbb893fba),
	.w7(32'hbbf85bce),
	.w8(32'h3c3ae67c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b9b52),
	.w1(32'hbc25b994),
	.w2(32'hbada3a49),
	.w3(32'h3c5fcf42),
	.w4(32'h3c1fdb6a),
	.w5(32'hbbb99cee),
	.w6(32'hba8e1e0a),
	.w7(32'hbb6150df),
	.w8(32'hba8ff751),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7f281),
	.w1(32'h3c5abc2e),
	.w2(32'h3bf4df93),
	.w3(32'hbc100c64),
	.w4(32'hbc27ce67),
	.w5(32'hb8d06ed6),
	.w6(32'hbb39413c),
	.w7(32'hbbc0ab36),
	.w8(32'hbbfb342b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380a36a9),
	.w1(32'h3c865658),
	.w2(32'h3c151e5b),
	.w3(32'h39cbc9b9),
	.w4(32'h3b1b2d0e),
	.w5(32'h3b2a163b),
	.w6(32'hbbd9be6c),
	.w7(32'h3b936b08),
	.w8(32'hbaa9215a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb83e45),
	.w1(32'hbbdb8c82),
	.w2(32'hbc3dc2da),
	.w3(32'h3b4aac45),
	.w4(32'h3ad67c3a),
	.w5(32'hbc0834d3),
	.w6(32'hbbaa8940),
	.w7(32'h3a0d0f07),
	.w8(32'hbb8b36bf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3887d4e7),
	.w1(32'h3c6e162d),
	.w2(32'hb85fe28e),
	.w3(32'hbc61129a),
	.w4(32'hbb67af0a),
	.w5(32'hbb42bc88),
	.w6(32'h39e65620),
	.w7(32'h3b59bbfc),
	.w8(32'hbbb1f3e2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c071513),
	.w1(32'h3c3e58f6),
	.w2(32'h3c896f14),
	.w3(32'hbb0c8cb5),
	.w4(32'h39b031cd),
	.w5(32'hbbdc9c68),
	.w6(32'hbafbcfde),
	.w7(32'h3b0b67fe),
	.w8(32'hb92ef5fa),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59ff01),
	.w1(32'hbc0ec77f),
	.w2(32'h3a0d5ad1),
	.w3(32'hba3aeab6),
	.w4(32'hbb212849),
	.w5(32'h3c777493),
	.w6(32'h3c87b4a6),
	.w7(32'h3a39cfd6),
	.w8(32'h3a391449),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde3a44),
	.w1(32'hbccf279d),
	.w2(32'hbcdc7e7b),
	.w3(32'h3d11232e),
	.w4(32'h3c15e82e),
	.w5(32'h3c0eb906),
	.w6(32'hbaab69b8),
	.w7(32'hbc9ba3c2),
	.w8(32'h3c197116),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49d46a),
	.w1(32'hbc8fab17),
	.w2(32'hbc32341c),
	.w3(32'h3cbf6d98),
	.w4(32'h3bd86a9b),
	.w5(32'hbcbb5edb),
	.w6(32'h3c0303de),
	.w7(32'h3be8666b),
	.w8(32'hbc817497),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96884e),
	.w1(32'h3cff5400),
	.w2(32'h3c6d86b8),
	.w3(32'hbd011ef3),
	.w4(32'hbca0a240),
	.w5(32'hbb9883eb),
	.w6(32'hbc2c2dc8),
	.w7(32'hbbb13f45),
	.w8(32'h3c1ebda3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0625a5),
	.w1(32'hbc0c6a91),
	.w2(32'h3c3df94b),
	.w3(32'h3c40bbe9),
	.w4(32'hbb8b86ba),
	.w5(32'h3c0b19e8),
	.w6(32'hbbe59e8a),
	.w7(32'hbb6cb8bf),
	.w8(32'hbbd13a8a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1de305),
	.w1(32'hbbf46a3a),
	.w2(32'hbbeab832),
	.w3(32'h3c7a49d4),
	.w4(32'h3b4f0435),
	.w5(32'h3c0646e8),
	.w6(32'hbc26f1fc),
	.w7(32'hbc2248bb),
	.w8(32'hbc01fa8d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafd1fe),
	.w1(32'h390acb94),
	.w2(32'hbbbea3df),
	.w3(32'hbbbb15c2),
	.w4(32'hbc2866cb),
	.w5(32'h3b195977),
	.w6(32'h3bb10636),
	.w7(32'hbb49afb8),
	.w8(32'hbbd288b6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe48fcf),
	.w1(32'h3c7f0a41),
	.w2(32'hba5aaafd),
	.w3(32'hbc657307),
	.w4(32'hbaa34b32),
	.w5(32'h3bbb1dbc),
	.w6(32'h3ae48bcb),
	.w7(32'h3bad1f4b),
	.w8(32'h390cec0c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49184d),
	.w1(32'h3affdcba),
	.w2(32'h3bbcf617),
	.w3(32'hbba8b37c),
	.w4(32'hbc00e9f8),
	.w5(32'h3bd25ee8),
	.w6(32'h3c85fa31),
	.w7(32'h3b261ed2),
	.w8(32'hbb505ec1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c006af8),
	.w1(32'h3b82290e),
	.w2(32'h3b00f091),
	.w3(32'h3b826650),
	.w4(32'h39cc6836),
	.w5(32'h3b45f448),
	.w6(32'h3b3550a1),
	.w7(32'h3c0d83b4),
	.w8(32'hbbc50ac2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba836baf),
	.w1(32'hbaf2da4a),
	.w2(32'hbbc35454),
	.w3(32'h3bc94713),
	.w4(32'h3b941c31),
	.w5(32'hbb627ed7),
	.w6(32'hbc0ece12),
	.w7(32'hbc16f5a5),
	.w8(32'hbc125022),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956b3ec),
	.w1(32'hba9a35b6),
	.w2(32'h3b8b0c60),
	.w3(32'hbbfe6e0e),
	.w4(32'hbc17489f),
	.w5(32'hbbe0f06e),
	.w6(32'h3bd5aea7),
	.w7(32'hbbff98b5),
	.w8(32'hbbba4707),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e1b01),
	.w1(32'h3c1af323),
	.w2(32'h3bd8b690),
	.w3(32'hbc246a1e),
	.w4(32'hbc00cc83),
	.w5(32'hbb43a37e),
	.w6(32'hbb82bcd1),
	.w7(32'h3bbe509d),
	.w8(32'hbbe71950),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac81915),
	.w1(32'h3cb27fca),
	.w2(32'h3b8e0118),
	.w3(32'hbca9598e),
	.w4(32'hbb803452),
	.w5(32'hbc52fe65),
	.w6(32'hba0876f9),
	.w7(32'h3bc5f1e8),
	.w8(32'hbc59a244),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe4401),
	.w1(32'h3cac0a74),
	.w2(32'h3bf2cdf4),
	.w3(32'hbc2253e6),
	.w4(32'hbb24054f),
	.w5(32'h3ca2e93a),
	.w6(32'hbaa9ed04),
	.w7(32'h3bd1f157),
	.w8(32'hbb046fbb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc27bb9),
	.w1(32'hbad88573),
	.w2(32'hbb452bde),
	.w3(32'h3bdc0824),
	.w4(32'hbaccb740),
	.w5(32'h3bbd0fdd),
	.w6(32'hbc1e7347),
	.w7(32'h3b439173),
	.w8(32'hba4db45e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f0b8c),
	.w1(32'hb953e69e),
	.w2(32'h3bbe5f63),
	.w3(32'h3c016251),
	.w4(32'h3b302ce4),
	.w5(32'hb9ea1dcc),
	.w6(32'hbc1d5c24),
	.w7(32'h3b876cab),
	.w8(32'hbc38772a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e78d1),
	.w1(32'hbc6bddbb),
	.w2(32'hbb25a840),
	.w3(32'h3ba7cd5d),
	.w4(32'h3bf0759f),
	.w5(32'hbb888380),
	.w6(32'hbc78488e),
	.w7(32'hbbe9aa15),
	.w8(32'h3b8c6b83),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af260f0),
	.w1(32'h3bd589b9),
	.w2(32'h3bf5797d),
	.w3(32'hba5338bd),
	.w4(32'hba6289d8),
	.w5(32'h3c040aaa),
	.w6(32'hba91ccde),
	.w7(32'hb9df71f5),
	.w8(32'h3954a0d4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73e7be),
	.w1(32'hbc7636f2),
	.w2(32'hbc38dc6b),
	.w3(32'h3c1a26ae),
	.w4(32'hbbc3ceeb),
	.w5(32'h3be5f2e7),
	.w6(32'hbc434c3a),
	.w7(32'hbc3b1f19),
	.w8(32'hb9296ca5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5562e8),
	.w1(32'hbcdd17fa),
	.w2(32'hbcaaa141),
	.w3(32'h3ce1b11d),
	.w4(32'h3c235575),
	.w5(32'hbb93a782),
	.w6(32'h3ac4a270),
	.w7(32'hbab4c70b),
	.w8(32'hbb89afff),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f738a),
	.w1(32'hbacfefe7),
	.w2(32'hbb869560),
	.w3(32'hbbdb969b),
	.w4(32'hba385242),
	.w5(32'hbaa3feeb),
	.w6(32'h3c207312),
	.w7(32'h3bd1e986),
	.w8(32'hbaf95fba),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e040e),
	.w1(32'h3a921df3),
	.w2(32'h3ad3737b),
	.w3(32'hb9a15ea6),
	.w4(32'h3a3afd28),
	.w5(32'hbb618e54),
	.w6(32'h381af325),
	.w7(32'h38c157f4),
	.w8(32'hbb8781ca),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cc333),
	.w1(32'hbb0966d5),
	.w2(32'hbb55572e),
	.w3(32'h3aaf50d9),
	.w4(32'hbb370979),
	.w5(32'h3b812c82),
	.w6(32'hba821ab0),
	.w7(32'hbb78ed06),
	.w8(32'h3b2c8353),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3850e59b),
	.w1(32'h3a8f7994),
	.w2(32'h3b8f5bb7),
	.w3(32'h3b236bf7),
	.w4(32'h3b98a016),
	.w5(32'h39a146b5),
	.w6(32'h3bac0256),
	.w7(32'h3be4a87f),
	.w8(32'hbc1b8713),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9355083),
	.w1(32'h39b86094),
	.w2(32'h3b374996),
	.w3(32'hbb41cbc2),
	.w4(32'h391e3561),
	.w5(32'h380d161f),
	.w6(32'hbbc83cd7),
	.w7(32'hbc2d5c96),
	.w8(32'h3b3609a9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d66a1),
	.w1(32'h3aaedda6),
	.w2(32'h3b144f9d),
	.w3(32'h3b46c3f8),
	.w4(32'h3b5e6e24),
	.w5(32'hbb814d90),
	.w6(32'h3b4f730a),
	.w7(32'h3aea736f),
	.w8(32'hbb81a818),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74b81c),
	.w1(32'hbb9edef1),
	.w2(32'hbb3ce0d5),
	.w3(32'hba95f1d6),
	.w4(32'hbb1ff61a),
	.w5(32'h3ab36bea),
	.w6(32'hbb4beb48),
	.w7(32'hbb5c066f),
	.w8(32'h3931a92d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbf986),
	.w1(32'hbac25764),
	.w2(32'h3b0facea),
	.w3(32'hb9c70415),
	.w4(32'h3a8d85bb),
	.w5(32'hbb1c379b),
	.w6(32'h3adfd9b5),
	.w7(32'h3bad4d07),
	.w8(32'h3ae6efdc),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bef3f),
	.w1(32'hb9b07366),
	.w2(32'h39f2cb75),
	.w3(32'hba1d4090),
	.w4(32'hbb873db5),
	.w5(32'hba879b02),
	.w6(32'h3add69b8),
	.w7(32'h3aa271b7),
	.w8(32'hbb78dfaf),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb921aae),
	.w1(32'h39b14e1e),
	.w2(32'hbb20b975),
	.w3(32'h3ac797f8),
	.w4(32'hb8eaa919),
	.w5(32'h3b3809fe),
	.w6(32'h388e1adc),
	.w7(32'hbb3301f9),
	.w8(32'h3afdbf72),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17c1c9),
	.w1(32'h3a8af0a0),
	.w2(32'h3a165adb),
	.w3(32'h3b411c64),
	.w4(32'h3758480f),
	.w5(32'hb8f89ea4),
	.w6(32'h3b19c2ee),
	.w7(32'h3988bec0),
	.w8(32'hb9bdb158),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f635c),
	.w1(32'h3aad9309),
	.w2(32'hba28f4c2),
	.w3(32'h3ad1bcaf),
	.w4(32'h3b44d0fc),
	.w5(32'hbab6e97c),
	.w6(32'h3b7312c0),
	.w7(32'h3add9832),
	.w8(32'h38a8c4b6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b296a5d),
	.w1(32'hb9e1a3ed),
	.w2(32'hbb873f54),
	.w3(32'hbaf05064),
	.w4(32'hbaa159e4),
	.w5(32'hba8e8090),
	.w6(32'hbafc937d),
	.w7(32'hbb6e5c93),
	.w8(32'hba93942d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd7004),
	.w1(32'hbacc05dc),
	.w2(32'h3aad812c),
	.w3(32'hb9afeb60),
	.w4(32'hb96097aa),
	.w5(32'hbb9148ac),
	.w6(32'h3aacf0dc),
	.w7(32'h3ae00d49),
	.w8(32'hba242088),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba927c00),
	.w1(32'hbb828909),
	.w2(32'hbaf126c6),
	.w3(32'hbb5039e6),
	.w4(32'hbb70f94e),
	.w5(32'hbb45a136),
	.w6(32'hbb8775b7),
	.w7(32'hbbc48342),
	.w8(32'h3ac68076),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b515fe7),
	.w1(32'h3b9bd297),
	.w2(32'h3ba2e01c),
	.w3(32'hbb05816c),
	.w4(32'hba1b73df),
	.w5(32'hbb3359a9),
	.w6(32'h3aa51c23),
	.w7(32'hba894a53),
	.w8(32'h3be3e507),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f25dc),
	.w1(32'hbb6e080b),
	.w2(32'hbaf45220),
	.w3(32'hbbc53ddc),
	.w4(32'hbb7bab9a),
	.w5(32'hbb13328d),
	.w6(32'h3bb56808),
	.w7(32'h3c1354f9),
	.w8(32'hbaf8e930),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7392c1),
	.w1(32'hba690a26),
	.w2(32'hbb6ee908),
	.w3(32'hbaf5a886),
	.w4(32'hbbc3203f),
	.w5(32'hbb1cf8e9),
	.w6(32'hbb46de9f),
	.w7(32'hbb4137e8),
	.w8(32'hba5287e2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d84c0),
	.w1(32'hba3693b3),
	.w2(32'h39ab8a9a),
	.w3(32'hbb0679a1),
	.w4(32'hba92a959),
	.w5(32'hbacb50b9),
	.w6(32'hbbd6e6ac),
	.w7(32'hbc08627f),
	.w8(32'hb9ce5cc4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd8185),
	.w1(32'hba1ddfc0),
	.w2(32'h3a5e9126),
	.w3(32'hbb257678),
	.w4(32'hbb263334),
	.w5(32'hb9f4d694),
	.w6(32'hbac90803),
	.w7(32'hbaa12540),
	.w8(32'hbb438220),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85d71b),
	.w1(32'hbb29aba2),
	.w2(32'hbac28c85),
	.w3(32'hb9c8d6cc),
	.w4(32'hba40ba77),
	.w5(32'h3b02a92c),
	.w6(32'h3ab6c082),
	.w7(32'hb991a354),
	.w8(32'h3c05335f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba25527),
	.w1(32'h3b557048),
	.w2(32'h3b032d0a),
	.w3(32'h3ae2d840),
	.w4(32'h380f6726),
	.w5(32'hbaf158ca),
	.w6(32'h3c32e773),
	.w7(32'h3c0cabe0),
	.w8(32'hbb404ca4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c7c4a),
	.w1(32'h3a57cd80),
	.w2(32'hbb0743cb),
	.w3(32'hbb6f9cbf),
	.w4(32'hb96bb75a),
	.w5(32'hbb4a3f2b),
	.w6(32'hbada0a49),
	.w7(32'hbb1adbdc),
	.w8(32'h3ad3ce0b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c218c),
	.w1(32'hbb320817),
	.w2(32'hbb8a4450),
	.w3(32'hbb62c715),
	.w4(32'hba4416b0),
	.w5(32'hbafc6d8b),
	.w6(32'h3a838b2f),
	.w7(32'hbae74321),
	.w8(32'hb9de32d3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53f9b9),
	.w1(32'hbb76fdf0),
	.w2(32'hbadad493),
	.w3(32'hb92fb127),
	.w4(32'hba941c10),
	.w5(32'hbb8fdaa7),
	.w6(32'hba6a9adb),
	.w7(32'hbaf14cc8),
	.w8(32'hbaabf70f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91a996),
	.w1(32'h3ba9b19c),
	.w2(32'h3a3f891c),
	.w3(32'hbb1f0a0b),
	.w4(32'hbb19b62a),
	.w5(32'hba1258aa),
	.w6(32'hbacdcb9d),
	.w7(32'hbaefeebd),
	.w8(32'hb9b207ac),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb5611),
	.w1(32'h39c478f9),
	.w2(32'hbaf98a3e),
	.w3(32'hbab488d7),
	.w4(32'h37c5335a),
	.w5(32'hbab2d8f6),
	.w6(32'h3a8661d9),
	.w7(32'h3a6ac9d5),
	.w8(32'hbb6c5c40),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d2265),
	.w1(32'h3a9663be),
	.w2(32'hb9cd7421),
	.w3(32'hba704ee7),
	.w4(32'hba9ecaa8),
	.w5(32'h3b395bf2),
	.w6(32'hbb71ae85),
	.w7(32'hbb6f7929),
	.w8(32'hbafeda48),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb990a82),
	.w1(32'hbbc1fb44),
	.w2(32'hbb85573f),
	.w3(32'h3b054891),
	.w4(32'h3b08f5e1),
	.w5(32'hbb1477dd),
	.w6(32'hb9a6ed8d),
	.w7(32'h3a0ceb61),
	.w8(32'h3b7ae7c5),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdab96),
	.w1(32'h3b17d156),
	.w2(32'hb9d28418),
	.w3(32'hbb0d002e),
	.w4(32'hbaa2b1f7),
	.w5(32'hbb45ff52),
	.w6(32'hbaceaec4),
	.w7(32'hbab68c15),
	.w8(32'h39120e5b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97b3e8),
	.w1(32'h3b7991a7),
	.w2(32'h3b6faa68),
	.w3(32'hbb28c45c),
	.w4(32'hbae99a77),
	.w5(32'hba96a731),
	.w6(32'hbad9676d),
	.w7(32'h39d2a4c4),
	.w8(32'hbb918837),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule