module layer_10_featuremap_390(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab5b21),
	.w1(32'hbbd076af),
	.w2(32'hbc91211a),
	.w3(32'h3b7016c5),
	.w4(32'h3ba15b04),
	.w5(32'h3b4c0e41),
	.w6(32'h3c541655),
	.w7(32'h3c14b933),
	.w8(32'h3cc9b77c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65dda8),
	.w1(32'h3b2134b8),
	.w2(32'hbbe0d3f8),
	.w3(32'h3ab15e22),
	.w4(32'hbbd62aed),
	.w5(32'h3a530170),
	.w6(32'h3c7e670a),
	.w7(32'hbc05744a),
	.w8(32'hbb81d75c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bded872),
	.w1(32'hbae4a1ba),
	.w2(32'hbc183375),
	.w3(32'h3c0b07ca),
	.w4(32'h3a6b8c3f),
	.w5(32'h389b28ab),
	.w6(32'hbb3607a2),
	.w7(32'hba169864),
	.w8(32'h3be7e0ac),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83e796),
	.w1(32'hbbe6866e),
	.w2(32'hbb98e46d),
	.w3(32'h38910915),
	.w4(32'hbc0e9b76),
	.w5(32'h3c1e3e37),
	.w6(32'h39b983d2),
	.w7(32'hb9f88b9f),
	.w8(32'h3bbc73bd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9279f),
	.w1(32'h38c5d79e),
	.w2(32'h3bc24c9b),
	.w3(32'hbbe9a697),
	.w4(32'h3b071ea4),
	.w5(32'hbb6b7064),
	.w6(32'hba32a088),
	.w7(32'hb9636b72),
	.w8(32'hba910b15),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b6f4b),
	.w1(32'h3c068fcf),
	.w2(32'h3c293043),
	.w3(32'h3a317440),
	.w4(32'hbb9c1211),
	.w5(32'h3b9c1baa),
	.w6(32'h3af92bea),
	.w7(32'hbc3dff96),
	.w8(32'hba9e2684),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43fe2d),
	.w1(32'hbbce506a),
	.w2(32'hbba24c90),
	.w3(32'h3c1a1430),
	.w4(32'hbc484c90),
	.w5(32'h3c316d98),
	.w6(32'hbc4ea21a),
	.w7(32'h3b04fe54),
	.w8(32'h3b6c0fe5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d6feb),
	.w1(32'h3bd7720b),
	.w2(32'h3bf3dd35),
	.w3(32'h3ca36df7),
	.w4(32'h3c4e2d8c),
	.w5(32'hbbf1fadb),
	.w6(32'h3c5801f0),
	.w7(32'h3c513d0c),
	.w8(32'h3bd846b6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4d9a1),
	.w1(32'hbaf945dc),
	.w2(32'hbbcd3a77),
	.w3(32'hbbb008dd),
	.w4(32'hba4feeb2),
	.w5(32'h3af73dac),
	.w6(32'hba3f965e),
	.w7(32'hbba51471),
	.w8(32'hbac6de26),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a06d3),
	.w1(32'h3c0b6bf7),
	.w2(32'h3c240469),
	.w3(32'hbbcb4b45),
	.w4(32'hbb914819),
	.w5(32'hbb3ac42f),
	.w6(32'hb898d3df),
	.w7(32'hbb4d0baf),
	.w8(32'h3c22aaf2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ccff9),
	.w1(32'h3b523a02),
	.w2(32'h3b597527),
	.w3(32'hbc15e66b),
	.w4(32'hb90672e1),
	.w5(32'h3c20ac1f),
	.w6(32'h3be2e680),
	.w7(32'h3bc60716),
	.w8(32'h3b0b9502),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc0231),
	.w1(32'h3c73a040),
	.w2(32'h3cb451ed),
	.w3(32'hbaa88e14),
	.w4(32'h3ac0cf66),
	.w5(32'hbaf5694a),
	.w6(32'hbc099bab),
	.w7(32'hbc070c27),
	.w8(32'hbc53e1b4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a80b0),
	.w1(32'h3bba3c9f),
	.w2(32'h3c9f4ba6),
	.w3(32'hbbce8029),
	.w4(32'hba9c2d7b),
	.w5(32'h3ba31899),
	.w6(32'hbcc25d10),
	.w7(32'hbc42dc6b),
	.w8(32'hbc8e2d2e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa9091),
	.w1(32'h3ac4d53f),
	.w2(32'hbbd580ad),
	.w3(32'hbb3983c2),
	.w4(32'h3c17d487),
	.w5(32'h3b7871ff),
	.w6(32'hbc08408b),
	.w7(32'h3c1662d0),
	.w8(32'h3ad5b0e8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdf6bf),
	.w1(32'hbc1cf4fd),
	.w2(32'h3a746cea),
	.w3(32'hbc357e6c),
	.w4(32'hbc29d97c),
	.w5(32'h3b87e609),
	.w6(32'hba640c32),
	.w7(32'hbbbfb35f),
	.w8(32'hbca64dfc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26b0b2),
	.w1(32'hbb463166),
	.w2(32'h3b3427cd),
	.w3(32'hbbac4930),
	.w4(32'hbbd04e3e),
	.w5(32'hbc132d34),
	.w6(32'hbab5700d),
	.w7(32'h3adddb03),
	.w8(32'hbc1746b8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b002588),
	.w1(32'hbb93e95e),
	.w2(32'hbb4265ea),
	.w3(32'hbbef82c7),
	.w4(32'hbc12e5e0),
	.w5(32'h3b51e8f5),
	.w6(32'hbbc16127),
	.w7(32'hb9abd16d),
	.w8(32'hbba463b8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74159c2),
	.w1(32'h3975fb7d),
	.w2(32'hbbe11f11),
	.w3(32'h3c1737bc),
	.w4(32'h3c55c288),
	.w5(32'h3c072b08),
	.w6(32'h3c3f7965),
	.w7(32'h3cdb432e),
	.w8(32'h3d34bd73),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22e332),
	.w1(32'h3add4e81),
	.w2(32'h3c5a0eb9),
	.w3(32'h3bfcada6),
	.w4(32'hbb9a55cf),
	.w5(32'h3bc7dc16),
	.w6(32'h3cd87352),
	.w7(32'hbbb5fc02),
	.w8(32'hbc1406f6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8b338),
	.w1(32'hbad7811d),
	.w2(32'hba0d4b36),
	.w3(32'hbbd810dd),
	.w4(32'hb9b8032b),
	.w5(32'h3bf955a0),
	.w6(32'hbc5155d1),
	.w7(32'h3c172f83),
	.w8(32'hbbad7d5c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94be1b),
	.w1(32'h3ca650a8),
	.w2(32'h3c9b7016),
	.w3(32'hbb254f3c),
	.w4(32'h3c1b0a83),
	.w5(32'h3b8c26a2),
	.w6(32'hbb3f17ed),
	.w7(32'hbbdc1958),
	.w8(32'hbc8e99e1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd76a2f),
	.w1(32'h3b377e78),
	.w2(32'hbba4e5d1),
	.w3(32'hbbe89a27),
	.w4(32'h3c0ca6ad),
	.w5(32'hbb31b132),
	.w6(32'hbcc40a60),
	.w7(32'h3b813823),
	.w8(32'hbc71a528),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab1fd9),
	.w1(32'h3c5711c7),
	.w2(32'h3c8858e4),
	.w3(32'h3bc1c302),
	.w4(32'hbc0099b8),
	.w5(32'h3b8111f6),
	.w6(32'h3cc2c27d),
	.w7(32'h3b93efc2),
	.w8(32'hbbdb66d8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd86a29),
	.w1(32'h3ac05e7a),
	.w2(32'h3b7d2e96),
	.w3(32'hbb41883c),
	.w4(32'hbc805337),
	.w5(32'hbbd35c75),
	.w6(32'hbc63a571),
	.w7(32'h38f1ad3f),
	.w8(32'h3b49ecbd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16cbeb),
	.w1(32'hbba5e677),
	.w2(32'hbc15666a),
	.w3(32'hbbf862dd),
	.w4(32'hbbe0628f),
	.w5(32'hba377a64),
	.w6(32'hba7ca03f),
	.w7(32'hbc31aeeb),
	.w8(32'hba6caa9c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d4876),
	.w1(32'h3aede188),
	.w2(32'hbab2cf49),
	.w3(32'hba909dfe),
	.w4(32'h3af8f29b),
	.w5(32'hb9316f7d),
	.w6(32'hb91fb6bf),
	.w7(32'hbbc59f4d),
	.w8(32'hba920a1c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc258dcf),
	.w1(32'h3c4b6011),
	.w2(32'hbb4b4442),
	.w3(32'hbad12eac),
	.w4(32'hbb9b0c8c),
	.w5(32'hbc0d5147),
	.w6(32'h3a09b76d),
	.w7(32'hbb55cea7),
	.w8(32'hbb18d192),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28b093),
	.w1(32'hbb128e62),
	.w2(32'hbbfd0e3f),
	.w3(32'hbbcd44fc),
	.w4(32'hbbb2b1f1),
	.w5(32'h3b5ff62f),
	.w6(32'h3b19b96d),
	.w7(32'h3a7caf68),
	.w8(32'h3a2a5aab),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3506),
	.w1(32'h3c1b2d12),
	.w2(32'h3bb7683e),
	.w3(32'hbbe226cb),
	.w4(32'hbbad1e6d),
	.w5(32'hbc69e079),
	.w6(32'hbbbee97b),
	.w7(32'hbc4bdf2e),
	.w8(32'hbbcd47c9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08c0fa),
	.w1(32'h3c8831a7),
	.w2(32'h3ce7bc25),
	.w3(32'hbc75dc02),
	.w4(32'hbb33431e),
	.w5(32'hbb8c9fe6),
	.w6(32'hbca34e7f),
	.w7(32'hbc704f5f),
	.w8(32'hbcc36f1a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce62d2e),
	.w1(32'hbb8ab338),
	.w2(32'hbbc48646),
	.w3(32'h3b7d82ee),
	.w4(32'hbc29de6f),
	.w5(32'hbae13545),
	.w6(32'hbc784489),
	.w7(32'h3bfba92a),
	.w8(32'h3b762d44),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39855d48),
	.w1(32'hbbc0d8e6),
	.w2(32'h3b721916),
	.w3(32'h3c5fec67),
	.w4(32'hbab0e19f),
	.w5(32'hbb2d77d7),
	.w6(32'h3b6d3a99),
	.w7(32'hbbc6e836),
	.w8(32'hbbcdc057),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984d48d),
	.w1(32'hbb3b651f),
	.w2(32'hba60c09f),
	.w3(32'hbbbadcc7),
	.w4(32'hbb1cf7f4),
	.w5(32'h3b95b979),
	.w6(32'hbb87ff35),
	.w7(32'h3a2d2747),
	.w8(32'h3b993602),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc8bc5),
	.w1(32'h3b0a70f1),
	.w2(32'hbb4a9819),
	.w3(32'h3ac6ba99),
	.w4(32'hbc28227c),
	.w5(32'h3b9b8794),
	.w6(32'h3c11d5ff),
	.w7(32'hba25da2a),
	.w8(32'h3b2d1c6e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0beabd),
	.w1(32'h3bd14e22),
	.w2(32'h3ad7aa0c),
	.w3(32'h3bda460c),
	.w4(32'h3bb6e459),
	.w5(32'h39ee2fab),
	.w6(32'h39ddbde9),
	.w7(32'h3be80143),
	.w8(32'h39e9c278),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1306ae),
	.w1(32'hbc6c621c),
	.w2(32'hbc04879e),
	.w3(32'h3c029851),
	.w4(32'hbbb0b415),
	.w5(32'h3c005a56),
	.w6(32'hb8d6628e),
	.w7(32'h3be017ce),
	.w8(32'h3cb4be9f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf6bc7),
	.w1(32'hbc2f0d64),
	.w2(32'h3b979e7b),
	.w3(32'h3bf7307c),
	.w4(32'hbc0ce7ce),
	.w5(32'h3ae73d1a),
	.w6(32'h3bd9e0fe),
	.w7(32'h3b84020b),
	.w8(32'h3b456909),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6efd80),
	.w1(32'hbc1ea07d),
	.w2(32'h3a860063),
	.w3(32'hbad14c26),
	.w4(32'hbc7f15c4),
	.w5(32'hbb15e474),
	.w6(32'hbc5055e4),
	.w7(32'hbc78985e),
	.w8(32'hbc56a9b1),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c584c),
	.w1(32'hbc82d53d),
	.w2(32'hbcf8a504),
	.w3(32'hbbe16639),
	.w4(32'hbc08f5f4),
	.w5(32'h3b97dcdf),
	.w6(32'hbcb7a859),
	.w7(32'h3a8da0ca),
	.w8(32'h3cc6bda2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6b983),
	.w1(32'hbc1dee8e),
	.w2(32'hbc1d2bbc),
	.w3(32'hbb88f885),
	.w4(32'hbba5344a),
	.w5(32'h3be26285),
	.w6(32'h3baccd39),
	.w7(32'h3b2b01e6),
	.w8(32'h3bb580d3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf224a6),
	.w1(32'h3a19c02e),
	.w2(32'h3a502bdd),
	.w3(32'hbc016eee),
	.w4(32'hbbc48a8e),
	.w5(32'hbc1d9136),
	.w6(32'h39bfd835),
	.w7(32'hbbb28f5e),
	.w8(32'h3af1026a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d6a47),
	.w1(32'h3b2f0c4a),
	.w2(32'h3bbdd63d),
	.w3(32'hbbdecb60),
	.w4(32'hb812dd98),
	.w5(32'h3b33f32f),
	.w6(32'hbc26d56a),
	.w7(32'hbb3c3bdc),
	.w8(32'hbc2a9a3d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafe50a),
	.w1(32'h3b31a954),
	.w2(32'h3c13d482),
	.w3(32'hba66ac1b),
	.w4(32'hbb040454),
	.w5(32'h3accb25a),
	.w6(32'h38cf9688),
	.w7(32'hbb673a9b),
	.w8(32'hbbd74a8f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35f7ab),
	.w1(32'hbbe25e2d),
	.w2(32'hbcf57887),
	.w3(32'h39d3f5aa),
	.w4(32'hba9e548c),
	.w5(32'h3c36d142),
	.w6(32'h3c2a72f6),
	.w7(32'h3c6414d0),
	.w8(32'h3d1f4067),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a0dd1),
	.w1(32'hbae3c64b),
	.w2(32'h3bb966ab),
	.w3(32'hb814a356),
	.w4(32'hbbd5fcb9),
	.w5(32'hbb975ecc),
	.w6(32'h3bee7e12),
	.w7(32'hbb9ebe42),
	.w8(32'hbb2d246a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be434b6),
	.w1(32'hba8a3698),
	.w2(32'hbb89a2c0),
	.w3(32'hbbc2fe0a),
	.w4(32'hbbc25ac0),
	.w5(32'hbc61ae15),
	.w6(32'h3b827626),
	.w7(32'h3a104298),
	.w8(32'hbacbe1d7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf0a9b),
	.w1(32'h3b678070),
	.w2(32'hbadab148),
	.w3(32'hbc0c97e4),
	.w4(32'hb973b150),
	.w5(32'h39e57a46),
	.w6(32'hbbffdf46),
	.w7(32'h3b5ae2cc),
	.w8(32'hbba68793),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d9917),
	.w1(32'h3c6f0cbb),
	.w2(32'h3c25a47c),
	.w3(32'h3ba0d88c),
	.w4(32'h3c1af58d),
	.w5(32'h3c9e5b62),
	.w6(32'h3bcf663b),
	.w7(32'h3c896177),
	.w8(32'h3cde6f61),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82e8000),
	.w1(32'hbb3869d8),
	.w2(32'h3bbd4ce8),
	.w3(32'h3a0deb90),
	.w4(32'hbbb421bd),
	.w5(32'hbbade79b),
	.w6(32'hbb85b5ee),
	.w7(32'hbbc0a38b),
	.w8(32'hba4f87c6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2abe5),
	.w1(32'hbb6c62d5),
	.w2(32'hbbbb29dd),
	.w3(32'hbad975f1),
	.w4(32'hbb323fec),
	.w5(32'hbbd11c9c),
	.w6(32'h3a1eef61),
	.w7(32'hbaf68a01),
	.w8(32'h3c40369e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb093e02),
	.w1(32'h3a257559),
	.w2(32'hbb6b9dcb),
	.w3(32'hbba22062),
	.w4(32'hbb2010a7),
	.w5(32'h3aea2e53),
	.w6(32'h3a3fc331),
	.w7(32'hbba85e0a),
	.w8(32'h3c062fb6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5bb5c),
	.w1(32'h3c68c805),
	.w2(32'hbc0790a6),
	.w3(32'hbb70e28c),
	.w4(32'h3ad0f4be),
	.w5(32'hba9432c2),
	.w6(32'hbc11736f),
	.w7(32'h3b89f379),
	.w8(32'h3ba332c2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe40f4e),
	.w1(32'hbaec11c5),
	.w2(32'h3b5c55ab),
	.w3(32'hbbc9f05d),
	.w4(32'hbb4672e2),
	.w5(32'h3b011337),
	.w6(32'hb9d9cd7e),
	.w7(32'hbb316884),
	.w8(32'h3bd1a9c9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dcb1c),
	.w1(32'h3c6ba331),
	.w2(32'h3c088e51),
	.w3(32'h3c3b007d),
	.w4(32'h3c8e4f30),
	.w5(32'hbb7c10f9),
	.w6(32'h3c94f711),
	.w7(32'h3c8b7f24),
	.w8(32'h3c34b54d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3256e),
	.w1(32'hba2e4777),
	.w2(32'hbba3d81f),
	.w3(32'hbc459cf4),
	.w4(32'hba8ac92c),
	.w5(32'h3af7eeef),
	.w6(32'hbb68329a),
	.w7(32'h3ba28b51),
	.w8(32'hb9930e76),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d4fbb),
	.w1(32'hbb51475a),
	.w2(32'hbba10c40),
	.w3(32'hb6183c66),
	.w4(32'hbb0c5e25),
	.w5(32'hbb3c5c31),
	.w6(32'h3bac493b),
	.w7(32'h3a054979),
	.w8(32'hbbb99145),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4472e3),
	.w1(32'hbad47cab),
	.w2(32'h3c233f22),
	.w3(32'h3a966636),
	.w4(32'h3acf6038),
	.w5(32'h3881a63c),
	.w6(32'hbb6e4a25),
	.w7(32'hbba8e1bf),
	.w8(32'hbc73bd90),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e4bff),
	.w1(32'hbab4abbf),
	.w2(32'hbbf02a64),
	.w3(32'hbafb4a18),
	.w4(32'h3bab076d),
	.w5(32'hbc8c2c30),
	.w6(32'hbc0d0fe0),
	.w7(32'hba2df963),
	.w8(32'hbc8abb0f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8edb9a),
	.w1(32'hbaae356d),
	.w2(32'hbb8a7450),
	.w3(32'hbb374cb0),
	.w4(32'hb9b12986),
	.w5(32'hba8e53d2),
	.w6(32'h3c313965),
	.w7(32'h3baf6b79),
	.w8(32'h3b91d369),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54feed),
	.w1(32'hbb9b565f),
	.w2(32'h3b86b3c5),
	.w3(32'hba8088f0),
	.w4(32'hbc830f73),
	.w5(32'hbbf2a30e),
	.w6(32'h3b5ded53),
	.w7(32'hbca92cc3),
	.w8(32'hbb91bddb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc733d5),
	.w1(32'hbaf438a6),
	.w2(32'hbba596c7),
	.w3(32'hb99d0f59),
	.w4(32'h3b784196),
	.w5(32'hbba8dc12),
	.w6(32'hbc142395),
	.w7(32'h3a11b338),
	.w8(32'h3c1c52ca),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fcef1),
	.w1(32'h3bd7d81f),
	.w2(32'h3b6a74e0),
	.w3(32'hbae2ea27),
	.w4(32'h3bb4440b),
	.w5(32'h3be2d660),
	.w6(32'h3c974dce),
	.w7(32'h3c2903da),
	.w8(32'h3b302261),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02cc3a),
	.w1(32'hbacfb629),
	.w2(32'hbc7dff4c),
	.w3(32'hbbaf7986),
	.w4(32'hbb1e0da9),
	.w5(32'h3ae01a84),
	.w6(32'h3a98f6fb),
	.w7(32'h3b8570f0),
	.w8(32'h3c35ee15),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44f9c3),
	.w1(32'h3bcdf82d),
	.w2(32'h3c104d0c),
	.w3(32'h3b21ce68),
	.w4(32'h3c2cf10b),
	.w5(32'hbc1a2174),
	.w6(32'h3b8e9ba8),
	.w7(32'hbb600672),
	.w8(32'hbc0cf2f9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b125fc4),
	.w1(32'h3c00d434),
	.w2(32'h3c2222c4),
	.w3(32'hbc147f17),
	.w4(32'h3c02681c),
	.w5(32'hba6baba4),
	.w6(32'hbbe919ac),
	.w7(32'h3c1a4284),
	.w8(32'h3bf1866c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b072c),
	.w1(32'hbb9113ed),
	.w2(32'hbbf88bbc),
	.w3(32'hbc08518a),
	.w4(32'hbaca0086),
	.w5(32'h3ad5fb38),
	.w6(32'h3a0786f4),
	.w7(32'h3bd7080d),
	.w8(32'h3c7da25d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe03133),
	.w1(32'h3ba8ce44),
	.w2(32'h3c0d409d),
	.w3(32'h3c151bec),
	.w4(32'h3c42769a),
	.w5(32'hbac6c3e4),
	.w6(32'h3c8765ab),
	.w7(32'h3a8550b8),
	.w8(32'hbb6f27f5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a924a75),
	.w1(32'hbba054af),
	.w2(32'hba70c08e),
	.w3(32'hbbeccd7c),
	.w4(32'hbb4ab8e3),
	.w5(32'h3b320d28),
	.w6(32'hbc093a0b),
	.w7(32'h393dc5cf),
	.w8(32'h3b89e0b1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30682a),
	.w1(32'h3bd0df89),
	.w2(32'hbc32337a),
	.w3(32'h3c54ca63),
	.w4(32'h3ba70e7a),
	.w5(32'h3bbed654),
	.w6(32'h3cb94c2b),
	.w7(32'h3c66b2a7),
	.w8(32'h3c9777d0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b571d9a),
	.w1(32'h3bf3a368),
	.w2(32'h3b1ee670),
	.w3(32'hbc431a94),
	.w4(32'h3c350342),
	.w5(32'h3b9f61c3),
	.w6(32'hbc0c8b52),
	.w7(32'h3badbe15),
	.w8(32'h3be62d5b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b693651),
	.w1(32'h3c1df24b),
	.w2(32'h3c4d1ae0),
	.w3(32'h3bde1e28),
	.w4(32'h3c14d6e4),
	.w5(32'h3a0e2460),
	.w6(32'h3b657c5e),
	.w7(32'hbb951792),
	.w8(32'hbc396459),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2434a),
	.w1(32'hbba9b537),
	.w2(32'hbb6eb955),
	.w3(32'hbc2b4fab),
	.w4(32'hbbec9db2),
	.w5(32'hbac31d96),
	.w6(32'hbc750574),
	.w7(32'hba6fb727),
	.w8(32'h3be44827),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd0218),
	.w1(32'h3c464e10),
	.w2(32'h3bc66848),
	.w3(32'h3a885f2a),
	.w4(32'h3cabcd28),
	.w5(32'h3c2c20f4),
	.w6(32'h3bc62f85),
	.w7(32'h3cc2b29b),
	.w8(32'h3bf2db45),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef64e3),
	.w1(32'h39651e81),
	.w2(32'hb81a392d),
	.w3(32'hbbb5abf7),
	.w4(32'h3a356134),
	.w5(32'h3a6073ed),
	.w6(32'hbc003d99),
	.w7(32'hbb119b85),
	.w8(32'hba088d04),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2b64e),
	.w1(32'h3c14b54c),
	.w2(32'h3c0965c4),
	.w3(32'hbae749f2),
	.w4(32'h3c0b8d36),
	.w5(32'h3c25683d),
	.w6(32'hbb512151),
	.w7(32'h3bc0c476),
	.w8(32'h3c114365),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad94725),
	.w1(32'h3c279004),
	.w2(32'h3c861ad9),
	.w3(32'h3b84d7f3),
	.w4(32'h3b3f4a60),
	.w5(32'hbb007a37),
	.w6(32'h3bf7eab5),
	.w7(32'h3a4c3a9a),
	.w8(32'hbabb6134),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb06b2e),
	.w1(32'h392278fb),
	.w2(32'h3be98bad),
	.w3(32'h3c7ccb8e),
	.w4(32'h3c40a595),
	.w5(32'h3c137304),
	.w6(32'h3bf0e1ee),
	.w7(32'h3bf8c561),
	.w8(32'h3bcaaa2e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07248c),
	.w1(32'hbbe99301),
	.w2(32'h3acc9450),
	.w3(32'hbbff3398),
	.w4(32'hb9f7e4ca),
	.w5(32'h3c09cf16),
	.w6(32'hbc2c81c5),
	.w7(32'h3b678e95),
	.w8(32'h3c04ccc6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf28af4),
	.w1(32'h3bb726b7),
	.w2(32'h3bc289a9),
	.w3(32'h3ac6432b),
	.w4(32'h3b07303c),
	.w5(32'h3a92a2af),
	.w6(32'hbaea0916),
	.w7(32'h3b40ae93),
	.w8(32'h3b7df9fb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ed3b),
	.w1(32'h3b8c95fa),
	.w2(32'h3bf01786),
	.w3(32'hbc76f6cd),
	.w4(32'h3b6eb05c),
	.w5(32'h3b1da734),
	.w6(32'hbc1a21d2),
	.w7(32'h3a3d7fad),
	.w8(32'h3b95c01b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c412bc1),
	.w1(32'hbc2a7be0),
	.w2(32'hbbacbe53),
	.w3(32'h3af4f3ef),
	.w4(32'hbbd24cc4),
	.w5(32'h3b30981f),
	.w6(32'h3b036bfc),
	.w7(32'hbbc0adae),
	.w8(32'hbbcbc061),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20af5b),
	.w1(32'h3b66a93a),
	.w2(32'h380c1f39),
	.w3(32'hbc0efcb4),
	.w4(32'h3bae607b),
	.w5(32'h3a7098c2),
	.w6(32'hbc48a671),
	.w7(32'h3ba5d2b9),
	.w8(32'h3b179a7b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46236c),
	.w1(32'h3a429612),
	.w2(32'h3b3f47ac),
	.w3(32'hbb043f40),
	.w4(32'hbb9977f2),
	.w5(32'h3997c796),
	.w6(32'hbb8ae617),
	.w7(32'hbba30d48),
	.w8(32'hbb984a2f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ad9751),
	.w1(32'h3c92722a),
	.w2(32'h3c621384),
	.w3(32'hba6e355b),
	.w4(32'h3bc5377b),
	.w5(32'hbb18b661),
	.w6(32'hb99bfcde),
	.w7(32'hbb8b6403),
	.w8(32'hbb93d017),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b593177),
	.w1(32'hbb994c34),
	.w2(32'hbc10efad),
	.w3(32'hbb46b62a),
	.w4(32'h3af3a221),
	.w5(32'hbbf68bbb),
	.w6(32'hbb07fecf),
	.w7(32'h3c4cd36b),
	.w8(32'h3a97f023),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eddf5),
	.w1(32'h3b568b32),
	.w2(32'hbbe35ddd),
	.w3(32'hbc13cd6a),
	.w4(32'hbbb9d5d6),
	.w5(32'hbc04d49a),
	.w6(32'hbb49bcbc),
	.w7(32'hbb9c10b0),
	.w8(32'h3b648c05),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dda90),
	.w1(32'hbb31ccf9),
	.w2(32'hbaea7aad),
	.w3(32'h3c1284de),
	.w4(32'hbbd8840c),
	.w5(32'hba9b250a),
	.w6(32'h3bb69760),
	.w7(32'hbb81ef09),
	.w8(32'hba1b2d3f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0570c5),
	.w1(32'hba306534),
	.w2(32'hbb35b080),
	.w3(32'hba5f4bc3),
	.w4(32'hb90b7d4c),
	.w5(32'h3b255833),
	.w6(32'hbaa6fcfc),
	.w7(32'h38e29bc6),
	.w8(32'h3bd7f2d9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942a653),
	.w1(32'h3c74984b),
	.w2(32'h3cae764c),
	.w3(32'h3b86ee08),
	.w4(32'h3beacbd3),
	.w5(32'h3b45c1bf),
	.w6(32'h3c176471),
	.w7(32'h3bd2e6ba),
	.w8(32'h3b394a97),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45b266),
	.w1(32'h3c5984f4),
	.w2(32'h3c23f3b5),
	.w3(32'h3c80c6a1),
	.w4(32'h3c538d02),
	.w5(32'h3b4011e8),
	.w6(32'h3c8f2cd6),
	.w7(32'h3c5d9b33),
	.w8(32'h3c023d68),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52a59f),
	.w1(32'h3afd3fad),
	.w2(32'hbbb2be56),
	.w3(32'h3bad0ab1),
	.w4(32'hbb021bf9),
	.w5(32'hbca86d1f),
	.w6(32'h3a899938),
	.w7(32'hbb299748),
	.w8(32'hbc55fb38),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a3f87),
	.w1(32'h3b5acf98),
	.w2(32'h3be5335e),
	.w3(32'h3a05115e),
	.w4(32'hbb3ac919),
	.w5(32'h3bcbc642),
	.w6(32'h3b22304b),
	.w7(32'h3a92056b),
	.w8(32'h3c25f4dd),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6cded),
	.w1(32'h3b7c31d9),
	.w2(32'h3b24e94a),
	.w3(32'hba62cac6),
	.w4(32'hbbc0fad9),
	.w5(32'hba5bc6a3),
	.w6(32'h3b850c5a),
	.w7(32'hbc1cc495),
	.w8(32'hbbebf363),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94e7ac),
	.w1(32'h3c6933f7),
	.w2(32'h3c24a3bc),
	.w3(32'hba502e25),
	.w4(32'h3aea4b7c),
	.w5(32'h3b463c1f),
	.w6(32'hbb2cc013),
	.w7(32'h3b63b924),
	.w8(32'h3ad0eec7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb60da7),
	.w1(32'h3c121122),
	.w2(32'h3ca02f4f),
	.w3(32'h3b2ad5a5),
	.w4(32'hbbb55910),
	.w5(32'hbb47bae6),
	.w6(32'hbb36f8b1),
	.w7(32'h3ad5c9a2),
	.w8(32'h3c1ec214),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96b15b),
	.w1(32'hbc02c850),
	.w2(32'hbb4d78bc),
	.w3(32'h3b3799ed),
	.w4(32'hbc222b98),
	.w5(32'h3a7659df),
	.w6(32'h3b864df8),
	.w7(32'hbc2c643e),
	.w8(32'hbbe98549),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab818d),
	.w1(32'hbb420eeb),
	.w2(32'hbb813016),
	.w3(32'h3be6ade2),
	.w4(32'hbb125da0),
	.w5(32'hbb248544),
	.w6(32'h3b54c0a8),
	.w7(32'hbaf99eb2),
	.w8(32'h3b4e4ed0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbee13a),
	.w1(32'hbbe4a116),
	.w2(32'h3c1bfb2c),
	.w3(32'h3b690b0f),
	.w4(32'hbc580076),
	.w5(32'h3b6ecbab),
	.w6(32'h3bc710fc),
	.w7(32'hbbd78fa4),
	.w8(32'h3c0445cb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca19fe6),
	.w1(32'h3b843045),
	.w2(32'h3bed9a9f),
	.w3(32'h3ca7d680),
	.w4(32'hbbf112f8),
	.w5(32'hbc0c470a),
	.w6(32'h3be0fb7d),
	.w7(32'hbc0e8d17),
	.w8(32'h3b7e73c7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b068bfe),
	.w1(32'h3c2b464c),
	.w2(32'h3cab2e4b),
	.w3(32'h3c42b72e),
	.w4(32'h3bbeefa8),
	.w5(32'h3bece814),
	.w6(32'h3baa73d8),
	.w7(32'h3c1a703a),
	.w8(32'h3b18bb90),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1029aa),
	.w1(32'h3c92e65e),
	.w2(32'h3c9eebbf),
	.w3(32'hbb8ff85e),
	.w4(32'hbc4012cd),
	.w5(32'hbbaf6dab),
	.w6(32'hbbcbc943),
	.w7(32'hbc63b9e5),
	.w8(32'hbc0cb68d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c164859),
	.w1(32'hbba4a381),
	.w2(32'hba8206f4),
	.w3(32'hbbc3c2b2),
	.w4(32'hbc3f38e6),
	.w5(32'h3b8173cf),
	.w6(32'hbbd1b5e6),
	.w7(32'hbbf2b7de),
	.w8(32'hbbcc478c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29e7a9),
	.w1(32'h3bb4ab79),
	.w2(32'h3c935672),
	.w3(32'h3bfa11c0),
	.w4(32'hbb48c810),
	.w5(32'h3c20c0bc),
	.w6(32'hb9a88195),
	.w7(32'hbb00a27b),
	.w8(32'h3b76eadc),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad69de7),
	.w1(32'h3ac59585),
	.w2(32'h3bbf8e8f),
	.w3(32'h3bfa89a3),
	.w4(32'h3bb4570c),
	.w5(32'h3bb7d668),
	.w6(32'h3bd6975f),
	.w7(32'hb9e950ed),
	.w8(32'h3b803b22),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68b3d8),
	.w1(32'h3c44439d),
	.w2(32'h3cc74168),
	.w3(32'h3c8fa4b8),
	.w4(32'h3a076d93),
	.w5(32'h3bd7c071),
	.w6(32'h3c4f8f26),
	.w7(32'h3ae69c96),
	.w8(32'h3c2a4fbe),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba179c14),
	.w1(32'hba641cfa),
	.w2(32'h3a127fc1),
	.w3(32'hbb50153a),
	.w4(32'hbbe1e90d),
	.w5(32'hb881bec4),
	.w6(32'hbb275a8f),
	.w7(32'hbba1a8d5),
	.w8(32'h3ac53966),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b099234),
	.w1(32'hbb6e3d22),
	.w2(32'hbbc0de76),
	.w3(32'h3adcab3a),
	.w4(32'hbaec0e16),
	.w5(32'hbab0f254),
	.w6(32'hbb609916),
	.w7(32'hbbaf5da1),
	.w8(32'hbb980f22),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73b233),
	.w1(32'hbb3d896f),
	.w2(32'hbb98617e),
	.w3(32'hbbb17e33),
	.w4(32'h3c3dac56),
	.w5(32'hbb4c49c8),
	.w6(32'hbb4ace87),
	.w7(32'h3c8c6f3d),
	.w8(32'h3bc5e8c4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55bfaa),
	.w1(32'h3b7619fc),
	.w2(32'h3c3fc41f),
	.w3(32'hbb641af5),
	.w4(32'hbc0742f8),
	.w5(32'h3afadba5),
	.w6(32'h3b4ea5e1),
	.w7(32'hbb9e8de3),
	.w8(32'hbb3dc6ab),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c598),
	.w1(32'hbb80988a),
	.w2(32'hba590950),
	.w3(32'hb8cbf8fb),
	.w4(32'hbc09fea2),
	.w5(32'hb984befb),
	.w6(32'hbbfdba8a),
	.w7(32'hbb9715a2),
	.w8(32'h3ad2f831),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11ae7f),
	.w1(32'h3baf09ff),
	.w2(32'hbc03a93b),
	.w3(32'h3b910e4a),
	.w4(32'hbbc39446),
	.w5(32'hbc6d9b6e),
	.w6(32'h3b51f006),
	.w7(32'h3bd8d523),
	.w8(32'h3b9c710d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb708f282),
	.w1(32'hba29e012),
	.w2(32'h3b362b96),
	.w3(32'hbb1a27e0),
	.w4(32'hbb8f7f69),
	.w5(32'hbb2d6de0),
	.w6(32'h3c87c012),
	.w7(32'hba118e2c),
	.w8(32'h3955297c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8af35),
	.w1(32'hbbb784ad),
	.w2(32'hbb84e96f),
	.w3(32'h3c32efcc),
	.w4(32'hb864b584),
	.w5(32'hbaa94113),
	.w6(32'hbabca4b2),
	.w7(32'hbb31d8cc),
	.w8(32'hbc087eae),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8beb6),
	.w1(32'h3b88e0bd),
	.w2(32'h399be9a5),
	.w3(32'h3a97090b),
	.w4(32'h3b445c03),
	.w5(32'h3b6cd9ac),
	.w6(32'h3b6a0364),
	.w7(32'h3a8d6c94),
	.w8(32'h3c4a3766),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba80e10),
	.w1(32'hb9f4d3d4),
	.w2(32'hbbd9e5af),
	.w3(32'h3b46ef86),
	.w4(32'hbc1ce96d),
	.w5(32'hbbd9c244),
	.w6(32'h3beff737),
	.w7(32'hbb9c3172),
	.w8(32'hbbc80e34),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb07311),
	.w1(32'h3be68e7a),
	.w2(32'h3be02abf),
	.w3(32'hbbe8527f),
	.w4(32'h3c8e843b),
	.w5(32'h3c281639),
	.w6(32'hbbc3e1e5),
	.w7(32'h3bef7476),
	.w8(32'h3a8f2413),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3398f),
	.w1(32'h3ac2916a),
	.w2(32'hb9987790),
	.w3(32'h3b0c50c3),
	.w4(32'hbb5f1415),
	.w5(32'hbb8ec9f7),
	.w6(32'hbbb12de9),
	.w7(32'h3a39c23b),
	.w8(32'hbb096527),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f4c08),
	.w1(32'h3b8e327c),
	.w2(32'hbafa312e),
	.w3(32'hba4fa098),
	.w4(32'hbc234ada),
	.w5(32'hbc08a1ca),
	.w6(32'h3a14cad1),
	.w7(32'hbbddce3c),
	.w8(32'hbc0fc1ec),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc93307),
	.w1(32'hbb837f8f),
	.w2(32'hbb4e4097),
	.w3(32'h3a7b3628),
	.w4(32'h3ac3d7d4),
	.w5(32'h3b9b53fb),
	.w6(32'hbc234187),
	.w7(32'hbb56e1ff),
	.w8(32'hba9cfd76),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab3529),
	.w1(32'hb892ce4d),
	.w2(32'h3b75f2ff),
	.w3(32'h399f8ebf),
	.w4(32'hbbfd1b86),
	.w5(32'hbba187e4),
	.w6(32'h3ab87ae3),
	.w7(32'hbb4982fe),
	.w8(32'h38e2be8b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c162345),
	.w1(32'h3bf0ecb6),
	.w2(32'h3c3c6e91),
	.w3(32'h3c2fa564),
	.w4(32'h3c84a23d),
	.w5(32'h3c8ee060),
	.w6(32'h3c11bbc7),
	.w7(32'h3c00fc80),
	.w8(32'h3c078d63),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afaa6a2),
	.w1(32'h3bbe6950),
	.w2(32'h3c8542fe),
	.w3(32'h3bbab22b),
	.w4(32'h3c0a674c),
	.w5(32'h3b44c4c1),
	.w6(32'h3accdd8c),
	.w7(32'h3b2a8f30),
	.w8(32'h3a854ed7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c345294),
	.w1(32'h3996b753),
	.w2(32'hba9a113b),
	.w3(32'h3b3d81ce),
	.w4(32'h3a8c75a1),
	.w5(32'h3b5987f2),
	.w6(32'hbb978c43),
	.w7(32'hb9cd6c08),
	.w8(32'hbac26351),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bb504),
	.w1(32'hb9e25cc6),
	.w2(32'h3acc387c),
	.w3(32'h3b24be70),
	.w4(32'hbb722c82),
	.w5(32'hb9c9a2fe),
	.w6(32'h3b1f303d),
	.w7(32'hbb4ef851),
	.w8(32'hbba98dcd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89fe876),
	.w1(32'h3b22ec68),
	.w2(32'h3bcb352f),
	.w3(32'hbb976657),
	.w4(32'h3acab772),
	.w5(32'h3be84c68),
	.w6(32'hbbfff71d),
	.w7(32'h3b3b8b3f),
	.w8(32'h3a40888e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc85d79),
	.w1(32'h3b7ed349),
	.w2(32'hba8258a5),
	.w3(32'h3bd4315f),
	.w4(32'h3abdaeef),
	.w5(32'h3bd14499),
	.w6(32'h39321bc6),
	.w7(32'hbb05b5ae),
	.w8(32'h3be63854),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5d55f),
	.w1(32'hbba117a6),
	.w2(32'hbb3db59e),
	.w3(32'h3a2238c8),
	.w4(32'hbb7f38a5),
	.w5(32'h3b024931),
	.w6(32'h3a4ae057),
	.w7(32'hbb95d2b7),
	.w8(32'hba40a8c3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25d847),
	.w1(32'h3c0e9b60),
	.w2(32'h3b8ae1fa),
	.w3(32'hbc0728d3),
	.w4(32'h3b23b570),
	.w5(32'h3af52b49),
	.w6(32'hbc19f6d0),
	.w7(32'hbab30944),
	.w8(32'h3ae0d125),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8188aa),
	.w1(32'h3ad3bb20),
	.w2(32'h3bfa7bdd),
	.w3(32'hbbbd65b5),
	.w4(32'hbbce5496),
	.w5(32'hb8bde341),
	.w6(32'h3a0b5d62),
	.w7(32'hbb2eb1c1),
	.w8(32'h39ac7fdf),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0cc4),
	.w1(32'h3b381b5b),
	.w2(32'h3a163953),
	.w3(32'hba0fb259),
	.w4(32'hbb0fef9f),
	.w5(32'hbb8e798e),
	.w6(32'hba09b3b6),
	.w7(32'hba80a536),
	.w8(32'h38985684),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41dc63),
	.w1(32'hba8ffb95),
	.w2(32'hbbf50c92),
	.w3(32'h3c2498b1),
	.w4(32'h3b154f63),
	.w5(32'hba4e80cc),
	.w6(32'h3c14d782),
	.w7(32'h38546251),
	.w8(32'h3aac7213),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e839ba),
	.w1(32'h3b491067),
	.w2(32'h3aa3ce27),
	.w3(32'h3bcf0b43),
	.w4(32'hbad0c5c7),
	.w5(32'h3a8a12d5),
	.w6(32'h3b91b4eb),
	.w7(32'h39c9ac4a),
	.w8(32'h3bcedab2),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae236e2),
	.w1(32'h3b11afc0),
	.w2(32'h3c253d1f),
	.w3(32'h3b8ce470),
	.w4(32'h380512f5),
	.w5(32'h3b956e69),
	.w6(32'h3b213278),
	.w7(32'hbaf15553),
	.w8(32'h3a899e20),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e0772),
	.w1(32'hbb1b49a3),
	.w2(32'hbb61c1c6),
	.w3(32'h3be6ac98),
	.w4(32'hbbfc6465),
	.w5(32'hbb6684a8),
	.w6(32'h3a78c013),
	.w7(32'hbb8cb0c9),
	.w8(32'hbb804b44),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1370fc),
	.w1(32'h3bc036fd),
	.w2(32'h3be532f7),
	.w3(32'h3c5b918d),
	.w4(32'hb8345764),
	.w5(32'h3759e97d),
	.w6(32'h3beb7403),
	.w7(32'h3af0dcac),
	.w8(32'h3bb0fb9a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb598d64),
	.w1(32'hbb864860),
	.w2(32'hbbfe29f6),
	.w3(32'hbbe2a46f),
	.w4(32'hbb9481e5),
	.w5(32'h39170ca7),
	.w6(32'hbc060022),
	.w7(32'h3a84cf48),
	.w8(32'hbb0627b6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb243876),
	.w1(32'h3aad60be),
	.w2(32'h3a9ed8a6),
	.w3(32'h3b402b04),
	.w4(32'hbb5611a1),
	.w5(32'hbbb04d13),
	.w6(32'h3aa655c5),
	.w7(32'h3af5adb2),
	.w8(32'h3a37c438),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad9a6f),
	.w1(32'h3cd00915),
	.w2(32'h3d0a8647),
	.w3(32'h3b436e2c),
	.w4(32'h3c5a68aa),
	.w5(32'h3c0992ea),
	.w6(32'h3b2057a8),
	.w7(32'h3b77b916),
	.w8(32'h3b117a77),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c402720),
	.w1(32'hbacee14b),
	.w2(32'h3b329619),
	.w3(32'hbb4b925e),
	.w4(32'hbc28ee1f),
	.w5(32'hbbeb242c),
	.w6(32'hbbd94883),
	.w7(32'hbb28f1c0),
	.w8(32'hba667047),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3c40f),
	.w1(32'h3a4f4a12),
	.w2(32'h3ac4b075),
	.w3(32'hbb28b9d2),
	.w4(32'h39807567),
	.w5(32'h3b644af8),
	.w6(32'h3a4c02dd),
	.w7(32'h3b27c075),
	.w8(32'h3b1b961f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a858fd9),
	.w1(32'h3b4146e8),
	.w2(32'h3b80a2bb),
	.w3(32'h3a28015f),
	.w4(32'h3c12c8f9),
	.w5(32'h3c81ffeb),
	.w6(32'hbb4132f1),
	.w7(32'h3a61fac8),
	.w8(32'h3bf7bfb0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9964d4),
	.w1(32'hbc03d81c),
	.w2(32'h3b1b0499),
	.w3(32'h3a532208),
	.w4(32'hbc681498),
	.w5(32'hbb6d95ac),
	.w6(32'hbb6857d2),
	.w7(32'h3b6a36e4),
	.w8(32'h3aaf75d6),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2c835),
	.w1(32'hbb585a5a),
	.w2(32'hb9a0a72c),
	.w3(32'hbb45251d),
	.w4(32'h3b8a9304),
	.w5(32'hbb2cc73c),
	.w6(32'h3aaf1545),
	.w7(32'h3bf27d98),
	.w8(32'hbbecc0d2),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b187581),
	.w1(32'hbbcd75c8),
	.w2(32'hbb7d276d),
	.w3(32'h3b8bc85f),
	.w4(32'h3be974ca),
	.w5(32'h3c0568c6),
	.w6(32'h396c596a),
	.w7(32'h3b837c18),
	.w8(32'h3aa6683b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b26e),
	.w1(32'hbc1b959d),
	.w2(32'hbc301cd4),
	.w3(32'h3b179f2f),
	.w4(32'h3a5f2a99),
	.w5(32'hbc314772),
	.w6(32'h3a3819b3),
	.w7(32'h3c22596e),
	.w8(32'h3a98bedb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f59d),
	.w1(32'h3b296d1c),
	.w2(32'hbb0ab22b),
	.w3(32'hbc05bcb1),
	.w4(32'hba63aca6),
	.w5(32'hbbf8411a),
	.w6(32'hbb2f60bb),
	.w7(32'h3906e323),
	.w8(32'hbbf04208),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6d2ea),
	.w1(32'hbb228832),
	.w2(32'h3bf109db),
	.w3(32'hbc8cfe10),
	.w4(32'h3ac2599a),
	.w5(32'h3bc67c58),
	.w6(32'hbc1e653e),
	.w7(32'h3be89400),
	.w8(32'h3c234851),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae24155),
	.w1(32'h3c1d16cb),
	.w2(32'h3bbcfcab),
	.w3(32'h3b3f57e2),
	.w4(32'h3c0c9a29),
	.w5(32'h3af96de1),
	.w6(32'h39b26d01),
	.w7(32'h3c70b078),
	.w8(32'h3c1f785b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb870166c),
	.w1(32'hbb9de642),
	.w2(32'hbbb1c092),
	.w3(32'h3b3793f3),
	.w4(32'hbbb5bf74),
	.w5(32'hbb6b25af),
	.w6(32'h3bfb6a15),
	.w7(32'hbb94c0d2),
	.w8(32'hbab582a2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b389f),
	.w1(32'h3a3b56b8),
	.w2(32'hba4d09d5),
	.w3(32'hbb8feb9f),
	.w4(32'hbb828a2c),
	.w5(32'hbb690893),
	.w6(32'hbaf39cb8),
	.w7(32'hb8a878a1),
	.w8(32'h3a2619f9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11146f),
	.w1(32'h3cb78dfa),
	.w2(32'h3c8def68),
	.w3(32'h3b89d0fd),
	.w4(32'h390f3bdc),
	.w5(32'h3bee9757),
	.w6(32'h3b324d88),
	.w7(32'hbb3f1163),
	.w8(32'hbaeac4f5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f781e),
	.w1(32'h3c24a0e9),
	.w2(32'h3cbfbe46),
	.w3(32'h3a7005df),
	.w4(32'h3c8c64b5),
	.w5(32'h3d11eeac),
	.w6(32'hbb8288e1),
	.w7(32'h3bb1537d),
	.w8(32'h3c7ff422),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7f144),
	.w1(32'h3b515857),
	.w2(32'hbb759e46),
	.w3(32'h3bdee7e6),
	.w4(32'hbbd0750a),
	.w5(32'hbc40f24f),
	.w6(32'hbc031723),
	.w7(32'h3b967097),
	.w8(32'hbb1237e7),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc22dd),
	.w1(32'hbbf58aaa),
	.w2(32'hbbe32977),
	.w3(32'hbc2e84dc),
	.w4(32'hbc246453),
	.w5(32'hbbad2f0f),
	.w6(32'hbc168190),
	.w7(32'hbbbf16f2),
	.w8(32'hbbcbde03),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab24590),
	.w1(32'hbc8a152f),
	.w2(32'hbc221162),
	.w3(32'hba890de2),
	.w4(32'hbc356134),
	.w5(32'h3b0d17a0),
	.w6(32'hbbc7e1cc),
	.w7(32'hba829bd9),
	.w8(32'h3c9878b3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb506df2),
	.w1(32'h3c1e8417),
	.w2(32'h3a4a08d0),
	.w3(32'h3c91b7c4),
	.w4(32'h3b750c77),
	.w5(32'hbbdc5475),
	.w6(32'h3cd7086c),
	.w7(32'hbab2d3e9),
	.w8(32'hbc3ef36f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c7c0b),
	.w1(32'h3ab8bc5b),
	.w2(32'hbb26166f),
	.w3(32'hbb823279),
	.w4(32'hbbad3757),
	.w5(32'hbbd522a4),
	.w6(32'hbc271205),
	.w7(32'hbc155bce),
	.w8(32'h3b4fbb02),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe29a0c),
	.w1(32'hba6c2f63),
	.w2(32'hbbe20bb6),
	.w3(32'hbbea0423),
	.w4(32'hb8d6e6e5),
	.w5(32'hbbcaefbd),
	.w6(32'h3c3f58ce),
	.w7(32'hba918e03),
	.w8(32'hbbd41f26),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a38b2),
	.w1(32'hb9954294),
	.w2(32'h3b3fbb1c),
	.w3(32'hbc23a415),
	.w4(32'h3c1e53fe),
	.w5(32'h3c02c0b1),
	.w6(32'hbc28828c),
	.w7(32'h3c2c24c0),
	.w8(32'h3c8d140d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16f900),
	.w1(32'h3a104cfa),
	.w2(32'hba90e239),
	.w3(32'h39fd8234),
	.w4(32'h3972daab),
	.w5(32'hbb470257),
	.w6(32'h3c05aa53),
	.w7(32'h3b26892f),
	.w8(32'hbb898d6f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aa4f0),
	.w1(32'h3c4ba7b3),
	.w2(32'h3cbc7019),
	.w3(32'h3b5d5594),
	.w4(32'hb8375636),
	.w5(32'hba92e638),
	.w6(32'h3b22d4b3),
	.w7(32'hbacd1bd0),
	.w8(32'h39079418),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ed841),
	.w1(32'h3a17514b),
	.w2(32'h3b794d0b),
	.w3(32'hba1e70e4),
	.w4(32'hbaaf112d),
	.w5(32'hbaaa8daa),
	.w6(32'hbc12ceb4),
	.w7(32'hbb026c78),
	.w8(32'hbbf0d535),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb8cb8),
	.w1(32'hbbd6a456),
	.w2(32'hbac6a365),
	.w3(32'h3a437b27),
	.w4(32'hbadc07aa),
	.w5(32'h398b53a5),
	.w6(32'hbbc5048b),
	.w7(32'hb99c1091),
	.w8(32'hbc18b90e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9890129),
	.w1(32'hbb1efc1b),
	.w2(32'h3b485d58),
	.w3(32'h3b807dc8),
	.w4(32'hbb5ee4d2),
	.w5(32'hba8357ef),
	.w6(32'hbbbdea39),
	.w7(32'hba890f0d),
	.w8(32'h3afa163f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a33d4),
	.w1(32'h3b8b60da),
	.w2(32'h3b3fa0b3),
	.w3(32'hbc7c674a),
	.w4(32'h3b2cab54),
	.w5(32'hbbbfa398),
	.w6(32'hbc4bca77),
	.w7(32'h3b926f80),
	.w8(32'h3b6a6dc3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39442c82),
	.w1(32'hbb8ce5f5),
	.w2(32'hbab85605),
	.w3(32'hbb1808dc),
	.w4(32'hbb8c849c),
	.w5(32'hba612d27),
	.w6(32'h3b110d0e),
	.w7(32'hbae1eafd),
	.w8(32'hbae6ca98),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6b62c),
	.w1(32'hbc029b8a),
	.w2(32'hb9c4c931),
	.w3(32'h3b130ce6),
	.w4(32'hbbafc443),
	.w5(32'h3adf28c7),
	.w6(32'hbaafdcd0),
	.w7(32'hbbb86060),
	.w8(32'hbb157dfc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae09c73),
	.w1(32'h3ae0901e),
	.w2(32'h37ca5467),
	.w3(32'hbb3a8f4b),
	.w4(32'hbad7956a),
	.w5(32'hbb10db31),
	.w6(32'hbba3251a),
	.w7(32'h3bc035ae),
	.w8(32'hba112f3f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd8605),
	.w1(32'hbc22ef91),
	.w2(32'h3adcfe7c),
	.w3(32'hbc090acf),
	.w4(32'hbc5ff11d),
	.w5(32'h3b3c09ad),
	.w6(32'h3a9db856),
	.w7(32'hba177850),
	.w8(32'h3a29a69f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc077990),
	.w1(32'hbb09f418),
	.w2(32'hbb8c8a24),
	.w3(32'hbc1e74a6),
	.w4(32'hbb834c96),
	.w5(32'hbb814db7),
	.w6(32'hbbfa007c),
	.w7(32'hbb9b3c94),
	.w8(32'hbb1a942c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd801ce),
	.w1(32'h3b94b2c1),
	.w2(32'h3b8a8cce),
	.w3(32'h3b72ba97),
	.w4(32'hbaff5ed2),
	.w5(32'h3bc49a15),
	.w6(32'h3b382185),
	.w7(32'hbbb38a33),
	.w8(32'h3bef4f18),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7fc56),
	.w1(32'hbb80e0d0),
	.w2(32'h3afb18d5),
	.w3(32'hbb147f36),
	.w4(32'hbb2b9d77),
	.w5(32'h3c078d9a),
	.w6(32'hb9506300),
	.w7(32'hbb943c78),
	.w8(32'h3b39d801),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b971676),
	.w1(32'h3c31ec3e),
	.w2(32'h3c6ae39e),
	.w3(32'h3bb3a00b),
	.w4(32'h3c32fba9),
	.w5(32'h3c054606),
	.w6(32'hbbcb47f4),
	.w7(32'h3bbfe71a),
	.w8(32'hbb833719),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4259c1),
	.w1(32'hbbdde534),
	.w2(32'h3afe847c),
	.w3(32'h38a82304),
	.w4(32'hba3b175a),
	.w5(32'h3a30eca6),
	.w6(32'hbbac2807),
	.w7(32'hbba925d9),
	.w8(32'hbb53596f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb639758),
	.w1(32'hbb5f00ce),
	.w2(32'hbba4addf),
	.w3(32'hbaefa639),
	.w4(32'hbbc3d3ea),
	.w5(32'h3ab88a8a),
	.w6(32'h3b459e60),
	.w7(32'h3b8e7199),
	.w8(32'h3c896d70),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc574757),
	.w1(32'hbb1bbf54),
	.w2(32'hbb82bae1),
	.w3(32'hba2c6138),
	.w4(32'hbb2fa02f),
	.w5(32'hbb8e5bdf),
	.w6(32'h3c0a6be3),
	.w7(32'hbb6f949b),
	.w8(32'hbb56ba4a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06cfb8),
	.w1(32'hbbc94fb0),
	.w2(32'hbb47966e),
	.w3(32'h3b5d71ea),
	.w4(32'hbc22d357),
	.w5(32'hbbf36d2d),
	.w6(32'h3b3bba17),
	.w7(32'hba383aed),
	.w8(32'h3ab420aa),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cdfd0),
	.w1(32'hbaff3e0c),
	.w2(32'h3aa534f5),
	.w3(32'hbc3d0e5e),
	.w4(32'hbb223317),
	.w5(32'hba3aaf73),
	.w6(32'hbb1f329b),
	.w7(32'h3a50de11),
	.w8(32'hbb29ad4c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7119f),
	.w1(32'h3aa02f86),
	.w2(32'hbaba2546),
	.w3(32'hbbf63d95),
	.w4(32'h3bb7609f),
	.w5(32'h3c24dba2),
	.w6(32'h394e7128),
	.w7(32'h3b12cbee),
	.w8(32'h3bda867e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34a30),
	.w1(32'hbc1a7fb3),
	.w2(32'hbb6b1684),
	.w3(32'h3c3e3b4d),
	.w4(32'hbc138e0b),
	.w5(32'hbbd6d784),
	.w6(32'h3bbf91fd),
	.w7(32'hbc382b4f),
	.w8(32'hbba0cad6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84a435),
	.w1(32'hbc12cbac),
	.w2(32'hbbcb0a5b),
	.w3(32'h3c3bce1b),
	.w4(32'hbc252f2a),
	.w5(32'hbb93a9df),
	.w6(32'h3bd79cc2),
	.w7(32'hbafb8fd8),
	.w8(32'hbb58c5db),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc015a7a),
	.w1(32'hbb2740ca),
	.w2(32'hba0ed1d2),
	.w3(32'hbc0b86ae),
	.w4(32'hbbbf9433),
	.w5(32'hbb74d9b1),
	.w6(32'hbbacd654),
	.w7(32'h3ba1930a),
	.w8(32'h3aa159ca),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f5a56),
	.w1(32'h3bbfc837),
	.w2(32'hbbecc58f),
	.w3(32'hbb138410),
	.w4(32'h3c41c463),
	.w5(32'hbbb313e3),
	.w6(32'hba006015),
	.w7(32'h3c8c4e24),
	.w8(32'hb6f751aa),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3becf2),
	.w1(32'hbb80f20d),
	.w2(32'hbacf6a1f),
	.w3(32'hbc55f50b),
	.w4(32'hbbc2a869),
	.w5(32'hbacd1806),
	.w6(32'hbc3609f5),
	.w7(32'hbbfa0d4b),
	.w8(32'hbb25068f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c4ac1),
	.w1(32'hbb305772),
	.w2(32'h3b9bb78d),
	.w3(32'hb982ddd5),
	.w4(32'hbb2bc676),
	.w5(32'h3c4edc43),
	.w6(32'hbb849991),
	.w7(32'hbbb1d0d8),
	.w8(32'h3c1f6786),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16c3ae),
	.w1(32'hbb2f1408),
	.w2(32'h3c0560e3),
	.w3(32'h3c4ff3e0),
	.w4(32'hbbddd616),
	.w5(32'hbb2b1cee),
	.w6(32'h3bcd71e9),
	.w7(32'hbc09de0a),
	.w8(32'hbbba72a1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e01e0),
	.w1(32'h3bef3156),
	.w2(32'h3b5c1c94),
	.w3(32'h3ba1ad33),
	.w4(32'h3b013b9d),
	.w5(32'h3c0f85fc),
	.w6(32'hbbda4db0),
	.w7(32'hbb81664f),
	.w8(32'hba56c99b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0491c),
	.w1(32'h3b61a7ad),
	.w2(32'h3b0d7d33),
	.w3(32'hbbf8ff28),
	.w4(32'h3c0d4e32),
	.w5(32'h3c473f8d),
	.w6(32'hbbc83628),
	.w7(32'h3cbe6dd5),
	.w8(32'h3cd54d73),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc382d88),
	.w1(32'hbc01b4e6),
	.w2(32'hbbd13ec2),
	.w3(32'hbc2a2370),
	.w4(32'hbbbf3854),
	.w5(32'h3b3aa76c),
	.w6(32'hbb8327b8),
	.w7(32'h3c0571d2),
	.w8(32'h3c7d73a7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3106fc),
	.w1(32'h3b5b9de0),
	.w2(32'h3af8b2fd),
	.w3(32'h3be22468),
	.w4(32'h3b29854b),
	.w5(32'hbb2c3647),
	.w6(32'h3c256c34),
	.w7(32'h3bd8d5b7),
	.w8(32'h3920b142),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980fef9),
	.w1(32'h3bcbe4d5),
	.w2(32'h3b700dca),
	.w3(32'h3a39e7e3),
	.w4(32'h3b703fb2),
	.w5(32'h3b8503d2),
	.w6(32'h3ac71f96),
	.w7(32'h3b0b82a3),
	.w8(32'hbaf94c1d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08de62),
	.w1(32'hbb207c01),
	.w2(32'h3b6a32ad),
	.w3(32'hba486536),
	.w4(32'h3b464fdd),
	.w5(32'h3c3bf502),
	.w6(32'h39cfa085),
	.w7(32'hbb640166),
	.w8(32'h3b2c70c5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950d2ac),
	.w1(32'hbc13ad7f),
	.w2(32'hbbb2a97e),
	.w3(32'h3bd6b4fb),
	.w4(32'hbbc31e1f),
	.w5(32'hb9889621),
	.w6(32'hba82c8ad),
	.w7(32'hbc075083),
	.w8(32'hbbd866bd),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74f683),
	.w1(32'hbbe14cd3),
	.w2(32'h3afad61c),
	.w3(32'hbc54c3db),
	.w4(32'hbc0d2335),
	.w5(32'hbabc7af7),
	.w6(32'hbc797b61),
	.w7(32'hbb6a3a11),
	.w8(32'hbb1f9402),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbec5f4),
	.w1(32'h3babd8f2),
	.w2(32'h3b0ee430),
	.w3(32'hbb2ff615),
	.w4(32'hbb657dba),
	.w5(32'hbbbe4287),
	.w6(32'hbb2ba699),
	.w7(32'h3b84569e),
	.w8(32'h3bd97e84),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ebdb8),
	.w1(32'hba220fbc),
	.w2(32'hbb9e2e4b),
	.w3(32'h3b0d2c23),
	.w4(32'hbbb604cd),
	.w5(32'hbc4fb623),
	.w6(32'hba8c38d3),
	.w7(32'hbb20159f),
	.w8(32'hbbdd7080),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9391b5),
	.w1(32'h3aaac38e),
	.w2(32'hbb494e85),
	.w3(32'h3ae2a5c8),
	.w4(32'hbad24768),
	.w5(32'hbc2fb14a),
	.w6(32'h3a913cc0),
	.w7(32'hbae7863e),
	.w8(32'hbae9631e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e0d30),
	.w1(32'h39c13079),
	.w2(32'h3b98a13f),
	.w3(32'h3b90c666),
	.w4(32'hbb3d04e2),
	.w5(32'h3b80f75a),
	.w6(32'h3bb659ec),
	.w7(32'hbab9a861),
	.w8(32'h3bac9005),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b103229),
	.w1(32'hbae904c5),
	.w2(32'hbaadf131),
	.w3(32'h38a237ba),
	.w4(32'hbaf4dd7e),
	.w5(32'h39c8e624),
	.w6(32'hbb08ad0a),
	.w7(32'hbb7459c6),
	.w8(32'hbb05472a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0eae),
	.w1(32'h3a5cd6cf),
	.w2(32'hba788261),
	.w3(32'hbab39cca),
	.w4(32'hba810d62),
	.w5(32'hbb0e0dad),
	.w6(32'hbafda9cd),
	.w7(32'hbad1049d),
	.w8(32'hbb3d9496),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d2c5c1),
	.w1(32'h3affeac4),
	.w2(32'h3b80c818),
	.w3(32'h3a9a2510),
	.w4(32'h3abaabc2),
	.w5(32'h3b02ede9),
	.w6(32'h3aeedb59),
	.w7(32'hbb20e301),
	.w8(32'h3a9a0711),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4a5a0),
	.w1(32'h3a9c2222),
	.w2(32'h39b96162),
	.w3(32'h3a09b027),
	.w4(32'hb939e7cc),
	.w5(32'hb93f46f0),
	.w6(32'h3a4c0355),
	.w7(32'h39720942),
	.w8(32'h3a943406),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a12db3),
	.w1(32'hbb7aeec4),
	.w2(32'hbb0f4686),
	.w3(32'h3b0404f9),
	.w4(32'hbb91242f),
	.w5(32'hbaabeaa4),
	.w6(32'h3b1fcc9f),
	.w7(32'hbb519fc8),
	.w8(32'hbac96a95),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0a73f),
	.w1(32'hba68360a),
	.w2(32'hbb458be6),
	.w3(32'hbb8597d2),
	.w4(32'hbb930388),
	.w5(32'hbb993790),
	.w6(32'hbb4afce3),
	.w7(32'hb9e191b9),
	.w8(32'h3afb5eae),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28e631),
	.w1(32'h3af8d174),
	.w2(32'h3b2d204c),
	.w3(32'hba83c5f8),
	.w4(32'hba11af02),
	.w5(32'h399c070f),
	.w6(32'hba33ecab),
	.w7(32'hba01834e),
	.w8(32'h3a4e536e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b650e),
	.w1(32'hba171c46),
	.w2(32'h36f1b729),
	.w3(32'h3a79a81f),
	.w4(32'hbaa7c007),
	.w5(32'hba0cd158),
	.w6(32'hb79cca79),
	.w7(32'h39e3f03d),
	.w8(32'h39bd2d20),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef53ee),
	.w1(32'hbae612cb),
	.w2(32'hbac4f87a),
	.w3(32'hbbd7724f),
	.w4(32'hbb7c3a22),
	.w5(32'hbb1657a6),
	.w6(32'hbbcf51a3),
	.w7(32'hbadb549a),
	.w8(32'hbb039f4e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa80723),
	.w1(32'hba18600b),
	.w2(32'h3a28910c),
	.w3(32'h3ac1947d),
	.w4(32'hbb5f0bfb),
	.w5(32'hbaaaab55),
	.w6(32'h3b8d1810),
	.w7(32'h3aa1621a),
	.w8(32'h3b46fb18),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bbb2b),
	.w1(32'h3b825abe),
	.w2(32'h3b32e72a),
	.w3(32'hbad33098),
	.w4(32'hba3938ea),
	.w5(32'h3b0a25f6),
	.w6(32'hbbc31b34),
	.w7(32'h3ad2eb6f),
	.w8(32'h3bbf3747),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b955910),
	.w1(32'h3a609b26),
	.w2(32'hb9100451),
	.w3(32'h3b6899ad),
	.w4(32'hb994289b),
	.w5(32'hb9e128b4),
	.w6(32'h3aa2cdad),
	.w7(32'hb90208e1),
	.w8(32'hba869b97),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a556ede),
	.w1(32'h3acd0ef3),
	.w2(32'h3a97bcee),
	.w3(32'h3a073935),
	.w4(32'h3b343fcc),
	.w5(32'h3a8085e9),
	.w6(32'h38922550),
	.w7(32'h3ab448a4),
	.w8(32'hb9eb5352),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaee211),
	.w1(32'hbb2cc5bf),
	.w2(32'hbae0bfa7),
	.w3(32'hbace4aab),
	.w4(32'hbb531f9c),
	.w5(32'h3b6ad718),
	.w6(32'hbaf2e94b),
	.w7(32'hbb4e5453),
	.w8(32'h3a26af39),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b981e76),
	.w1(32'h3b95042a),
	.w2(32'h3b9bf161),
	.w3(32'h3a6ef7fd),
	.w4(32'hbb195a1d),
	.w5(32'h386ab7cf),
	.w6(32'h3c31ff3b),
	.w7(32'h3bf6d978),
	.w8(32'h3c06e024),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec1256),
	.w1(32'hbb32745e),
	.w2(32'hbb57801c),
	.w3(32'hbb5b9879),
	.w4(32'hbbaa837e),
	.w5(32'hbb4a829a),
	.w6(32'hbb08245f),
	.w7(32'hbb6813e1),
	.w8(32'h371287e3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6cc4b),
	.w1(32'hbb5b67ea),
	.w2(32'hbace940e),
	.w3(32'hbaa38b04),
	.w4(32'hbbd23854),
	.w5(32'hbba6c14e),
	.w6(32'hbb756740),
	.w7(32'hbacfc6eb),
	.w8(32'hba375489),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2fa26),
	.w1(32'h39fb0b43),
	.w2(32'h3a0a449b),
	.w3(32'h394109ac),
	.w4(32'h39820cb2),
	.w5(32'hb758626c),
	.w6(32'hbb160c54),
	.w7(32'hb9e19bd2),
	.w8(32'hbaa5b6a0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f6da7),
	.w1(32'hb9c99ee4),
	.w2(32'h39edcdc8),
	.w3(32'h3b12f67a),
	.w4(32'h3a128ee5),
	.w5(32'hb8e08e06),
	.w6(32'hb981a49b),
	.w7(32'h3a75ef2b),
	.w8(32'h3b07fc84),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae63414),
	.w1(32'hbc056971),
	.w2(32'hba375216),
	.w3(32'h3b527518),
	.w4(32'hbb974565),
	.w5(32'h3b538214),
	.w6(32'h3abd9e56),
	.w7(32'hbb1e4399),
	.w8(32'h3b1465f6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fdb97),
	.w1(32'h3c350308),
	.w2(32'h3be00813),
	.w3(32'h3c123c99),
	.w4(32'h3bc8239b),
	.w5(32'h3ba91189),
	.w6(32'h3c0ef069),
	.w7(32'h3c0b1b28),
	.w8(32'h3c09b1cd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8271ef),
	.w1(32'hb9bd463b),
	.w2(32'h3b81c78f),
	.w3(32'h3b0777fa),
	.w4(32'h3a8b581f),
	.w5(32'h3ae63d54),
	.w6(32'h3b569814),
	.w7(32'h3a87abcc),
	.w8(32'h3b0b7582),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bce729),
	.w1(32'h39e74d63),
	.w2(32'h38bb5019),
	.w3(32'hbaabd6fa),
	.w4(32'hb9fab4d6),
	.w5(32'hbb0b9e65),
	.w6(32'hbb4131a7),
	.w7(32'hba345b75),
	.w8(32'hbb054cd4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081514),
	.w1(32'hba9275a0),
	.w2(32'hbb01f83e),
	.w3(32'hbaf1ccd0),
	.w4(32'hbbaf30fd),
	.w5(32'hbb804041),
	.w6(32'hba1984e8),
	.w7(32'hbb414864),
	.w8(32'hba45e293),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae73f52),
	.w1(32'hbb3226ea),
	.w2(32'hbb3f4d61),
	.w3(32'h395e969f),
	.w4(32'hbb18ef2d),
	.w5(32'hbab240d6),
	.w6(32'h3a5c62ee),
	.w7(32'hba83f823),
	.w8(32'h3a434369),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd01e7),
	.w1(32'hbaa9c6df),
	.w2(32'hbb901fa7),
	.w3(32'hba9aee6c),
	.w4(32'hba81b352),
	.w5(32'hba15f84e),
	.w6(32'hb660bbba),
	.w7(32'hbb0502d4),
	.w8(32'h3a064569),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaccc5e),
	.w1(32'hb9356ddc),
	.w2(32'hbb0bdf91),
	.w3(32'hbb2bfbbc),
	.w4(32'hbaf0a0ff),
	.w5(32'hb8c9c6b5),
	.w6(32'hbb5aae9c),
	.w7(32'hbb22ce30),
	.w8(32'h3a064b39),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9490a3),
	.w1(32'hba9bf765),
	.w2(32'hb9738a15),
	.w3(32'hb9ec6e5d),
	.w4(32'hbb07d27d),
	.w5(32'h39707964),
	.w6(32'h3a0ac608),
	.w7(32'hbad7cb3f),
	.w8(32'hb9ef8f2f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb388659),
	.w1(32'hbab05d31),
	.w2(32'hbaded1bc),
	.w3(32'hbb1124f9),
	.w4(32'hbb55c299),
	.w5(32'hbb17a728),
	.w6(32'hbb678cb0),
	.w7(32'hba9b10ac),
	.w8(32'hb9e8cf2e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77df25),
	.w1(32'h394cac10),
	.w2(32'h3b933328),
	.w3(32'hb9a8bdd9),
	.w4(32'hbb891245),
	.w5(32'h389bad73),
	.w6(32'h3b9a411c),
	.w7(32'h3ae5073f),
	.w8(32'h3b4b8f02),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8240c),
	.w1(32'hb81fb1d7),
	.w2(32'hbb1e9d3b),
	.w3(32'hbb2aa06a),
	.w4(32'hbb754a20),
	.w5(32'hbb12a462),
	.w6(32'hbaf36992),
	.w7(32'hbb88bcc6),
	.w8(32'h39b3cc88),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1782c),
	.w1(32'h39f34f66),
	.w2(32'hbade43d9),
	.w3(32'hb92f45bf),
	.w4(32'h3a0d3508),
	.w5(32'hba5f6f36),
	.w6(32'hba21660c),
	.w7(32'h39b60bfa),
	.w8(32'h38597d22),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3168aa),
	.w1(32'h3aaabd07),
	.w2(32'h3c0be387),
	.w3(32'h3b7d6776),
	.w4(32'h3ab280b0),
	.w5(32'h3b554137),
	.w6(32'h3b146f94),
	.w7(32'h3abae108),
	.w8(32'h3bc69a9a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb9fec),
	.w1(32'hba968043),
	.w2(32'hba26c6a9),
	.w3(32'hb88dbaad),
	.w4(32'hbb2a50aa),
	.w5(32'h3ab42ecc),
	.w6(32'h3a2d946f),
	.w7(32'h3b04dc60),
	.w8(32'h3b387a4b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac85b4),
	.w1(32'h3a4e91b9),
	.w2(32'h3a80554b),
	.w3(32'hba38c7c9),
	.w4(32'h39cd82d8),
	.w5(32'h3aa000f2),
	.w6(32'hba53e666),
	.w7(32'h3839a258),
	.w8(32'h3a24638c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25a175),
	.w1(32'h3b9b216f),
	.w2(32'h3b85a9ad),
	.w3(32'h3bbf1b95),
	.w4(32'h3b3dfde9),
	.w5(32'h3b76d0d9),
	.w6(32'h3b46ab70),
	.w7(32'h3b4545f0),
	.w8(32'h3b9da3ee),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a218eb),
	.w1(32'hb8e65405),
	.w2(32'hb95cadf2),
	.w3(32'h3a0d6de5),
	.w4(32'h3aaa4da3),
	.w5(32'h378e3393),
	.w6(32'h3a49d89e),
	.w7(32'h3a27de2c),
	.w8(32'hba8b3b6c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b4219),
	.w1(32'hbaaef627),
	.w2(32'hbaec8d11),
	.w3(32'hbb0c0517),
	.w4(32'hbb072cbe),
	.w5(32'hbabe2e5d),
	.w6(32'hbadef29b),
	.w7(32'hba610b53),
	.w8(32'hb9909914),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8fb22),
	.w1(32'h3a021538),
	.w2(32'hb8f2c14b),
	.w3(32'hba62bf07),
	.w4(32'hba078d54),
	.w5(32'h3986c022),
	.w6(32'hbad3dad3),
	.w7(32'h39cd36b8),
	.w8(32'hb74f424a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac594bd),
	.w1(32'hba8d0d67),
	.w2(32'hba282efd),
	.w3(32'hb9a3bafd),
	.w4(32'hbad7038d),
	.w5(32'hba914a72),
	.w6(32'hba581905),
	.w7(32'hba8cdc08),
	.w8(32'hb9f04839),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c9cdf),
	.w1(32'hba6103e5),
	.w2(32'hbb900cb8),
	.w3(32'h3a8b6383),
	.w4(32'hba832c85),
	.w5(32'h39fc37cf),
	.w6(32'hbb28cf81),
	.w7(32'hba9249ab),
	.w8(32'hbadb57a1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1858f6),
	.w1(32'h3af4ee07),
	.w2(32'hba067549),
	.w3(32'hbb5b7d07),
	.w4(32'hbbbd3eda),
	.w5(32'hbb7c32ba),
	.w6(32'h3b2993e3),
	.w7(32'h3b39f31e),
	.w8(32'h3b89e7bf),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b936f27),
	.w1(32'h3b9e6133),
	.w2(32'h3bb0b2a2),
	.w3(32'h3b940743),
	.w4(32'h3ade7da9),
	.w5(32'h3b664763),
	.w6(32'h3b1671b6),
	.w7(32'h3b2107ff),
	.w8(32'h3bb9bcd7),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6923ec),
	.w1(32'h39226326),
	.w2(32'h3aa6cddf),
	.w3(32'h39c2fa3f),
	.w4(32'h39b1779a),
	.w5(32'hbad3f8cc),
	.w6(32'h3a8ab372),
	.w7(32'h3b97b178),
	.w8(32'h3ba6e221),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeee6a5),
	.w1(32'hb9ac5cd7),
	.w2(32'h39d7461d),
	.w3(32'h3a4b6494),
	.w4(32'h3a288720),
	.w5(32'h38816e13),
	.w6(32'h3a8b86db),
	.w7(32'hb9934f1c),
	.w8(32'hba7a8457),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68046b),
	.w1(32'hba5a5a32),
	.w2(32'hbb107c6c),
	.w3(32'hb7d93e0b),
	.w4(32'hb914e583),
	.w5(32'hb99204db),
	.w6(32'hba1ef245),
	.w7(32'hba3f5060),
	.w8(32'h39df8930),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93ee40),
	.w1(32'hba3f99dc),
	.w2(32'hb9e1b532),
	.w3(32'h3ae05fa2),
	.w4(32'h38e0ca43),
	.w5(32'hb994f292),
	.w6(32'h3b07048f),
	.w7(32'hbabcc5aa),
	.w8(32'hba640b2c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ba7fd),
	.w1(32'h3b04a45d),
	.w2(32'h3ac8fee2),
	.w3(32'hba20ab12),
	.w4(32'h3a95125a),
	.w5(32'hba8bbd9e),
	.w6(32'hbaad56c3),
	.w7(32'hba372c8a),
	.w8(32'hb9d64e9d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b24c0),
	.w1(32'h3b353499),
	.w2(32'h3baa8e10),
	.w3(32'h39d53c0f),
	.w4(32'h3ad5c042),
	.w5(32'h3b11c2f7),
	.w6(32'h3ab379ed),
	.w7(32'h3b1d98fc),
	.w8(32'h3b0e03f6),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f28545),
	.w1(32'hbaf4de06),
	.w2(32'h3a026d01),
	.w3(32'h3a6bfcf0),
	.w4(32'hb9e69c57),
	.w5(32'h3b0890c1),
	.w6(32'h3a93ec4f),
	.w7(32'hb85dd521),
	.w8(32'h3acc565b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa80f5e),
	.w1(32'hb9567d58),
	.w2(32'h3aae983c),
	.w3(32'h3a93cdf6),
	.w4(32'h386c0b18),
	.w5(32'h3a92c452),
	.w6(32'h3ae31c3b),
	.w7(32'h3a1d6737),
	.w8(32'h3b3ee438),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe0e86),
	.w1(32'hb91d66b8),
	.w2(32'hb9f081d8),
	.w3(32'h3b5ebfe2),
	.w4(32'hba31ce29),
	.w5(32'hb9120c4b),
	.w6(32'h3b238389),
	.w7(32'hba1a4fca),
	.w8(32'h3b0ed6bd),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ac90d),
	.w1(32'h397a2548),
	.w2(32'hba9d169c),
	.w3(32'h3ab090f3),
	.w4(32'hb8d51647),
	.w5(32'h3a652e0d),
	.w6(32'hba94125e),
	.w7(32'hba9d49f2),
	.w8(32'hba4a493e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99aca00),
	.w1(32'h3a64c61a),
	.w2(32'h3a8b910f),
	.w3(32'hbaa17311),
	.w4(32'hb9f723c3),
	.w5(32'h3ae95cad),
	.w6(32'hbae9c858),
	.w7(32'h36a5bfbd),
	.w8(32'h3b85ee67),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39583be4),
	.w1(32'hb8e69a0a),
	.w2(32'h38bbcac5),
	.w3(32'hba673fa6),
	.w4(32'hbabde3e4),
	.w5(32'hbb067004),
	.w6(32'hba1aa370),
	.w7(32'hba0cefad),
	.w8(32'h39966ce1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f1665),
	.w1(32'h3c1e4d12),
	.w2(32'h3c0a5603),
	.w3(32'h3a5c2cc3),
	.w4(32'h3bab0bcb),
	.w5(32'h3ba21ee2),
	.w6(32'h3bcb8838),
	.w7(32'h3c08dcff),
	.w8(32'h3b5abd71),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefe2a5),
	.w1(32'hbb200b7f),
	.w2(32'hba39bed6),
	.w3(32'hba6ecf30),
	.w4(32'hbae3e9ce),
	.w5(32'h3b07b32e),
	.w6(32'h3a071b30),
	.w7(32'hbaf36198),
	.w8(32'hba495734),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ef374),
	.w1(32'h3a83269f),
	.w2(32'hbb23e30f),
	.w3(32'h3af8aaf3),
	.w4(32'hbb225560),
	.w5(32'hbb403fc3),
	.w6(32'h3b8047e2),
	.w7(32'hbb1d6b46),
	.w8(32'hbb15c634),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule