module layer_10_featuremap_258(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf71d9b),
	.w1(32'h3b81e71c),
	.w2(32'h3be5db7f),
	.w3(32'hbba8bde6),
	.w4(32'h3ab7548b),
	.w5(32'hbaca228c),
	.w6(32'hbb1fd0c6),
	.w7(32'h3b1264b9),
	.w8(32'hba10d8b3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb432bec),
	.w1(32'h3a53541d),
	.w2(32'h36a6ce7c),
	.w3(32'hbc4e98e9),
	.w4(32'hbbdbf9b6),
	.w5(32'h3b0e00d1),
	.w6(32'hbc2bf685),
	.w7(32'hbc15b7c5),
	.w8(32'hbb9025cb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d3cb),
	.w1(32'h394bfea4),
	.w2(32'h3a839ea7),
	.w3(32'h3ad4fb9c),
	.w4(32'h3a92fa7e),
	.w5(32'h3a1516b9),
	.w6(32'h3a22f990),
	.w7(32'hbb6a6ce0),
	.w8(32'h3b1aee67),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8ff52),
	.w1(32'h3a317a25),
	.w2(32'hbba9e3be),
	.w3(32'hba7f8b66),
	.w4(32'h3a08b92c),
	.w5(32'h39de08cf),
	.w6(32'hb9f6a200),
	.w7(32'h398e870c),
	.w8(32'hbb65e228),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1638bb),
	.w1(32'hbb56c205),
	.w2(32'hbadfb33f),
	.w3(32'hbbdee269),
	.w4(32'hbb032f8a),
	.w5(32'hba5c82f7),
	.w6(32'hbc217ade),
	.w7(32'hbb890314),
	.w8(32'hbb43f1d9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b060145),
	.w1(32'h39790d83),
	.w2(32'h3a1d0e17),
	.w3(32'hbbb08426),
	.w4(32'hb8c998b9),
	.w5(32'h3a36d129),
	.w6(32'hbb9fd32b),
	.w7(32'h3afd40ab),
	.w8(32'hba33a5b8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb124081),
	.w1(32'hbc931ac6),
	.w2(32'hba22a0bd),
	.w3(32'hbb4417b2),
	.w4(32'hbc06cbba),
	.w5(32'h3c2b68d0),
	.w6(32'h3b50025d),
	.w7(32'h3aa2a969),
	.w8(32'h3b777f25),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a910999),
	.w1(32'h3c801680),
	.w2(32'h3cd01ca1),
	.w3(32'h3b743c05),
	.w4(32'h3ca7f58c),
	.w5(32'h3c4aa2d6),
	.w6(32'h3d413b79),
	.w7(32'h3c769864),
	.w8(32'h3baf3f63),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b411cb5),
	.w1(32'h3aaa9b54),
	.w2(32'h3b7b977c),
	.w3(32'hbb38d053),
	.w4(32'h3aa9c05f),
	.w5(32'hba6ebba9),
	.w6(32'hbb660201),
	.w7(32'h3b0c0e88),
	.w8(32'hbb06794f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab5ee3),
	.w1(32'hbb7cf09c),
	.w2(32'hbb87a3dd),
	.w3(32'hbc469c99),
	.w4(32'hbbe4e629),
	.w5(32'hbb2a1568),
	.w6(32'hbb03f767),
	.w7(32'h3a53c11a),
	.w8(32'hbbd1c2a1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6600d9),
	.w1(32'h3b1ebbd1),
	.w2(32'h3977497b),
	.w3(32'hbc0173a1),
	.w4(32'hbab7f63a),
	.w5(32'h3b14d055),
	.w6(32'hbbb8d6da),
	.w7(32'hb9e717d1),
	.w8(32'h3b8b45ad),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c170d47),
	.w1(32'hbccadef8),
	.w2(32'hbc6a68bb),
	.w3(32'h3ba7514b),
	.w4(32'hbba66e49),
	.w5(32'hbbb38ac3),
	.w6(32'h3cda17e7),
	.w7(32'h3c38783b),
	.w8(32'hbb9b772c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0e5d3),
	.w1(32'hba02e260),
	.w2(32'hbb03d5d8),
	.w3(32'h3a923edf),
	.w4(32'hbc120a14),
	.w5(32'hbb833fa1),
	.w6(32'h3c381e8d),
	.w7(32'h3b3c7e70),
	.w8(32'hbbdd88fb),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099192),
	.w1(32'hbbf9f6ad),
	.w2(32'h3bc9919c),
	.w3(32'hbbd4af0e),
	.w4(32'h39bc16d7),
	.w5(32'h3bfb494e),
	.w6(32'hbaabc6c0),
	.w7(32'hba6dcedf),
	.w8(32'h3b9fbc31),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e1cbe),
	.w1(32'h3ba45c1b),
	.w2(32'hbb0d5ed6),
	.w3(32'hbc2503dc),
	.w4(32'hbb4eb30a),
	.w5(32'hba9501bc),
	.w6(32'hbbfc1a7a),
	.w7(32'hbadacc49),
	.w8(32'h3b7400ad),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66cde5),
	.w1(32'hbc414f49),
	.w2(32'h3b91a0e5),
	.w3(32'hbc93cd1a),
	.w4(32'hbbf08d20),
	.w5(32'hbaa8a562),
	.w6(32'hbbde5147),
	.w7(32'h3a80a0db),
	.w8(32'h3b066aaf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba431e5a),
	.w1(32'h3a7c64a3),
	.w2(32'hbb06ffca),
	.w3(32'hbad7a373),
	.w4(32'h3b13c6e7),
	.w5(32'h3965b4d3),
	.w6(32'hbad35aeb),
	.w7(32'h387ee8c5),
	.w8(32'hb9cb18cd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c7358),
	.w1(32'hbbed8cfb),
	.w2(32'h3bb8f5c3),
	.w3(32'h3b801ba7),
	.w4(32'h396789f8),
	.w5(32'h3c3e1eff),
	.w6(32'h3c24b90f),
	.w7(32'hbb8b41f9),
	.w8(32'hbc61b945),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48a7c7),
	.w1(32'hbbd0b358),
	.w2(32'hbb0cc5bd),
	.w3(32'h3b74c005),
	.w4(32'hbb1f353e),
	.w5(32'hbb97be19),
	.w6(32'h3bef6a90),
	.w7(32'hba2aeddd),
	.w8(32'hbc4f6aca),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8b6e1),
	.w1(32'hbaa82631),
	.w2(32'hbb44386d),
	.w3(32'hba3e441a),
	.w4(32'hbaea9be9),
	.w5(32'h3afbd6e0),
	.w6(32'hba7df2f9),
	.w7(32'hbba73450),
	.w8(32'hba0f74b2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff7c49),
	.w1(32'hbbeb6ecf),
	.w2(32'hba9844e4),
	.w3(32'hbc0bec2b),
	.w4(32'hbba95e19),
	.w5(32'hba182e28),
	.w6(32'hbb5ca282),
	.w7(32'hba11e207),
	.w8(32'h3b63ca24),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06be6e),
	.w1(32'h3b9e13e0),
	.w2(32'h3aef77ed),
	.w3(32'hbaad3bdd),
	.w4(32'h3a9d32a2),
	.w5(32'hbb333dca),
	.w6(32'hbae7672c),
	.w7(32'h3b73c635),
	.w8(32'h3b1402ad),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad92023),
	.w1(32'hbb828545),
	.w2(32'h3c0d1ee5),
	.w3(32'hbb8616ae),
	.w4(32'hbb32ef4c),
	.w5(32'h3c369d46),
	.w6(32'hbb6a3d20),
	.w7(32'h3b53009f),
	.w8(32'hbc402946),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc139632),
	.w1(32'hbbc4d062),
	.w2(32'h3c34bd63),
	.w3(32'hbc667ce2),
	.w4(32'hbbcd8c92),
	.w5(32'hb7ac390c),
	.w6(32'hbc48f641),
	.w7(32'h3c17d74a),
	.w8(32'hbb54b660),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b7ff4),
	.w1(32'h3c9ce121),
	.w2(32'h3c26e2a8),
	.w3(32'hbc2c8f10),
	.w4(32'hb93207b0),
	.w5(32'hbbbdd6bb),
	.w6(32'hbcc8f1e9),
	.w7(32'hbba9a2f8),
	.w8(32'h3bca56c4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383d0569),
	.w1(32'hbb39a1d2),
	.w2(32'hb9eaa643),
	.w3(32'hbb631b69),
	.w4(32'hbadedc0e),
	.w5(32'hbacbc20a),
	.w6(32'h3af1c518),
	.w7(32'h3aaf0fef),
	.w8(32'hbb1c8dbf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77cb8b),
	.w1(32'hbab97513),
	.w2(32'hbac21f93),
	.w3(32'hbad108e8),
	.w4(32'hbaf535d1),
	.w5(32'h3a1eee04),
	.w6(32'hbacd63f7),
	.w7(32'hbab496d2),
	.w8(32'hbb5de7ab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b538fb3),
	.w1(32'h3c3b2a27),
	.w2(32'hbb3bf503),
	.w3(32'hbc74a0f9),
	.w4(32'h3b99e930),
	.w5(32'h3b22f9bb),
	.w6(32'hbbf5bf2f),
	.w7(32'h3badcb59),
	.w8(32'hbaacc74a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a968b77),
	.w1(32'hba87292c),
	.w2(32'hbbadafbb),
	.w3(32'h3a5e1850),
	.w4(32'hbb5fccc3),
	.w5(32'hbaed7d79),
	.w6(32'hbb6eb8ea),
	.w7(32'hbbf29e93),
	.w8(32'hbaf7338f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf684c),
	.w1(32'h3b041661),
	.w2(32'hbbbfeacf),
	.w3(32'hbcefbdbe),
	.w4(32'hbb273d8a),
	.w5(32'h3b3686cd),
	.w6(32'hbcc334b8),
	.w7(32'hbbe50650),
	.w8(32'h3c0dd1f9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd3e63),
	.w1(32'h3b454bd8),
	.w2(32'h3b8b2452),
	.w3(32'h3c1b462b),
	.w4(32'h3b674963),
	.w5(32'hbb0b4d4a),
	.w6(32'h3afe84b5),
	.w7(32'h3bb9267e),
	.w8(32'hbbf8fec1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0e68),
	.w1(32'hbb57df2f),
	.w2(32'hbbaec915),
	.w3(32'hbb8e80a5),
	.w4(32'h39cf4134),
	.w5(32'hb8ba9d90),
	.w6(32'hbb6b7953),
	.w7(32'hbb573860),
	.w8(32'hbb40852d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924e1e1),
	.w1(32'hbb7f3fe0),
	.w2(32'hbb0f88a1),
	.w3(32'hbb211514),
	.w4(32'hbbb824f5),
	.w5(32'hba45129e),
	.w6(32'h3b1c60d6),
	.w7(32'hbad674a4),
	.w8(32'h3b17aa87),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bfa8b),
	.w1(32'h39dbc7fd),
	.w2(32'h3b0a03bc),
	.w3(32'hbbcd63fa),
	.w4(32'hbbfe9fd4),
	.w5(32'hbbffb722),
	.w6(32'hbc0aa7ec),
	.w7(32'hbba8393f),
	.w8(32'h3b6141b5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26056f),
	.w1(32'h3c118a5c),
	.w2(32'h3b211b4d),
	.w3(32'hbbf5754a),
	.w4(32'hbbcef658),
	.w5(32'h3b3aee75),
	.w6(32'h3ad78405),
	.w7(32'hba897db3),
	.w8(32'h3b11b427),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15266e),
	.w1(32'h3b4a6b80),
	.w2(32'h3bbe0fa2),
	.w3(32'h3c427e9c),
	.w4(32'hbb22e546),
	.w5(32'hbb11526d),
	.w6(32'h3ba1fb4b),
	.w7(32'h3b8d9802),
	.w8(32'hbbd71977),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d256c2c),
	.w1(32'hbcc5f570),
	.w2(32'hbc85917b),
	.w3(32'hbb23ca48),
	.w4(32'hbd2c8073),
	.w5(32'hbbec092d),
	.w6(32'hbbc8c523),
	.w7(32'hbcac3c34),
	.w8(32'hbc6bae35),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c4fa3),
	.w1(32'h3c915361),
	.w2(32'h3ba5934f),
	.w3(32'hbd0104bd),
	.w4(32'hbb3d80d3),
	.w5(32'h3aa2495b),
	.w6(32'hbd099966),
	.w7(32'h3b8c3d5d),
	.w8(32'h3cab1321),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e68bc),
	.w1(32'h3d12b4b5),
	.w2(32'h3c946b40),
	.w3(32'hbae88dce),
	.w4(32'h3c5ef4b5),
	.w5(32'h3bedb04a),
	.w6(32'hbcefd5a4),
	.w7(32'h3a6a3a80),
	.w8(32'h3cf03909),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac10952),
	.w1(32'h3b35a60c),
	.w2(32'h3b647c60),
	.w3(32'hba9ef31a),
	.w4(32'hba455865),
	.w5(32'hbab995f9),
	.w6(32'hbb058be0),
	.w7(32'h3b08c087),
	.w8(32'h3b82765d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d6ec4),
	.w1(32'hb8b68636),
	.w2(32'hbb8b3b85),
	.w3(32'h3ac46c20),
	.w4(32'h3b85f168),
	.w5(32'h3a53f540),
	.w6(32'h3be7c7d2),
	.w7(32'h3b24abd5),
	.w8(32'h3aa4b7d4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d790b6),
	.w1(32'hba4bd455),
	.w2(32'hbaa2f590),
	.w3(32'hbaf445ea),
	.w4(32'h3a5e105d),
	.w5(32'h3a2f33c4),
	.w6(32'h3a6ebdf9),
	.w7(32'hbadae9df),
	.w8(32'hbb0336fa),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaabbad),
	.w1(32'hba3b0bf0),
	.w2(32'h3a3bad9b),
	.w3(32'h3b4fa327),
	.w4(32'h3b23354e),
	.w5(32'h39d71f93),
	.w6(32'hbaccdf98),
	.w7(32'h3b31a48b),
	.w8(32'hbac2ddf4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd68778),
	.w1(32'hb9de4245),
	.w2(32'h3bc54217),
	.w3(32'h3b942e87),
	.w4(32'h3af6edad),
	.w5(32'h3aade9fc),
	.w6(32'h3bf5053b),
	.w7(32'h3a8e3bed),
	.w8(32'hbc4a76c9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b096),
	.w1(32'h3bd5dfcc),
	.w2(32'h3a1348bf),
	.w3(32'hbc16a18c),
	.w4(32'hbab2a070),
	.w5(32'hbbbf6eae),
	.w6(32'hbc22bdb7),
	.w7(32'h378154f8),
	.w8(32'h3bf3dc5b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4557e9),
	.w1(32'h3b2fe381),
	.w2(32'h3ae93be0),
	.w3(32'h3a932118),
	.w4(32'hb8f819c2),
	.w5(32'hbc479c92),
	.w6(32'h3b03a292),
	.w7(32'hb9caa6a8),
	.w8(32'hbbcdf6a3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0968ea),
	.w1(32'hbb1659f0),
	.w2(32'hbb6b409d),
	.w3(32'hbc3eb76d),
	.w4(32'hbb18b745),
	.w5(32'hbb2b65bb),
	.w6(32'hbb6b830c),
	.w7(32'hba7d4e24),
	.w8(32'h3accf407),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02404d),
	.w1(32'hbb327c48),
	.w2(32'h39148dd8),
	.w3(32'h3be94f0e),
	.w4(32'hbaef8d27),
	.w5(32'h3b11f438),
	.w6(32'h3cbc5560),
	.w7(32'h3ada7690),
	.w8(32'hbc504a6c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1c5e5),
	.w1(32'h3b0238ee),
	.w2(32'h3b80d9d5),
	.w3(32'h3a6b7718),
	.w4(32'h3a1c2aa4),
	.w5(32'hbab8e0b4),
	.w6(32'h3b39ebc6),
	.w7(32'h3b5c710c),
	.w8(32'h3acb7f09),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fc7ec),
	.w1(32'h3adf0ff8),
	.w2(32'h38e8a0fc),
	.w3(32'hbaf15695),
	.w4(32'hb8693bc0),
	.w5(32'h3bcad93d),
	.w6(32'h3a581cc2),
	.w7(32'h3a3a05f5),
	.w8(32'h3b0b21a3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd446e9),
	.w1(32'h3ad5c694),
	.w2(32'h3bc3e6e9),
	.w3(32'hba069ba7),
	.w4(32'hba6a94c7),
	.w5(32'h3993face),
	.w6(32'hbb1f3151),
	.w7(32'h3a4234a3),
	.w8(32'hb86227d9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6da379),
	.w1(32'hbaf352c7),
	.w2(32'h3b6868ba),
	.w3(32'h3b1ae909),
	.w4(32'h3b80dd9a),
	.w5(32'h395a2aa6),
	.w6(32'hbbd7c21f),
	.w7(32'h3b627862),
	.w8(32'hbb6130ad),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb911a2e),
	.w1(32'hbb9864a4),
	.w2(32'hbb916ad2),
	.w3(32'h39da6212),
	.w4(32'hbb6d3571),
	.w5(32'hbae4f503),
	.w6(32'hbaa4bfd1),
	.w7(32'hbb8d94bb),
	.w8(32'h3a26d020),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb812c708),
	.w1(32'hbc58fec1),
	.w2(32'hbc138ccd),
	.w3(32'hbc3c8ceb),
	.w4(32'hbbd3e850),
	.w5(32'hba2f296b),
	.w6(32'h3ca64172),
	.w7(32'hbbebc816),
	.w8(32'hbc642bc7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5acbb7),
	.w1(32'hbb43446f),
	.w2(32'hbb81d418),
	.w3(32'h3a88dcb0),
	.w4(32'hb849aaa6),
	.w5(32'hba855be4),
	.w6(32'h3b825570),
	.w7(32'hbb4ad84e),
	.w8(32'hba8b4b30),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac620de),
	.w1(32'h3b72dbc2),
	.w2(32'h3b015463),
	.w3(32'hbb4bf283),
	.w4(32'hbbaad477),
	.w5(32'h3a1d76d2),
	.w6(32'hb983df00),
	.w7(32'hbb56551d),
	.w8(32'h3b4b55ca),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b969c7d),
	.w1(32'h3a2a9221),
	.w2(32'hbac9592c),
	.w3(32'h3a5391e8),
	.w4(32'h3b20bf3e),
	.w5(32'hba8670db),
	.w6(32'h3b5f6cf8),
	.w7(32'h3ac99fa0),
	.w8(32'hbb2bd372),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc60658),
	.w1(32'hbbb24b04),
	.w2(32'hbba84d08),
	.w3(32'hbb7d43c4),
	.w4(32'hbb1b7fe3),
	.w5(32'h3b043b7e),
	.w6(32'hba9b7e6c),
	.w7(32'hbb20c0f2),
	.w8(32'h3ad31e32),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa07c2),
	.w1(32'h3a244c44),
	.w2(32'h3a5b75ac),
	.w3(32'hbb5d01ee),
	.w4(32'h3a8186c9),
	.w5(32'hbba48f6c),
	.w6(32'hbaa7517a),
	.w7(32'h3b2b0796),
	.w8(32'hbbeb83bf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae7165),
	.w1(32'hbc01340e),
	.w2(32'hbbe97bd5),
	.w3(32'hbb521cd7),
	.w4(32'hbb488e3e),
	.w5(32'h3b9680de),
	.w6(32'hbace690f),
	.w7(32'hbbc73aac),
	.w8(32'h3c02fc71),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8406e),
	.w1(32'h3c44f652),
	.w2(32'h3bec97e0),
	.w3(32'h3c6ef0ef),
	.w4(32'h3c2a4efd),
	.w5(32'h3b863818),
	.w6(32'hbb2e6462),
	.w7(32'hbbffcb91),
	.w8(32'hbb2d7356),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4d511),
	.w1(32'h3bb782e3),
	.w2(32'hb90956a7),
	.w3(32'h3baa86b6),
	.w4(32'h3ca32e9a),
	.w5(32'hbaccfd17),
	.w6(32'hba54bf98),
	.w7(32'h3b04ee35),
	.w8(32'hbc429493),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b2724),
	.w1(32'h3ba0fe8c),
	.w2(32'h3b57da44),
	.w3(32'hb8ca8b66),
	.w4(32'hbb1764dd),
	.w5(32'hbb4e9dd3),
	.w6(32'hbac1f982),
	.w7(32'hbaeb2274),
	.w8(32'h39c44b6a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e3b0c),
	.w1(32'h3b04523d),
	.w2(32'hbae33c22),
	.w3(32'hbb8efb93),
	.w4(32'hbac0ea63),
	.w5(32'hbb1d9719),
	.w6(32'h3a44ec0c),
	.w7(32'hbb217cf7),
	.w8(32'hbb12a214),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a15a8),
	.w1(32'hbb8b9ea9),
	.w2(32'hbb6bb786),
	.w3(32'hbb63e9b5),
	.w4(32'h3a25679e),
	.w5(32'h3a75f287),
	.w6(32'hbb838466),
	.w7(32'hbb303666),
	.w8(32'hbb15294d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73adc6),
	.w1(32'hbbbdbf1d),
	.w2(32'hbba16fde),
	.w3(32'h3b58e9ae),
	.w4(32'h3aeb21c5),
	.w5(32'h3b58b8aa),
	.w6(32'h3a9d8ee6),
	.w7(32'hbaae0c24),
	.w8(32'hbb59885c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2964fd),
	.w1(32'hbc1f16f4),
	.w2(32'hbc7e253d),
	.w3(32'hbcefce9d),
	.w4(32'hbad9e9b4),
	.w5(32'h3b76d4d0),
	.w6(32'h3cc416c2),
	.w7(32'hba9553b0),
	.w8(32'hbb604806),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80717e),
	.w1(32'hbbd9fb8b),
	.w2(32'hba48779c),
	.w3(32'h3c1f0568),
	.w4(32'hbb5a8baf),
	.w5(32'h3a9e29f5),
	.w6(32'h3bce7fa0),
	.w7(32'hb98bae08),
	.w8(32'h3a5fbd10),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2546e),
	.w1(32'hbb627a07),
	.w2(32'h3c05f865),
	.w3(32'h3b503571),
	.w4(32'h3bd0cb92),
	.w5(32'hb91c54f3),
	.w6(32'hbb637657),
	.w7(32'hb98a4b0a),
	.w8(32'hbbf415ef),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99c86e),
	.w1(32'h3c11f9a7),
	.w2(32'hbbe66511),
	.w3(32'hbc7a512e),
	.w4(32'hb9f5080c),
	.w5(32'hbc68a27d),
	.w6(32'hbce8cea8),
	.w7(32'h39fe05f7),
	.w8(32'h3b03e0ea),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c227d),
	.w1(32'hbb4f6516),
	.w2(32'hbabc9535),
	.w3(32'hba148275),
	.w4(32'h372dfe56),
	.w5(32'h3c2b4193),
	.w6(32'hbb006963),
	.w7(32'h3a5788a2),
	.w8(32'h3cb40352),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8ad17),
	.w1(32'hbbdbcb43),
	.w2(32'h3bf5e700),
	.w3(32'h3c6d724a),
	.w4(32'h3b4b1403),
	.w5(32'h3c8d315d),
	.w6(32'hbbc14461),
	.w7(32'hbc11edf0),
	.w8(32'h3b41c144),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb504e0a),
	.w1(32'h3a254e68),
	.w2(32'h3b6254a4),
	.w3(32'h3ce95315),
	.w4(32'h3c7d4f8d),
	.w5(32'hbac696e2),
	.w6(32'hbbf83a84),
	.w7(32'hbb2a42a6),
	.w8(32'h3999d0ca),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c0e9b),
	.w1(32'hbb6d2044),
	.w2(32'hbb1ad0d2),
	.w3(32'h3b4b695d),
	.w4(32'h3ab3b9ef),
	.w5(32'h3b0c09ad),
	.w6(32'h3bac199b),
	.w7(32'hbb90869f),
	.w8(32'hbb861745),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a840c25),
	.w1(32'h3a29b113),
	.w2(32'hb5a7d590),
	.w3(32'hbc13139e),
	.w4(32'h3a9e9444),
	.w5(32'h3b606525),
	.w6(32'h3ae3fd9e),
	.w7(32'h3a351d81),
	.w8(32'h3ae70fbd),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199c55),
	.w1(32'hbb2fb186),
	.w2(32'hbb58f632),
	.w3(32'h3b6b54f5),
	.w4(32'hbb59fc70),
	.w5(32'hba8d6f30),
	.w6(32'h3c6df0c6),
	.w7(32'h3a74c737),
	.w8(32'hbbf24618),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0508fa),
	.w1(32'h39b0b5cb),
	.w2(32'hbb19bc23),
	.w3(32'h3c08d815),
	.w4(32'h3b48104d),
	.w5(32'h3ba12155),
	.w6(32'h3cbccbe2),
	.w7(32'h3b35d621),
	.w8(32'hbb3ede94),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0541be),
	.w1(32'h3bc621ac),
	.w2(32'h3b143596),
	.w3(32'hbc4f0723),
	.w4(32'hbb07c101),
	.w5(32'hbb9fa43b),
	.w6(32'hbc7425bd),
	.w7(32'hba0c021e),
	.w8(32'h3ab79234),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86065e),
	.w1(32'hb99a8872),
	.w2(32'hb8b09f6d),
	.w3(32'hbbe97c4c),
	.w4(32'hbb058042),
	.w5(32'h3b2d437a),
	.w6(32'h3b5cf248),
	.w7(32'hbb2f3873),
	.w8(32'hbaaad6f1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f6505),
	.w1(32'hbbcba7ba),
	.w2(32'hbc231dc6),
	.w3(32'hbc43e903),
	.w4(32'hbb53e73c),
	.w5(32'hbb44bc18),
	.w6(32'h3a594ef8),
	.w7(32'hbba5030d),
	.w8(32'h3b075c4e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2210f),
	.w1(32'hbb2389a1),
	.w2(32'hbb930d3e),
	.w3(32'hbc20d502),
	.w4(32'hbb9b3d01),
	.w5(32'hba0d0585),
	.w6(32'hbb875db9),
	.w7(32'hbba64a96),
	.w8(32'hbb38a169),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951eaff),
	.w1(32'hbb7e9177),
	.w2(32'hbadd7920),
	.w3(32'h3bf9bcee),
	.w4(32'hbae42ecd),
	.w5(32'h3b92a25a),
	.w6(32'h3bca0d77),
	.w7(32'h37ee001a),
	.w8(32'hbbe4d88b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9883e78),
	.w1(32'hbab5a2d9),
	.w2(32'hb97cc5aa),
	.w3(32'hbb1c4817),
	.w4(32'hba5108bd),
	.w5(32'hba7a27fd),
	.w6(32'hbba73059),
	.w7(32'hbb58fa64),
	.w8(32'h3aa567de),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafaefeb),
	.w1(32'hb81e6c5e),
	.w2(32'hba477ecf),
	.w3(32'hbb5c2459),
	.w4(32'hbb0fdecb),
	.w5(32'h3b715101),
	.w6(32'h3b0e5d51),
	.w7(32'h3b2dc23e),
	.w8(32'hbac991d4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76e2a7),
	.w1(32'hbada3767),
	.w2(32'hba546eed),
	.w3(32'h3af2b0c6),
	.w4(32'h3ab206c7),
	.w5(32'h3ae67926),
	.w6(32'hbb772198),
	.w7(32'hbb3ee043),
	.w8(32'hbbf32e67),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb215475),
	.w1(32'h3b881eaa),
	.w2(32'h3ae44e1c),
	.w3(32'hbb1b6819),
	.w4(32'h3abf78db),
	.w5(32'h3bd05001),
	.w6(32'hbb2d655b),
	.w7(32'hba4ac036),
	.w8(32'h3bfb3341),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0d88),
	.w1(32'h3acc1c39),
	.w2(32'hb7571bd2),
	.w3(32'hbc095071),
	.w4(32'hbb57f21c),
	.w5(32'hbc4ca3f4),
	.w6(32'hbbcab42c),
	.w7(32'hbb054603),
	.w8(32'hbbacf348),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07be2c),
	.w1(32'hba469c96),
	.w2(32'hbb06c843),
	.w3(32'hbadb9bb7),
	.w4(32'hba7c000a),
	.w5(32'h3a67eb41),
	.w6(32'hbbc2f61b),
	.w7(32'hbbaeae33),
	.w8(32'h3b1b52d5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c330d),
	.w1(32'h3bae3b19),
	.w2(32'h3b95ff0d),
	.w3(32'h395d7d24),
	.w4(32'h3a65e056),
	.w5(32'hbc1ef9b2),
	.w6(32'hbbb2e41a),
	.w7(32'hba352202),
	.w8(32'hbac73179),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf394bd),
	.w1(32'hbbac533a),
	.w2(32'hbba17daf),
	.w3(32'hbb3d9b8a),
	.w4(32'h39ff1dc7),
	.w5(32'h3b4e0c08),
	.w6(32'h3c99f57c),
	.w7(32'h3b151d68),
	.w8(32'hbbd26db9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80a5e2),
	.w1(32'h3b85e24e),
	.w2(32'hba425e80),
	.w3(32'hbc88eed3),
	.w4(32'hbb027658),
	.w5(32'h3af43ebf),
	.w6(32'hbb94bda3),
	.w7(32'hbb489dde),
	.w8(32'h3b960073),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c046ebc),
	.w1(32'hbc2058a6),
	.w2(32'hbc649d20),
	.w3(32'hbb9d3dc3),
	.w4(32'hbc73d614),
	.w5(32'hbc2dea82),
	.w6(32'h3c038f02),
	.w7(32'h3ae85b1e),
	.w8(32'hbbc6cc0d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc498d53),
	.w1(32'hba8a28c0),
	.w2(32'hbadf488f),
	.w3(32'hbc62d16a),
	.w4(32'hbc167664),
	.w5(32'hbb469df4),
	.w6(32'hbc1dcf7b),
	.w7(32'hba10983b),
	.w8(32'hb9525182),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39e8f3),
	.w1(32'hbba20dfc),
	.w2(32'h3b0911e7),
	.w3(32'hbc47c915),
	.w4(32'hba08bfac),
	.w5(32'hba26b9bc),
	.w6(32'h3996e634),
	.w7(32'hbb55847c),
	.w8(32'hbb4d0e67),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8156c1),
	.w1(32'hbc044eb6),
	.w2(32'hbb6361de),
	.w3(32'hbc771970),
	.w4(32'hbc12b265),
	.w5(32'hbb868ea2),
	.w6(32'hbbb72777),
	.w7(32'hbc0fe595),
	.w8(32'hbaa74a79),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1103fe),
	.w1(32'h3b8fa512),
	.w2(32'h3a0c8a43),
	.w3(32'hbc838525),
	.w4(32'h3bbefd44),
	.w5(32'h38767bcf),
	.w6(32'hbc7c37a2),
	.w7(32'h395d2bc7),
	.w8(32'h3c5cbe40),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b338237),
	.w1(32'h3b3c370b),
	.w2(32'hbaa17747),
	.w3(32'hbb179120),
	.w4(32'hbb36c15c),
	.w5(32'hbb8232da),
	.w6(32'h39a16bdd),
	.w7(32'hbb567c69),
	.w8(32'hba4b2ed2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8378c1),
	.w1(32'hbbccc5c2),
	.w2(32'h3b890361),
	.w3(32'hbbb15b62),
	.w4(32'hbbc7e5b1),
	.w5(32'hbc05c85c),
	.w6(32'h3ba319e9),
	.w7(32'h39a48a81),
	.w8(32'hbc439f8b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca99660),
	.w1(32'hbc440d50),
	.w2(32'hbcb529fe),
	.w3(32'hbc4f34ce),
	.w4(32'hbca7d0c4),
	.w5(32'h3c394ebb),
	.w6(32'h3c0205aa),
	.w7(32'hbc041be8),
	.w8(32'hbc1cf5a9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca22e74),
	.w1(32'hbd1b1d6a),
	.w2(32'h3ccb7df6),
	.w3(32'h3d93ed0b),
	.w4(32'h3b8af670),
	.w5(32'h3c5c2a56),
	.w6(32'hbb05a37b),
	.w7(32'h3ca603aa),
	.w8(32'hb9deded8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f9830),
	.w1(32'h3b219fcc),
	.w2(32'hbbd84aac),
	.w3(32'hbc2cb138),
	.w4(32'h3c456048),
	.w5(32'h3b88224d),
	.w6(32'hbc44f40b),
	.w7(32'h3c6b7bbf),
	.w8(32'h3c6869a2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcbc51),
	.w1(32'hbbd0fb63),
	.w2(32'hbba18696),
	.w3(32'hb9e73e69),
	.w4(32'hbc091fa2),
	.w5(32'hbbcbc64d),
	.w6(32'hbced02e2),
	.w7(32'hbca2fb9d),
	.w8(32'h3b9f2ca5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a0666),
	.w1(32'hbc6682c2),
	.w2(32'hbb977ff1),
	.w3(32'hbb9e7ff2),
	.w4(32'hbcbd010f),
	.w5(32'h3c803870),
	.w6(32'h3bf4cb1a),
	.w7(32'hbc02ce06),
	.w8(32'hbcfbac5a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3725cd),
	.w1(32'hbc933316),
	.w2(32'hbbe32833),
	.w3(32'h3d678a96),
	.w4(32'h3d14f4b4),
	.w5(32'h3b2959d2),
	.w6(32'hba37bb4a),
	.w7(32'hba164f6b),
	.w8(32'hbc33df61),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d315dc1),
	.w1(32'h3b5d1453),
	.w2(32'hbc201b62),
	.w3(32'h3acb9d5c),
	.w4(32'hbcc8fdf3),
	.w5(32'h3ce97f00),
	.w6(32'h3c48ce48),
	.w7(32'hbc959824),
	.w8(32'h3a19e4bc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42e3f2),
	.w1(32'hbcfef192),
	.w2(32'hbccb350b),
	.w3(32'h3d1deecd),
	.w4(32'h3cbaf0e3),
	.w5(32'h3ab8c807),
	.w6(32'h3b65bfb2),
	.w7(32'h3b9c0acb),
	.w8(32'hbb350cc0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0e02d),
	.w1(32'hbc722b41),
	.w2(32'h3b1ab5c1),
	.w3(32'h3c688694),
	.w4(32'h3c572607),
	.w5(32'hb9cbbe24),
	.w6(32'hbcd87260),
	.w7(32'hba48798c),
	.w8(32'h3bb199f9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b020de9),
	.w1(32'hbc18895e),
	.w2(32'h3adb0bcd),
	.w3(32'hbc06268c),
	.w4(32'hbc14a192),
	.w5(32'hbc1d49d5),
	.w6(32'hbb9ad4d3),
	.w7(32'hb95d0897),
	.w8(32'hba5bab65),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5124c),
	.w1(32'hbc1d796f),
	.w2(32'hbbbb99e3),
	.w3(32'hbc221a52),
	.w4(32'hbc41b819),
	.w5(32'hbd0f582c),
	.w6(32'h3ab1d9aa),
	.w7(32'hbbbd5a1a),
	.w8(32'hbc153222),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c8bc7),
	.w1(32'h3c98a486),
	.w2(32'h3bc05dba),
	.w3(32'hbd5036be),
	.w4(32'hbd1aaf86),
	.w5(32'h3b82fc63),
	.w6(32'hbcc791f7),
	.w7(32'hbc571094),
	.w8(32'h3c20b0bd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb356154),
	.w1(32'h3c20fc9f),
	.w2(32'h3ba3810e),
	.w3(32'hbb883929),
	.w4(32'h36b03a94),
	.w5(32'h3bb178f3),
	.w6(32'hbaf7d344),
	.w7(32'h3c27529d),
	.w8(32'h3c4068b3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba2b85),
	.w1(32'hbaeed08d),
	.w2(32'hbb3a6019),
	.w3(32'hbc165d95),
	.w4(32'hbc1d0add),
	.w5(32'hbc944bd5),
	.w6(32'hbbabd060),
	.w7(32'hbb5bff06),
	.w8(32'h39b4bb04),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c107e72),
	.w1(32'h3cd4c3a6),
	.w2(32'h3ba81cb1),
	.w3(32'hbc5cd529),
	.w4(32'hbc5a3091),
	.w5(32'hbc128173),
	.w6(32'h3bdc4046),
	.w7(32'hb9e8b7c7),
	.w8(32'hbc1fc0c5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc886020),
	.w1(32'hbc15e2b8),
	.w2(32'h3b5cf322),
	.w3(32'hbc14085e),
	.w4(32'hbb096ff8),
	.w5(32'h3c876443),
	.w6(32'hbc18d68d),
	.w7(32'hbc14360f),
	.w8(32'h3849c5cc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ade3),
	.w1(32'hbc60d4d8),
	.w2(32'hbbcbc981),
	.w3(32'h3ba91d25),
	.w4(32'h3c593279),
	.w5(32'h3c41875d),
	.w6(32'hbc997bca),
	.w7(32'hbb675a13),
	.w8(32'h3bb23395),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb238458),
	.w1(32'hbbbe03aa),
	.w2(32'hbb64015b),
	.w3(32'h3c2827c9),
	.w4(32'hbba3c0a0),
	.w5(32'hbc912ff2),
	.w6(32'h3aa8a29b),
	.w7(32'hbb88984d),
	.w8(32'h3b4c797f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0de59a),
	.w1(32'h3c416af9),
	.w2(32'h3bc538a1),
	.w3(32'hbcb63550),
	.w4(32'hbcd40f42),
	.w5(32'hbc316c77),
	.w6(32'hb81c3107),
	.w7(32'hbbb01400),
	.w8(32'hbc005b49),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4000f),
	.w1(32'hbc10aee5),
	.w2(32'hbc03fb9d),
	.w3(32'h3b9e7e8c),
	.w4(32'h3bf43b25),
	.w5(32'hbb020d2e),
	.w6(32'hb9c41f33),
	.w7(32'hbbe3090e),
	.w8(32'hbb9e9b87),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a4d15),
	.w1(32'hbc5c514c),
	.w2(32'hbb953a22),
	.w3(32'hbc3a1078),
	.w4(32'hbb88dafb),
	.w5(32'h3bbb9ee8),
	.w6(32'hbc5a450b),
	.w7(32'hbbcac897),
	.w8(32'hbc6a8c87),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a7ee7),
	.w1(32'hbd2675a4),
	.w2(32'hbcdf93d1),
	.w3(32'h3ca2b696),
	.w4(32'h3c0639ea),
	.w5(32'h3a58f86e),
	.w6(32'hbced8613),
	.w7(32'hbc8b8a5a),
	.w8(32'h3aa56e6d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3773d7),
	.w1(32'hbc42da11),
	.w2(32'hbc4b0158),
	.w3(32'h3af066cf),
	.w4(32'hbba7f673),
	.w5(32'h3bbbdb3a),
	.w6(32'h3b2172dd),
	.w7(32'h3a563b08),
	.w8(32'hba079a2c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc83312),
	.w1(32'h3bd47b82),
	.w2(32'h3b9a0651),
	.w3(32'h3ade3184),
	.w4(32'hbc0c1107),
	.w5(32'h3c1d944d),
	.w6(32'h3cb86634),
	.w7(32'h3c43493e),
	.w8(32'h3b35aa53),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bef70),
	.w1(32'h3c827e49),
	.w2(32'h3c19b23d),
	.w3(32'hbbe227aa),
	.w4(32'h3c51cc78),
	.w5(32'hbbc48906),
	.w6(32'hbcbe3cf2),
	.w7(32'hbb8ef343),
	.w8(32'h3c376773),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b605828),
	.w1(32'h3c52bcb3),
	.w2(32'h3a7b8d26),
	.w3(32'hb928b589),
	.w4(32'h3bbbdeda),
	.w5(32'h3b8d2eb7),
	.w6(32'hba49d20d),
	.w7(32'h3b8418e0),
	.w8(32'h3b9af3d2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7a133),
	.w1(32'h3c2282a4),
	.w2(32'h3bf19244),
	.w3(32'h3a3d54d5),
	.w4(32'h3b66cf6c),
	.w5(32'h3982a680),
	.w6(32'hbc0d0895),
	.w7(32'hbb22b887),
	.w8(32'hbbe95142),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c6a3f),
	.w1(32'hbb3f03f0),
	.w2(32'hbaac5425),
	.w3(32'h3b32c024),
	.w4(32'h3b3cd522),
	.w5(32'hbc3fe8f6),
	.w6(32'h3b35ffec),
	.w7(32'hb98544eb),
	.w8(32'h3bb53911),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8279bf),
	.w1(32'h3c15e6b4),
	.w2(32'hbb1f8016),
	.w3(32'hbcbca5b5),
	.w4(32'hbc44821b),
	.w5(32'h3c2a06a7),
	.w6(32'hbab755b2),
	.w7(32'hbbf69a49),
	.w8(32'hbb0625ee),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc621581),
	.w1(32'hbcea57e1),
	.w2(32'h3c4861a5),
	.w3(32'h3d045555),
	.w4(32'h3c835418),
	.w5(32'hbba3f373),
	.w6(32'hbbf983ac),
	.w7(32'h3c607dc9),
	.w8(32'hbb6fad45),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a322cf2),
	.w1(32'h3b606a17),
	.w2(32'hbbc19327),
	.w3(32'hbc82c436),
	.w4(32'hbca73080),
	.w5(32'h3c1502e7),
	.w6(32'h3c784d3b),
	.w7(32'hbc038836),
	.w8(32'h3b5feca2),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c148ecd),
	.w1(32'h3c531d40),
	.w2(32'h3bc004e6),
	.w3(32'hbaef0f92),
	.w4(32'h3bd1fba3),
	.w5(32'h3c697abd),
	.w6(32'h3c0ae075),
	.w7(32'hbb83b93b),
	.w8(32'hbb3425d9),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2907cd),
	.w1(32'hbb7c12a3),
	.w2(32'h3aeb4570),
	.w3(32'h3b42ae73),
	.w4(32'h3a3e6c46),
	.w5(32'hbb554574),
	.w6(32'hbc3daa4f),
	.w7(32'hbb67aa34),
	.w8(32'h3befe76d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc50b33),
	.w1(32'h3c53630d),
	.w2(32'h3a767890),
	.w3(32'hbc60b847),
	.w4(32'hbbcabec7),
	.w5(32'hbc59addd),
	.w6(32'h3b9902eb),
	.w7(32'hba800854),
	.w8(32'hbd10de31),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc071b24),
	.w1(32'h3bad2b48),
	.w2(32'h3c3a7d1b),
	.w3(32'h3c72ea26),
	.w4(32'h3c43210d),
	.w5(32'hbc88186b),
	.w6(32'hbccb4c76),
	.w7(32'hbc91e9ed),
	.w8(32'h3b34b059),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c424768),
	.w1(32'h3cf8ffe7),
	.w2(32'h3c471b7d),
	.w3(32'hbd231862),
	.w4(32'hbce60d00),
	.w5(32'hbc081edb),
	.w6(32'hbbd0d949),
	.w7(32'hbb966c8a),
	.w8(32'h3c1b6540),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64377b),
	.w1(32'h3c353cbd),
	.w2(32'h3c15b0ad),
	.w3(32'hbc8a8ff2),
	.w4(32'hbc888dd4),
	.w5(32'hbc35e8ee),
	.w6(32'h3cc7070d),
	.w7(32'h3b60a94c),
	.w8(32'hbc9089c2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae85f6a),
	.w1(32'h3c1db738),
	.w2(32'h3bc4751a),
	.w3(32'hbcd5a5c9),
	.w4(32'hbcf087f2),
	.w5(32'hbc87b167),
	.w6(32'hbc0e30e5),
	.w7(32'h3b456f65),
	.w8(32'h3c0482f9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca31a96),
	.w1(32'h3cd28b32),
	.w2(32'h3c4c7137),
	.w3(32'hbcf6d889),
	.w4(32'hbd003314),
	.w5(32'hbcb6382d),
	.w6(32'hbba492f0),
	.w7(32'hbbedeb52),
	.w8(32'hbbadc36e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e8fb6),
	.w1(32'h3bc4f9c6),
	.w2(32'h3b37aab6),
	.w3(32'hbcdf2591),
	.w4(32'hbd1461ac),
	.w5(32'hbb51325a),
	.w6(32'h3b98e5d9),
	.w7(32'hbc351101),
	.w8(32'hba8597ea),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcbc8b),
	.w1(32'h3c986fb6),
	.w2(32'h3bb68199),
	.w3(32'hbc31607b),
	.w4(32'hbc77f8cf),
	.w5(32'h3ba3f7ca),
	.w6(32'h3c2e4241),
	.w7(32'h3ba5a83c),
	.w8(32'hbc0656aa),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17dd22),
	.w1(32'hbc879a03),
	.w2(32'hbc29769c),
	.w3(32'h3bc6e672),
	.w4(32'hb95724eb),
	.w5(32'h3bc1fee7),
	.w6(32'hbc79dd99),
	.w7(32'hbc0fc01a),
	.w8(32'hbcb4ca0b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca186ed),
	.w1(32'h3a845060),
	.w2(32'hbc118f50),
	.w3(32'h3ce215e6),
	.w4(32'h3c890784),
	.w5(32'h3b0c4e12),
	.w6(32'hbaabccc0),
	.w7(32'hbb58dc9a),
	.w8(32'hba5f2657),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1cf49),
	.w1(32'h3bab5f9a),
	.w2(32'hbaf3aa97),
	.w3(32'hbc52ce20),
	.w4(32'h3c6dedbc),
	.w5(32'h3c1a0125),
	.w6(32'hbc958e56),
	.w7(32'h3c13b642),
	.w8(32'h3ca1bc3b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01987e),
	.w1(32'h3c8ca039),
	.w2(32'h3c3c407c),
	.w3(32'hbbe42cce),
	.w4(32'hbb2de8e5),
	.w5(32'hbba01dd2),
	.w6(32'h3c48aae6),
	.w7(32'h3c397f01),
	.w8(32'hba3b1007),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6049c7),
	.w1(32'h3c1b32af),
	.w2(32'h3ba3fc0e),
	.w3(32'hbc501bed),
	.w4(32'h3a27aac5),
	.w5(32'hbbe5e40e),
	.w6(32'h3b8178c4),
	.w7(32'h392695d2),
	.w8(32'h3b6d863d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c055757),
	.w1(32'h3c934aa5),
	.w2(32'h3c294da5),
	.w3(32'hbc8dea5a),
	.w4(32'hbc9aa003),
	.w5(32'h3c1a1ab2),
	.w6(32'hb9c7f1be),
	.w7(32'hbb0bf2b9),
	.w8(32'hbbb1cb0f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f1878),
	.w1(32'hbc620b0c),
	.w2(32'hbc28fcab),
	.w3(32'h3c798de6),
	.w4(32'h3c9b94b5),
	.w5(32'hbbd5a1ac),
	.w6(32'hbb7bfd2c),
	.w7(32'h3b00f31f),
	.w8(32'hbc5ae3ff),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02245d),
	.w1(32'hbc3c23e0),
	.w2(32'hbc647ab6),
	.w3(32'h3ab6f8f0),
	.w4(32'hba759f84),
	.w5(32'hbbf7ac42),
	.w6(32'hbc65367b),
	.w7(32'hbc6b0b15),
	.w8(32'hbbc06f84),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ddd74),
	.w1(32'h3ae10fc9),
	.w2(32'hbbcb1ed5),
	.w3(32'hbb4c02eb),
	.w4(32'hba9b0629),
	.w5(32'hbb28a8a3),
	.w6(32'hba17a7e2),
	.w7(32'hbc08aa43),
	.w8(32'hbb8cf841),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a9cd7),
	.w1(32'h3bbd0c23),
	.w2(32'h3bdeeeba),
	.w3(32'h3b911b2a),
	.w4(32'h3bc6ecdc),
	.w5(32'hbc2044c8),
	.w6(32'h3bc940ba),
	.w7(32'h3bb17b06),
	.w8(32'h3bbf6dc1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca19855),
	.w1(32'h3c7a61a4),
	.w2(32'h3bdc36cd),
	.w3(32'hbcc73da4),
	.w4(32'hbce3d4f4),
	.w5(32'hba375cc3),
	.w6(32'h3c476ccd),
	.w7(32'hbb1bd342),
	.w8(32'h3b3fe8bc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0e4a9),
	.w1(32'hbaa72295),
	.w2(32'h39a0c644),
	.w3(32'h3b9962d1),
	.w4(32'h3bddb7ba),
	.w5(32'hbba188fc),
	.w6(32'h3b9f9927),
	.w7(32'h3b824b9d),
	.w8(32'h3ba601e6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8862cd),
	.w1(32'h3b5888cb),
	.w2(32'hbab27245),
	.w3(32'h3abe8c3c),
	.w4(32'hbb582198),
	.w5(32'hbb810980),
	.w6(32'h3ca46f4a),
	.w7(32'h3ba8c9c2),
	.w8(32'hbba8813a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53575d),
	.w1(32'h3b558a38),
	.w2(32'hbc67a108),
	.w3(32'hbc05b4a0),
	.w4(32'hbc1454aa),
	.w5(32'hbc20b962),
	.w6(32'hbcbceeba),
	.w7(32'hbc2a5e51),
	.w8(32'h3bba200a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8744a),
	.w1(32'h3beb9e93),
	.w2(32'h3bab2975),
	.w3(32'hbc7f5e9b),
	.w4(32'hbc9833e3),
	.w5(32'hbbc19395),
	.w6(32'h3b71c222),
	.w7(32'hbaf7f1b1),
	.w8(32'h3c0fbc60),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20714a),
	.w1(32'hba7306fc),
	.w2(32'h3acdb611),
	.w3(32'hbc5a6c4a),
	.w4(32'hbb7f686b),
	.w5(32'hbcd24314),
	.w6(32'h3b851720),
	.w7(32'hb8c32eb9),
	.w8(32'hbbc6c005),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a9fe2),
	.w1(32'h3ca0c960),
	.w2(32'h3b8691fb),
	.w3(32'hbd1e60ab),
	.w4(32'hbd0d9a7a),
	.w5(32'hbc7c4d3e),
	.w6(32'hbcae1146),
	.w7(32'hbc9878ba),
	.w8(32'hbc0f7fe5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb91ee3),
	.w1(32'hba83844b),
	.w2(32'hb94764ff),
	.w3(32'hbc0f03bb),
	.w4(32'h3c5390ca),
	.w5(32'hbbb80c62),
	.w6(32'hbc571f42),
	.w7(32'h3b51c140),
	.w8(32'hbb2f6953),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba810462),
	.w1(32'h3b96e199),
	.w2(32'h3b736fc4),
	.w3(32'hbb9105e7),
	.w4(32'hbbac5b4a),
	.w5(32'hbc1981ee),
	.w6(32'hbb035cc8),
	.w7(32'h3c072bfb),
	.w8(32'hba70e51c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50a229),
	.w1(32'hbca1911e),
	.w2(32'hbc1d4caa),
	.w3(32'hbb8f10de),
	.w4(32'hbc515b11),
	.w5(32'h3ba86b3c),
	.w6(32'hbae2fcd5),
	.w7(32'hbc61ff3b),
	.w8(32'hbc1beb8e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc538c98),
	.w1(32'hbb364f86),
	.w2(32'hbc75433e),
	.w3(32'h3ada1507),
	.w4(32'h3a182d4a),
	.w5(32'h3bd8d678),
	.w6(32'hbcbad3a1),
	.w7(32'hbba741e0),
	.w8(32'hbb59ec43),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88f3f9),
	.w1(32'hbc1f8cb4),
	.w2(32'h3b9f95e3),
	.w3(32'h3beba222),
	.w4(32'hbc4cb6cf),
	.w5(32'h3befef02),
	.w6(32'h3c1fe555),
	.w7(32'hbb81c92e),
	.w8(32'hbc6389c2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d9d04),
	.w1(32'hbcc20c8f),
	.w2(32'hbc81c694),
	.w3(32'h3ca03175),
	.w4(32'h3c4aa7d0),
	.w5(32'h3b80f25e),
	.w6(32'hbc173203),
	.w7(32'hba5ec821),
	.w8(32'h3b3ac576),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5787),
	.w1(32'h3bdf8e2c),
	.w2(32'hbb834e60),
	.w3(32'h3b60564f),
	.w4(32'h3c41c2fe),
	.w5(32'h3bf14e4c),
	.w6(32'hbbb7a726),
	.w7(32'hba12f6fe),
	.w8(32'h3c0ec381),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe03a92),
	.w1(32'hbc848469),
	.w2(32'hbbe5aee2),
	.w3(32'h3c9f58cb),
	.w4(32'h3c2d3fc8),
	.w5(32'hbb5e33f2),
	.w6(32'hbaeee6ef),
	.w7(32'h3aadcb51),
	.w8(32'hbc2edca1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc960a22),
	.w1(32'hbcd18dfa),
	.w2(32'hbc6991af),
	.w3(32'hbb2b35f6),
	.w4(32'h3ad9d6d9),
	.w5(32'hbbc5b9da),
	.w6(32'hbb336c35),
	.w7(32'hbc18ea6e),
	.w8(32'h3c1ae370),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88aaec),
	.w1(32'h3ca91dca),
	.w2(32'h3c1f8da1),
	.w3(32'hbc94d0cf),
	.w4(32'hbca17a79),
	.w5(32'h3c354e0c),
	.w6(32'h3c9047da),
	.w7(32'hba8b653e),
	.w8(32'h3ba06881),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0be7f8),
	.w1(32'h3c5135bb),
	.w2(32'h3bb87dee),
	.w3(32'h3b970191),
	.w4(32'h3abf7461),
	.w5(32'hbc717887),
	.w6(32'h3a02fd0a),
	.w7(32'h3ae8916b),
	.w8(32'hba05ecee),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5266b4),
	.w1(32'h3c96b870),
	.w2(32'h3bb1e591),
	.w3(32'hbc4a80ee),
	.w4(32'hbca4aa25),
	.w5(32'h3b86402c),
	.w6(32'h3c2231d7),
	.w7(32'hbc070bfd),
	.w8(32'h3b6cb7a3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad33a90),
	.w1(32'hbc0adcaf),
	.w2(32'hbc19a4b5),
	.w3(32'h3cbdf976),
	.w4(32'h3c0c6b40),
	.w5(32'hbb3760cd),
	.w6(32'h3c934f84),
	.w7(32'h3c0435ef),
	.w8(32'h3ba67c40),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50b8b9),
	.w1(32'h3b43b11a),
	.w2(32'hbb2f4097),
	.w3(32'hbc88b4a2),
	.w4(32'hbc246d51),
	.w5(32'h3c11bc95),
	.w6(32'h3c00e345),
	.w7(32'h3a064863),
	.w8(32'hbb1df043),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ef055),
	.w1(32'hbc3297b0),
	.w2(32'hbc598b74),
	.w3(32'h3c19226a),
	.w4(32'h3c6c59d5),
	.w5(32'h3c30e756),
	.w6(32'hbc11f838),
	.w7(32'hbbd1e0ab),
	.w8(32'h3c5be98f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092ab5),
	.w1(32'h3c1568dd),
	.w2(32'h3c2b8fe2),
	.w3(32'hbc10c047),
	.w4(32'h3c108da4),
	.w5(32'h39d9b5ce),
	.w6(32'hbb9c06eb),
	.w7(32'h3beb99e7),
	.w8(32'hbb516ca3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4a2c6),
	.w1(32'hbc489088),
	.w2(32'hbbeba196),
	.w3(32'hbaf1c396),
	.w4(32'hbac78b85),
	.w5(32'h3bbd13a9),
	.w6(32'hbbbc592e),
	.w7(32'hbb32e5f6),
	.w8(32'hbbbad598),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0135d5),
	.w1(32'hbc476f20),
	.w2(32'hbbd514e7),
	.w3(32'hbba83f66),
	.w4(32'hbb16de3a),
	.w5(32'h3c843580),
	.w6(32'h3a24148c),
	.w7(32'hbb73e13e),
	.w8(32'h3bbda7b0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4afd),
	.w1(32'hbc8e4fd6),
	.w2(32'hb956c607),
	.w3(32'h3c8a6f36),
	.w4(32'h3c5a3a51),
	.w5(32'hbca201b3),
	.w6(32'h3b5be6b4),
	.w7(32'hba6c3fbf),
	.w8(32'hbbc1b5a8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb55ba2),
	.w1(32'h3d14cc67),
	.w2(32'h3c5a4db0),
	.w3(32'hbd10394e),
	.w4(32'hbcfdb5d8),
	.w5(32'hbbc0dd6f),
	.w6(32'h3b8ad45f),
	.w7(32'hbbf3ccd4),
	.w8(32'hbbbbf6e1),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81f5d7),
	.w1(32'hbb06edc3),
	.w2(32'hbc12fbb6),
	.w3(32'hbbe84bd2),
	.w4(32'h3c1920ad),
	.w5(32'hbc31dab3),
	.w6(32'h3b93abbd),
	.w7(32'h3ba0af55),
	.w8(32'h3b2ccc03),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca65130),
	.w1(32'h3cac979c),
	.w2(32'h3bfa4cb1),
	.w3(32'hbca65d24),
	.w4(32'hbcdee42f),
	.w5(32'h3b37f801),
	.w6(32'h3c2f30d5),
	.w7(32'hbb90e21b),
	.w8(32'hbb29b078),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ee85d),
	.w1(32'hbaee82f0),
	.w2(32'h3b64a82d),
	.w3(32'h3c6e7032),
	.w4(32'hbc16346e),
	.w5(32'h3bc21418),
	.w6(32'h390e4738),
	.w7(32'hbc2013ff),
	.w8(32'hbafa6f03),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc093c0b),
	.w1(32'hbbdd042f),
	.w2(32'hbb8f49bd),
	.w3(32'h3c43ad62),
	.w4(32'h3c290f25),
	.w5(32'h3ba0a77d),
	.w6(32'hbbade891),
	.w7(32'hbbaf009f),
	.w8(32'h3bcef3f8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4cfc2),
	.w1(32'hbbad47ec),
	.w2(32'h3b12bd93),
	.w3(32'hbb7b7b4e),
	.w4(32'hbb86edcd),
	.w5(32'hbbecf39f),
	.w6(32'h3befb7ce),
	.w7(32'h3b95c085),
	.w8(32'hbc11a069),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe438f6),
	.w1(32'hbc4379c4),
	.w2(32'hbc2b6f3b),
	.w3(32'hbb64933f),
	.w4(32'h3c7b9c3e),
	.w5(32'h3bb3a40c),
	.w6(32'h3b955872),
	.w7(32'hbb20792d),
	.w8(32'hbbd4a315),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05582c),
	.w1(32'hba83a485),
	.w2(32'hbb7f156b),
	.w3(32'h3c08bb6b),
	.w4(32'h3c2a3f12),
	.w5(32'hbbd7d2d5),
	.w6(32'hbb86d96b),
	.w7(32'hba13adaa),
	.w8(32'hbb9fb51d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0b67),
	.w1(32'h3b373fc8),
	.w2(32'hbbb613c1),
	.w3(32'h3a21c308),
	.w4(32'h3bcc8a33),
	.w5(32'hbc3c20f8),
	.w6(32'hbc48a0fb),
	.w7(32'hbbfbb79f),
	.w8(32'hbb6cdeb0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9ecd3),
	.w1(32'hbc75565d),
	.w2(32'hbc305d04),
	.w3(32'hbba6627c),
	.w4(32'hbc319db1),
	.w5(32'hbc1103e3),
	.w6(32'hbc731f64),
	.w7(32'hbc7a875f),
	.w8(32'hbc7858e6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6ab40),
	.w1(32'h3bc341a1),
	.w2(32'hbc184847),
	.w3(32'h3bf8af10),
	.w4(32'hbadb58cd),
	.w5(32'hbc65be70),
	.w6(32'h3c91e476),
	.w7(32'h3c0730d1),
	.w8(32'h3be5f473),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c990c19),
	.w1(32'h3c9f9db1),
	.w2(32'h3bd5c0c1),
	.w3(32'hbc9acbca),
	.w4(32'hbcbded25),
	.w5(32'hbb809a01),
	.w6(32'h3c50b3b0),
	.w7(32'hbaf8adfd),
	.w8(32'hbb5acdce),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4560c9),
	.w1(32'hbc074b8a),
	.w2(32'h3aaeb89d),
	.w3(32'h3c25db76),
	.w4(32'hbc97d0f6),
	.w5(32'h3a4f5b72),
	.w6(32'h3c72b0ac),
	.w7(32'hbbcfb047),
	.w8(32'hbbf3f180),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd42a6d),
	.w1(32'h3cbbfde0),
	.w2(32'hb9123b28),
	.w3(32'hbd02cebc),
	.w4(32'hbc36bbf7),
	.w5(32'hbc81e112),
	.w6(32'hbba9cf53),
	.w7(32'hbb83658e),
	.w8(32'h3c30eccb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a3b6d),
	.w1(32'h3c28e8a7),
	.w2(32'hbbcf34a7),
	.w3(32'hbc6c7c2b),
	.w4(32'hbc0f0a13),
	.w5(32'hbad7bd55),
	.w6(32'h3c2fbacb),
	.w7(32'h3b5c9bc1),
	.w8(32'hbc1fe850),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf59a3),
	.w1(32'hbc0486ac),
	.w2(32'hbc08f72f),
	.w3(32'h3c45567c),
	.w4(32'h3b73d8a9),
	.w5(32'hbb19075b),
	.w6(32'hbbeffe9c),
	.w7(32'hbbf621a9),
	.w8(32'h3b0d39eb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c6299),
	.w1(32'h3b05b24e),
	.w2(32'hba8f065f),
	.w3(32'h3c3a809f),
	.w4(32'h3c81c70d),
	.w5(32'h3ad7fc66),
	.w6(32'h3bc811af),
	.w7(32'h3b41f626),
	.w8(32'hbb3e2211),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98cb77),
	.w1(32'h3a43bf81),
	.w2(32'hbbb1670b),
	.w3(32'h3ba95287),
	.w4(32'h3bf17ca7),
	.w5(32'h3b8a9117),
	.w6(32'hb8eb6d7c),
	.w7(32'h3b27bf1b),
	.w8(32'hbaf7a04a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb5152),
	.w1(32'hbca0ac2b),
	.w2(32'hbc2207b0),
	.w3(32'h3c99f223),
	.w4(32'hbab57405),
	.w5(32'hbb6ecdfc),
	.w6(32'hbb884f75),
	.w7(32'hbba8bcc2),
	.w8(32'hba3f5578),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4cfa),
	.w1(32'h3c78ed02),
	.w2(32'h3c5749ab),
	.w3(32'hbc8ed3a2),
	.w4(32'hbc6de3e4),
	.w5(32'hbbef6980),
	.w6(32'h3bf6167e),
	.w7(32'h3be35b9a),
	.w8(32'hbbdebb98),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d07a6),
	.w1(32'h3c6c81dd),
	.w2(32'h3c2ddea4),
	.w3(32'hbca6526c),
	.w4(32'h3a75d813),
	.w5(32'h3b65651b),
	.w6(32'hbc84706c),
	.w7(32'hb9da82ea),
	.w8(32'h3c163883),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63487e),
	.w1(32'hbafbe1d5),
	.w2(32'h3ad1a418),
	.w3(32'hbb3b926d),
	.w4(32'hbbd75f00),
	.w5(32'h3c4c275a),
	.w6(32'hb96d4a22),
	.w7(32'h3b0882ec),
	.w8(32'h3b8b0289),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7524fa),
	.w1(32'hbca0da25),
	.w2(32'hbc0bf594),
	.w3(32'h3c32cf53),
	.w4(32'h3bb31cf5),
	.w5(32'h398b216f),
	.w6(32'h3b4fc60c),
	.w7(32'h399109df),
	.w8(32'hbc2a71a3),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe1d15),
	.w1(32'hbb9cd48e),
	.w2(32'hbc253bdf),
	.w3(32'h3c24cb9a),
	.w4(32'hbb79d431),
	.w5(32'hbc387982),
	.w6(32'hbaa23b8b),
	.w7(32'hbc3f6ea5),
	.w8(32'hbc339526),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2140d0),
	.w1(32'h3bb65ecc),
	.w2(32'hb9db96f8),
	.w3(32'h3b2bd833),
	.w4(32'hbc0120dd),
	.w5(32'h3ac9c535),
	.w6(32'h3b44116c),
	.w7(32'hba137942),
	.w8(32'h3bac96a9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c037540),
	.w1(32'h3c719547),
	.w2(32'h3bd8dfde),
	.w3(32'hbc14f99f),
	.w4(32'hbb53239b),
	.w5(32'h3b9beb7d),
	.w6(32'h38e253a0),
	.w7(32'h3bbab9c7),
	.w8(32'hbc83cc8d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce0bc5e),
	.w1(32'hbcc74a36),
	.w2(32'hbca30608),
	.w3(32'h3ca03732),
	.w4(32'h3af6658a),
	.w5(32'hbbd2bf7e),
	.w6(32'h3b8e3d0d),
	.w7(32'hbbac1d03),
	.w8(32'h3ba0bfc4),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06bca5),
	.w1(32'h3c9fc99b),
	.w2(32'h3c16128d),
	.w3(32'hbc78d892),
	.w4(32'hbbdfc3ce),
	.w5(32'h3c22c76f),
	.w6(32'h3ca2ec33),
	.w7(32'h3c1564b1),
	.w8(32'hbcba3fe8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd132771),
	.w1(32'hbca6bbc1),
	.w2(32'hbcb240a6),
	.w3(32'h3cfa2649),
	.w4(32'h3d06ba01),
	.w5(32'hbae6c047),
	.w6(32'hbcbfc483),
	.w7(32'hbbdf5aa1),
	.w8(32'h3bb672da),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4f374),
	.w1(32'hbb32d384),
	.w2(32'hbb6e8f91),
	.w3(32'h3be7f598),
	.w4(32'hbb17dd97),
	.w5(32'h3c0b920f),
	.w6(32'hbb5b3cb7),
	.w7(32'hbc210137),
	.w8(32'hbc60e234),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06cc9f),
	.w1(32'hbc878e0f),
	.w2(32'hbc3a3391),
	.w3(32'h3cef72c8),
	.w4(32'h3cafc351),
	.w5(32'hbc09f223),
	.w6(32'hbcb05352),
	.w7(32'hbc09dff8),
	.w8(32'hbc3e4c79),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc5c3f),
	.w1(32'h3c14074f),
	.w2(32'hbbac730d),
	.w3(32'hbc78ef22),
	.w4(32'hbb2f24ec),
	.w5(32'hbc9e0025),
	.w6(32'hbbf3afab),
	.w7(32'hbc01a8e0),
	.w8(32'h3b0b323d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e1e87),
	.w1(32'h3cc8ca9b),
	.w2(32'h3c36c9cc),
	.w3(32'hbcee5f6a),
	.w4(32'hbcb4919e),
	.w5(32'hbae98b32),
	.w6(32'hbb9a9b80),
	.w7(32'hbc2714b5),
	.w8(32'hbb1f9c99),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9201c1),
	.w1(32'hbb42ae08),
	.w2(32'hba8cc2c8),
	.w3(32'h3c148d0d),
	.w4(32'h3ac4d8c8),
	.w5(32'hbae9ba3d),
	.w6(32'h3cd13eb2),
	.w7(32'h3c8a7bc6),
	.w8(32'hbc679966),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdcd80a),
	.w1(32'hbce9d85e),
	.w2(32'hbcce69ab),
	.w3(32'h3c94f6f6),
	.w4(32'h3c80fe74),
	.w5(32'h3bf20f72),
	.w6(32'hbb18771e),
	.w7(32'hbb130f08),
	.w8(32'h3c19d903),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef4fa4),
	.w1(32'hbc40cf3d),
	.w2(32'hbc1a5048),
	.w3(32'h3bdd7beb),
	.w4(32'hbbffa33d),
	.w5(32'hbad41e20),
	.w6(32'h3b0926af),
	.w7(32'hbc2c8e5c),
	.w8(32'h3bad637a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94f72f),
	.w1(32'h3be66a7e),
	.w2(32'hbc343b2a),
	.w3(32'hbb16a949),
	.w4(32'hbc122eee),
	.w5(32'hbbaac15a),
	.w6(32'h3cafd4a3),
	.w7(32'h3c0b1c90),
	.w8(32'hbacd2865),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d01e6),
	.w1(32'hbc57f887),
	.w2(32'hbbeaadf0),
	.w3(32'h3c2e24b7),
	.w4(32'hba569ce9),
	.w5(32'hbb0c8abe),
	.w6(32'h3c264e96),
	.w7(32'hbae63ed6),
	.w8(32'h3c124051),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab9742),
	.w1(32'hba4ce3f4),
	.w2(32'h3b14fcd7),
	.w3(32'hbc43d3a7),
	.w4(32'hbc1af64b),
	.w5(32'h3b65a758),
	.w6(32'hbc2c2548),
	.w7(32'hb910f15c),
	.w8(32'h3b94e6d0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9d5b9),
	.w1(32'hbca6682a),
	.w2(32'hbcaeb014),
	.w3(32'hbca6d648),
	.w4(32'hbbd8985d),
	.w5(32'hbb907daf),
	.w6(32'hbb37b9ef),
	.w7(32'hbc0a8d58),
	.w8(32'hbc594b97),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38d28b),
	.w1(32'hbb765c37),
	.w2(32'h3aea67ca),
	.w3(32'h3bc8c25e),
	.w4(32'h3aadec9b),
	.w5(32'hbbe43e32),
	.w6(32'hbc37a8de),
	.w7(32'hbbae863e),
	.w8(32'h3c14cab7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c781549),
	.w1(32'h3cd939b8),
	.w2(32'h3c6ff23e),
	.w3(32'hbccd568d),
	.w4(32'hbcbc8652),
	.w5(32'hbc098377),
	.w6(32'h3c007994),
	.w7(32'hbbd25dde),
	.w8(32'hba5eea4e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d040e8d),
	.w1(32'hbc189de3),
	.w2(32'hbc2e2232),
	.w3(32'h3d0cc03d),
	.w4(32'hbc6058a5),
	.w5(32'hbc3faad6),
	.w6(32'h3cd48e7a),
	.w7(32'h3c834eb5),
	.w8(32'hbb98a2b8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cf2a8),
	.w1(32'h3a6ec296),
	.w2(32'hba57a5a4),
	.w3(32'h3bd4afae),
	.w4(32'h3b71bc8c),
	.w5(32'h3886da32),
	.w6(32'h3c7578ac),
	.w7(32'hb91011cf),
	.w8(32'hbc6d1feb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a96c4),
	.w1(32'hbc326872),
	.w2(32'h3ba0b69e),
	.w3(32'h3c8e3b3d),
	.w4(32'h3bf88477),
	.w5(32'h3c556170),
	.w6(32'h3c1ff780),
	.w7(32'h3ca40336),
	.w8(32'hbc334dbb),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7febaa),
	.w1(32'hbb0ee2d0),
	.w2(32'hbc117ece),
	.w3(32'hbbbc287f),
	.w4(32'h3ccb3b1b),
	.w5(32'h3a764e4c),
	.w6(32'hbd01af25),
	.w7(32'hbbcde3f3),
	.w8(32'h3c786a3c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b2080),
	.w1(32'h3aaccb1e),
	.w2(32'h3c0fbd9a),
	.w3(32'hbcef9273),
	.w4(32'h3b1f7a0d),
	.w5(32'hbca49bf9),
	.w6(32'hbcb31ae9),
	.w7(32'h3bd013ac),
	.w8(32'h3b64b020),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dca1b),
	.w1(32'h3c10b562),
	.w2(32'h3b8d0982),
	.w3(32'hbc6fe896),
	.w4(32'hbc803e56),
	.w5(32'h3c0c9e5b),
	.w6(32'h3ba1c991),
	.w7(32'hba7fd39f),
	.w8(32'hbc328838),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b3ed7),
	.w1(32'hbc14b6c1),
	.w2(32'hbbade8a9),
	.w3(32'hb87f79cc),
	.w4(32'hbaedb26f),
	.w5(32'hbb21a7d5),
	.w6(32'hbc9df6c1),
	.w7(32'hbbb3467d),
	.w8(32'h3a307617),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fa71a),
	.w1(32'h3b78268f),
	.w2(32'hbb5ca718),
	.w3(32'h3c451156),
	.w4(32'h3bbd0e6e),
	.w5(32'h3918b130),
	.w6(32'h3c27f53c),
	.w7(32'hbba2b2ec),
	.w8(32'hbaad7532),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11db96),
	.w1(32'hba81d4a8),
	.w2(32'h3bcdb6aa),
	.w3(32'h3b5b4427),
	.w4(32'hbc7b636e),
	.w5(32'hbb2b1d2f),
	.w6(32'h3c0509a6),
	.w7(32'hbc11c4fc),
	.w8(32'hba9212d5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd2b23),
	.w1(32'hbbfbfc64),
	.w2(32'hbb56d9f0),
	.w3(32'h3abb2a81),
	.w4(32'hb9bf060a),
	.w5(32'h3bebd8e9),
	.w6(32'h3b368ae6),
	.w7(32'h3b067459),
	.w8(32'h3bb3841b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6caa6b),
	.w1(32'h3b335ece),
	.w2(32'h3bda2fe7),
	.w3(32'h3c8be04a),
	.w4(32'hbba4c1bf),
	.w5(32'h3b891f9a),
	.w6(32'h3c429e55),
	.w7(32'hbb406aea),
	.w8(32'h3b4bcfba),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02348b),
	.w1(32'hbb2151f2),
	.w2(32'hbbc4d4f7),
	.w3(32'hbb81924f),
	.w4(32'hbb94cb64),
	.w5(32'hbc0b6850),
	.w6(32'hbc1da131),
	.w7(32'hbb671f6d),
	.w8(32'hbbb9f475),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d8ad3),
	.w1(32'hbbf2124b),
	.w2(32'hbbb50d26),
	.w3(32'hbb6f3842),
	.w4(32'hbacac1d5),
	.w5(32'h3bee213b),
	.w6(32'h3b089748),
	.w7(32'hbb9068da),
	.w8(32'h3b6ee1ef),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73295e),
	.w1(32'hbbc774fe),
	.w2(32'hb9a69b21),
	.w3(32'h3ce9a0e8),
	.w4(32'h3a4ec2fb),
	.w5(32'h3ad80f95),
	.w6(32'h3d23b9f6),
	.w7(32'h3c0bb9d6),
	.w8(32'hbbea8e9b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67afef),
	.w1(32'hba4b546d),
	.w2(32'h3bbfff6d),
	.w3(32'hb9b92549),
	.w4(32'h3b82faa2),
	.w5(32'h3a211ebd),
	.w6(32'h3b8c7676),
	.w7(32'h3b049ffd),
	.w8(32'hbbe052ef),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19868f),
	.w1(32'hbbe817d7),
	.w2(32'hbaf5c79b),
	.w3(32'h38193009),
	.w4(32'hbba8f342),
	.w5(32'hbb8d0f73),
	.w6(32'h3bdf9893),
	.w7(32'h3be3af77),
	.w8(32'hbb2c7f24),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9988bc),
	.w1(32'hbbfafc39),
	.w2(32'hbba09742),
	.w3(32'hbb4a886c),
	.w4(32'hbb3426ef),
	.w5(32'hb9d8549a),
	.w6(32'hbbd52b09),
	.w7(32'h3b422fee),
	.w8(32'hbaeb39c6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81bc9e),
	.w1(32'hbbc313a8),
	.w2(32'hbbb14091),
	.w3(32'hb9dc3339),
	.w4(32'h3a5cbacb),
	.w5(32'h3b9dff4b),
	.w6(32'h3a6e7842),
	.w7(32'hbba2b3f9),
	.w8(32'h3a10243f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c78ef),
	.w1(32'h3bce03c0),
	.w2(32'h3b70a424),
	.w3(32'hba002738),
	.w4(32'hba29decc),
	.w5(32'h3a963e27),
	.w6(32'h3a3c0070),
	.w7(32'hbb260039),
	.w8(32'h3ba5ccf5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b816ec8),
	.w1(32'h3b4666a1),
	.w2(32'hbc042629),
	.w3(32'h3bf10ffb),
	.w4(32'hb93cdb5e),
	.w5(32'hbae22f12),
	.w6(32'h3b85a4c0),
	.w7(32'hbb2b34de),
	.w8(32'hbb9c816d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd94729),
	.w1(32'hbbd5dd4a),
	.w2(32'h3b0ede50),
	.w3(32'h3b22b977),
	.w4(32'h3af0594c),
	.w5(32'hbbac8076),
	.w6(32'h3a9e89ed),
	.w7(32'h3b11b696),
	.w8(32'hbbbb5158),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf83757),
	.w1(32'hbbc540aa),
	.w2(32'hbbad93df),
	.w3(32'hbbae36bc),
	.w4(32'hbb2f086f),
	.w5(32'hba2824c5),
	.w6(32'hbbe9f7e3),
	.w7(32'hbb19bd90),
	.w8(32'h3b916fd8),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfbaba),
	.w1(32'hbbbad67f),
	.w2(32'hbb625095),
	.w3(32'hbbd34fb8),
	.w4(32'h3af03f42),
	.w5(32'hbbcfab36),
	.w6(32'h3ca80fc4),
	.w7(32'h3c03e6c3),
	.w8(32'hbc19bc99),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8758),
	.w1(32'hbbbbf183),
	.w2(32'hbb28878b),
	.w3(32'h3aff870c),
	.w4(32'hbbac5f63),
	.w5(32'hbba5da3b),
	.w6(32'h3c1f1736),
	.w7(32'hbb5d19cc),
	.w8(32'hbc33f122),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd98731),
	.w1(32'hbb93b40a),
	.w2(32'hbb747abc),
	.w3(32'hbbb887ba),
	.w4(32'hbba935fd),
	.w5(32'h3bf0d3f6),
	.w6(32'h3b2504ea),
	.w7(32'h3a102ff8),
	.w8(32'hbb2b3b09),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7feee5),
	.w1(32'h3c4d2141),
	.w2(32'hbb880f0d),
	.w3(32'h3b1a8497),
	.w4(32'h3990dce1),
	.w5(32'hbc3d2fbd),
	.w6(32'h3c296fa4),
	.w7(32'hbba253bb),
	.w8(32'hbc489408),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb771242),
	.w1(32'h3a0ddfac),
	.w2(32'hbb40c3b6),
	.w3(32'h3a2519fb),
	.w4(32'h3ba81f50),
	.w5(32'h3c0395c5),
	.w6(32'h3c2c5a79),
	.w7(32'h3aa89b3d),
	.w8(32'h3bb61e84),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb9d89),
	.w1(32'h3b2c04ac),
	.w2(32'h3adf5351),
	.w3(32'hb96def73),
	.w4(32'h3a224165),
	.w5(32'h3b4237e9),
	.w6(32'hbaf02b84),
	.w7(32'hbb3fa626),
	.w8(32'hbb0196e7),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb717034),
	.w1(32'hbbec4467),
	.w2(32'hbc25388e),
	.w3(32'hbc4e36bc),
	.w4(32'hbc0fb5f4),
	.w5(32'h39ea6ace),
	.w6(32'hbb7f3a6d),
	.w7(32'hbbf7d130),
	.w8(32'hbae4d5a7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1197a0),
	.w1(32'h3b2f8fe4),
	.w2(32'hbb4d93b7),
	.w3(32'hbb9172fc),
	.w4(32'hb938c651),
	.w5(32'h3bbc1e53),
	.w6(32'h3b1d33de),
	.w7(32'hbb6fb943),
	.w8(32'hbbede87e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb774bd0),
	.w1(32'hbb76b6fb),
	.w2(32'h39c902e9),
	.w3(32'h3afafd70),
	.w4(32'h3adb9114),
	.w5(32'hbb60c073),
	.w6(32'h39944c12),
	.w7(32'h3b025f50),
	.w8(32'hba499852),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8701817),
	.w1(32'h3b96166d),
	.w2(32'h3c2942ac),
	.w3(32'h3a821352),
	.w4(32'h3bcb91f6),
	.w5(32'h3b67bff4),
	.w6(32'h3b652282),
	.w7(32'h3c27bd7a),
	.w8(32'h3a87b109),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4e231),
	.w1(32'h3c2c58c1),
	.w2(32'h3c7a732f),
	.w3(32'h3c8c661b),
	.w4(32'h3caee860),
	.w5(32'hbc94e1c9),
	.w6(32'h3c7b1ce0),
	.w7(32'h3caae784),
	.w8(32'hbba60296),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d5794),
	.w1(32'hbac1f995),
	.w2(32'hbc9d26ab),
	.w3(32'h3a2d915c),
	.w4(32'h3c1d8a2b),
	.w5(32'h3c548f08),
	.w6(32'hbb28fb84),
	.w7(32'hbbdb107e),
	.w8(32'h3c44611a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a52f4),
	.w1(32'h3aa6b8ae),
	.w2(32'h3c6e8f28),
	.w3(32'h3bf88af7),
	.w4(32'hbc0c8a2b),
	.w5(32'hbc578f0e),
	.w6(32'h3c9cb1e4),
	.w7(32'h3b3f4cec),
	.w8(32'hbc51552a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c180a89),
	.w1(32'hbb5f3614),
	.w2(32'hbc87c588),
	.w3(32'hbb7fd407),
	.w4(32'h39e5679a),
	.w5(32'h3ab05c57),
	.w6(32'hba8494e2),
	.w7(32'h3b8e91f4),
	.w8(32'hbabbb380),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45b4bf),
	.w1(32'h3c1b17a4),
	.w2(32'h3c411980),
	.w3(32'hbc8d5fb6),
	.w4(32'h3c0fb191),
	.w5(32'h3bd3379a),
	.w6(32'h3c6aa681),
	.w7(32'h3c1d4b5a),
	.w8(32'hbc0759b6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61e84e),
	.w1(32'hbb33c6ee),
	.w2(32'h3b07066a),
	.w3(32'h3969f168),
	.w4(32'h3b1c3efe),
	.w5(32'h3b2ba67f),
	.w6(32'hba859215),
	.w7(32'hbb1b8534),
	.w8(32'h3bff4c05),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1597fa),
	.w1(32'h3b3055f4),
	.w2(32'hb6fd58ee),
	.w3(32'h3b4e1860),
	.w4(32'h3b494bcb),
	.w5(32'hbc144dda),
	.w6(32'hbc49fc1f),
	.w7(32'hbb53b8d5),
	.w8(32'hbba42c86),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule