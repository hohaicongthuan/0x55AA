module layer_10_featuremap_314(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813039),
	.w1(32'h3a49dd48),
	.w2(32'hba31b9d9),
	.w3(32'h3b835981),
	.w4(32'h3b4e9007),
	.w5(32'h3aab52ef),
	.w6(32'h3aa3cbb2),
	.w7(32'h3b2e2388),
	.w8(32'h3b3cab51),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae21b6),
	.w1(32'h3b143727),
	.w2(32'h3a4d9ccc),
	.w3(32'hb9538e9c),
	.w4(32'hba83e6c6),
	.w5(32'h3b929b40),
	.w6(32'h38c7af93),
	.w7(32'h3ad4739c),
	.w8(32'h3aa5d9a4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab76df1),
	.w1(32'h3a74f59b),
	.w2(32'hb9770f45),
	.w3(32'h3bb2fe76),
	.w4(32'hbaf6edc9),
	.w5(32'h3b9cfde8),
	.w6(32'h3ba26460),
	.w7(32'h3be80979),
	.w8(32'h3a8f2db6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a49d7),
	.w1(32'h3b4ffd92),
	.w2(32'h3b75f139),
	.w3(32'h3bd7e03e),
	.w4(32'h3b90caca),
	.w5(32'h3bab1789),
	.w6(32'h3bfb9a65),
	.w7(32'h3bd006ce),
	.w8(32'hbac2defe),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97a326),
	.w1(32'hbb60f0ed),
	.w2(32'hbba0f9b9),
	.w3(32'hbb3dc4a3),
	.w4(32'hbba1c6a4),
	.w5(32'hbad0479b),
	.w6(32'hbb9a41da),
	.w7(32'hbbfcfb6a),
	.w8(32'hbb30b5dd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84c84a),
	.w1(32'hbabbca33),
	.w2(32'hbb183a60),
	.w3(32'h3a82c036),
	.w4(32'h3a8903c1),
	.w5(32'h3a55f139),
	.w6(32'h3a36a0eb),
	.w7(32'h3ab8cd55),
	.w8(32'hba8b54da),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ddd4d),
	.w1(32'hbad6e451),
	.w2(32'h391ac6d8),
	.w3(32'h3ad11dbf),
	.w4(32'h3a01fba2),
	.w5(32'h3baed94e),
	.w6(32'h3ad4e9d9),
	.w7(32'h39b21c66),
	.w8(32'h3b72ddfe),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395045c0),
	.w1(32'h3b353d3d),
	.w2(32'h3b3c4dd3),
	.w3(32'h3be2e9ff),
	.w4(32'h3bb6b6b8),
	.w5(32'hba8caca1),
	.w6(32'h3b36f8be),
	.w7(32'h3ba2cd42),
	.w8(32'hbac7ea1e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc9185),
	.w1(32'hbaa38376),
	.w2(32'hbb13f964),
	.w3(32'hb80df36a),
	.w4(32'hbb07581e),
	.w5(32'hbae395b2),
	.w6(32'hba1903a7),
	.w7(32'hbac667e2),
	.w8(32'hbb090a43),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90612e),
	.w1(32'h3b10a334),
	.w2(32'h3aa310dd),
	.w3(32'h3b6ecfbf),
	.w4(32'h3b54f0f9),
	.w5(32'h3b61d4f4),
	.w6(32'h3b84e261),
	.w7(32'h3b7117e9),
	.w8(32'h39df5ded),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1d473),
	.w1(32'hb83b8b33),
	.w2(32'hb99e8203),
	.w3(32'h3b0207b1),
	.w4(32'hba7cda87),
	.w5(32'hbac6a487),
	.w6(32'h3ae9fbe3),
	.w7(32'h39a02dd5),
	.w8(32'hbb77bfad),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04032f),
	.w1(32'hbbbe4d07),
	.w2(32'hbb7728e9),
	.w3(32'hba4d44ca),
	.w4(32'hbb8fb6cf),
	.w5(32'h3b8a30aa),
	.w6(32'hbb564863),
	.w7(32'hba987dcc),
	.w8(32'h3ab05cdf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1711fc),
	.w1(32'h3ba75240),
	.w2(32'h3b9f4e81),
	.w3(32'h3ac336ec),
	.w4(32'h3b82bd99),
	.w5(32'h3c30a6e0),
	.w6(32'h3ac5462a),
	.w7(32'h3b0b8d6f),
	.w8(32'h3be3fee1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8fd6d),
	.w1(32'h38ab3d82),
	.w2(32'h3a73725d),
	.w3(32'h3a603f62),
	.w4(32'hbafa1a70),
	.w5(32'h3ac158ec),
	.w6(32'h3aeaad45),
	.w7(32'hb9904d13),
	.w8(32'hbad54409),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9683e9),
	.w1(32'hba125537),
	.w2(32'h3b607c85),
	.w3(32'h3ae478e4),
	.w4(32'h3b3d1a70),
	.w5(32'hbb887272),
	.w6(32'h39e21ef7),
	.w7(32'h3a506a3a),
	.w8(32'hbb2a5c03),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad2453),
	.w1(32'h398cb547),
	.w2(32'h3a087222),
	.w3(32'hbbb9eb28),
	.w4(32'hba85e77e),
	.w5(32'hbb8bd034),
	.w6(32'hbb75b1c0),
	.w7(32'hbaff4c4b),
	.w8(32'hbbb7f7e2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc61eed),
	.w1(32'hbbd77606),
	.w2(32'hbb8dc531),
	.w3(32'hbba99326),
	.w4(32'hbad24b35),
	.w5(32'hbb6d7724),
	.w6(32'hbb862e39),
	.w7(32'hbb22092c),
	.w8(32'hbb48b9ce),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e75d4),
	.w1(32'h37efdd12),
	.w2(32'hbb8ed120),
	.w3(32'hba65b585),
	.w4(32'hbb420d97),
	.w5(32'hbbb31d4d),
	.w6(32'h3a2a6052),
	.w7(32'hbb0ceba0),
	.w8(32'hbbb0c251),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54e0c1),
	.w1(32'h3b1c0b79),
	.w2(32'h3b98b4fd),
	.w3(32'hb992b8c0),
	.w4(32'hba04dad7),
	.w5(32'hbb001624),
	.w6(32'h3aea4b67),
	.w7(32'hbb028e52),
	.w8(32'h3aca1451),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88c9f0),
	.w1(32'hbac08bab),
	.w2(32'hbb6f7745),
	.w3(32'hbb47772d),
	.w4(32'hba95eb84),
	.w5(32'hba3680c8),
	.w6(32'hb9f5f1e9),
	.w7(32'hbb5bf212),
	.w8(32'hba054f6c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991d01a),
	.w1(32'hba007da0),
	.w2(32'h3ab27fcd),
	.w3(32'hbb859269),
	.w4(32'hbacc2aa8),
	.w5(32'h3b12edbd),
	.w6(32'hb9d44452),
	.w7(32'hba317db8),
	.w8(32'h3a9cc1d1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6de0e),
	.w1(32'h3add9a6f),
	.w2(32'h3b02319f),
	.w3(32'h3adf9537),
	.w4(32'h3b242df6),
	.w5(32'h38bff9f6),
	.w6(32'h36c02856),
	.w7(32'h3aeb5ec0),
	.w8(32'h3986746d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4e9f7),
	.w1(32'hb933d501),
	.w2(32'hba58c708),
	.w3(32'hbad869a3),
	.w4(32'h3a1da573),
	.w5(32'h3b77168b),
	.w6(32'hbb451f13),
	.w7(32'h38587cf0),
	.w8(32'h3b31c58e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaae6bc),
	.w1(32'h3ba713ec),
	.w2(32'h3bae6e35),
	.w3(32'h3b1f05db),
	.w4(32'h3a2133e5),
	.w5(32'hbacfd97a),
	.w6(32'h39c84088),
	.w7(32'h3aa2f166),
	.w8(32'h387ba0bb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81ca2c),
	.w1(32'h3b9dc2a2),
	.w2(32'h3b49ca1f),
	.w3(32'h3995a1e7),
	.w4(32'hbaf29aa5),
	.w5(32'hbb4be897),
	.w6(32'h39b9c10d),
	.w7(32'hbb09b87c),
	.w8(32'hbba3ba2f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3fc80),
	.w1(32'hbbb61861),
	.w2(32'hba91fbc0),
	.w3(32'hbafb3fcc),
	.w4(32'hba72afb6),
	.w5(32'h3b1dd6a6),
	.w6(32'hbb7db793),
	.w7(32'hbb05321f),
	.w8(32'h3b1d5917),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c7cdd),
	.w1(32'hbb12c523),
	.w2(32'h3b10711a),
	.w3(32'h3b52bbd1),
	.w4(32'h3bb41ea3),
	.w5(32'h392a56e6),
	.w6(32'h3aad1523),
	.w7(32'h3c0406e5),
	.w8(32'hba0d052b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cdb38),
	.w1(32'hbaa8093e),
	.w2(32'hbb6d5b11),
	.w3(32'h3a911910),
	.w4(32'hb80cc7ae),
	.w5(32'h3b801da3),
	.w6(32'hb8bc66b1),
	.w7(32'hba55d225),
	.w8(32'h3bb8e705),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b16ab),
	.w1(32'h3ae9b14b),
	.w2(32'h3a0da618),
	.w3(32'h3a007206),
	.w4(32'h39dc5b54),
	.w5(32'h3b4baa08),
	.w6(32'h3bd3cd1f),
	.w7(32'h39908d7a),
	.w8(32'h3b4527c7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51ab71),
	.w1(32'hbb07ec95),
	.w2(32'h3b7da28d),
	.w3(32'h3abd89ca),
	.w4(32'h3b1f5c68),
	.w5(32'hba249e46),
	.w6(32'hb86f20ad),
	.w7(32'h3bb5170a),
	.w8(32'h3b58a4f5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5acfc9),
	.w1(32'h3c1dc052),
	.w2(32'h3b1c727d),
	.w3(32'hb9c0d430),
	.w4(32'hbb695ca1),
	.w5(32'hbb928877),
	.w6(32'hbaeb1dc7),
	.w7(32'hba2e3f73),
	.w8(32'hbb859a3c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38d4f1),
	.w1(32'hbb9c103d),
	.w2(32'hbc1e5786),
	.w3(32'hbb9039bb),
	.w4(32'hb9d7a3e1),
	.w5(32'hbbf4f79a),
	.w6(32'h3a529597),
	.w7(32'hbb5c6286),
	.w8(32'hbb9acc2e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b850b),
	.w1(32'hbb1fbc38),
	.w2(32'h3a2705fb),
	.w3(32'hba27969e),
	.w4(32'hb9c36055),
	.w5(32'hbad7ee1d),
	.w6(32'hbb5ddcd7),
	.w7(32'hba9037d5),
	.w8(32'h3ac57827),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820f89),
	.w1(32'hba29dc2e),
	.w2(32'hbb88ca9f),
	.w3(32'hbb0c7fde),
	.w4(32'hba15db95),
	.w5(32'hb8d88eba),
	.w6(32'hba942799),
	.w7(32'h3a31b23d),
	.w8(32'h3af27257),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d0b08),
	.w1(32'hba3c8061),
	.w2(32'hbb29f9a4),
	.w3(32'h3a456cad),
	.w4(32'h3b9b1e00),
	.w5(32'h3b19684f),
	.w6(32'h39898b37),
	.w7(32'hba9e1800),
	.w8(32'h3a66c9d3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb009e4a),
	.w1(32'hbb28d65a),
	.w2(32'hbb10e087),
	.w3(32'hbbb7659f),
	.w4(32'hba4bb6be),
	.w5(32'hbc23f3bc),
	.w6(32'hbaddb2c7),
	.w7(32'h3a91b3e1),
	.w8(32'hb8d20e14),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f1145),
	.w1(32'hb9de2b14),
	.w2(32'hbb81fe4d),
	.w3(32'hbaa7605a),
	.w4(32'h3b7478bd),
	.w5(32'hb93a3480),
	.w6(32'hbc1dcfb7),
	.w7(32'hbc043e25),
	.w8(32'hb9c2bf3a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3acb3),
	.w1(32'h3acae39a),
	.w2(32'h3ad52a11),
	.w3(32'h3b6d7053),
	.w4(32'h393b3e0b),
	.w5(32'hbbf8cf06),
	.w6(32'h3b8459a1),
	.w7(32'h3c012118),
	.w8(32'hbba75a49),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65fe0a),
	.w1(32'hbad0b195),
	.w2(32'hbb136a6e),
	.w3(32'hbbfd192e),
	.w4(32'hbbbbf48b),
	.w5(32'h3a09e917),
	.w6(32'hbbaca576),
	.w7(32'hbbc22659),
	.w8(32'h3b4d3b04),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06ed7b),
	.w1(32'h3ae49db7),
	.w2(32'hbb58fdff),
	.w3(32'h3b793dd4),
	.w4(32'h3b8ce7a5),
	.w5(32'h3adb4eaf),
	.w6(32'h3b63823d),
	.w7(32'h3abea5ec),
	.w8(32'h3ba914f5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca0161),
	.w1(32'hbaa4b8c4),
	.w2(32'h39027963),
	.w3(32'hbb0b32d0),
	.w4(32'hbb295b0b),
	.w5(32'hb9c1d31f),
	.w6(32'hbb7746f3),
	.w7(32'h3940478c),
	.w8(32'hbaaf6f44),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc88839),
	.w1(32'hbbb2f442),
	.w2(32'h39864f7a),
	.w3(32'h3b4a64e1),
	.w4(32'h3a926efb),
	.w5(32'h3b3c1a9a),
	.w6(32'h3b734c41),
	.w7(32'h3b8a417c),
	.w8(32'h3a6ce5cb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82c1b8),
	.w1(32'h3b073819),
	.w2(32'h397a7669),
	.w3(32'h3c078409),
	.w4(32'h3aba8a96),
	.w5(32'hbba13211),
	.w6(32'h3c12df37),
	.w7(32'h3c17c46e),
	.w8(32'hbab80a87),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52447),
	.w1(32'hbb4726ec),
	.w2(32'hbb993e5b),
	.w3(32'h3aa6d901),
	.w4(32'hbba8008a),
	.w5(32'hb821c9aa),
	.w6(32'h3c813494),
	.w7(32'h3bf2c276),
	.w8(32'h3a37e208),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b003a),
	.w1(32'h3b406ef6),
	.w2(32'h3bd72f60),
	.w3(32'h3c8b1c75),
	.w4(32'h3c59e58a),
	.w5(32'h3c19b777),
	.w6(32'h3c74ebc5),
	.w7(32'h3c3c2a8b),
	.w8(32'hb9f67ea2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921da93),
	.w1(32'h39fd7ecc),
	.w2(32'h3a152dd3),
	.w3(32'h3c3e13c3),
	.w4(32'h3b97598d),
	.w5(32'h3c370e44),
	.w6(32'h3b9d4971),
	.w7(32'h3b80f4dd),
	.w8(32'h3befae86),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eb419),
	.w1(32'h3ad7bd18),
	.w2(32'h3b25b186),
	.w3(32'h3c84c914),
	.w4(32'h3bfae875),
	.w5(32'hba5d83f4),
	.w6(32'h3c1aa0d9),
	.w7(32'h3be08b8d),
	.w8(32'hba406914),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a2424),
	.w1(32'h3b3ac027),
	.w2(32'h3b5e1c45),
	.w3(32'hbb2481f5),
	.w4(32'h38d118b4),
	.w5(32'h3ba051bf),
	.w6(32'hbadf6403),
	.w7(32'hbaced37f),
	.w8(32'h3ba087ba),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd99c86),
	.w1(32'h3bb1e471),
	.w2(32'h3b7925e5),
	.w3(32'h3b21dce0),
	.w4(32'h3b936f54),
	.w5(32'h3a6739a2),
	.w6(32'h3b195edd),
	.w7(32'h3b88ddf3),
	.w8(32'hba086305),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7a057),
	.w1(32'hba079783),
	.w2(32'h3b04d698),
	.w3(32'h3b18cb76),
	.w4(32'h3b8732cd),
	.w5(32'hbb40738f),
	.w6(32'hbabc07c9),
	.w7(32'h3a27b8fe),
	.w8(32'hbb3e27a7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3c366),
	.w1(32'hbc11c9f8),
	.w2(32'hbb9bb5aa),
	.w3(32'hbaf12aaa),
	.w4(32'hbb6420bd),
	.w5(32'h3b15212c),
	.w6(32'hbc03a5fd),
	.w7(32'hbaebc695),
	.w8(32'h3c0bd159),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc09e00),
	.w1(32'h3becd473),
	.w2(32'h3b211423),
	.w3(32'h3bfe790d),
	.w4(32'h3ae442d6),
	.w5(32'h3c0da1cb),
	.w6(32'h3c83fcc3),
	.w7(32'h3c5f1d31),
	.w8(32'h3b455b6b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c1e30),
	.w1(32'hbb0d57e1),
	.w2(32'h3b1035c3),
	.w3(32'h3bbe0f8c),
	.w4(32'hba39551a),
	.w5(32'h3a4d80f8),
	.w6(32'hbb3a9907),
	.w7(32'hb8df2f90),
	.w8(32'h3b84c9ba),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb645769),
	.w1(32'hb8dac64d),
	.w2(32'h3b4ede47),
	.w3(32'hbaa686dc),
	.w4(32'h3c026e52),
	.w5(32'hbb93f748),
	.w6(32'hbb81adaf),
	.w7(32'h3baa56cb),
	.w8(32'hbb11fd96),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb1043),
	.w1(32'h39cb9e7a),
	.w2(32'hbb812df0),
	.w3(32'hbb2a62b9),
	.w4(32'h3b31318d),
	.w5(32'h3b7b7f77),
	.w6(32'hba70bc78),
	.w7(32'hbb8143e8),
	.w8(32'h3af68eb0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a23a7),
	.w1(32'h3977030d),
	.w2(32'hb8cd31c7),
	.w3(32'h3b520d60),
	.w4(32'h3b74481a),
	.w5(32'hbb1a6818),
	.w6(32'h3c134181),
	.w7(32'h3b497f36),
	.w8(32'h3a4c7cee),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9fb3a),
	.w1(32'h3aafa36e),
	.w2(32'h394694a1),
	.w3(32'hba26299c),
	.w4(32'h3b084f03),
	.w5(32'h3bbdd93a),
	.w6(32'h3ad1f33e),
	.w7(32'h3b2042ec),
	.w8(32'h3c0f5895),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6ba37),
	.w1(32'h3b019198),
	.w2(32'hba83442b),
	.w3(32'h3a2f4944),
	.w4(32'h3b94a26b),
	.w5(32'hba5a2fe6),
	.w6(32'hba577ac8),
	.w7(32'h3be2a870),
	.w8(32'hbb242bdf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb698089),
	.w1(32'hbb47a778),
	.w2(32'h3a1dfd39),
	.w3(32'hba9b4156),
	.w4(32'h3a4415e0),
	.w5(32'h3a9a8959),
	.w6(32'hbb3f6263),
	.w7(32'hba9c4792),
	.w8(32'h3a506192),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39417c77),
	.w1(32'h3bccd747),
	.w2(32'h3bef04d7),
	.w3(32'h3c055c09),
	.w4(32'h3b0b1882),
	.w5(32'h3ab3df16),
	.w6(32'h3be16436),
	.w7(32'h3be43f35),
	.w8(32'hba0fe5c2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67e753),
	.w1(32'hba646b5e),
	.w2(32'h39f05aa6),
	.w3(32'h3a72fc6c),
	.w4(32'hb8d017aa),
	.w5(32'h3ad04132),
	.w6(32'h3a980c6a),
	.w7(32'h3a40525f),
	.w8(32'hbb19259f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb853f84),
	.w1(32'hbb9db3a6),
	.w2(32'hba5ebbb7),
	.w3(32'h3a75553c),
	.w4(32'hb974d017),
	.w5(32'h3a8b8f1e),
	.w6(32'h3aed12a9),
	.w7(32'hbb249797),
	.w8(32'h3aeb6b70),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71ecc8),
	.w1(32'h3b066f17),
	.w2(32'hba59c28f),
	.w3(32'hbad5e8ee),
	.w4(32'h3ab2f77a),
	.w5(32'h38815a6f),
	.w6(32'hbad248fe),
	.w7(32'hbb3e0cad),
	.w8(32'h3b0e794e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf27a7),
	.w1(32'hbb809b6d),
	.w2(32'hbaf20d5c),
	.w3(32'hbb4ec795),
	.w4(32'h3a8a04f0),
	.w5(32'h378162bb),
	.w6(32'hbaf9a555),
	.w7(32'hba1a3e10),
	.w8(32'hbaabb6fb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395aec11),
	.w1(32'hb74908e7),
	.w2(32'h3b1a1e8d),
	.w3(32'hbab23004),
	.w4(32'h3b729d08),
	.w5(32'hbb1a57cf),
	.w6(32'h3a082232),
	.w7(32'h3b6fd8ed),
	.w8(32'hbae86ff2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b123423),
	.w1(32'h3aab7587),
	.w2(32'hbabec964),
	.w3(32'hbab5b9c4),
	.w4(32'hbb00280c),
	.w5(32'h3b7b978a),
	.w6(32'hbacb8e32),
	.w7(32'hbb033150),
	.w8(32'h3af5b080),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea310a),
	.w1(32'h3aeeda58),
	.w2(32'h3a9bc7f4),
	.w3(32'h3b378b6c),
	.w4(32'h3b2a0f6b),
	.w5(32'hbb6126c6),
	.w6(32'h3acd1416),
	.w7(32'h3857ea0b),
	.w8(32'hbb6ba943),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b189a09),
	.w1(32'hbab1b729),
	.w2(32'hbadb22cd),
	.w3(32'hbbdf257a),
	.w4(32'hbb62ca83),
	.w5(32'hbacccde9),
	.w6(32'hbbb75f23),
	.w7(32'hbb805f81),
	.w8(32'hbabb4246),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab615d9),
	.w1(32'hbbaa5238),
	.w2(32'h39a6bfdc),
	.w3(32'hbb40d037),
	.w4(32'h3b448399),
	.w5(32'h3b4c0cd0),
	.w6(32'hb8cb6fbf),
	.w7(32'h3b562eae),
	.w8(32'h3b9c110f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21fb85),
	.w1(32'h3c178d91),
	.w2(32'h3befa6c5),
	.w3(32'h3c16d867),
	.w4(32'h3c00f252),
	.w5(32'h3af45ea8),
	.w6(32'h3c85ba4f),
	.w7(32'h3c6bea0f),
	.w8(32'h3b8d87e6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f2e5a),
	.w1(32'h3b652525),
	.w2(32'h3be69614),
	.w3(32'h3c0df78f),
	.w4(32'h3bc43633),
	.w5(32'hb9e6c57e),
	.w6(32'h3b9fc3cd),
	.w7(32'h3bd4d554),
	.w8(32'h3b04ebd2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b144a4f),
	.w1(32'hba2f94f2),
	.w2(32'hba850aba),
	.w3(32'hbb79a1be),
	.w4(32'hbaea72b2),
	.w5(32'hbbd34087),
	.w6(32'hbb9d81ba),
	.w7(32'hbb0f7f11),
	.w8(32'hbb8f8ba9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb099608),
	.w1(32'hbb38588e),
	.w2(32'hbb5f5957),
	.w3(32'hbbd9f53a),
	.w4(32'hbb54b067),
	.w5(32'h3ad71321),
	.w6(32'hbba8629f),
	.w7(32'hbb80ddae),
	.w8(32'h3b8692dd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71f4b3),
	.w1(32'h398dc38e),
	.w2(32'hbb17056e),
	.w3(32'h3a8bd6b0),
	.w4(32'h3b2510fb),
	.w5(32'hbae4a8c1),
	.w6(32'h3a83fa9d),
	.w7(32'h3bc517e6),
	.w8(32'hba38f9dc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a941),
	.w1(32'hba230345),
	.w2(32'hbb54e14e),
	.w3(32'hba5c13e3),
	.w4(32'hb9716f78),
	.w5(32'hba13bb19),
	.w6(32'h3a01e49b),
	.w7(32'hb9a84f7f),
	.w8(32'hba1ec6e4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b81d2),
	.w1(32'h3b1559ee),
	.w2(32'hb97f93ec),
	.w3(32'hbb6cede3),
	.w4(32'hbb969f5e),
	.w5(32'hba2c5335),
	.w6(32'h39e9d98f),
	.w7(32'hbaea1a31),
	.w8(32'hbb369fe6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2239c),
	.w1(32'h3a5bd2df),
	.w2(32'h3b934b8a),
	.w3(32'hbacb4842),
	.w4(32'hbb460585),
	.w5(32'hbb882b7e),
	.w6(32'hbbda3632),
	.w7(32'h389c7e0a),
	.w8(32'hbb782d2f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46b504),
	.w1(32'h38fadf07),
	.w2(32'hbb5b688d),
	.w3(32'h3c06ca85),
	.w4(32'h3b7590b0),
	.w5(32'h3b1ebcfc),
	.w6(32'h3c019f97),
	.w7(32'h3be22872),
	.w8(32'h39d2c42b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7edf5),
	.w1(32'hba519290),
	.w2(32'hb9467e07),
	.w3(32'h3af34380),
	.w4(32'hba8d8be0),
	.w5(32'h39bd81cd),
	.w6(32'hbaaacf94),
	.w7(32'h39190e47),
	.w8(32'hbac59f31),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3fa4a),
	.w1(32'hba2a9351),
	.w2(32'hbb32819f),
	.w3(32'hbaa7a2ce),
	.w4(32'h3ac69524),
	.w5(32'h3bb6a8e7),
	.w6(32'hba9c9646),
	.w7(32'hba5ed1a1),
	.w8(32'h3b1b6b30),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b484e61),
	.w1(32'hbae54266),
	.w2(32'h3b19d26d),
	.w3(32'h3b0e722e),
	.w4(32'h3a57cfb7),
	.w5(32'hba18e36d),
	.w6(32'hbb02c1e2),
	.w7(32'h3b2c6548),
	.w8(32'hba839024),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50e0f0),
	.w1(32'hb77fad6c),
	.w2(32'hba2d2a56),
	.w3(32'hbb4aa8e0),
	.w4(32'hbabb60d2),
	.w5(32'hbaa44087),
	.w6(32'hbae99d69),
	.w7(32'hbb205178),
	.w8(32'hba5fdfb1),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34affb),
	.w1(32'h3a17c48f),
	.w2(32'h3ba8deff),
	.w3(32'hbab4ed6e),
	.w4(32'h3addbcf2),
	.w5(32'hbb8e6883),
	.w6(32'hbb9c0bb4),
	.w7(32'h3b91d63d),
	.w8(32'hbb59268e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4610b4),
	.w1(32'hbba57c01),
	.w2(32'hbaf4470a),
	.w3(32'hbbf69302),
	.w4(32'hbb8bb39d),
	.w5(32'h3af28025),
	.w6(32'hbbd99f1f),
	.w7(32'hbb59245b),
	.w8(32'hba172ae7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926189e),
	.w1(32'hb8563d98),
	.w2(32'hb9999e07),
	.w3(32'hbae67aad),
	.w4(32'hba3e0659),
	.w5(32'h382f6c8e),
	.w6(32'hbb87ce9f),
	.w7(32'hb9b81187),
	.w8(32'h3a1768ac),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a41ad9),
	.w1(32'hba7de1ab),
	.w2(32'hbad0b5ab),
	.w3(32'h3b300d9e),
	.w4(32'hba7f1003),
	.w5(32'hb90a1fa2),
	.w6(32'h3b9e3442),
	.w7(32'h3b7f3262),
	.w8(32'hbaaa89e6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e3aa3),
	.w1(32'hbb845612),
	.w2(32'hb9bf26e1),
	.w3(32'h397f1ae9),
	.w4(32'h3b8cff1a),
	.w5(32'hbb804b94),
	.w6(32'h3a8896f7),
	.w7(32'h3c2c76f6),
	.w8(32'hbb29b816),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9095be),
	.w1(32'hbb0bb044),
	.w2(32'hbbccf8da),
	.w3(32'hbb84b161),
	.w4(32'hbaaa56c7),
	.w5(32'hbb2a2901),
	.w6(32'hb9fc4661),
	.w7(32'hbb635c1e),
	.w8(32'hbb8e7704),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb82ccc),
	.w1(32'hbb06e086),
	.w2(32'hba9810e6),
	.w3(32'h3aa58bcc),
	.w4(32'h3a33f1b2),
	.w5(32'h3b8c6623),
	.w6(32'hba2abb40),
	.w7(32'hb89fbcd0),
	.w8(32'h3aace7f2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e80b1),
	.w1(32'hbb18704d),
	.w2(32'hbb6f33e3),
	.w3(32'h39a8f396),
	.w4(32'h3adf012f),
	.w5(32'h3a620677),
	.w6(32'hbb9296ff),
	.w7(32'hbb28dc4e),
	.w8(32'h3a4545fe),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5a182),
	.w1(32'hbaac4950),
	.w2(32'hbb0eeef0),
	.w3(32'hbb1f79dd),
	.w4(32'h39d3f8e5),
	.w5(32'h3c23e615),
	.w6(32'hbb38e7a4),
	.w7(32'hbba28c82),
	.w8(32'h3bd2ad6d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b780aa5),
	.w1(32'hbb0ff642),
	.w2(32'h3ac2ceef),
	.w3(32'h3b46b92b),
	.w4(32'hbbacdb92),
	.w5(32'h3b91ed15),
	.w6(32'h3bec4578),
	.w7(32'hba1db0d2),
	.w8(32'h3aeb4731),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a597),
	.w1(32'h3a0d9345),
	.w2(32'h3b02256b),
	.w3(32'hbb0b834c),
	.w4(32'h3aa46d1a),
	.w5(32'h3b576545),
	.w6(32'h3c87d06b),
	.w7(32'hbb00dc75),
	.w8(32'h3be7f319),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acafe68),
	.w1(32'hba318599),
	.w2(32'hbc132655),
	.w3(32'hba8dddc2),
	.w4(32'hbc06d17f),
	.w5(32'h3aaad7b4),
	.w6(32'h3bb456b2),
	.w7(32'hbb0d7890),
	.w8(32'h3a9a4471),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898bf72),
	.w1(32'hb9fc6eb2),
	.w2(32'h3afd6db9),
	.w3(32'h3b318ca3),
	.w4(32'h3a7b352a),
	.w5(32'hbb014c44),
	.w6(32'h3a6e5d69),
	.w7(32'h3b156bdf),
	.w8(32'hbb402f02),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91799c1),
	.w1(32'hb99c958d),
	.w2(32'hbab75159),
	.w3(32'h3b9ba3bc),
	.w4(32'h3b86f74e),
	.w5(32'hbad17eb0),
	.w6(32'h3c58b2b8),
	.w7(32'h3c86e4ea),
	.w8(32'hbb48a649),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860cfd),
	.w1(32'hb9fd8c6b),
	.w2(32'hbac0489d),
	.w3(32'h3a0c8514),
	.w4(32'hbada1d7b),
	.w5(32'hbb992f61),
	.w6(32'hbac14efb),
	.w7(32'hbbac57c2),
	.w8(32'hbbe796e9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedda1a),
	.w1(32'h3b9d8603),
	.w2(32'h3be8cda6),
	.w3(32'h3ae0a8b6),
	.w4(32'h3b5eead9),
	.w5(32'h3ac5b436),
	.w6(32'hbb12a444),
	.w7(32'h3b1a206c),
	.w8(32'h3aa09851),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3943dd60),
	.w1(32'h3a7b84d8),
	.w2(32'hbaf37da7),
	.w3(32'hb7b96f7b),
	.w4(32'hbaef269e),
	.w5(32'h39d74e83),
	.w6(32'h3a454e46),
	.w7(32'hba92a34b),
	.w8(32'hb8cb6e74),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11ddc8),
	.w1(32'hbae19089),
	.w2(32'hbb7dc78b),
	.w3(32'hbae8b4f7),
	.w4(32'hbb296654),
	.w5(32'h3b8aabb1),
	.w6(32'hbbd9313b),
	.w7(32'hbb1d7fc6),
	.w8(32'h3bb2b9cf),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6131c3),
	.w1(32'h3b90ae2c),
	.w2(32'h3b5dfc55),
	.w3(32'h3b57446a),
	.w4(32'h39c75e5e),
	.w5(32'hbbadb9fb),
	.w6(32'h3b98a29f),
	.w7(32'h3ae6a819),
	.w8(32'hbb3138d6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aef21),
	.w1(32'hbb8a0752),
	.w2(32'hbb120770),
	.w3(32'hb55ea2e6),
	.w4(32'h39e57389),
	.w5(32'h3b93ce63),
	.w6(32'hba749cb9),
	.w7(32'h399b24bd),
	.w8(32'h3b288940),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49d097),
	.w1(32'h3ac73c36),
	.w2(32'h3abba9ea),
	.w3(32'h3b3b9439),
	.w4(32'h3b1e96bd),
	.w5(32'hbb5267c6),
	.w6(32'h3adfb210),
	.w7(32'h3b0735ed),
	.w8(32'hbba8c0fe),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffd3bf),
	.w1(32'hbae412e8),
	.w2(32'hbb119b82),
	.w3(32'hbb7efedc),
	.w4(32'hbae143d7),
	.w5(32'h3b2680c4),
	.w6(32'hbb087036),
	.w7(32'hbaadba1c),
	.w8(32'h3ba74858),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f41ee),
	.w1(32'hbadcdf17),
	.w2(32'hbb35a61b),
	.w3(32'h3a0a3f68),
	.w4(32'h3aee8088),
	.w5(32'hbb197ee6),
	.w6(32'h3a4d8712),
	.w7(32'hbaad0a96),
	.w8(32'hbb4b89c1),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d5474),
	.w1(32'hbb505bb2),
	.w2(32'hbb3fc763),
	.w3(32'hbabe91a2),
	.w4(32'hbb59828c),
	.w5(32'h3b5e0c92),
	.w6(32'hbb3c5c39),
	.w7(32'hbb5bd699),
	.w8(32'h3b2a5dd6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5ab30),
	.w1(32'h3ab0f457),
	.w2(32'h3a9cfd6c),
	.w3(32'h3b37582d),
	.w4(32'h3b0b4058),
	.w5(32'h3b34805e),
	.w6(32'h3b06ab67),
	.w7(32'hba34d8c3),
	.w8(32'h3b511f74),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3354bd),
	.w1(32'h3a091ef9),
	.w2(32'hbb0afabe),
	.w3(32'h3a9761a6),
	.w4(32'hbad21d3a),
	.w5(32'hbb841afa),
	.w6(32'hbae66abe),
	.w7(32'hbb3d990c),
	.w8(32'hbb89e46b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59297e),
	.w1(32'hba8c7b6e),
	.w2(32'hbb9e7668),
	.w3(32'hba3b8d89),
	.w4(32'hbbb4f85e),
	.w5(32'h3b852a44),
	.w6(32'hbb0f36fb),
	.w7(32'hbbdb8639),
	.w8(32'h3b91424e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62bf83),
	.w1(32'h3b8c5ff9),
	.w2(32'h3addc21f),
	.w3(32'h3b4430fe),
	.w4(32'h39f5fd88),
	.w5(32'h3b0c5497),
	.w6(32'h3b7cd8bf),
	.w7(32'h3a57324c),
	.w8(32'hb982c1e9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1854e),
	.w1(32'hbbc301bb),
	.w2(32'hbb778d64),
	.w3(32'h3a306af5),
	.w4(32'hbbad6702),
	.w5(32'h3b1d5a77),
	.w6(32'hbb7fd531),
	.w7(32'hbbaeee6d),
	.w8(32'h3aef2789),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03a1b6),
	.w1(32'h38bdd414),
	.w2(32'hbb021009),
	.w3(32'h3a9b4eb2),
	.w4(32'hba7d3894),
	.w5(32'h3a97e23f),
	.w6(32'hb905984f),
	.w7(32'hba8effc1),
	.w8(32'h3ab897e3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7e035),
	.w1(32'h3a804e57),
	.w2(32'h3b029d32),
	.w3(32'h3b05ae45),
	.w4(32'h3aef5f6e),
	.w5(32'h3b181420),
	.w6(32'h3a9960e7),
	.w7(32'h3aa8c5db),
	.w8(32'hba22cce8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a146417),
	.w1(32'hbabc651d),
	.w2(32'hba83fa26),
	.w3(32'h3b1b6b2d),
	.w4(32'h3ace235b),
	.w5(32'hba1821b6),
	.w6(32'h3a72ccd7),
	.w7(32'h3af5a6b4),
	.w8(32'hbab40ef6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b5934),
	.w1(32'h39e17c78),
	.w2(32'hba97a972),
	.w3(32'h389905ae),
	.w4(32'hba3dd8d3),
	.w5(32'h3a116343),
	.w6(32'hbb3fba83),
	.w7(32'hba9e169e),
	.w8(32'h3a7072c0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd5390),
	.w1(32'hbb0f31f4),
	.w2(32'hbb461c47),
	.w3(32'hba072db8),
	.w4(32'hba87a20c),
	.w5(32'hb9cbb5e5),
	.w6(32'hbaba3292),
	.w7(32'hba2c681e),
	.w8(32'h39ce50cb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b131356),
	.w1(32'h3ae792e3),
	.w2(32'h3b55cde3),
	.w3(32'h3a5aac43),
	.w4(32'h3ad22c9e),
	.w5(32'hb925582b),
	.w6(32'h3a05df37),
	.w7(32'h39c7d18e),
	.w8(32'h3c0315ab),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d887d),
	.w1(32'h3abb059f),
	.w2(32'hbb028974),
	.w3(32'hb92db827),
	.w4(32'h39f7955a),
	.w5(32'hba817031),
	.w6(32'h3a0c065c),
	.w7(32'hb91c5dd0),
	.w8(32'hbb0253f4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a82d8),
	.w1(32'hbb0eb808),
	.w2(32'hbb1f3a5c),
	.w3(32'hba3926fb),
	.w4(32'hbaced8ca),
	.w5(32'h3a9d6ad6),
	.w6(32'hbae190e7),
	.w7(32'hba9a683a),
	.w8(32'h3b693c39),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831d5b),
	.w1(32'h3bc9acd2),
	.w2(32'h3a6f8035),
	.w3(32'h3ba60143),
	.w4(32'h39a6ace1),
	.w5(32'h3b1c542a),
	.w6(32'h3bfc0ccd),
	.w7(32'h3a913e6d),
	.w8(32'hb885ed62),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa35301),
	.w1(32'hba59663e),
	.w2(32'h394035e9),
	.w3(32'hb9f4ef64),
	.w4(32'hba81d3ec),
	.w5(32'hba8e200d),
	.w6(32'hbab8eadc),
	.w7(32'hbaa226ac),
	.w8(32'hbadeb948),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d94a4),
	.w1(32'hbba078c8),
	.w2(32'hbbf4c71d),
	.w3(32'hbb89a7f6),
	.w4(32'hbbbc2f3e),
	.w5(32'h3b5b8ae5),
	.w6(32'hbb989d26),
	.w7(32'hbbd18d74),
	.w8(32'h3b5a1ee4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a5cea),
	.w1(32'hbad1ff60),
	.w2(32'hbb55d152),
	.w3(32'h3b7d1c5b),
	.w4(32'h3b2c8b5c),
	.w5(32'hbabc5579),
	.w6(32'hb9294009),
	.w7(32'h3ac6048b),
	.w8(32'h3995ee19),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad324f4),
	.w1(32'h3a2e4846),
	.w2(32'hbb267aac),
	.w3(32'hbb72474e),
	.w4(32'hbad35668),
	.w5(32'h3a5a2c1e),
	.w6(32'hbaf865b1),
	.w7(32'hbaff424c),
	.w8(32'hba489f95),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b23325),
	.w1(32'hb99073ae),
	.w2(32'hbaf57bfe),
	.w3(32'h3b27e85d),
	.w4(32'h3a80bb92),
	.w5(32'h3a0200e2),
	.w6(32'hba5d45ca),
	.w7(32'hb993a461),
	.w8(32'h39d68c5d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5d216),
	.w1(32'hb9eaf600),
	.w2(32'hbb330ce9),
	.w3(32'h3b29427c),
	.w4(32'h3b2569ae),
	.w5(32'h3b67894c),
	.w6(32'hba0ebb09),
	.w7(32'hb9f24f6d),
	.w8(32'h3c02f213),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07236b),
	.w1(32'h3b821bf9),
	.w2(32'hbb4127a5),
	.w3(32'hba8d5c33),
	.w4(32'hbab7c4bd),
	.w5(32'h3a3b94c0),
	.w6(32'h39a64286),
	.w7(32'hbaf2f0de),
	.w8(32'hbb0d9657),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42e6da),
	.w1(32'hbaf20586),
	.w2(32'hbb0b876a),
	.w3(32'h3a47d017),
	.w4(32'h39cbb6cd),
	.w5(32'h3ba757a7),
	.w6(32'h3a70c7c0),
	.w7(32'hbaa6a784),
	.w8(32'h3b62f195),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36628f),
	.w1(32'h3aec436a),
	.w2(32'h3b4fe950),
	.w3(32'h3b5b5e06),
	.w4(32'h3991016a),
	.w5(32'h3aa9a199),
	.w6(32'h3bb874a4),
	.w7(32'h3b0920b9),
	.w8(32'h3b125f26),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56905a),
	.w1(32'h3ba02aa7),
	.w2(32'hbab67630),
	.w3(32'hba4a69c4),
	.w4(32'h3af0d978),
	.w5(32'hbaac9737),
	.w6(32'h389f23d2),
	.w7(32'h3aaa3e0e),
	.w8(32'h3a524111),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5cf8e),
	.w1(32'hbb39f16e),
	.w2(32'hbb892ead),
	.w3(32'hbb2642d6),
	.w4(32'hbb77051c),
	.w5(32'hb87ef06c),
	.w6(32'hbae505db),
	.w7(32'hba8e22bf),
	.w8(32'h3aae430e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b004053),
	.w1(32'hbaa28790),
	.w2(32'hbb6e833e),
	.w3(32'hbb1a3eb1),
	.w4(32'hbb6d8c15),
	.w5(32'h390b03bf),
	.w6(32'hbb8be790),
	.w7(32'hbb8e1bef),
	.w8(32'h3b8280bb),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f3a60),
	.w1(32'h3b824372),
	.w2(32'hbafcd56e),
	.w3(32'h3bbd313d),
	.w4(32'h3b383911),
	.w5(32'h3b0caccd),
	.w6(32'h3bd83d3c),
	.w7(32'h39dbec69),
	.w8(32'h3b463441),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59da91),
	.w1(32'hba6aad4e),
	.w2(32'hbb6a67b1),
	.w3(32'hba8ccfea),
	.w4(32'hbb85a25f),
	.w5(32'h39aed5b3),
	.w6(32'hbb336478),
	.w7(32'hbb921bf8),
	.w8(32'h3b28f230),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52f449),
	.w1(32'h3b3f7d4d),
	.w2(32'hba201b03),
	.w3(32'h3a782137),
	.w4(32'hb8bc3bc2),
	.w5(32'h3b8f1829),
	.w6(32'h3990a5e8),
	.w7(32'hba998112),
	.w8(32'h3b5e73c2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ef2fb),
	.w1(32'hbb7cf9f5),
	.w2(32'h3b9e02e8),
	.w3(32'h3b535a0d),
	.w4(32'hb9885d40),
	.w5(32'h3a4f4d13),
	.w6(32'hbaaab624),
	.w7(32'hba832619),
	.w8(32'h3a9fcab0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab02e5e),
	.w1(32'h3a66c29e),
	.w2(32'h3a17674c),
	.w3(32'h3af36e40),
	.w4(32'h398f11c0),
	.w5(32'h3a2877ba),
	.w6(32'h3a645dbf),
	.w7(32'hba12f006),
	.w8(32'h3afb0906),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa96fa5),
	.w1(32'hb9bb3414),
	.w2(32'hbb807c0b),
	.w3(32'hba9c53a5),
	.w4(32'hbb5232e4),
	.w5(32'h3af33050),
	.w6(32'hbb227856),
	.w7(32'hbb987acf),
	.w8(32'h3ab11272),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e5ad0),
	.w1(32'hbb118f69),
	.w2(32'hbb9665a5),
	.w3(32'hbae4490a),
	.w4(32'hbba7f609),
	.w5(32'h3b0d1201),
	.w6(32'hbba4195f),
	.w7(32'hbbc50cc6),
	.w8(32'h3aa6678b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc096e),
	.w1(32'hbb8dc92b),
	.w2(32'hbb7a04fd),
	.w3(32'hba6fd097),
	.w4(32'hbb18b4db),
	.w5(32'h3aa6d53a),
	.w6(32'hbb167c8e),
	.w7(32'hbab10c70),
	.w8(32'h398ebec3),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7616a3),
	.w1(32'h3b07ce53),
	.w2(32'h3b3a2e17),
	.w3(32'h3b8c127d),
	.w4(32'h3b84ec19),
	.w5(32'h3b3ae754),
	.w6(32'h3b4d1bee),
	.w7(32'h3b9bc67b),
	.w8(32'h3a5dae71),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0723db),
	.w1(32'h3b844af9),
	.w2(32'h3a26822b),
	.w3(32'h3b42cd33),
	.w4(32'h3a267750),
	.w5(32'hba1580ec),
	.w6(32'h3b4fab9e),
	.w7(32'h3a98c968),
	.w8(32'hba9179c0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ff87),
	.w1(32'hbbd9cf72),
	.w2(32'hbbbc5a2b),
	.w3(32'hbaf9a9bb),
	.w4(32'hbbea559e),
	.w5(32'hbb11d794),
	.w6(32'hbbd49c87),
	.w7(32'hbbe2db1a),
	.w8(32'hbb826e74),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb489d07),
	.w1(32'hb91241c8),
	.w2(32'hba78bfa3),
	.w3(32'hba2fa4ed),
	.w4(32'hba362c24),
	.w5(32'h3baeb56c),
	.w6(32'hbab7ec00),
	.w7(32'hba0c786f),
	.w8(32'h3b4989eb),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b010a7f),
	.w1(32'hbb119aff),
	.w2(32'hbafd366d),
	.w3(32'h3a0f787f),
	.w4(32'hbaaed81b),
	.w5(32'hba6af478),
	.w6(32'hbb335077),
	.w7(32'h37989697),
	.w8(32'hbb0559d6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa23f08),
	.w1(32'hbb133dee),
	.w2(32'hbb2ffc30),
	.w3(32'hbadea264),
	.w4(32'hbae388d3),
	.w5(32'h38cc7a4a),
	.w6(32'hbb31c7c6),
	.w7(32'hbb538214),
	.w8(32'hba6c7c57),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a104f),
	.w1(32'hbb4eed19),
	.w2(32'hbb30d112),
	.w3(32'hb9e93780),
	.w4(32'hba9a1ccb),
	.w5(32'h3b292740),
	.w6(32'hbaca937d),
	.w7(32'hbade4546),
	.w8(32'h3b407122),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5fc5),
	.w1(32'h3b0b58b8),
	.w2(32'hba590338),
	.w3(32'h3a4007a5),
	.w4(32'h3b014f0c),
	.w5(32'hba2ff6d0),
	.w6(32'hb9ffcc86),
	.w7(32'hba3c9a46),
	.w8(32'hbb3823a6),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8b1e8),
	.w1(32'h3a8840b9),
	.w2(32'hb92bd530),
	.w3(32'h3aac552e),
	.w4(32'h399ba172),
	.w5(32'h3a984827),
	.w6(32'hb906a25d),
	.w7(32'h3899de2a),
	.w8(32'h3acd0bfc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8242fc),
	.w1(32'h3aea6fbb),
	.w2(32'h3b49ea56),
	.w3(32'h3a1b661f),
	.w4(32'h3afd064e),
	.w5(32'h3bac7dd7),
	.w6(32'h3a31d16f),
	.w7(32'h3afdd6c5),
	.w8(32'h3b58edb7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08fcae),
	.w1(32'h3b074773),
	.w2(32'h3b72efdf),
	.w3(32'h3b35a9d7),
	.w4(32'h3ba0d8c5),
	.w5(32'hbb31ddfe),
	.w6(32'h3b1ffd8c),
	.w7(32'h3bc037ec),
	.w8(32'hbbaaffe3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb808d4b),
	.w1(32'h3ae08e4c),
	.w2(32'h3afdc61d),
	.w3(32'h3a8bb647),
	.w4(32'h3950c75f),
	.w5(32'hbb7618b1),
	.w6(32'h3ab15940),
	.w7(32'h3a378191),
	.w8(32'hba4e639e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41e3e1),
	.w1(32'hbaa1c59b),
	.w2(32'hbace8654),
	.w3(32'hbb00ca12),
	.w4(32'hbb470f6d),
	.w5(32'h3b0a69b8),
	.w6(32'hbac1f1d1),
	.w7(32'hba14e47f),
	.w8(32'h3a9197ff),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab44e91),
	.w1(32'hbb5268f7),
	.w2(32'hbb8c46ea),
	.w3(32'h3a1e0b55),
	.w4(32'hbbb43529),
	.w5(32'h3ac2cb86),
	.w6(32'hbb291934),
	.w7(32'hbba2ea2d),
	.w8(32'h3afcebb4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dab883),
	.w1(32'h3b2a228c),
	.w2(32'hba86ef4b),
	.w3(32'h3b8d6f9c),
	.w4(32'hbafa863f),
	.w5(32'h3b8525e6),
	.w6(32'h3b0f80b6),
	.w7(32'hbb03d238),
	.w8(32'h3b98c30a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbab4e2),
	.w1(32'h3bf11a62),
	.w2(32'h3b9d12b2),
	.w3(32'h3bcc17eb),
	.w4(32'h3b8340c2),
	.w5(32'hbb4d97bb),
	.w6(32'h3c0baa94),
	.w7(32'h3b9ce345),
	.w8(32'h39fa5f57),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9949916),
	.w1(32'hbb3fc3dd),
	.w2(32'hbb82df8c),
	.w3(32'hbbb0c304),
	.w4(32'hbb83d216),
	.w5(32'hbabc32ce),
	.w6(32'hbb9b3f23),
	.w7(32'hbb935c87),
	.w8(32'hbb05c5ec),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab566da),
	.w1(32'hbb899fea),
	.w2(32'hbbb23e15),
	.w3(32'hbb86d90a),
	.w4(32'hbb5e9b7f),
	.w5(32'hbb84de14),
	.w6(32'hbb904006),
	.w7(32'hbb78628c),
	.w8(32'h3a5d030f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34372a),
	.w1(32'h3b93824f),
	.w2(32'h3bb9eaf2),
	.w3(32'hbace70e4),
	.w4(32'hb9a41e1c),
	.w5(32'h3a7c6701),
	.w6(32'h3b55b7f3),
	.w7(32'hba68cad0),
	.w8(32'h3a0d95e3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6941bd),
	.w1(32'hbb4b2284),
	.w2(32'hba96680c),
	.w3(32'hba74c923),
	.w4(32'h3a82a437),
	.w5(32'hbaf305de),
	.w6(32'h3ae7d1f7),
	.w7(32'h3abc648c),
	.w8(32'hbb806f5b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb887601),
	.w1(32'hbb3ad232),
	.w2(32'hbb87e05e),
	.w3(32'hbb854d23),
	.w4(32'hbb21d90d),
	.w5(32'hba33c60b),
	.w6(32'h3a2dc32e),
	.w7(32'hbb7787ee),
	.w8(32'hbad3a69b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89fba2),
	.w1(32'hbae021ee),
	.w2(32'hbb9f4695),
	.w3(32'hbad92acc),
	.w4(32'hbb81f70f),
	.w5(32'hb9ca7ca1),
	.w6(32'hbb85a718),
	.w7(32'hbbbe7ee2),
	.w8(32'h3b0ac10f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa18380),
	.w1(32'hb9d57288),
	.w2(32'h3ae53e2a),
	.w3(32'h3ac50671),
	.w4(32'h3a097516),
	.w5(32'h3a8037d9),
	.w6(32'h3aa861cb),
	.w7(32'h3b4f2257),
	.w8(32'hba6f5032),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80f8f88),
	.w1(32'hba048748),
	.w2(32'h37893af2),
	.w3(32'hba9dc16d),
	.w4(32'hbb17f2cc),
	.w5(32'hb98a592b),
	.w6(32'hbb929e5f),
	.w7(32'hbac1c4e5),
	.w8(32'h3bc6c3ec),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad38e0f),
	.w1(32'h39fabc75),
	.w2(32'h3abba03d),
	.w3(32'hbb2728d7),
	.w4(32'hb9a69d4a),
	.w5(32'h3a43a8c1),
	.w6(32'h3b79064a),
	.w7(32'hba21921d),
	.w8(32'h3acfa58c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2abdfc),
	.w1(32'h3b7400aa),
	.w2(32'h39d4ba55),
	.w3(32'h3ba056b0),
	.w4(32'h3a83b521),
	.w5(32'hbaf63c4d),
	.w6(32'h3b581dd6),
	.w7(32'h3a047eda),
	.w8(32'hb9599fbb),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432c91),
	.w1(32'h3b69c07f),
	.w2(32'h3b5d08b5),
	.w3(32'hbba9cc48),
	.w4(32'hbac0fef4),
	.w5(32'h377dfc5f),
	.w6(32'hba8a896c),
	.w7(32'h3ad787b2),
	.w8(32'hbb061b69),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1492f7),
	.w1(32'hbafcc3ff),
	.w2(32'hba289054),
	.w3(32'hbb1c5c8c),
	.w4(32'h3984cb12),
	.w5(32'hbafc4e04),
	.w6(32'hbbad93f0),
	.w7(32'hbb3deb0d),
	.w8(32'hbb579cac),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f2da3),
	.w1(32'hbb10a1cf),
	.w2(32'hba503ca4),
	.w3(32'hbac2fc72),
	.w4(32'hba71beb6),
	.w5(32'h3bd55ee4),
	.w6(32'hbad92214),
	.w7(32'hba0434e8),
	.w8(32'h3c0480fb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6da37),
	.w1(32'h3b0dd0d7),
	.w2(32'hb9b9f757),
	.w3(32'h3b3f5c6b),
	.w4(32'hbada780b),
	.w5(32'hbb2f88fc),
	.w6(32'h39cfaac5),
	.w7(32'hb99e158c),
	.w8(32'hbb150665),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2eb86e),
	.w1(32'h3b820de2),
	.w2(32'h3b561c1c),
	.w3(32'h3b82e7fb),
	.w4(32'h3bc1d6e9),
	.w5(32'hb932b2ad),
	.w6(32'h3a7b7619),
	.w7(32'h3ac81cf4),
	.w8(32'hb893503d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0730f),
	.w1(32'h39aa156b),
	.w2(32'hbb1efad3),
	.w3(32'h3afdd4b4),
	.w4(32'hba1f7f18),
	.w5(32'h3b19ae2e),
	.w6(32'hbbe2d806),
	.w7(32'hbb740ff3),
	.w8(32'h3b6a4796),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b276c67),
	.w1(32'h3b9f20f6),
	.w2(32'h3b6f6dab),
	.w3(32'h3b7258f3),
	.w4(32'h3b3d6278),
	.w5(32'h3c04b760),
	.w6(32'h3bdb070a),
	.w7(32'h3b5caf49),
	.w8(32'h3c20c7a7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26a1e0),
	.w1(32'h3c0cc8d0),
	.w2(32'h3b53a511),
	.w3(32'h3b17832d),
	.w4(32'h39ebb8ac),
	.w5(32'hbb057de7),
	.w6(32'h3ba6927c),
	.w7(32'h3b950730),
	.w8(32'h389a1c16),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1339c0),
	.w1(32'h3b652690),
	.w2(32'hb9b8f114),
	.w3(32'h3af2e5d7),
	.w4(32'h39037c73),
	.w5(32'h3b2b2f49),
	.w6(32'h3ab499bf),
	.w7(32'hba8027f4),
	.w8(32'h3b1878ab),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0359e6),
	.w1(32'h3b46b46b),
	.w2(32'h3b8b4bb2),
	.w3(32'h3b11d808),
	.w4(32'h3b25f490),
	.w5(32'hbb61878c),
	.w6(32'h3b50aa78),
	.w7(32'h3b779d8d),
	.w8(32'hbbaf362e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96dd13),
	.w1(32'hbae0cc68),
	.w2(32'hbaa09d8a),
	.w3(32'h391f8166),
	.w4(32'hbb77574f),
	.w5(32'h3b23db2a),
	.w6(32'hbab4ab25),
	.w7(32'hbb4ae825),
	.w8(32'h3b533e33),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af23b48),
	.w1(32'h39f5d68e),
	.w2(32'h39792e84),
	.w3(32'h39dda575),
	.w4(32'hba3c9a0f),
	.w5(32'h3b776371),
	.w6(32'h3b033c57),
	.w7(32'h3a05a5c0),
	.w8(32'h3b27e891),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b578f23),
	.w1(32'h3b1ffc71),
	.w2(32'hbaac426e),
	.w3(32'h3b6e47d9),
	.w4(32'hb8313f87),
	.w5(32'hba2860ba),
	.w6(32'hb9836cfa),
	.w7(32'hbab548d6),
	.w8(32'h3a5247c8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acae614),
	.w1(32'h399c60b4),
	.w2(32'hbb1777a2),
	.w3(32'hb91d60dd),
	.w4(32'hbab9a294),
	.w5(32'h39bd492d),
	.w6(32'hbb3e28a8),
	.w7(32'hba0a51bd),
	.w8(32'hba32edb1),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a69ca),
	.w1(32'hbb7c4d86),
	.w2(32'hbb3322a3),
	.w3(32'hbb16eaa1),
	.w4(32'hbb8343f6),
	.w5(32'h3bcb101d),
	.w6(32'hbba97eff),
	.w7(32'hbb4f0267),
	.w8(32'h3bd8f825),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d3a4b),
	.w1(32'hbaa73e85),
	.w2(32'h3b0149d7),
	.w3(32'h3aa771dc),
	.w4(32'h38f8bf3f),
	.w5(32'hbad9499d),
	.w6(32'hbaf38c08),
	.w7(32'hbb0acecc),
	.w8(32'hbb0b8ea0),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cfaff),
	.w1(32'hbb657fbe),
	.w2(32'hbb599151),
	.w3(32'hbb2af295),
	.w4(32'hbb0eadaf),
	.w5(32'hbab23f52),
	.w6(32'hbb747d77),
	.w7(32'hbb3be443),
	.w8(32'h3a731931),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2f397),
	.w1(32'h3a915262),
	.w2(32'hbabceb99),
	.w3(32'hb7d8a772),
	.w4(32'hbae4cc73),
	.w5(32'hbb1ff75d),
	.w6(32'h3981ffe1),
	.w7(32'hbad27427),
	.w8(32'hbaf5e91f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec3220),
	.w1(32'h3a9ca266),
	.w2(32'h3a6d96f5),
	.w3(32'hba7cde99),
	.w4(32'hbaac93b5),
	.w5(32'h3b7b6244),
	.w6(32'hba7cb8a0),
	.w7(32'hbaca8e8c),
	.w8(32'h3b9ebd27),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9057f4),
	.w1(32'h3aed404a),
	.w2(32'h3b4b3176),
	.w3(32'h3aabf5df),
	.w4(32'h3b71ed6e),
	.w5(32'h3abec4fd),
	.w6(32'h3a8fd044),
	.w7(32'h3a966991),
	.w8(32'h3b32285f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d169a),
	.w1(32'h3a8b851c),
	.w2(32'hba2a0451),
	.w3(32'h3aaf5974),
	.w4(32'hbae83182),
	.w5(32'hbb836f8b),
	.w6(32'h3b227f11),
	.w7(32'hbac0e7c5),
	.w8(32'hbb8bce33),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956d7fc),
	.w1(32'h3bc42920),
	.w2(32'h3c0128b1),
	.w3(32'h3b25ac5e),
	.w4(32'h3bbd4c47),
	.w5(32'h3b02c809),
	.w6(32'hb826ea60),
	.w7(32'h3bcf921b),
	.w8(32'h3aa2e55b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3df003),
	.w1(32'hb9bb84df),
	.w2(32'hbaabc0fa),
	.w3(32'hbbadfa09),
	.w4(32'hbb8ecbce),
	.w5(32'h3b99b534),
	.w6(32'hbb719556),
	.w7(32'hbb6e0904),
	.w8(32'h3bbbe28b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b960858),
	.w1(32'h3ad1fc29),
	.w2(32'hba9040cb),
	.w3(32'h3aa672d7),
	.w4(32'hbade8dcb),
	.w5(32'h38be2241),
	.w6(32'h39c8a060),
	.w7(32'hbaabac84),
	.w8(32'h3a1b7f80),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb053970),
	.w1(32'hb9a14993),
	.w2(32'h3a1b9834),
	.w3(32'h3a57b700),
	.w4(32'hba9c7099),
	.w5(32'hba1ccdfd),
	.w6(32'h3ad6b4bb),
	.w7(32'h3acac27d),
	.w8(32'h3a4f701b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986c072),
	.w1(32'h3b10139d),
	.w2(32'h3ada0e3b),
	.w3(32'h3ac2c8b2),
	.w4(32'h3a036b22),
	.w5(32'h3ad67d10),
	.w6(32'h3ae3d021),
	.w7(32'h3a846a5a),
	.w8(32'h3b4fa6c8),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b268a6c),
	.w1(32'h3af4c22c),
	.w2(32'hb7c71e65),
	.w3(32'h39d44873),
	.w4(32'h3a94ec30),
	.w5(32'hb942cfea),
	.w6(32'h3b17b330),
	.w7(32'hb8ea94f0),
	.w8(32'hbb0cb820),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f2162),
	.w1(32'hbb87f825),
	.w2(32'hbb964c38),
	.w3(32'hbaa8a785),
	.w4(32'hbb76c50f),
	.w5(32'h3bc4db2b),
	.w6(32'hbb9fca29),
	.w7(32'hbb9c1899),
	.w8(32'h3be3cc9b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b8d04),
	.w1(32'hbb9ad0a9),
	.w2(32'hba676efb),
	.w3(32'h39b282e9),
	.w4(32'hbb2aa20a),
	.w5(32'hbb587cf6),
	.w6(32'hbb46067c),
	.w7(32'hba22f75a),
	.w8(32'hbb400102),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39939ab4),
	.w1(32'h3c16460d),
	.w2(32'h3bb9a82e),
	.w3(32'h3bf367c4),
	.w4(32'h3b6f7ac3),
	.w5(32'hba9960c3),
	.w6(32'h3bcc7a7f),
	.w7(32'h3b487090),
	.w8(32'hbb65c60c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb451b1a),
	.w1(32'h36034bd1),
	.w2(32'hbb46837a),
	.w3(32'hba93f811),
	.w4(32'hbaf78c04),
	.w5(32'hb9281576),
	.w6(32'h3a7976eb),
	.w7(32'hbb50317d),
	.w8(32'hbb09bb9b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a3a65),
	.w1(32'hba812b7a),
	.w2(32'hbaf39808),
	.w3(32'h38ad23fb),
	.w4(32'hbb18bd5a),
	.w5(32'h3b00fb08),
	.w6(32'hbbd9d38e),
	.w7(32'hbbc37737),
	.w8(32'h3b6f5990),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933230f),
	.w1(32'h3af65493),
	.w2(32'h3b1cfbd8),
	.w3(32'h3b43a5b3),
	.w4(32'h3b3d32a0),
	.w5(32'hbaa5d407),
	.w6(32'h3b74e3a7),
	.w7(32'h3b28a6b3),
	.w8(32'hbb4cc3ef),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5eacee),
	.w1(32'hba0220d4),
	.w2(32'h3a35b723),
	.w3(32'hb9d3e122),
	.w4(32'hbb28550c),
	.w5(32'hbb923f36),
	.w6(32'hbaadbe11),
	.w7(32'h3a867f42),
	.w8(32'hbbb8e3e6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf08c22),
	.w1(32'h3af0b00a),
	.w2(32'hba197053),
	.w3(32'hbb09ac86),
	.w4(32'hbaf5d5f5),
	.w5(32'hbadfae54),
	.w6(32'hba5ab93e),
	.w7(32'hba99216a),
	.w8(32'hba27f357),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb929b140),
	.w1(32'h3a03ec21),
	.w2(32'hbb4b107b),
	.w3(32'hbb2d8bdf),
	.w4(32'hbadafe17),
	.w5(32'h3b80b97a),
	.w6(32'hbb27ed06),
	.w7(32'hbb6f7c6a),
	.w8(32'h3b3f4569),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5177d),
	.w1(32'hb8c53f9a),
	.w2(32'hbafe6282),
	.w3(32'h3aa9cd4b),
	.w4(32'hba8f5397),
	.w5(32'hbb9094b0),
	.w6(32'hba4430b5),
	.w7(32'hbac0914c),
	.w8(32'hbbc6c97b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66f325),
	.w1(32'hba461076),
	.w2(32'hbb2fcd22),
	.w3(32'hbac0deac),
	.w4(32'hbb1d9654),
	.w5(32'hbabc9449),
	.w6(32'hbb2a5563),
	.w7(32'hbb00ca34),
	.w8(32'hbb3609d6),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafad037),
	.w1(32'hb897c9d9),
	.w2(32'hba53255e),
	.w3(32'h39697d1c),
	.w4(32'hba8b21ee),
	.w5(32'hb96cb0fc),
	.w6(32'hb9dd66f2),
	.w7(32'hb931b4b0),
	.w8(32'hb9d5d5d5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38399840),
	.w1(32'h391d2053),
	.w2(32'hbb0b40c4),
	.w3(32'hb90e845f),
	.w4(32'hbaca21fd),
	.w5(32'h3ac79c2a),
	.w6(32'hbb0a6878),
	.w7(32'hbb02fdc9),
	.w8(32'h398a251b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39939125),
	.w1(32'hba8521bd),
	.w2(32'h393e12af),
	.w3(32'hb965625a),
	.w4(32'hbb23b84e),
	.w5(32'h3b8f8113),
	.w6(32'hbb1e619a),
	.w7(32'hbb29bb45),
	.w8(32'h3bbcc1c4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93bc77),
	.w1(32'h3aca6ae4),
	.w2(32'h3a6ade14),
	.w3(32'h3b11de95),
	.w4(32'hba57ece4),
	.w5(32'hbb86663f),
	.w6(32'h3a55927d),
	.w7(32'h3a167549),
	.w8(32'hbbc9f635),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1f908),
	.w1(32'hbb8bd152),
	.w2(32'h3a9dee91),
	.w3(32'h3a3390c4),
	.w4(32'h3a12f284),
	.w5(32'hbae4139b),
	.w6(32'hbb3b96ae),
	.w7(32'hbaed8ba5),
	.w8(32'hbb2dbe6c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4336fa),
	.w1(32'hbb1ac2b5),
	.w2(32'hbb197991),
	.w3(32'hbab5f387),
	.w4(32'hbb0dedde),
	.w5(32'h3b5ece57),
	.w6(32'hbb1f1898),
	.w7(32'hbb61304d),
	.w8(32'h3ae58523),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941b982),
	.w1(32'hb9f3149d),
	.w2(32'h3a6ea40b),
	.w3(32'h3ab0b64f),
	.w4(32'h3aab4894),
	.w5(32'hbb62a63d),
	.w6(32'h3ab4ee75),
	.w7(32'h3a81f3dd),
	.w8(32'hbbea5c12),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbded4cd),
	.w1(32'hbc1296be),
	.w2(32'hbc247289),
	.w3(32'hbbbe1b94),
	.w4(32'hbbd3bc83),
	.w5(32'h3b7a2cab),
	.w6(32'hbc4caac1),
	.w7(32'hbc14353e),
	.w8(32'h3b339dd5),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c8992),
	.w1(32'hb9b38b81),
	.w2(32'h3a2147ac),
	.w3(32'h3b8e4a5f),
	.w4(32'h3b81c00b),
	.w5(32'h3b8704a7),
	.w6(32'h3b1cfc25),
	.w7(32'h3b3f82bb),
	.w8(32'h3bd95479),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbace63),
	.w1(32'h3bd05a33),
	.w2(32'h3ae82deb),
	.w3(32'h3ba216f5),
	.w4(32'hbabc69e4),
	.w5(32'h3b855f38),
	.w6(32'h3b579f01),
	.w7(32'hbad6e1f0),
	.w8(32'h3b9f692c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19d121),
	.w1(32'h3a0c3027),
	.w2(32'h3a477499),
	.w3(32'h3b7a610a),
	.w4(32'h3a24329d),
	.w5(32'h3a4b8af4),
	.w6(32'hba569572),
	.w7(32'h39b54bb9),
	.w8(32'h3a7d8ad6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4a7de),
	.w1(32'h3a4b65b0),
	.w2(32'hbac82786),
	.w3(32'h3acf926c),
	.w4(32'h3ad60b81),
	.w5(32'h3b11ecab),
	.w6(32'hba058a72),
	.w7(32'hb9180447),
	.w8(32'h3b59e638),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbfcb4),
	.w1(32'h38cf11e5),
	.w2(32'hba99f664),
	.w3(32'h39c79bf2),
	.w4(32'hbaae5763),
	.w5(32'h3aa34953),
	.w6(32'hb8cf8d01),
	.w7(32'hba9df583),
	.w8(32'hb9a29595),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf777f1),
	.w1(32'hbb91e0a8),
	.w2(32'hbbc07a9d),
	.w3(32'hbb4ab067),
	.w4(32'hbbdb5a79),
	.w5(32'hba0ba98d),
	.w6(32'hbb44698d),
	.w7(32'hbbc602a7),
	.w8(32'hba9cf6fe),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9326f3),
	.w1(32'h3a396385),
	.w2(32'hbb082fab),
	.w3(32'h3a8b2b49),
	.w4(32'h3a8c0d65),
	.w5(32'h3aa396e7),
	.w6(32'h3b3ac1c2),
	.w7(32'h3b1d1c04),
	.w8(32'h39c7a3c1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4508c5),
	.w1(32'hba209ca6),
	.w2(32'hbb705994),
	.w3(32'hbb172cd2),
	.w4(32'hbb4ec314),
	.w5(32'h3b7e60a8),
	.w6(32'hba718196),
	.w7(32'hbb899c14),
	.w8(32'h3b264cdb),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0d35e),
	.w1(32'h3ac0d11e),
	.w2(32'hbb261d16),
	.w3(32'h3b89e2f0),
	.w4(32'h3a1c47f3),
	.w5(32'hb9c0f2d6),
	.w6(32'h3bb86fe8),
	.w7(32'hba8cffe2),
	.w8(32'hba0e2e11),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07657f),
	.w1(32'hbb20b7a7),
	.w2(32'hbb313274),
	.w3(32'hba1db21a),
	.w4(32'hbaf4036a),
	.w5(32'hb9658d9a),
	.w6(32'hba998b54),
	.w7(32'hba3b0c66),
	.w8(32'hbac1018a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ccb9a),
	.w1(32'hba918da2),
	.w2(32'hbb03c50d),
	.w3(32'hba0e61af),
	.w4(32'hbb4d61c7),
	.w5(32'h3b183916),
	.w6(32'h3a3cfb54),
	.w7(32'hbae1b1f2),
	.w8(32'hba2fdf70),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba931c4e),
	.w1(32'h39479f2e),
	.w2(32'h3a5f364b),
	.w3(32'h39ec160c),
	.w4(32'hba9ef32c),
	.w5(32'hbb648e67),
	.w6(32'h3a91ea2c),
	.w7(32'h39982e98),
	.w8(32'hbb4146cb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13b1ca),
	.w1(32'h3b686670),
	.w2(32'hb8f6bb7b),
	.w3(32'hbb5bf9f2),
	.w4(32'h3a845107),
	.w5(32'hbab1d629),
	.w6(32'hbad7d77b),
	.w7(32'hb6f55d29),
	.w8(32'hbae977ce),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb697f7d),
	.w1(32'h3a4378f7),
	.w2(32'h39c632f9),
	.w3(32'h3a4e5108),
	.w4(32'h3a28d29f),
	.w5(32'hba0e53e9),
	.w6(32'h3b8521ba),
	.w7(32'hbb43a728),
	.w8(32'hba10b6dc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95768f0),
	.w1(32'hba71c5d2),
	.w2(32'hba2dc254),
	.w3(32'hba1f9979),
	.w4(32'hb9dc54cd),
	.w5(32'hbaa2a201),
	.w6(32'hba9a6572),
	.w7(32'hba817b18),
	.w8(32'hbae6c443),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa10df8),
	.w1(32'hba70eb36),
	.w2(32'hb9a511d5),
	.w3(32'hb8d18dce),
	.w4(32'hba763a59),
	.w5(32'hba6186fe),
	.w6(32'hbac8a75f),
	.w7(32'hba0e00cb),
	.w8(32'hbabac602),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99938da),
	.w1(32'hba2845c9),
	.w2(32'hbacccfa1),
	.w3(32'hba8567fe),
	.w4(32'hb927c0f5),
	.w5(32'hba9e0890),
	.w6(32'hba2fee86),
	.w7(32'hbaa40de8),
	.w8(32'hba3c1dc6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e6cba),
	.w1(32'h3a88874f),
	.w2(32'h3a93b13a),
	.w3(32'hbabfc19c),
	.w4(32'hbaaf3eae),
	.w5(32'h3a34b28a),
	.w6(32'hba2e2198),
	.w7(32'hb9db14ad),
	.w8(32'h39df012f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f179a),
	.w1(32'h39e30c0b),
	.w2(32'h39cb018f),
	.w3(32'hba57780d),
	.w4(32'h39e07213),
	.w5(32'hbabe3137),
	.w6(32'hb9e8bd3f),
	.w7(32'h39312802),
	.w8(32'hbb14e103),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb164e96),
	.w1(32'hbaec7527),
	.w2(32'hbb037a86),
	.w3(32'hb9838a17),
	.w4(32'hba8c56dc),
	.w5(32'hba7dff9f),
	.w6(32'hbb069756),
	.w7(32'hbaf40e33),
	.w8(32'hb814e566),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba922040),
	.w1(32'hbaeac3bc),
	.w2(32'hbafe137d),
	.w3(32'hbae63264),
	.w4(32'hbaafa76f),
	.w5(32'hbaa00adb),
	.w6(32'hbb1e2051),
	.w7(32'hbaef6691),
	.w8(32'hbb16cc80),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6f57a),
	.w1(32'hbabbba3d),
	.w2(32'hba99c766),
	.w3(32'hba33b284),
	.w4(32'hba863ea8),
	.w5(32'h3a4ff49e),
	.w6(32'hbab04732),
	.w7(32'hba97cc4e),
	.w8(32'h3a5228c1),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3f601),
	.w1(32'hb9fb4198),
	.w2(32'hb93da828),
	.w3(32'h39c4aaff),
	.w4(32'hbb016904),
	.w5(32'h3a28fc23),
	.w6(32'h3a0a05db),
	.w7(32'hba67aece),
	.w8(32'h39c13759),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df438a),
	.w1(32'hb9df955a),
	.w2(32'hb7cd3f36),
	.w3(32'h39aed533),
	.w4(32'h39b3d6c5),
	.w5(32'hbad29157),
	.w6(32'hb91af73f),
	.w7(32'h38afc50d),
	.w8(32'hbae0f570),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafb8e7),
	.w1(32'hbac083ea),
	.w2(32'hba7b3298),
	.w3(32'hba59769c),
	.w4(32'hba1c92ef),
	.w5(32'hb9cc6680),
	.w6(32'hbae2f6dc),
	.w7(32'hbabcfa29),
	.w8(32'hb7ce4ce7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9be09),
	.w1(32'hba0e119e),
	.w2(32'h3a15914b),
	.w3(32'hb9f703d2),
	.w4(32'h3a760ecb),
	.w5(32'hba582d6a),
	.w6(32'hb9e9184a),
	.w7(32'h398ed549),
	.w8(32'hb9fc894b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a616dd),
	.w1(32'hb9a50574),
	.w2(32'hba8732ec),
	.w3(32'hbad1b1d0),
	.w4(32'hba8a6e99),
	.w5(32'hbac42688),
	.w6(32'hba85e480),
	.w7(32'hb8cbf46d),
	.w8(32'hbb3d99cb),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0476b7),
	.w1(32'hba5d4379),
	.w2(32'h3a838be6),
	.w3(32'h38a46904),
	.w4(32'h3a9e79cc),
	.w5(32'h3b3d489c),
	.w6(32'hb9cc0e4f),
	.w7(32'h392542a2),
	.w8(32'h3b2b0d1b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e3bd9),
	.w1(32'h3af636ea),
	.w2(32'h3b2af712),
	.w3(32'h3ae31ebf),
	.w4(32'h3b3cb900),
	.w5(32'h3abe54c0),
	.w6(32'h3a4a7725),
	.w7(32'h3b005ca6),
	.w8(32'h3a8efa09),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e4c390),
	.w1(32'h3a66882c),
	.w2(32'h3a01e028),
	.w3(32'h3ad4e5d3),
	.w4(32'h3a2d35b6),
	.w5(32'h39f54e6d),
	.w6(32'h3a86b7b5),
	.w7(32'h39ab63f0),
	.w8(32'hb9807175),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394716f1),
	.w1(32'h390e8d8e),
	.w2(32'hba0d3574),
	.w3(32'hb95bc8e2),
	.w4(32'hbac2d4ce),
	.w5(32'hba3c06be),
	.w6(32'hba25aae1),
	.w7(32'hbaab7146),
	.w8(32'hbadf31e3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa27af),
	.w1(32'hba988b75),
	.w2(32'h3a5e045d),
	.w3(32'hba88b257),
	.w4(32'h399b1f99),
	.w5(32'h3acfa90d),
	.w6(32'hbab9e789),
	.w7(32'hb908e3e1),
	.w8(32'h3a87bd7b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78b3a5),
	.w1(32'h3a8f3ec0),
	.w2(32'h3a76375f),
	.w3(32'h3ab7b09d),
	.w4(32'h3ac01030),
	.w5(32'hba9342e2),
	.w6(32'h3a644ac6),
	.w7(32'h3a87da25),
	.w8(32'h39e36148),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77ca5b),
	.w1(32'hb7a67b23),
	.w2(32'h388ad145),
	.w3(32'h39cbfe75),
	.w4(32'h3a2fd976),
	.w5(32'hba851092),
	.w6(32'h3a1316e4),
	.w7(32'h3a0f3b4a),
	.w8(32'hba04a88f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3b4f9),
	.w1(32'hb9bdbca2),
	.w2(32'h397b687b),
	.w3(32'hba94ff1e),
	.w4(32'hb72ab656),
	.w5(32'hbaec89dd),
	.w6(32'hba9fb4ea),
	.w7(32'hba806cbe),
	.w8(32'hbb03db1b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa337c4),
	.w1(32'hba727a75),
	.w2(32'hba839585),
	.w3(32'hbaea7fae),
	.w4(32'hba93de76),
	.w5(32'h3a692870),
	.w6(32'hba9c8685),
	.w7(32'hba86b7f0),
	.w8(32'hb75bf96e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eb15de),
	.w1(32'hb9ab9d36),
	.w2(32'hb97d66c9),
	.w3(32'h3895a796),
	.w4(32'h3a0b5098),
	.w5(32'hba778f56),
	.w6(32'hb9b8ed30),
	.w7(32'hb9810b19),
	.w8(32'hba867820),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52240c),
	.w1(32'hbac2621b),
	.w2(32'hbaa4ccce),
	.w3(32'hbae88435),
	.w4(32'hba7e74f3),
	.w5(32'hb93d1215),
	.w6(32'hba839771),
	.w7(32'hbaa3e40d),
	.w8(32'hb8e2a52c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6e85c),
	.w1(32'h39a84b9c),
	.w2(32'h399d526d),
	.w3(32'h3a084733),
	.w4(32'hba556625),
	.w5(32'h392465cb),
	.w6(32'h39d0c63f),
	.w7(32'hb84ef10e),
	.w8(32'h39cf3f0e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a508f97),
	.w1(32'h3982fe23),
	.w2(32'hba20d3ea),
	.w3(32'hb9dacdb6),
	.w4(32'h3a401ce2),
	.w5(32'h3a1b4607),
	.w6(32'hba81637a),
	.w7(32'hb96c4691),
	.w8(32'h38dcf539),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b6b4c),
	.w1(32'h39a949d3),
	.w2(32'h3a857d7a),
	.w3(32'h398a8ae5),
	.w4(32'h3960690c),
	.w5(32'hb73f1b46),
	.w6(32'h39a4cc0e),
	.w7(32'h39136ebe),
	.w8(32'h3a0b2a16),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c479f),
	.w1(32'h3ab60c3c),
	.w2(32'h3a9d5088),
	.w3(32'hba1984d1),
	.w4(32'hbab88abb),
	.w5(32'hb93b2759),
	.w6(32'hb7febeef),
	.w7(32'hb951fba0),
	.w8(32'h39fd0370),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b1e9b),
	.w1(32'h388f01b7),
	.w2(32'h39e8796c),
	.w3(32'h3a087bf8),
	.w4(32'h3a40aff2),
	.w5(32'h3a5fe7a0),
	.w6(32'h38f24285),
	.w7(32'h3996c9f9),
	.w8(32'h3923dfea),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c628f1),
	.w1(32'h3b1e3f95),
	.w2(32'h3b04cdc4),
	.w3(32'hba3a36e5),
	.w4(32'h3ab46ece),
	.w5(32'h3b1d4796),
	.w6(32'hb97e9825),
	.w7(32'hb934b743),
	.w8(32'h3ad869da),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule