module layer_8_featuremap_206(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3107d),
	.w1(32'h3a42d733),
	.w2(32'h3b2dad92),
	.w3(32'h3b1f4ff5),
	.w4(32'h3c78ffd0),
	.w5(32'h3c0b1d4a),
	.w6(32'h3c1771e9),
	.w7(32'h3c6bd5a5),
	.w8(32'h3ccb7d09),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbee21b),
	.w1(32'hba18a306),
	.w2(32'hbb7e97e8),
	.w3(32'h3c2579b7),
	.w4(32'hbb2c6a89),
	.w5(32'hbbc673c6),
	.w6(32'h3a9741f4),
	.w7(32'hbb90e64f),
	.w8(32'hbbe7c860),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af57e3e),
	.w1(32'h3bb4beb7),
	.w2(32'h3be74308),
	.w3(32'h3b92edca),
	.w4(32'h3b056d53),
	.w5(32'h3b92b1ec),
	.w6(32'h3cb012e9),
	.w7(32'h3c1a7049),
	.w8(32'h3bdacc6d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7529b9),
	.w1(32'h3be29e71),
	.w2(32'h3b925cf5),
	.w3(32'h3c3f7528),
	.w4(32'h39cac2ad),
	.w5(32'hbc06e3b9),
	.w6(32'h3c67c5d7),
	.w7(32'h3ca066db),
	.w8(32'h3c948024),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4bc3d),
	.w1(32'h3baa0223),
	.w2(32'h3ba04242),
	.w3(32'hbb9da3d4),
	.w4(32'h3b51b76a),
	.w5(32'h3b0dab48),
	.w6(32'h3bc934a5),
	.w7(32'h3ba87c08),
	.w8(32'h3b9e6db9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68fc02),
	.w1(32'h3b9fde53),
	.w2(32'hbb6d8d57),
	.w3(32'hba70b8a8),
	.w4(32'hbba3651b),
	.w5(32'hbc1130c3),
	.w6(32'h3b1ad1c6),
	.w7(32'hbad2ddda),
	.w8(32'hb988f906),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3019e5),
	.w1(32'h3ad2d0c5),
	.w2(32'h3b95946d),
	.w3(32'h3b43bb18),
	.w4(32'hb988439a),
	.w5(32'h3b68d052),
	.w6(32'h39ee9741),
	.w7(32'h3b18420b),
	.w8(32'h3a2ecacd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f6c75),
	.w1(32'h3b9a788d),
	.w2(32'h3b904567),
	.w3(32'h3c213643),
	.w4(32'h3cc982dc),
	.w5(32'h3c4daaac),
	.w6(32'hbb890ad6),
	.w7(32'h3c2a303c),
	.w8(32'h3c37d08b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a0c59),
	.w1(32'h3be3864f),
	.w2(32'hbb0b92ba),
	.w3(32'hba074798),
	.w4(32'h3bc5e5a2),
	.w5(32'hbbb1e143),
	.w6(32'h3bfbbd68),
	.w7(32'hbb373b8a),
	.w8(32'hbc0a6509),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b978cde),
	.w1(32'hbba9ac1b),
	.w2(32'hbbca381b),
	.w3(32'h3bfd34f3),
	.w4(32'hbb0a1e8d),
	.w5(32'hbc079d4e),
	.w6(32'h3bb30471),
	.w7(32'hbc0b419f),
	.w8(32'hbc52078a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38917b),
	.w1(32'h3b32a22a),
	.w2(32'h3c34d840),
	.w3(32'h3b47b695),
	.w4(32'h3c0a747f),
	.w5(32'h39cec0a3),
	.w6(32'h3acedf83),
	.w7(32'h3c2481d6),
	.w8(32'h3b93775b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb72d2d),
	.w1(32'h3a440d39),
	.w2(32'hbaf6e3e0),
	.w3(32'h3c274dea),
	.w4(32'hba0f6d34),
	.w5(32'hbbb88dc6),
	.w6(32'h3bac6e2a),
	.w7(32'h3723d0a4),
	.w8(32'h3bdc3c8c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c8c0a),
	.w1(32'h3b12c206),
	.w2(32'hbbf6bcc9),
	.w3(32'h3b7d9948),
	.w4(32'hbc065507),
	.w5(32'h3a57161e),
	.w6(32'h3baefe65),
	.w7(32'hbc450d9b),
	.w8(32'hbbbdcdc6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa97e8c),
	.w1(32'hbaa3eb51),
	.w2(32'hbc06ccaa),
	.w3(32'h3c2d9312),
	.w4(32'h3a4fb253),
	.w5(32'hbbdd0392),
	.w6(32'h3bb61cee),
	.w7(32'h3b5834b7),
	.w8(32'h3b0d05cd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc385b5e),
	.w1(32'hb9c69674),
	.w2(32'hb972f0f3),
	.w3(32'hbb862978),
	.w4(32'hba473b3a),
	.w5(32'hba2ef712),
	.w6(32'hbac6f079),
	.w7(32'hbb298155),
	.w8(32'hbbd2fd33),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bc391),
	.w1(32'h3b9ef4c7),
	.w2(32'h3bb56f75),
	.w3(32'hbb10bafc),
	.w4(32'h3a69528b),
	.w5(32'h3c02e5d4),
	.w6(32'h3ae89ad4),
	.w7(32'h3ba3acc9),
	.w8(32'h3c8e5f01),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf88892),
	.w1(32'h3bd9fdfd),
	.w2(32'h3c5f584c),
	.w3(32'h3cb5d9ba),
	.w4(32'h3c105bba),
	.w5(32'hbc0c7b7b),
	.w6(32'h3c1d4608),
	.w7(32'h3c9f8714),
	.w8(32'h3c9b3a85),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2358a),
	.w1(32'hbbb9d5d2),
	.w2(32'hbc801643),
	.w3(32'h3c50d050),
	.w4(32'h3ae45c96),
	.w5(32'hbc2e423b),
	.w6(32'h38ed18f6),
	.w7(32'hbbebe152),
	.w8(32'hba4b8f66),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992eaf5),
	.w1(32'hba09b9c0),
	.w2(32'hbc931df8),
	.w3(32'h3c4be594),
	.w4(32'h3c43dc8c),
	.w5(32'hbc789507),
	.w6(32'h3c8d00a0),
	.w7(32'h3a3ce87c),
	.w8(32'hbcc1b7c7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae9fa8),
	.w1(32'hbb88a33d),
	.w2(32'hbaa38391),
	.w3(32'hbc2ceed1),
	.w4(32'hbacd8386),
	.w5(32'h3b46486c),
	.w6(32'h3afc8dd5),
	.w7(32'hba8dfc1a),
	.w8(32'h3b6aeb1b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d5470),
	.w1(32'hbaf38783),
	.w2(32'hbc1b91a3),
	.w3(32'hbb733e10),
	.w4(32'hbb81ddd6),
	.w5(32'hbbf73c6f),
	.w6(32'hba74972e),
	.w7(32'hbbe1ef1b),
	.w8(32'hbb871ea7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea6e36),
	.w1(32'h3a06497d),
	.w2(32'h3c159cfe),
	.w3(32'h3a80fc7d),
	.w4(32'h3ca2ecd1),
	.w5(32'h3c7649b4),
	.w6(32'h3b4d9ce0),
	.w7(32'hbbb289e1),
	.w8(32'hbb7220b1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fe583),
	.w1(32'hbbf6c8a1),
	.w2(32'hbc56f630),
	.w3(32'h3c4031f1),
	.w4(32'h3a6bef54),
	.w5(32'hbc7d0e75),
	.w6(32'hbbbff067),
	.w7(32'hbb727d5c),
	.w8(32'hbcbd63f9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c2f05),
	.w1(32'h3c70d2d4),
	.w2(32'h3c534fbf),
	.w3(32'h3a6e5d36),
	.w4(32'h3c42d4b0),
	.w5(32'h3ce0a480),
	.w6(32'h3ba3ae2c),
	.w7(32'hbb8f78b2),
	.w8(32'hbb1ae66f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c351a15),
	.w1(32'hbbab6513),
	.w2(32'hbb878fa3),
	.w3(32'h3c806c74),
	.w4(32'hbbbe7474),
	.w5(32'hba056ca1),
	.w6(32'h3b908c3b),
	.w7(32'h3acf765d),
	.w8(32'h3bbd2a82),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24ca69),
	.w1(32'hbb474389),
	.w2(32'hbc0e6585),
	.w3(32'h3b13dce8),
	.w4(32'h3c65973c),
	.w5(32'h3baafa13),
	.w6(32'h3bfa955f),
	.w7(32'hbc1d97c9),
	.w8(32'h3af71a83),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0246dc),
	.w1(32'h3c165445),
	.w2(32'h3c6095bd),
	.w3(32'h3c1f8252),
	.w4(32'hb9ede6bb),
	.w5(32'hbbf72686),
	.w6(32'h3c511ccc),
	.w7(32'h3cb811bb),
	.w8(32'h3d01d1f2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3da96d56),
	.w1(32'h3cae640c),
	.w2(32'hbca9a49d),
	.w3(32'h3d359a22),
	.w4(32'h3bd2f9be),
	.w5(32'h3ca3284b),
	.w6(32'h3d6dd4ab),
	.w7(32'h3ce72e5d),
	.w8(32'hbc6105ae),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d7efd),
	.w1(32'h3bb02340),
	.w2(32'hbb4cbaa0),
	.w3(32'hba3fb69b),
	.w4(32'h3b7b2d16),
	.w5(32'hbc0cc22f),
	.w6(32'h3bb3db5a),
	.w7(32'h3b7c0121),
	.w8(32'hbbb00d26),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb691076),
	.w1(32'h3a14f9c3),
	.w2(32'h3a572382),
	.w3(32'hbab867d2),
	.w4(32'hbb8fd175),
	.w5(32'hbbb02801),
	.w6(32'h3b92d133),
	.w7(32'h3b69bfd2),
	.w8(32'h3c105e45),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a7b62),
	.w1(32'h3acc1096),
	.w2(32'hbaa4ebe7),
	.w3(32'h3b4d49a7),
	.w4(32'h3aa09592),
	.w5(32'hba75a274),
	.w6(32'h3a35374f),
	.w7(32'hbb7bb16e),
	.w8(32'hbb6d84ff),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1111ee),
	.w1(32'hba4a1b18),
	.w2(32'h39323ecf),
	.w3(32'h3a4f56ef),
	.w4(32'hbba1ebef),
	.w5(32'h3b73c8aa),
	.w6(32'hbad3e9ba),
	.w7(32'hbb91105d),
	.w8(32'hbb0ffcd2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc296b30),
	.w1(32'hbb337643),
	.w2(32'hbbd7d191),
	.w3(32'hbbc056a8),
	.w4(32'hb9c28b08),
	.w5(32'hbc2a20ee),
	.w6(32'h3c5ef730),
	.w7(32'hba124118),
	.w8(32'h39844d4c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd49931),
	.w1(32'hbab8c64f),
	.w2(32'h3bf9f3b9),
	.w3(32'hbbe7a0e0),
	.w4(32'hbba08ecd),
	.w5(32'hbb94875e),
	.w6(32'h3b34f630),
	.w7(32'h3bb10d44),
	.w8(32'h3c9b9144),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b582a),
	.w1(32'hbbafd6b8),
	.w2(32'hbb968f3c),
	.w3(32'hbb990019),
	.w4(32'hbb716598),
	.w5(32'hba6bdd55),
	.w6(32'h3b901be7),
	.w7(32'hbafa6037),
	.w8(32'h39d051fd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5feeaf),
	.w1(32'h3cd06488),
	.w2(32'h3c4b4a09),
	.w3(32'h3c111df0),
	.w4(32'hbb30ea63),
	.w5(32'hbbf7ee24),
	.w6(32'h3c4f0cb0),
	.w7(32'h3c65c678),
	.w8(32'h3ba7051a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dcefe),
	.w1(32'h3b376e5f),
	.w2(32'h3afa8dc8),
	.w3(32'hbca652eb),
	.w4(32'h3b2af435),
	.w5(32'hbaaf649c),
	.w6(32'h3b00b205),
	.w7(32'h3b3707af),
	.w8(32'hbac2bc23),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d44a7),
	.w1(32'h3bcdb6ec),
	.w2(32'h3b71aeb2),
	.w3(32'hba303fbf),
	.w4(32'h3b9fa05f),
	.w5(32'h3b54cef5),
	.w6(32'h3b6a992e),
	.w7(32'hbab34d0e),
	.w8(32'hbbfcd529),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acaf944),
	.w1(32'hbc2f1ec6),
	.w2(32'hbbd9ba7f),
	.w3(32'h3ba9b9b1),
	.w4(32'h3b1c42ae),
	.w5(32'h3c174fa9),
	.w6(32'hbbc84200),
	.w7(32'hbbda4d31),
	.w8(32'hbc1cb661),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22c8c0),
	.w1(32'h3c4b87f3),
	.w2(32'h3c85115b),
	.w3(32'h3c730b0b),
	.w4(32'h3c58bf77),
	.w5(32'h3c90c815),
	.w6(32'hbbb78c38),
	.w7(32'hbbae223c),
	.w8(32'hbc0bf762),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba7689),
	.w1(32'h3ab511a2),
	.w2(32'hbb01e179),
	.w3(32'h3c9dc5a4),
	.w4(32'h3c1a61b2),
	.w5(32'hb9040a17),
	.w6(32'h3cb6d988),
	.w7(32'h3be15477),
	.w8(32'h3bbf52e9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04c795),
	.w1(32'h3b59b50f),
	.w2(32'h3a4254f1),
	.w3(32'hb99ca182),
	.w4(32'h3c10551b),
	.w5(32'h3b591f23),
	.w6(32'h3be035af),
	.w7(32'hba7152c0),
	.w8(32'hbba8724e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8794ae),
	.w1(32'hbbaedf62),
	.w2(32'hbabc99bd),
	.w3(32'hbb904b15),
	.w4(32'hbba0fc9f),
	.w5(32'hbc242379),
	.w6(32'h3b10eb9e),
	.w7(32'h3bf5d5f1),
	.w8(32'hbb0482c5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb233d),
	.w1(32'hbbe2ac0f),
	.w2(32'hbbddb07c),
	.w3(32'hbb32cd31),
	.w4(32'hbba5bcdd),
	.w5(32'hbc67ca5c),
	.w6(32'hbbd52590),
	.w7(32'hbc2e795a),
	.w8(32'hbb8b556e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ec678),
	.w1(32'h3c82cc12),
	.w2(32'hbbb22965),
	.w3(32'h3bc90b9b),
	.w4(32'hbb3b5a2c),
	.w5(32'hbcafe860),
	.w6(32'h3cdee30a),
	.w7(32'h3c8fcc49),
	.w8(32'hbc4cb225),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06ea73),
	.w1(32'h3bb2f491),
	.w2(32'hbb40a446),
	.w3(32'hbcdaf5bf),
	.w4(32'h38a7b4e0),
	.w5(32'hbbc89f75),
	.w6(32'h3bd975dd),
	.w7(32'hba57724e),
	.w8(32'hbbe7b3ab),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8546dc),
	.w1(32'hba853c04),
	.w2(32'h3ad16c2c),
	.w3(32'hba8253a7),
	.w4(32'hb8a96661),
	.w5(32'h3b1459d7),
	.w6(32'h397b5daf),
	.w7(32'h3a80a035),
	.w8(32'h3c071f18),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b066),
	.w1(32'h3c3a42e3),
	.w2(32'h3c34b1d0),
	.w3(32'hbae04604),
	.w4(32'h3b71183d),
	.w5(32'hbb6d5573),
	.w6(32'hbaa65667),
	.w7(32'hbb57b608),
	.w8(32'hbc5cd5f2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3e420),
	.w1(32'h3c5d8821),
	.w2(32'h3c26fdf3),
	.w3(32'h3ad9fcaf),
	.w4(32'h3b0e108e),
	.w5(32'h3aa49fd5),
	.w6(32'h3bb857f7),
	.w7(32'h3c3a80cb),
	.w8(32'hbac719d8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913881b),
	.w1(32'h3ad39b8a),
	.w2(32'hbc5d35d0),
	.w3(32'h3bbbe3a2),
	.w4(32'h3bdb9d80),
	.w5(32'hbbb8297b),
	.w6(32'hbb55226c),
	.w7(32'hbc2e6e72),
	.w8(32'hbba3feeb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81a329),
	.w1(32'hbc1467fa),
	.w2(32'hbc25d96a),
	.w3(32'hbc327071),
	.w4(32'hbc1b5bc4),
	.w5(32'hbc240c4f),
	.w6(32'hbb04142b),
	.w7(32'hbc48629c),
	.w8(32'hbc1ca636),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b49dd),
	.w1(32'h3c4044ce),
	.w2(32'hba458612),
	.w3(32'h3c744994),
	.w4(32'h3c872f63),
	.w5(32'hbb054f61),
	.w6(32'h3caf7079),
	.w7(32'h3c39875a),
	.w8(32'hbc1549fe),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c5151),
	.w1(32'h3b3a370a),
	.w2(32'h3b11c0f7),
	.w3(32'hbc08451a),
	.w4(32'h3b3ddca8),
	.w5(32'h3ad29e0b),
	.w6(32'h3b90fa96),
	.w7(32'h3a875a7b),
	.w8(32'hbb95c460),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5082e2),
	.w1(32'hbc047109),
	.w2(32'hbcf1e661),
	.w3(32'h3bd09834),
	.w4(32'hbbce075c),
	.w5(32'hbcaa96ad),
	.w6(32'hbbcf8b78),
	.w7(32'hbca93a24),
	.w8(32'hbce90004),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc817d6),
	.w1(32'hb9c59750),
	.w2(32'hbb413d16),
	.w3(32'hbc473d28),
	.w4(32'hbbb3e816),
	.w5(32'hbb7a128f),
	.w6(32'h3a9bfc04),
	.w7(32'hbbd01dae),
	.w8(32'hbbaf9d34),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b571e9b),
	.w1(32'hbb4d05ce),
	.w2(32'h39d33f37),
	.w3(32'hbaab2566),
	.w4(32'h3b1381db),
	.w5(32'hbabedb47),
	.w6(32'hb801b2b9),
	.w7(32'hbc43a156),
	.w8(32'hbbdde302),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96c3fc),
	.w1(32'h3b0b62e8),
	.w2(32'hbb46d726),
	.w3(32'h3c66a9a1),
	.w4(32'h3a8ecdd7),
	.w5(32'hbbc436dc),
	.w6(32'h3bbf918c),
	.w7(32'h3ba8da66),
	.w8(32'h3bd86acb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9871bf),
	.w1(32'h3bd0b3ca),
	.w2(32'hbb3a4196),
	.w3(32'h3c6bd426),
	.w4(32'h3bd5216d),
	.w5(32'hbc29dfa0),
	.w6(32'h3c65a99f),
	.w7(32'h3b32acfb),
	.w8(32'hbc034fa5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9b9bd),
	.w1(32'hb873b72b),
	.w2(32'h3a7904a6),
	.w3(32'hbc086e0d),
	.w4(32'h3b14fe3f),
	.w5(32'h3baaa719),
	.w6(32'hbb12d510),
	.w7(32'hbb0fabab),
	.w8(32'hbb8bbefa),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a65a9),
	.w1(32'h3c780a4b),
	.w2(32'h3c33f5eb),
	.w3(32'h3bd7abb5),
	.w4(32'h3c9090e5),
	.w5(32'h3cc3c1b2),
	.w6(32'h3baea3eb),
	.w7(32'h3b8b9eb2),
	.w8(32'hbbf94106),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8710f9),
	.w1(32'hbb48b263),
	.w2(32'h3a2fa3e8),
	.w3(32'h3c4ff9b8),
	.w4(32'h3af131de),
	.w5(32'h3c120abe),
	.w6(32'hbba0be44),
	.w7(32'hbbf51ce6),
	.w8(32'hbc046d6e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baee5e1),
	.w1(32'hbb28bf52),
	.w2(32'h3ad95dac),
	.w3(32'h3c8f93aa),
	.w4(32'hbb495ce5),
	.w5(32'hbb04f3fd),
	.w6(32'hbb2f0937),
	.w7(32'h3a07afae),
	.w8(32'hba5021fe),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5189b2),
	.w1(32'h3ab93b9d),
	.w2(32'h3b5943fd),
	.w3(32'h3c2520f0),
	.w4(32'h3b25bdf1),
	.w5(32'hba6617a8),
	.w6(32'h3b604e84),
	.w7(32'hbb6d6cec),
	.w8(32'hbac3b363),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c85b0),
	.w1(32'hbb242c6a),
	.w2(32'hba8a0aef),
	.w3(32'h3bad8ef0),
	.w4(32'h3ad24afa),
	.w5(32'h3a1bc50c),
	.w6(32'h3ba27099),
	.w7(32'h3bb3fb58),
	.w8(32'h3b696c5d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb465c6c),
	.w1(32'hbb889826),
	.w2(32'hbb33edb0),
	.w3(32'hbb082e9b),
	.w4(32'hbaf170f9),
	.w5(32'hb9d7fce3),
	.w6(32'hbc0befa3),
	.w7(32'hbbf6f9df),
	.w8(32'hbbe29023),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae39b41),
	.w1(32'h3bfd9899),
	.w2(32'h3beccd84),
	.w3(32'h3ba7bc2d),
	.w4(32'h3cb3f665),
	.w5(32'h3c9ea903),
	.w6(32'hbaec44ef),
	.w7(32'hbbaf5f60),
	.w8(32'hbbd936af),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba31e3b),
	.w1(32'hbc43e6e6),
	.w2(32'hbc7ae544),
	.w3(32'h3c0f395f),
	.w4(32'hbcabc1d8),
	.w5(32'hbc868564),
	.w6(32'hbb8189ad),
	.w7(32'hbbf909cf),
	.w8(32'hbc844f24),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc067ca4),
	.w1(32'hba283439),
	.w2(32'h3b22fda2),
	.w3(32'hbb30dcca),
	.w4(32'h3b967536),
	.w5(32'h3b660968),
	.w6(32'h3a223d92),
	.w7(32'hbc383344),
	.w8(32'h3c202cef),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c006e98),
	.w1(32'h3b63d05b),
	.w2(32'hba313ab9),
	.w3(32'h3c0e8a0c),
	.w4(32'h3b20cad8),
	.w5(32'h3b302574),
	.w6(32'hbb4a3298),
	.w7(32'hbb92edcc),
	.w8(32'h3b1b13d2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ee06c),
	.w1(32'h3c38acff),
	.w2(32'h3c8385c2),
	.w3(32'hbbd79c6e),
	.w4(32'h3c717e77),
	.w5(32'h3bfff221),
	.w6(32'h3c3fbcf5),
	.w7(32'h3ca527c5),
	.w8(32'hbca4609d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f176ef),
	.w1(32'h3b1f9efc),
	.w2(32'hbb1caa3e),
	.w3(32'h3c2a7a39),
	.w4(32'h3a182e86),
	.w5(32'hbb8e9d03),
	.w6(32'h3abc3d6f),
	.w7(32'hbbeaa642),
	.w8(32'hbb8f942e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfe2af),
	.w1(32'h3b47a9eb),
	.w2(32'h399c118c),
	.w3(32'h3afccd02),
	.w4(32'hbba28de7),
	.w5(32'hbc59b6ec),
	.w6(32'h3ccef00c),
	.w7(32'h3cccc8a7),
	.w8(32'h3c79e836),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1737d5),
	.w1(32'h3c27a34b),
	.w2(32'h3ad0e816),
	.w3(32'hbc1ff840),
	.w4(32'hbc1df8b9),
	.w5(32'hbc4f81fb),
	.w6(32'h3c3335ed),
	.w7(32'h3c8d3881),
	.w8(32'h3bc95c3b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d16b),
	.w1(32'hbbb87762),
	.w2(32'hbc02605f),
	.w3(32'hbc048a7c),
	.w4(32'hbb615359),
	.w5(32'hbc0ff533),
	.w6(32'hbada3387),
	.w7(32'hbbf96856),
	.w8(32'hbbef61cc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a35840),
	.w1(32'h3b7b7382),
	.w2(32'hbb8a41bd),
	.w3(32'hbb8f4d9a),
	.w4(32'hbbdd147e),
	.w5(32'hbc064931),
	.w6(32'h3c01f6b8),
	.w7(32'h3bb51aae),
	.w8(32'hbac73d53),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccf890),
	.w1(32'h3c3925b3),
	.w2(32'h3c4071b9),
	.w3(32'hbc1ca85e),
	.w4(32'h3c063233),
	.w5(32'h3b627b80),
	.w6(32'h3c214524),
	.w7(32'h3c11ee36),
	.w8(32'hba1a1d8e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4a6d4),
	.w1(32'h3b69c82e),
	.w2(32'hbab4353c),
	.w3(32'h3b3669d6),
	.w4(32'h39426ef3),
	.w5(32'hbbe0f738),
	.w6(32'h3b57d8fe),
	.w7(32'hb9df318f),
	.w8(32'hba7c5b40),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85caa7),
	.w1(32'h3a32e60b),
	.w2(32'hbb604d19),
	.w3(32'hbb0eb684),
	.w4(32'h3bdaf854),
	.w5(32'hbb89dbaf),
	.w6(32'h3c016183),
	.w7(32'h3b80d2ce),
	.w8(32'hbb0b3e37),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8e1fa),
	.w1(32'hba406514),
	.w2(32'hbc233ade),
	.w3(32'h3bc8589f),
	.w4(32'h3bebdbd1),
	.w5(32'hbb98e60c),
	.w6(32'h3c39e8ff),
	.w7(32'h3aacf2e5),
	.w8(32'hbbd8172f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc336b7e),
	.w1(32'hbc57f659),
	.w2(32'h3bd775e8),
	.w3(32'hbb9fefa1),
	.w4(32'hbb0b98ec),
	.w5(32'h3a8f5b3d),
	.w6(32'hbc1795ec),
	.w7(32'hbb127297),
	.w8(32'h3c3370c2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c8cda),
	.w1(32'h3b347a7a),
	.w2(32'h3b8b9ad2),
	.w3(32'h3c1906cf),
	.w4(32'hba3a9f95),
	.w5(32'h3ab94219),
	.w6(32'h3be3b299),
	.w7(32'h3c0a0525),
	.w8(32'hb87a1b1f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e9fd6),
	.w1(32'h3c18f207),
	.w2(32'h3bcad80e),
	.w3(32'h3c16feec),
	.w4(32'h3c50eda4),
	.w5(32'h3a94f480),
	.w6(32'h3c2a395b),
	.w7(32'h3b5255b6),
	.w8(32'h3c8fd40a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33a8ab),
	.w1(32'hbc109eb3),
	.w2(32'hbc094334),
	.w3(32'h3b39fff6),
	.w4(32'hbb32bc68),
	.w5(32'hbc6c0621),
	.w6(32'h3c06d695),
	.w7(32'hbbece211),
	.w8(32'hbbf00c18),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f3a3d),
	.w1(32'hbb3ef3f6),
	.w2(32'hbb94a23b),
	.w3(32'h3c8ab694),
	.w4(32'hba2e6175),
	.w5(32'h3aa68f96),
	.w6(32'h3c95f869),
	.w7(32'h3c59eb79),
	.w8(32'h3adaef0d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d7892),
	.w1(32'hbb91bd73),
	.w2(32'hbc5fd048),
	.w3(32'h3a91c26d),
	.w4(32'h3ac70739),
	.w5(32'hbc9125cb),
	.w6(32'h3c93dcb5),
	.w7(32'h3bfeb76f),
	.w8(32'hbbf0bf28),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96b71b),
	.w1(32'h3c06a6e8),
	.w2(32'h3c309b60),
	.w3(32'hbc9604ac),
	.w4(32'h3b133527),
	.w5(32'h3c15ae17),
	.w6(32'h3bf9b018),
	.w7(32'h3c82dead),
	.w8(32'h3ca06625),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14753c),
	.w1(32'hbb1c6774),
	.w2(32'hbb172742),
	.w3(32'h3c01575d),
	.w4(32'h3b4994d3),
	.w5(32'h3beade29),
	.w6(32'hbbada615),
	.w7(32'hbbcf1898),
	.w8(32'hbaa041bd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d5cfd),
	.w1(32'hbaf4855b),
	.w2(32'h3a9c957a),
	.w3(32'h3c0f1272),
	.w4(32'h39c7c234),
	.w5(32'h39e79b49),
	.w6(32'hbbfc584e),
	.w7(32'hbbc55645),
	.w8(32'h3b00c476),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a439c),
	.w1(32'hba79bdbe),
	.w2(32'hb83341b3),
	.w3(32'hbb866393),
	.w4(32'hbaf4a305),
	.w5(32'h3a974f21),
	.w6(32'h393ad2eb),
	.w7(32'hbb21be6b),
	.w8(32'h3ac4bb8d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a664a),
	.w1(32'h3c48af1f),
	.w2(32'h3c4221c4),
	.w3(32'h3bb12558),
	.w4(32'h3b587b03),
	.w5(32'h3b6ecf80),
	.w6(32'h3af75457),
	.w7(32'h3c794450),
	.w8(32'h3c051491),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19bf31),
	.w1(32'h3a6343d4),
	.w2(32'h3b9f749c),
	.w3(32'h3c028c33),
	.w4(32'hbbc836a0),
	.w5(32'hbc28b5ed),
	.w6(32'h3c3dd34d),
	.w7(32'h3cc77764),
	.w8(32'h3c57e44d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18e7c5),
	.w1(32'h39c2fd01),
	.w2(32'h3b528b0c),
	.w3(32'hbcb099e2),
	.w4(32'hbb02f7cf),
	.w5(32'h3a8e579b),
	.w6(32'h3bbc71da),
	.w7(32'h3b3ed691),
	.w8(32'h3c1e3f22),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2547bc),
	.w1(32'hbadeb724),
	.w2(32'hbafec635),
	.w3(32'h3ba28583),
	.w4(32'h3a495aa7),
	.w5(32'h3b2776e9),
	.w6(32'h3bba8756),
	.w7(32'hba4948d9),
	.w8(32'hbb668f48),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee289),
	.w1(32'hbbbb4108),
	.w2(32'hbb725b4d),
	.w3(32'h3a1378e6),
	.w4(32'hbb245188),
	.w5(32'h3918dc26),
	.w6(32'hbb5b830b),
	.w7(32'hbbbadc73),
	.w8(32'hbb3a0037),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56d9d3),
	.w1(32'hba90d9f1),
	.w2(32'hbc6aa06a),
	.w3(32'h3b49c9a8),
	.w4(32'h3b0f01ec),
	.w5(32'hbc9f3d80),
	.w6(32'h3b9e3785),
	.w7(32'h3b892035),
	.w8(32'hbc0fe597),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88e9bb),
	.w1(32'hbb035971),
	.w2(32'hbb881ea7),
	.w3(32'hbcab0dbe),
	.w4(32'hbb787c6d),
	.w5(32'hbc048630),
	.w6(32'hbaad9cf3),
	.w7(32'hbb47dbfb),
	.w8(32'hbbca2bac),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6f2bf),
	.w1(32'h3bd9a32d),
	.w2(32'h3beb42f7),
	.w3(32'h3a8a98df),
	.w4(32'h3bf1d7a1),
	.w5(32'hbb589a53),
	.w6(32'h3c98cab4),
	.w7(32'h3cacfd2b),
	.w8(32'hbb8f7170),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8625b),
	.w1(32'hbc0efc3d),
	.w2(32'hbbec692a),
	.w3(32'hbacf587a),
	.w4(32'hbc00dcc7),
	.w5(32'hba252fa4),
	.w6(32'hb887e236),
	.w7(32'hbb98029b),
	.w8(32'hbbf79b69),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13b712),
	.w1(32'hbc9651f3),
	.w2(32'hbc2cce26),
	.w3(32'h3bc3de1a),
	.w4(32'hbc25d05c),
	.w5(32'h39e65b73),
	.w6(32'hbc53a030),
	.w7(32'hbc9d0031),
	.w8(32'hbb5568a4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e3944),
	.w1(32'hbb783821),
	.w2(32'hbb8202cf),
	.w3(32'h3c792a19),
	.w4(32'h3a8a00e6),
	.w5(32'hbb40acd7),
	.w6(32'h3b38c275),
	.w7(32'h3c2b23be),
	.w8(32'h3bd44ce8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44f73c),
	.w1(32'hbc669543),
	.w2(32'hbc8fdab6),
	.w3(32'hba0bafc9),
	.w4(32'hbc9449c6),
	.w5(32'hbcb6f3ed),
	.w6(32'h3b208e43),
	.w7(32'hbbb0d7f7),
	.w8(32'hbc71152b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd5903b),
	.w1(32'h3beec7d6),
	.w2(32'hbb2fcc9b),
	.w3(32'hbc533bb8),
	.w4(32'hbc52bc63),
	.w5(32'hbc8747fa),
	.w6(32'h3c3ba572),
	.w7(32'h3c6a4e28),
	.w8(32'h3a87bf96),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1f75f),
	.w1(32'hbb18686b),
	.w2(32'h3aabdebb),
	.w3(32'hbcbb4938),
	.w4(32'hbb1b9982),
	.w5(32'hbbcc7cff),
	.w6(32'h3b450a69),
	.w7(32'h3bfd2076),
	.w8(32'h3b213cd4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb4bf0),
	.w1(32'h3b30a78b),
	.w2(32'hba97df79),
	.w3(32'hbac5c6ac),
	.w4(32'h3b1fc657),
	.w5(32'h3a0a87ba),
	.w6(32'h3c532292),
	.w7(32'h3c0592f9),
	.w8(32'hbb6d875a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6aad4),
	.w1(32'hbc4af98c),
	.w2(32'h3b86ac2c),
	.w3(32'h3aa2ea2e),
	.w4(32'hbc52e2e4),
	.w5(32'hbb52fb06),
	.w6(32'hbc02a837),
	.w7(32'h3b96bea1),
	.w8(32'h3c2a1847),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd64c80),
	.w1(32'h3b7a709e),
	.w2(32'hb93f8791),
	.w3(32'h3a9f4bd8),
	.w4(32'h3bfcf9b7),
	.w5(32'h3b3881e4),
	.w6(32'h3b7d443f),
	.w7(32'hbb3ec33a),
	.w8(32'hbc27c4e8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a6ba4),
	.w1(32'hbb7bb7d7),
	.w2(32'hbbaf9bd3),
	.w3(32'hba37f172),
	.w4(32'h3b38dac0),
	.w5(32'h3bf3f689),
	.w6(32'hba932c51),
	.w7(32'hbba797ab),
	.w8(32'h3a129677),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59cbf),
	.w1(32'h3a33fe66),
	.w2(32'hb892979a),
	.w3(32'h3c52917c),
	.w4(32'h3b2a73ec),
	.w5(32'hbbbf8df7),
	.w6(32'h3bc14bd1),
	.w7(32'h3a95e110),
	.w8(32'h3ba9718d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3edf08),
	.w1(32'h3bfe6050),
	.w2(32'h3cb82243),
	.w3(32'hbb993042),
	.w4(32'h3b9391c8),
	.w5(32'h3ca3c055),
	.w6(32'h3c07493c),
	.w7(32'h3c7ac908),
	.w8(32'h3cc00a79),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce88754),
	.w1(32'h3b952781),
	.w2(32'h3b1ad997),
	.w3(32'h3ca647ec),
	.w4(32'h3ba0cfb6),
	.w5(32'h3afa9ca2),
	.w6(32'h3b62748b),
	.w7(32'h3a8bf660),
	.w8(32'hba27cbae),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18bfe1),
	.w1(32'h3b29272a),
	.w2(32'hbb9f8afc),
	.w3(32'h3c065239),
	.w4(32'hbb392d7d),
	.w5(32'hbbf34e24),
	.w6(32'h3c783731),
	.w7(32'h3c402907),
	.w8(32'h3c31fc8a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baedde3),
	.w1(32'hbb89daeb),
	.w2(32'hba7c0238),
	.w3(32'hbc5c4b5c),
	.w4(32'hbb765e66),
	.w5(32'h3902812e),
	.w6(32'h395c7282),
	.w7(32'hbbb1bd19),
	.w8(32'h3a3c5d89),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d038e),
	.w1(32'h3a792e50),
	.w2(32'h3bf4fe84),
	.w3(32'h39e8d92a),
	.w4(32'h3a1393a4),
	.w5(32'h3bda5330),
	.w6(32'h3bcfd4ca),
	.w7(32'h3a2583ff),
	.w8(32'h3b557cf5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a888bfe),
	.w1(32'hbc6d03fb),
	.w2(32'hbc7cc893),
	.w3(32'h3c188205),
	.w4(32'hbca2795d),
	.w5(32'hbc92bcd2),
	.w6(32'h3a5918ed),
	.w7(32'h3a9c8121),
	.w8(32'hbc15d4d5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9c300),
	.w1(32'h3aab3361),
	.w2(32'h397471d9),
	.w3(32'hbb2d91ac),
	.w4(32'h3baa562d),
	.w5(32'h3b9913bb),
	.w6(32'hbb0c1e00),
	.w7(32'hb99cae22),
	.w8(32'hb9aa753a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9730fb),
	.w1(32'h3a9794de),
	.w2(32'h3affd300),
	.w3(32'h3b0d834d),
	.w4(32'h3b0fec92),
	.w5(32'h3b8b417f),
	.w6(32'hbb17b73a),
	.w7(32'hbb3dc0fc),
	.w8(32'hbb2a5943),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5e143),
	.w1(32'h3a6ce67c),
	.w2(32'hbafcc14f),
	.w3(32'h3ba15d49),
	.w4(32'hbb21c3d6),
	.w5(32'h3b286e87),
	.w6(32'h3b5b2564),
	.w7(32'hbb45d96f),
	.w8(32'h3b2ffbc2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5844b),
	.w1(32'h3b52c890),
	.w2(32'h3ab431d3),
	.w3(32'h3c19d27d),
	.w4(32'h3b9d1e48),
	.w5(32'h3b9fdc32),
	.w6(32'h3bc32028),
	.w7(32'hbb62cee6),
	.w8(32'h3bb228d0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa80eb),
	.w1(32'hbc0fe30d),
	.w2(32'hbc755bb7),
	.w3(32'hb98950a1),
	.w4(32'hbc476467),
	.w5(32'hbc3e3e88),
	.w6(32'hbbdafdc0),
	.w7(32'hbc36f27f),
	.w8(32'hbbff6b7c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f802a),
	.w1(32'h3b926152),
	.w2(32'h3abfee50),
	.w3(32'hbc2abc35),
	.w4(32'hbbbd5cd1),
	.w5(32'hbba86bd8),
	.w6(32'h3bd201a6),
	.w7(32'h3ba842a3),
	.w8(32'h3bb8ab26),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cce941),
	.w1(32'h3b06d7d9),
	.w2(32'h3c4d0104),
	.w3(32'hbb0a801c),
	.w4(32'hba957a2c),
	.w5(32'hbbaa0478),
	.w6(32'h3a379e5b),
	.w7(32'hbb8701a0),
	.w8(32'h3bd3d07b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2375e7),
	.w1(32'h3ba65294),
	.w2(32'hbaa63b2a),
	.w3(32'h3bf056ef),
	.w4(32'h3b6d7066),
	.w5(32'h3902662f),
	.w6(32'h3a6a19a6),
	.w7(32'hbaea8e89),
	.w8(32'h3b3f85a8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ffe73),
	.w1(32'hbb384c19),
	.w2(32'hbb513936),
	.w3(32'hbb3676f7),
	.w4(32'hbb69d269),
	.w5(32'hbb828591),
	.w6(32'h3b05d04e),
	.w7(32'hb94042aa),
	.w8(32'h38038546),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad79b34),
	.w1(32'h3c17053e),
	.w2(32'h3c5c3956),
	.w3(32'hba7a8a93),
	.w4(32'h3be0b775),
	.w5(32'h3c3368a4),
	.w6(32'h39027f8b),
	.w7(32'hbbe8d5f6),
	.w8(32'h3afe0ae4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1fa4d),
	.w1(32'hbc683646),
	.w2(32'hbc9424d2),
	.w3(32'hb93d00e8),
	.w4(32'hbbf7600e),
	.w5(32'hbcb50266),
	.w6(32'hbbcb54c2),
	.w7(32'hbc6f9e69),
	.w8(32'hbc3ae06d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0f7af),
	.w1(32'h3c406421),
	.w2(32'h3c08e19d),
	.w3(32'hbb858c56),
	.w4(32'h3c140bf4),
	.w5(32'h3bd92ce9),
	.w6(32'hba9b3875),
	.w7(32'hbaf2b87f),
	.w8(32'hbbb998d0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5880f7),
	.w1(32'h3b175616),
	.w2(32'hbb3dfd1f),
	.w3(32'h3c3200a0),
	.w4(32'h3a8b7aa2),
	.w5(32'hbb3ccad4),
	.w6(32'h3b2c0d7a),
	.w7(32'hbb2a7a93),
	.w8(32'h3a2d4e8e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a980abe),
	.w1(32'hbc304dce),
	.w2(32'h3c1f0fda),
	.w3(32'h3ab63aa9),
	.w4(32'hbbeb4264),
	.w5(32'h3bb9cd46),
	.w6(32'hbbd52aed),
	.w7(32'h3c33f7bf),
	.w8(32'hbb8ec7e1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule