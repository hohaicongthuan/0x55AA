module layer_10_featuremap_144(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938cd51),
	.w1(32'hbc71b105),
	.w2(32'hbbc37c33),
	.w3(32'hba302971),
	.w4(32'hbc60e131),
	.w5(32'hbbd18068),
	.w6(32'hbbe24b19),
	.w7(32'h3b3214bd),
	.w8(32'h3c03bc96),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa904bd),
	.w1(32'hb9ff0b1d),
	.w2(32'hbb6d63af),
	.w3(32'hbb875e1e),
	.w4(32'h3b0fd855),
	.w5(32'hbab51581),
	.w6(32'hbb1c7b14),
	.w7(32'h3a7d1da4),
	.w8(32'hbb02085b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c14c22),
	.w1(32'hbaf7fae3),
	.w2(32'hbb2044d1),
	.w3(32'hb9b8c13f),
	.w4(32'hba8c3edf),
	.w5(32'hbb0e84b8),
	.w6(32'hba96917f),
	.w7(32'hbb1f85b6),
	.w8(32'hbadd3e25),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e123c),
	.w1(32'h3b830ca1),
	.w2(32'h3b939402),
	.w3(32'hbae2e162),
	.w4(32'h3a987857),
	.w5(32'h3b551f89),
	.w6(32'hba8c3821),
	.w7(32'h3b0d226b),
	.w8(32'h3b1a8b31),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab7d10),
	.w1(32'h3b7b3ab1),
	.w2(32'h3b0cae4d),
	.w3(32'h3bfa347c),
	.w4(32'h3b90e4a3),
	.w5(32'h3b086981),
	.w6(32'h3affc031),
	.w7(32'hbaa049a9),
	.w8(32'hbb633ba5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76fd74),
	.w1(32'h3bca9371),
	.w2(32'h3c0ecbe6),
	.w3(32'hbaafd161),
	.w4(32'h3b92d7b3),
	.w5(32'h3be8d51a),
	.w6(32'h3b725fdd),
	.w7(32'h3c0b5001),
	.w8(32'h3bcd522d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5c508),
	.w1(32'hbc129c9b),
	.w2(32'hbc454cbc),
	.w3(32'h3b6dbd15),
	.w4(32'hbc1d51dd),
	.w5(32'hbc476658),
	.w6(32'hbb577716),
	.w7(32'hbc127d7b),
	.w8(32'hbc1364c3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc441ead),
	.w1(32'hbb8288a2),
	.w2(32'hbad677f2),
	.w3(32'hbc6d3561),
	.w4(32'hbc1e3589),
	.w5(32'hba3d9afe),
	.w6(32'hbc2f41e7),
	.w7(32'hba3eaeee),
	.w8(32'hbb836a66),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2307dd),
	.w1(32'hba728eac),
	.w2(32'h3a2d431c),
	.w3(32'h3a985fc6),
	.w4(32'hbaec03e1),
	.w5(32'h3a867b22),
	.w6(32'hbb732679),
	.w7(32'h38e34b20),
	.w8(32'hbb4227b5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b34cc),
	.w1(32'hbc0fda85),
	.w2(32'hbcab4c88),
	.w3(32'hbbaccc60),
	.w4(32'hbbb307ba),
	.w5(32'hbc935ff1),
	.w6(32'hbc558c7a),
	.w7(32'hbc3beb4c),
	.w8(32'hbc89f83a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c0d68),
	.w1(32'h3bbe2fde),
	.w2(32'h3bd3fa34),
	.w3(32'hbbea1110),
	.w4(32'h3b1d7b0f),
	.w5(32'h3b4e80b6),
	.w6(32'h3b8500de),
	.w7(32'h3bb47ada),
	.w8(32'h3bc5ed07),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd71f0),
	.w1(32'h3bc47131),
	.w2(32'h39af8e7f),
	.w3(32'hb984fa18),
	.w4(32'hb8a81752),
	.w5(32'hbb35789c),
	.w6(32'hbbcfe530),
	.w7(32'h3b3adc57),
	.w8(32'hbbe724af),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942ce5),
	.w1(32'hbb3821e2),
	.w2(32'hbc2c87ac),
	.w3(32'hba51c4b5),
	.w4(32'hba82e805),
	.w5(32'hbc14eadb),
	.w6(32'hbb62c83c),
	.w7(32'hba96186a),
	.w8(32'hbbec7f41),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bee7f),
	.w1(32'hbbeb21aa),
	.w2(32'hbaeb6023),
	.w3(32'hbb166641),
	.w4(32'hbbb63550),
	.w5(32'h3aca174d),
	.w6(32'hbc02709d),
	.w7(32'h3a35aa07),
	.w8(32'hba584304),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f6cc1),
	.w1(32'h3bb90c39),
	.w2(32'hba52e756),
	.w3(32'h3ba012a9),
	.w4(32'h3b9940be),
	.w5(32'h3a7d4594),
	.w6(32'hbbe199ac),
	.w7(32'hbab9d4af),
	.w8(32'hbc09ad78),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020ccd),
	.w1(32'hbb8a363b),
	.w2(32'hbc088dbf),
	.w3(32'hbbf42013),
	.w4(32'hb92594ff),
	.w5(32'hbb0fe60f),
	.w6(32'hbc1464c5),
	.w7(32'hbb251b76),
	.w8(32'hbc0ec9a8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba493e8d),
	.w1(32'h3addd1e8),
	.w2(32'h3b5d049e),
	.w3(32'h3990709e),
	.w4(32'h3a08da49),
	.w5(32'h3af8fb61),
	.w6(32'h3b3e1c9b),
	.w7(32'h3b35f3ad),
	.w8(32'h3b896537),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc31ed2),
	.w1(32'hbc6ef7b1),
	.w2(32'hbca964c0),
	.w3(32'hbc13aa7a),
	.w4(32'hbc5eff4c),
	.w5(32'hbca9f5e2),
	.w6(32'hbc6d7dbe),
	.w7(32'hbc70a9a8),
	.w8(32'hbc849119),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc763b0b),
	.w1(32'hbb4f77fd),
	.w2(32'hbbe7b620),
	.w3(32'hbc58a3cd),
	.w4(32'hbb9b29ac),
	.w5(32'hbc0863eb),
	.w6(32'hbb8506aa),
	.w7(32'hbb99e198),
	.w8(32'hbbe589da),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c650a),
	.w1(32'hbb6f8344),
	.w2(32'hb9cc39df),
	.w3(32'hb9f91057),
	.w4(32'hbb8a1826),
	.w5(32'hb973f9e2),
	.w6(32'hbb9cbe44),
	.w7(32'hba523783),
	.w8(32'hbb4dd4e3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15ad1b),
	.w1(32'h3ae91a32),
	.w2(32'h3ba5d5ec),
	.w3(32'hbb279a4b),
	.w4(32'h3a381983),
	.w5(32'h3b961db0),
	.w6(32'hb944ba15),
	.w7(32'h3bb1ee6c),
	.w8(32'h3a4d708c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62a47e),
	.w1(32'hb8c31442),
	.w2(32'hb9264df4),
	.w3(32'h3b7a740e),
	.w4(32'h3bcc196f),
	.w5(32'h3baa6283),
	.w6(32'hbb33282b),
	.w7(32'h3b0d6814),
	.w8(32'h3b27b620),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc235104),
	.w1(32'hbaefab91),
	.w2(32'hbc46d45b),
	.w3(32'hbbd30291),
	.w4(32'h3a5ef3b3),
	.w5(32'hbc1d1412),
	.w6(32'hbc5f4043),
	.w7(32'hbbd50c19),
	.w8(32'hbca58e9c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfffbea),
	.w1(32'h396555d4),
	.w2(32'hbbe9a9f1),
	.w3(32'h3a9093ec),
	.w4(32'h3b701261),
	.w5(32'hbb72832f),
	.w6(32'hbc106d66),
	.w7(32'h3b7fe942),
	.w8(32'hbc19a125),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22a63a),
	.w1(32'h3bc7b1ff),
	.w2(32'hbb7b00e9),
	.w3(32'hbbf04261),
	.w4(32'h3c038adf),
	.w5(32'hbab0b31f),
	.w6(32'hbc44a4c4),
	.w7(32'h3b93ee43),
	.w8(32'hbb576db3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f73dd),
	.w1(32'h3bb00907),
	.w2(32'h3bf574f9),
	.w3(32'h3b1e4059),
	.w4(32'h3bbeeba2),
	.w5(32'h3ba50fe4),
	.w6(32'h3907b592),
	.w7(32'hb99662d5),
	.w8(32'hba1ca4d5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe7405),
	.w1(32'hbb344ab3),
	.w2(32'h38ce7165),
	.w3(32'h3b383660),
	.w4(32'hbb50a761),
	.w5(32'hb9722eac),
	.w6(32'hbb92761f),
	.w7(32'hbabf2706),
	.w8(32'hbb526141),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48edc7),
	.w1(32'h3bf30804),
	.w2(32'hba096aa7),
	.w3(32'hbb54c1e5),
	.w4(32'h3bc3eee5),
	.w5(32'h3b1bad65),
	.w6(32'hb9a686a7),
	.w7(32'h3b9726f9),
	.w8(32'h3b15e41b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6976f4),
	.w1(32'h3b8fb8fb),
	.w2(32'h3afba724),
	.w3(32'h39d201e7),
	.w4(32'h3b72d436),
	.w5(32'h3ac9f604),
	.w6(32'hb86c46df),
	.w7(32'h3be0409c),
	.w8(32'h3973ff5d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c3dda),
	.w1(32'h3bdf7307),
	.w2(32'hbb6ab21a),
	.w3(32'hbb195eaa),
	.w4(32'h3bddc7bd),
	.w5(32'hbb18f763),
	.w6(32'hbb83cdc6),
	.w7(32'h3b4fbf72),
	.w8(32'hba973d29),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9831d0),
	.w1(32'hb7c69a0a),
	.w2(32'h3aca56db),
	.w3(32'h3a706592),
	.w4(32'hbaa55f62),
	.w5(32'h39b310e2),
	.w6(32'hb9cd8454),
	.w7(32'h3b127037),
	.w8(32'hbb191f6c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf66e95),
	.w1(32'hbad37fd0),
	.w2(32'hba6afcc4),
	.w3(32'hbb29c5de),
	.w4(32'hba93aed7),
	.w5(32'hba050acd),
	.w6(32'hbb2c9eeb),
	.w7(32'hbabf3db7),
	.w8(32'hbb64c7f0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc07bce),
	.w1(32'h3b3b4599),
	.w2(32'h3bd0d6ae),
	.w3(32'hbb72125b),
	.w4(32'h3b5881ab),
	.w5(32'h3bb22c5a),
	.w6(32'h3a31c65c),
	.w7(32'h3c17de1b),
	.w8(32'hb994c66c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab79a5c),
	.w1(32'hba3974c3),
	.w2(32'h3a231d68),
	.w3(32'h3a927dde),
	.w4(32'h3b332758),
	.w5(32'h39219b51),
	.w6(32'hbbb729db),
	.w7(32'hba3b6861),
	.w8(32'hbaad1eb5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9433f6),
	.w1(32'hbba17561),
	.w2(32'hbbe88ccf),
	.w3(32'hbaa8f397),
	.w4(32'hbbb86503),
	.w5(32'hbc04fe71),
	.w6(32'hbb5ae08a),
	.w7(32'hbbd09299),
	.w8(32'hbb6c83a5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce7d5e),
	.w1(32'hbaa18d7f),
	.w2(32'hbab2ca41),
	.w3(32'hbba2c460),
	.w4(32'hbb6a5a1b),
	.w5(32'hbb2087d4),
	.w6(32'hbaa7775d),
	.w7(32'hba79ee4b),
	.w8(32'hbbe606c6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22e3e9),
	.w1(32'h3a4a39e2),
	.w2(32'hbc14da0f),
	.w3(32'hbb75b07e),
	.w4(32'h3a8a6db3),
	.w5(32'hbc034a72),
	.w6(32'h3bd935a4),
	.w7(32'h3bcd75b2),
	.w8(32'hbb5debef),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc028733),
	.w1(32'h3c25b1e0),
	.w2(32'hbbaf2401),
	.w3(32'hbbb5b42e),
	.w4(32'h3c71ac6f),
	.w5(32'h39e1b72b),
	.w6(32'hbca2a7a8),
	.w7(32'h3bbcbf92),
	.w8(32'hbc01465a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77ecf7),
	.w1(32'h3c81b475),
	.w2(32'h3a823ac3),
	.w3(32'hbc064168),
	.w4(32'h3c3e1ecf),
	.w5(32'hb94c026b),
	.w6(32'hbc986b03),
	.w7(32'h3be47534),
	.w8(32'hbc07fdc5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833a2a),
	.w1(32'h3940981b),
	.w2(32'hb8c105cb),
	.w3(32'hbb812f77),
	.w4(32'h3a76e092),
	.w5(32'h39dfce77),
	.w6(32'hbb85efcd),
	.w7(32'hba84d403),
	.w8(32'hbaae2ccc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba117837),
	.w1(32'hba908157),
	.w2(32'hbab62381),
	.w3(32'hba01d054),
	.w4(32'hba534672),
	.w5(32'hba3f9488),
	.w6(32'h393fc629),
	.w7(32'h3a3cd08b),
	.w8(32'h3b225328),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab070de),
	.w1(32'h3b893a1a),
	.w2(32'h3b8f6332),
	.w3(32'h3ae78c37),
	.w4(32'hb8954f8e),
	.w5(32'hb9281d54),
	.w6(32'h3b990a78),
	.w7(32'h3ba620d1),
	.w8(32'h3bb65668),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd623a),
	.w1(32'h3ae04f6f),
	.w2(32'h3a9b6f8f),
	.w3(32'hbae5d381),
	.w4(32'h3b6298e4),
	.w5(32'h3b12771f),
	.w6(32'hba2b76a7),
	.w7(32'h3b927614),
	.w8(32'h383902b2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1528df),
	.w1(32'hbbf7e7ac),
	.w2(32'hbc7371fa),
	.w3(32'hbc0acb35),
	.w4(32'hbb96c4f2),
	.w5(32'hbc48b6b0),
	.w6(32'hbc6e137c),
	.w7(32'hbc78a411),
	.w8(32'hbc4e799c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a0a4f),
	.w1(32'hbc7148e4),
	.w2(32'hbcc9acf1),
	.w3(32'hba7d2823),
	.w4(32'hbbd8a54d),
	.w5(32'hbc923161),
	.w6(32'hbcad72c3),
	.w7(32'hbc569947),
	.w8(32'hbcbecac7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce3a601),
	.w1(32'hbbb8f297),
	.w2(32'hbc7df954),
	.w3(32'hbc938368),
	.w4(32'h3a088c37),
	.w5(32'hbc35511a),
	.w6(32'hbc586c63),
	.w7(32'hbb9afff3),
	.w8(32'hbc662c3a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc565b94),
	.w1(32'h3b6b3313),
	.w2(32'hbb019cbb),
	.w3(32'hbc2af416),
	.w4(32'h396b940f),
	.w5(32'hbb4e24ce),
	.w6(32'hbc1fa743),
	.w7(32'hb99e97b2),
	.w8(32'hbc1c9503),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9c3de),
	.w1(32'hbc07713c),
	.w2(32'hbc7bf3e3),
	.w3(32'hbc0323a4),
	.w4(32'hbc47f980),
	.w5(32'hbc804c79),
	.w6(32'hbbc12a3a),
	.w7(32'hbc58cf3c),
	.w8(32'hbc3ef316),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae00c98),
	.w1(32'hbae45310),
	.w2(32'h39de1c60),
	.w3(32'hbacf1a86),
	.w4(32'hba9ed0b5),
	.w5(32'h3958041a),
	.w6(32'hbb1641fb),
	.w7(32'hb9f66f6f),
	.w8(32'hbadb9e76),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87341f),
	.w1(32'h3a87f897),
	.w2(32'h3b824918),
	.w3(32'hbae4ac21),
	.w4(32'hba409eac),
	.w5(32'h3b45fc6e),
	.w6(32'hbb19c8ae),
	.w7(32'h3adfad12),
	.w8(32'hb8d3ff31),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d0823),
	.w1(32'hbc631ea4),
	.w2(32'hbc5f1152),
	.w3(32'h3a556428),
	.w4(32'hbc50e4b8),
	.w5(32'hbc5870af),
	.w6(32'hbc3f8faf),
	.w7(32'hbc5bfe94),
	.w8(32'hbc2ce3f7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84f7ff),
	.w1(32'hbc411707),
	.w2(32'hbbc5c158),
	.w3(32'hbc4288b3),
	.w4(32'hbc132c10),
	.w5(32'hb8020094),
	.w6(32'hbc7fb443),
	.w7(32'hb7779e40),
	.w8(32'hbadf13fc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97dc7d),
	.w1(32'h3b61893c),
	.w2(32'h3bb2d162),
	.w3(32'h3c1f297f),
	.w4(32'h3a88bf26),
	.w5(32'h3b2a57d2),
	.w6(32'h3a8e10e5),
	.w7(32'h3bed7b45),
	.w8(32'h3b4d1387),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb87ce7),
	.w1(32'h39cccb46),
	.w2(32'hbc239953),
	.w3(32'hbbdbd283),
	.w4(32'hbaa7b9c4),
	.w5(32'hbc2800ce),
	.w6(32'hbb806609),
	.w7(32'hbbaa7796),
	.w8(32'hbc330ec1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3d028),
	.w1(32'h3b99536e),
	.w2(32'h3b211f18),
	.w3(32'hbbd711e0),
	.w4(32'h3b3e82aa),
	.w5(32'h3a6756a4),
	.w6(32'h3b30b90e),
	.w7(32'h3b448d81),
	.w8(32'h3b443c10),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48349e),
	.w1(32'h375ebf85),
	.w2(32'hbb13536b),
	.w3(32'h3b412b13),
	.w4(32'hbab8c6e2),
	.w5(32'hba62abc8),
	.w6(32'h391900da),
	.w7(32'h3ace717a),
	.w8(32'hbacfce03),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84388f),
	.w1(32'hbb9e93d9),
	.w2(32'hbb8f4143),
	.w3(32'hbb2b5309),
	.w4(32'hbb88231b),
	.w5(32'hbb8ae9f9),
	.w6(32'hbb5066b5),
	.w7(32'hbb5c0199),
	.w8(32'hba3ae4e6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba78ed7d),
	.w1(32'h3abe4ad8),
	.w2(32'h3ac15e8d),
	.w3(32'hbae7f5cd),
	.w4(32'h3b65e555),
	.w5(32'h3a9cdbce),
	.w6(32'h389f4b20),
	.w7(32'hbae5d455),
	.w8(32'h3b07bfaf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf16b4e),
	.w1(32'hbaa6d71c),
	.w2(32'hbb6c4320),
	.w3(32'h3b79d520),
	.w4(32'hba2c06fe),
	.w5(32'hbb5ab2cf),
	.w6(32'hbb31bda7),
	.w7(32'hbb03c8a3),
	.w8(32'hbb4cbcd3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90b60b),
	.w1(32'hbb1526c6),
	.w2(32'hb90ca9e2),
	.w3(32'hbb6f4e55),
	.w4(32'hbb5ab62d),
	.w5(32'hb9b89c0b),
	.w6(32'hbb62e41d),
	.w7(32'h39d0a1c4),
	.w8(32'hbb003b48),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb98aaa),
	.w1(32'hbb27b4a7),
	.w2(32'hbbdd561b),
	.w3(32'hbbbfa04e),
	.w4(32'hbb1b329b),
	.w5(32'hbbc80913),
	.w6(32'hbb823961),
	.w7(32'hbb5fb2b8),
	.w8(32'hbb76f83a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08ffd6),
	.w1(32'hbb252084),
	.w2(32'hb8b715ff),
	.w3(32'hbbd22151),
	.w4(32'hbba67e8d),
	.w5(32'h39c7fdb6),
	.w6(32'hbb38094d),
	.w7(32'h3ae1ca41),
	.w8(32'h3a7b2134),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b748c5e),
	.w1(32'hbabc6378),
	.w2(32'h3b8d78fd),
	.w3(32'h3aa17a99),
	.w4(32'hbb8261a1),
	.w5(32'h3b849166),
	.w6(32'hb949dcfe),
	.w7(32'h3b8a7efb),
	.w8(32'hbae44916),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed0b5b),
	.w1(32'hbb41cc33),
	.w2(32'hbb84d83c),
	.w3(32'hbb15f6c9),
	.w4(32'hbacd0b6e),
	.w5(32'hbb7b137c),
	.w6(32'hba7be632),
	.w7(32'hbba18b5c),
	.w8(32'hba8014ff),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134168),
	.w1(32'hbb074014),
	.w2(32'hbafa916f),
	.w3(32'hba3573a4),
	.w4(32'hbb2cfbf7),
	.w5(32'hbb347161),
	.w6(32'hba71422f),
	.w7(32'hbad71696),
	.w8(32'h398ce628),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a54f61),
	.w1(32'hbbb46bc4),
	.w2(32'hbb9fe274),
	.w3(32'hb9a5d6a6),
	.w4(32'hbb6b0810),
	.w5(32'hbb8360f5),
	.w6(32'hbb8f7d52),
	.w7(32'hbbd2f81b),
	.w8(32'hba53e568),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993f51),
	.w1(32'hbb82d83f),
	.w2(32'hbbf47e2b),
	.w3(32'hbc1d602d),
	.w4(32'hbbe8e9ea),
	.w5(32'hbba9d32b),
	.w6(32'hbbb6a025),
	.w7(32'hbba156ce),
	.w8(32'hbb80e81e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23d20a),
	.w1(32'hb94fbbf6),
	.w2(32'hbc2b08fa),
	.w3(32'hbbfa4669),
	.w4(32'h3af87713),
	.w5(32'hbc265b02),
	.w6(32'hbbfe43a5),
	.w7(32'hb990b1e8),
	.w8(32'hbc3414c6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc076c34),
	.w1(32'h3b674d0b),
	.w2(32'hbb67e03a),
	.w3(32'hbb73e09f),
	.w4(32'h3b57d6be),
	.w5(32'hbb60b77a),
	.w6(32'hbc4aab2d),
	.w7(32'h3b3fc657),
	.w8(32'hbbd0b7a3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe74182),
	.w1(32'hbc0de1c5),
	.w2(32'hbcfa0675),
	.w3(32'hbb2bd02f),
	.w4(32'h3a849e82),
	.w5(32'hbcb27096),
	.w6(32'hbd01dcd4),
	.w7(32'hbc2ef5cf),
	.w8(32'hbcc6b843),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc806bae),
	.w1(32'hbb91c930),
	.w2(32'hbba7b332),
	.w3(32'hbc88840d),
	.w4(32'hbb6c744f),
	.w5(32'hbb9a811f),
	.w6(32'hbb235074),
	.w7(32'hbb922973),
	.w8(32'hbb4dd390),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d956),
	.w1(32'hb92235f3),
	.w2(32'h3950ca2a),
	.w3(32'hbb621b45),
	.w4(32'hbb10a3ad),
	.w5(32'hba863f99),
	.w6(32'hba934baa),
	.w7(32'h3a068092),
	.w8(32'hba660083),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11108e),
	.w1(32'hbaa4ecae),
	.w2(32'h3a4ed7fe),
	.w3(32'hbb17687c),
	.w4(32'hbb3fd6d0),
	.w5(32'h39522875),
	.w6(32'hbb2c5ecd),
	.w7(32'h3a570262),
	.w8(32'hba7b0edc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7118c),
	.w1(32'h39a7b904),
	.w2(32'h3af3ea98),
	.w3(32'hbb2f0d66),
	.w4(32'hba56b3a0),
	.w5(32'hb9a1b121),
	.w6(32'hbb93fe05),
	.w7(32'h3a5eb325),
	.w8(32'hbb4f92e8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab69bfd),
	.w1(32'h3929cddd),
	.w2(32'h39cdd38d),
	.w3(32'hbb4322db),
	.w4(32'hba46bfab),
	.w5(32'hba3b419b),
	.w6(32'h3a8d5d2c),
	.w7(32'h3a07b1a5),
	.w8(32'h3a8df2cb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb204e77),
	.w1(32'h3b844581),
	.w2(32'h3bd764c3),
	.w3(32'hbbb70d15),
	.w4(32'hbbdf8ab3),
	.w5(32'hbac93bb5),
	.w6(32'hbba1822a),
	.w7(32'h3a70d753),
	.w8(32'h3aa904e0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef5b5d),
	.w1(32'hbb501dcf),
	.w2(32'hba9cebe9),
	.w3(32'hbbd18574),
	.w4(32'hbb2f9562),
	.w5(32'hba3953cc),
	.w6(32'hbc248ac6),
	.w7(32'h39b97e7b),
	.w8(32'hbb297884),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb345591),
	.w1(32'hbb87ac71),
	.w2(32'hbc1a9a83),
	.w3(32'hbb694990),
	.w4(32'hba73d97d),
	.w5(32'hbbd1e2a7),
	.w6(32'hbc138206),
	.w7(32'hbb405067),
	.w8(32'hbc022b3d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17bbe6),
	.w1(32'hb9b1d1bc),
	.w2(32'hbb66ccf4),
	.w3(32'hbbedf96a),
	.w4(32'h3ac22dca),
	.w5(32'hbb4ea4c6),
	.w6(32'hbba9d66a),
	.w7(32'hb9befcea),
	.w8(32'hbb3754eb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba090481),
	.w1(32'hbae28e44),
	.w2(32'h38233185),
	.w3(32'hbb56f8c3),
	.w4(32'hbb9b4c27),
	.w5(32'hbaff78fe),
	.w6(32'hba8dad20),
	.w7(32'h3b781b16),
	.w8(32'hbbbc313c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e123b),
	.w1(32'h3a942915),
	.w2(32'hbb8bc1d2),
	.w3(32'hbb162413),
	.w4(32'h3b471acf),
	.w5(32'hbaa74a48),
	.w6(32'h392702bd),
	.w7(32'h3b402760),
	.w8(32'hba7330b0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c973b),
	.w1(32'h3a85e380),
	.w2(32'hb8ebedd1),
	.w3(32'hbb81a2b8),
	.w4(32'hba465182),
	.w5(32'hbb3ae725),
	.w6(32'h3aff785a),
	.w7(32'h3b05b822),
	.w8(32'h39b675e5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6d628),
	.w1(32'h3ac4349c),
	.w2(32'h3ae8271a),
	.w3(32'h3b858c39),
	.w4(32'hba357979),
	.w5(32'hb9fd47de),
	.w6(32'h3ac168f5),
	.w7(32'h3b00e8a5),
	.w8(32'h3b18216b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad96192),
	.w1(32'hba9596e5),
	.w2(32'hba98e07a),
	.w3(32'h398bb882),
	.w4(32'hba7a1c71),
	.w5(32'hbaa941a2),
	.w6(32'hb9d23b0d),
	.w7(32'hbaa1f9a8),
	.w8(32'hbaa0e164),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb1233),
	.w1(32'h3a9837e6),
	.w2(32'hbb1ac293),
	.w3(32'hbad3de30),
	.w4(32'h3a9dee85),
	.w5(32'hbb477ad3),
	.w6(32'h3b87e261),
	.w7(32'h3a4dee2e),
	.w8(32'hbace19c5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80a68c),
	.w1(32'h39b44db5),
	.w2(32'hb8d81205),
	.w3(32'hbb9e7b2d),
	.w4(32'h39ba92a2),
	.w5(32'hb9b1a40c),
	.w6(32'h39a4ac59),
	.w7(32'h39424ec0),
	.w8(32'h3916c628),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf391f8),
	.w1(32'hbaca996f),
	.w2(32'hbb4873f9),
	.w3(32'hbbd828c8),
	.w4(32'h3a74817a),
	.w5(32'hb9d8ff0b),
	.w6(32'hbc4ef529),
	.w7(32'hba55b09d),
	.w8(32'hbb86037a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6871b),
	.w1(32'h3a70010a),
	.w2(32'h3b003062),
	.w3(32'hbb860da7),
	.w4(32'h39110923),
	.w5(32'h3aa93316),
	.w6(32'hbb0c8705),
	.w7(32'h3b362560),
	.w8(32'hba9df527),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb92f7d),
	.w1(32'h3ba530c9),
	.w2(32'h3a4f7768),
	.w3(32'hbb5a8f7b),
	.w4(32'h3bcee1a2),
	.w5(32'h3a71c929),
	.w6(32'h3b430b99),
	.w7(32'h3ba46650),
	.w8(32'h3a17997f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fee45),
	.w1(32'hbbb1fcef),
	.w2(32'hbba16a9a),
	.w3(32'hbc0c287f),
	.w4(32'hbbe8b848),
	.w5(32'hbbb0be86),
	.w6(32'hbc84312b),
	.w7(32'hbbb331ca),
	.w8(32'hbc099715),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba846f8f),
	.w1(32'h3c285d46),
	.w2(32'h3b7e6148),
	.w3(32'hbb82c6af),
	.w4(32'h3c029280),
	.w5(32'h3b5d859b),
	.w6(32'hbb0d5322),
	.w7(32'h3c0bd48b),
	.w8(32'hba8002d1),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23d236),
	.w1(32'hbc3e5f39),
	.w2(32'hbc8a02d7),
	.w3(32'hbafa727e),
	.w4(32'hbbfa0079),
	.w5(32'hbc58f0c6),
	.w6(32'hbc15a3db),
	.w7(32'hbc6a5d9e),
	.w8(32'hbc873b6f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14cbf0),
	.w1(32'h3be7de0b),
	.w2(32'h3a3d740c),
	.w3(32'hbbf03c18),
	.w4(32'h3bca7267),
	.w5(32'hb9fb25d4),
	.w6(32'h3b71a03c),
	.w7(32'h3bd99c1f),
	.w8(32'h3b3ff8ce),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0bd80),
	.w1(32'hbb1c3ac6),
	.w2(32'hbbeb4491),
	.w3(32'hbb734d74),
	.w4(32'h3a8691cb),
	.w5(32'hbb13d4bf),
	.w6(32'hbbbf1008),
	.w7(32'h3b156da6),
	.w8(32'hbba07a87),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb30d17),
	.w1(32'hb9271ac4),
	.w2(32'hbb7613ca),
	.w3(32'hbb82f772),
	.w4(32'h3af2afb4),
	.w5(32'hba4dc560),
	.w6(32'hbb654ede),
	.w7(32'hba8b76cf),
	.w8(32'hbb1f8909),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5cc2),
	.w1(32'h3b5984b2),
	.w2(32'hbb0bb4d1),
	.w3(32'hbbca174e),
	.w4(32'h3b35abf8),
	.w5(32'hbb90927b),
	.w6(32'hba3831c2),
	.w7(32'h3c1ecf69),
	.w8(32'h39a2cb2f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb659036),
	.w1(32'h39fb5a10),
	.w2(32'hbb27a0ec),
	.w3(32'hbc04fe6e),
	.w4(32'h3aff3050),
	.w5(32'hb9e3cc6f),
	.w6(32'h39aee979),
	.w7(32'hbb1d1889),
	.w8(32'h38ea0881),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec3af3),
	.w1(32'hbbabdc8d),
	.w2(32'hbc105c00),
	.w3(32'hba205257),
	.w4(32'hbb2362b9),
	.w5(32'hbbdcc9a1),
	.w6(32'hbc3c8d81),
	.w7(32'hbac39bf9),
	.w8(32'hbc1a60b8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb079b16),
	.w1(32'h3b7b6d30),
	.w2(32'hbb531a6e),
	.w3(32'hbb185066),
	.w4(32'h3b45b8ff),
	.w5(32'hbb1913be),
	.w6(32'hba6b9290),
	.w7(32'h3ae65d19),
	.w8(32'hbb8b997f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaefbe0),
	.w1(32'h3a3516d1),
	.w2(32'hbc221117),
	.w3(32'hba07ac99),
	.w4(32'h3adfc4c7),
	.w5(32'hbc04a311),
	.w6(32'hbabd359b),
	.w7(32'h3a45468d),
	.w8(32'hbc1dc92c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf2945),
	.w1(32'h3c35b37a),
	.w2(32'h3a8a170c),
	.w3(32'hbb9cc1ac),
	.w4(32'h3cbc793d),
	.w5(32'h3bf7dbb7),
	.w6(32'hbc6595a8),
	.w7(32'h3c0b4e5c),
	.w8(32'h3a27c419),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5e8a7),
	.w1(32'h3ac264dc),
	.w2(32'hbc0ce8f9),
	.w3(32'h3b2b7c7c),
	.w4(32'h3b9e6d89),
	.w5(32'hbbeb1a1b),
	.w6(32'hba678a55),
	.w7(32'h3ac1dc24),
	.w8(32'hbbb5284d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7eab7),
	.w1(32'hbb538c75),
	.w2(32'hba680504),
	.w3(32'hbbe70543),
	.w4(32'hbb694070),
	.w5(32'h3a50d93d),
	.w6(32'hba9f1c11),
	.w7(32'h3bbe387a),
	.w8(32'hbb8c7466),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef768a),
	.w1(32'hb88d6737),
	.w2(32'h3aaa9cda),
	.w3(32'h3b9dd5a2),
	.w4(32'hbb1ff21d),
	.w5(32'hb9cad768),
	.w6(32'hbb23acb5),
	.w7(32'h39467cff),
	.w8(32'hbb1117c9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc710c39),
	.w1(32'hbba0ae3e),
	.w2(32'hbb90652a),
	.w3(32'hbc37121e),
	.w4(32'hb9a0cace),
	.w5(32'hbaf92553),
	.w6(32'hbb43833a),
	.w7(32'h3c059ee1),
	.w8(32'h378d6834),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb724d),
	.w1(32'hbaf3b238),
	.w2(32'hbb1b248a),
	.w3(32'hba2f845a),
	.w4(32'hbb2a9f98),
	.w5(32'hbb5b2f59),
	.w6(32'hbbb99855),
	.w7(32'hb95f61eb),
	.w8(32'hbbb161f0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dda7a2),
	.w1(32'hbac5c591),
	.w2(32'hbb00b742),
	.w3(32'hb9a531dd),
	.w4(32'hb9e52d66),
	.w5(32'hbaa970d4),
	.w6(32'hba4b75b5),
	.w7(32'hba9c0a7c),
	.w8(32'hba91c205),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68092b),
	.w1(32'h3ac77590),
	.w2(32'h3b6f0ffa),
	.w3(32'hbb0c4e4d),
	.w4(32'h3a5d2031),
	.w5(32'h3b38fffd),
	.w6(32'hbabe3c94),
	.w7(32'h3ba226c2),
	.w8(32'hba2ebf11),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eadfe),
	.w1(32'hbb48f794),
	.w2(32'hbb01a5d9),
	.w3(32'hbbbd029c),
	.w4(32'hbb8d05b4),
	.w5(32'hbb184255),
	.w6(32'hbbfa1127),
	.w7(32'hbb7206d4),
	.w8(32'hbbeb95d0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdc7ba),
	.w1(32'hbc1076b2),
	.w2(32'hbc5a5e2e),
	.w3(32'h3ae99d35),
	.w4(32'hbbe3ba2a),
	.w5(32'hbc3adbee),
	.w6(32'hbc538623),
	.w7(32'hbbf55439),
	.w8(32'hbc3f2604),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eb70a),
	.w1(32'h3a7504ef),
	.w2(32'h3a737a0e),
	.w3(32'hbc4cea54),
	.w4(32'h39cac435),
	.w5(32'h3b10bd5f),
	.w6(32'hbc1410da),
	.w7(32'h3ae6e412),
	.w8(32'hbbbef0bf),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93c46c),
	.w1(32'hbb615e66),
	.w2(32'hbaeb904d),
	.w3(32'h3a8a446d),
	.w4(32'hbb05aa41),
	.w5(32'h3ad89344),
	.w6(32'hbbf0ed95),
	.w7(32'h3b69f4a3),
	.w8(32'hbb9f5da7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fc20b),
	.w1(32'h3b7a5f0c),
	.w2(32'h3b672afc),
	.w3(32'hbb105913),
	.w4(32'h3b383f58),
	.w5(32'h3b7b372f),
	.w6(32'hbbafef3f),
	.w7(32'h3ba37a61),
	.w8(32'hbab0488f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb688257),
	.w1(32'hbbdd515c),
	.w2(32'hbc2236f1),
	.w3(32'hb9709671),
	.w4(32'hbb4c757e),
	.w5(32'hbbf565c1),
	.w6(32'hbbb60951),
	.w7(32'hbb9f4c7a),
	.w8(32'hbbc2fd5d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf537bb),
	.w1(32'hba7c6c52),
	.w2(32'h39ed8337),
	.w3(32'hbbcdac13),
	.w4(32'hb9c1adf3),
	.w5(32'h38b2bb88),
	.w6(32'hbbba3590),
	.w7(32'h3a4cff8d),
	.w8(32'hbb336075),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2befbf),
	.w1(32'h3a3440ee),
	.w2(32'h3ba91953),
	.w3(32'h3a4490bc),
	.w4(32'hba018e21),
	.w5(32'h3ba5825e),
	.w6(32'hbb24ee1b),
	.w7(32'h3b7622d4),
	.w8(32'h3b052b26),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aee07),
	.w1(32'h3a02db25),
	.w2(32'h3aea674b),
	.w3(32'h3b4d26ed),
	.w4(32'hb9c5aba3),
	.w5(32'h3acd892e),
	.w6(32'hba9932df),
	.w7(32'h3b2839d2),
	.w8(32'h3a2d44ec),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4bece),
	.w1(32'h3b19726b),
	.w2(32'h3b767b53),
	.w3(32'hb9215d65),
	.w4(32'h3a3a6667),
	.w5(32'h3b4f250b),
	.w6(32'h395b204c),
	.w7(32'h3b81cb82),
	.w8(32'h3affe435),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3566ec),
	.w1(32'hbb751d2a),
	.w2(32'hba148b38),
	.w3(32'h3a9c1d69),
	.w4(32'hbae6f398),
	.w5(32'h3b35509f),
	.w6(32'hb9a6bca3),
	.w7(32'h3aca58c2),
	.w8(32'h3b8f9db4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb354404),
	.w1(32'hbaf0b6bf),
	.w2(32'hbc1192da),
	.w3(32'h397de794),
	.w4(32'h3a95ba26),
	.w5(32'hbbf51652),
	.w6(32'hbbb91182),
	.w7(32'hbb5585a7),
	.w8(32'hbb7f3af5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada3adc),
	.w1(32'h39d32f18),
	.w2(32'hbb3b4f6c),
	.w3(32'hba421e65),
	.w4(32'h39a7e0d7),
	.w5(32'hbb52b1ca),
	.w6(32'hbaf55e9f),
	.w7(32'hbb064b32),
	.w8(32'hbc2122cf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc294d28),
	.w1(32'hbbc4a838),
	.w2(32'hbc105dfb),
	.w3(32'hbc33b0d3),
	.w4(32'hbc05e6b0),
	.w5(32'hbc079619),
	.w6(32'hbb9aeea4),
	.w7(32'hbb84056b),
	.w8(32'hbbd79587),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4540b3),
	.w1(32'hba6c2316),
	.w2(32'hbac08f03),
	.w3(32'hbc33f793),
	.w4(32'h3aee7ea9),
	.w5(32'h3ab7ee0c),
	.w6(32'hbc32d646),
	.w7(32'h3b0bea53),
	.w8(32'hbbd715f6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a522adf),
	.w1(32'hbbfc4e8c),
	.w2(32'hbb711242),
	.w3(32'hba14d558),
	.w4(32'hbbd4b7e0),
	.w5(32'hbb672c03),
	.w6(32'hbace850d),
	.w7(32'hba5b0859),
	.w8(32'h3b23da46),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6eeb4b),
	.w1(32'h3be3eee1),
	.w2(32'h3bd7156b),
	.w3(32'hbb0fe684),
	.w4(32'h3b8644ee),
	.w5(32'h3b7b68d7),
	.w6(32'h3c01796e),
	.w7(32'h3c2bb37b),
	.w8(32'h3bc1abbb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b667f46),
	.w1(32'h3a9f9698),
	.w2(32'h3b8a9585),
	.w3(32'hba17fdb8),
	.w4(32'hba558980),
	.w5(32'h3b3855c3),
	.w6(32'hba8aff58),
	.w7(32'h3b830743),
	.w8(32'hbae6a1dd),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacee681),
	.w1(32'hb945f0e1),
	.w2(32'hb90dd49f),
	.w3(32'hbb5bf61d),
	.w4(32'hba015ee2),
	.w5(32'h3900d1aa),
	.w6(32'hbaed9454),
	.w7(32'hbacdd983),
	.w8(32'hbaefdd61),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62af60),
	.w1(32'hbbbb2399),
	.w2(32'hbb9f841b),
	.w3(32'hbaa34a25),
	.w4(32'hbba98527),
	.w5(32'hbbde951b),
	.w6(32'hba66ef4c),
	.w7(32'hbb89af6c),
	.w8(32'hbbbaac5b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd6ccd),
	.w1(32'hbb25c141),
	.w2(32'hbbebd943),
	.w3(32'hbba0337c),
	.w4(32'hbb24ed9d),
	.w5(32'hbbd5972c),
	.w6(32'hbb856753),
	.w7(32'hbb384577),
	.w8(32'hbc03ca92),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba202142),
	.w1(32'hba471100),
	.w2(32'hba3f55eb),
	.w3(32'hb9c0f369),
	.w4(32'hba060f1b),
	.w5(32'hb973b2c8),
	.w6(32'h39b32ac9),
	.w7(32'h37dcfbab),
	.w8(32'hb936a7c9),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee08ed),
	.w1(32'h39d205a0),
	.w2(32'hbabee837),
	.w3(32'hbad7c0c1),
	.w4(32'h3860ee85),
	.w5(32'hba86be31),
	.w6(32'hbb618d97),
	.w7(32'hba000f3b),
	.w8(32'hbb1665f2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb1af7),
	.w1(32'h3a0bc9b0),
	.w2(32'hbab50397),
	.w3(32'hbadb4781),
	.w4(32'h3abdbdb0),
	.w5(32'hba05eb82),
	.w6(32'hbabd6ac4),
	.w7(32'h3aa396e2),
	.w8(32'hbae0cdae),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb357e76),
	.w1(32'hb7910cf4),
	.w2(32'hbb212b96),
	.w3(32'hba8220d3),
	.w4(32'h3a22892f),
	.w5(32'hba9ce204),
	.w6(32'hbb073594),
	.w7(32'hb8e74d2f),
	.w8(32'hbb01d4fe),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0a48b),
	.w1(32'hba272653),
	.w2(32'hbb87a2b4),
	.w3(32'hbb3d0cbf),
	.w4(32'h3b37ce90),
	.w5(32'h399d4d96),
	.w6(32'hbb3fa209),
	.w7(32'h3ae9999a),
	.w8(32'hb9f850e7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac603c),
	.w1(32'hbb44f172),
	.w2(32'hbbf861d7),
	.w3(32'hbbc58316),
	.w4(32'hbb8c8ea0),
	.w5(32'hbc02bbe0),
	.w6(32'hbb803b3e),
	.w7(32'hbb8c31ba),
	.w8(32'hbc10caa9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941935),
	.w1(32'h3a38eb9a),
	.w2(32'hbafb86ba),
	.w3(32'hbb16b0b3),
	.w4(32'h3b57ebe7),
	.w5(32'h393fbf9a),
	.w6(32'hbb87265b),
	.w7(32'h3a9a8b28),
	.w8(32'hbb5cbe6c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb881462),
	.w1(32'hba9499b7),
	.w2(32'hbb858919),
	.w3(32'hbace7802),
	.w4(32'h3b074e89),
	.w5(32'hba3a55f7),
	.w6(32'hbb30f1d9),
	.w7(32'hba5ff1f7),
	.w8(32'hbbb33f19),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02f163),
	.w1(32'hbb91179e),
	.w2(32'hbbed21b6),
	.w3(32'hbbaa6d1f),
	.w4(32'hbb933b7a),
	.w5(32'hbc00c07b),
	.w6(32'hbb28029f),
	.w7(32'hbaedeb84),
	.w8(32'hbbb304ae),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcd8db),
	.w1(32'hb98e9f41),
	.w2(32'hba60f5eb),
	.w3(32'hbb48aadd),
	.w4(32'h3ae4fcf5),
	.w5(32'h3a089ef6),
	.w6(32'hbbaab586),
	.w7(32'h38889c42),
	.w8(32'hbb0e6bc6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cbc7d),
	.w1(32'hbabf7bd8),
	.w2(32'hbb8c0c50),
	.w3(32'hbb200f0f),
	.w4(32'hba50a10f),
	.w5(32'hbb807614),
	.w6(32'hbae159dd),
	.w7(32'hbae2f42d),
	.w8(32'hbbae1c99),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a4fb5),
	.w1(32'h39e46be3),
	.w2(32'hba9baf64),
	.w3(32'hb904fcd9),
	.w4(32'h3a8bfc52),
	.w5(32'hba3f08f6),
	.w6(32'hba734560),
	.w7(32'h39b2b5dd),
	.w8(32'hbab2d63e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89558d),
	.w1(32'h3c042f28),
	.w2(32'h38b516a9),
	.w3(32'hbbe13f0d),
	.w4(32'h3bc26d1d),
	.w5(32'hbaa2d9cd),
	.w6(32'hbbf62cc0),
	.w7(32'h3b9074bf),
	.w8(32'hbb9d33df),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77995d),
	.w1(32'h3aef40f4),
	.w2(32'h3b18142f),
	.w3(32'hbb7d344e),
	.w4(32'h39fe148e),
	.w5(32'h3aa5f7fb),
	.w6(32'hbba751c6),
	.w7(32'hb8939271),
	.w8(32'hba9d0ab4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb817a825),
	.w1(32'hb83fa4e5),
	.w2(32'hb82e0b8b),
	.w3(32'hb8c5673f),
	.w4(32'hb8e9259f),
	.w5(32'hb8c41c01),
	.w6(32'hb81338ed),
	.w7(32'hb8483423),
	.w8(32'hb79dda02),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382b6c08),
	.w1(32'h38b0ca40),
	.w2(32'h382eeda8),
	.w3(32'hb6d53905),
	.w4(32'h364e2c76),
	.w5(32'h35c97876),
	.w6(32'h38c36ec7),
	.w7(32'h390ea930),
	.w8(32'h39025abc),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18c9a1),
	.w1(32'hba175c70),
	.w2(32'hbab19a91),
	.w3(32'hbb2332d9),
	.w4(32'h38e513cf),
	.w5(32'h39c248fc),
	.w6(32'hbb34507e),
	.w7(32'hb8f857ef),
	.w8(32'hba785216),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe90439),
	.w1(32'h3a0c6586),
	.w2(32'hba0c8748),
	.w3(32'hbb87b3cb),
	.w4(32'h3b831a43),
	.w5(32'h3a692d5b),
	.w6(32'hbbbeb936),
	.w7(32'h3b191520),
	.w8(32'hbb5e4ebf),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb8b15),
	.w1(32'h384633a7),
	.w2(32'hbb896504),
	.w3(32'hbbee3fcf),
	.w4(32'h3b01974f),
	.w5(32'hbb4043b7),
	.w6(32'hbbff2214),
	.w7(32'hba6f46d6),
	.w8(32'hbba6ba94),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aea2a0),
	.w1(32'h35ca4822),
	.w2(32'h3784e583),
	.w3(32'h382e79bf),
	.w4(32'h378e0f1d),
	.w5(32'h380ab812),
	.w6(32'h38808049),
	.w7(32'h37fcff7c),
	.w8(32'h38846527),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca1e50),
	.w1(32'hbab3824c),
	.w2(32'hbbdeebe4),
	.w3(32'hbb9c235f),
	.w4(32'hb9bed2cb),
	.w5(32'hbbb92caf),
	.w6(32'hbbbc84a9),
	.w7(32'hbaebdbe5),
	.w8(32'hbbdf6823),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dc351),
	.w1(32'hb9164e10),
	.w2(32'hbb19bb7d),
	.w3(32'hbb2ebe7a),
	.w4(32'h3710ebce),
	.w5(32'hbadc9f06),
	.w6(32'hbb861a6f),
	.w7(32'hbaf6e3a6),
	.w8(32'hbb90baeb),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb620586),
	.w1(32'hbb8bc7fd),
	.w2(32'hbc12ccea),
	.w3(32'hbb8ef543),
	.w4(32'hbb548dc6),
	.w5(32'hbbd11c16),
	.w6(32'hba4792be),
	.w7(32'hbb2154a8),
	.w8(32'hbbbc7178),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82a011),
	.w1(32'h3c00325d),
	.w2(32'hbb400e5d),
	.w3(32'h39f41318),
	.w4(32'h3c1fc7e3),
	.w5(32'hba71d0a8),
	.w6(32'hbb721b73),
	.w7(32'h3bd336db),
	.w8(32'hba31eecf),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb191377),
	.w1(32'h3a0dc7fb),
	.w2(32'h39dfb312),
	.w3(32'hbaff3585),
	.w4(32'h3a96a28c),
	.w5(32'h39a8e897),
	.w6(32'hbb791c5d),
	.w7(32'h39e09e4a),
	.w8(32'hbad04d72),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cc5f6),
	.w1(32'h3a8caad3),
	.w2(32'h3a906112),
	.w3(32'h3a69651a),
	.w4(32'h3a49a185),
	.w5(32'h3a5b809d),
	.w6(32'h3a816999),
	.w7(32'h3a808788),
	.w8(32'h3a7a007e),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb159d7a),
	.w1(32'h3b96b80d),
	.w2(32'h3aa3cd9a),
	.w3(32'h39449711),
	.w4(32'h3bcad20d),
	.w5(32'h3b1c0f9f),
	.w6(32'hbb54fc73),
	.w7(32'h3b89b936),
	.w8(32'h3a19317f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb971054),
	.w1(32'h3baa0471),
	.w2(32'h3a065431),
	.w3(32'hbb8dd4de),
	.w4(32'h3bdcba2e),
	.w5(32'h3af2ee7b),
	.w6(32'hbbe8db30),
	.w7(32'h3b8ed12d),
	.w8(32'hbb3877ee),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e8d29),
	.w1(32'h3bc03ad0),
	.w2(32'h38d452fe),
	.w3(32'hb9d5e791),
	.w4(32'h3bc5ee0f),
	.w5(32'h3a8e43a5),
	.w6(32'hbb45adf4),
	.w7(32'h3b996445),
	.w8(32'hb9d8f549),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b7685),
	.w1(32'hba649393),
	.w2(32'hba8497f1),
	.w3(32'hbb08d4c8),
	.w4(32'hbae9a47d),
	.w5(32'hba9a8a3b),
	.w6(32'hba731e2a),
	.w7(32'hba80450c),
	.w8(32'hba9452a1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986f4b1),
	.w1(32'hb9e4b393),
	.w2(32'hb9bc8386),
	.w3(32'hb9b0554d),
	.w4(32'hb94e4513),
	.w5(32'hb8bb64a6),
	.w6(32'hba1324f8),
	.w7(32'hb9eec409),
	.w8(32'hb9ee406e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc32898),
	.w1(32'hbb119747),
	.w2(32'hbba7d81c),
	.w3(32'hbb8e11ff),
	.w4(32'hbaa645d5),
	.w5(32'hbb945eba),
	.w6(32'hbb8c99cc),
	.w7(32'hbb11ea5a),
	.w8(32'hbbad1834),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b272a8),
	.w1(32'hb932efbe),
	.w2(32'hba2aeebc),
	.w3(32'hb94ce035),
	.w4(32'hb9bcc64c),
	.w5(32'hba2688c1),
	.w6(32'h3a09a617),
	.w7(32'h39a2004a),
	.w8(32'hb95b3281),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc27b0),
	.w1(32'h3b11d225),
	.w2(32'hba516696),
	.w3(32'h3a1e5934),
	.w4(32'h3b56714f),
	.w5(32'h39d53e57),
	.w6(32'hb9f9f968),
	.w7(32'h3b4e7930),
	.w8(32'h3865c8ed),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39354590),
	.w1(32'hb84a4747),
	.w2(32'hb9a846f6),
	.w3(32'h393d3702),
	.w4(32'h397b7226),
	.w5(32'h37c23a32),
	.w6(32'h3932ea65),
	.w7(32'h3a0244d5),
	.w8(32'h392c1448),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea440f),
	.w1(32'h39fdb317),
	.w2(32'hbba91a74),
	.w3(32'hbb596146),
	.w4(32'hbac93f23),
	.w5(32'hbbe44c56),
	.w6(32'hbb229cad),
	.w7(32'hbab91241),
	.w8(32'hbbe1f845),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4c070),
	.w1(32'h3663d98d),
	.w2(32'h392da100),
	.w3(32'h38b26b10),
	.w4(32'h3675759c),
	.w5(32'h3909558d),
	.w6(32'h39411022),
	.w7(32'h38d227f1),
	.w8(32'h39347b72),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ce906),
	.w1(32'hb72401e5),
	.w2(32'hb9631a3a),
	.w3(32'hb946de16),
	.w4(32'hb88e8a7a),
	.w5(32'hb981a33d),
	.w6(32'hb8b6fbab),
	.w7(32'hb898ac1b),
	.w8(32'hb99a21a2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3198ca),
	.w1(32'h3aceae92),
	.w2(32'h398d55c0),
	.w3(32'hba770825),
	.w4(32'h3b5ca7b6),
	.w5(32'h3adddbed),
	.w6(32'hbb2bf1e7),
	.w7(32'h3adc9ec7),
	.w8(32'hbab53995),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf54520),
	.w1(32'hba138783),
	.w2(32'hbbca1e6c),
	.w3(32'hbbda28ca),
	.w4(32'hbb0cbf5a),
	.w5(32'hbc4572b7),
	.w6(32'hbbd23e9a),
	.w7(32'hbb0ff77d),
	.w8(32'hbc5bbe8a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96178a6),
	.w1(32'h3b27d1a1),
	.w2(32'hba9a0d41),
	.w3(32'hba64b5b7),
	.w4(32'h3ad354cd),
	.w5(32'hbad7bb36),
	.w6(32'hbb2a15f0),
	.w7(32'h3a78624e),
	.w8(32'hbb08a881),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9796f6),
	.w1(32'hba387406),
	.w2(32'hbb9b2143),
	.w3(32'hbae1cbf0),
	.w4(32'h3a42f3fa),
	.w5(32'hbb7ca065),
	.w6(32'hbb7ad8e0),
	.w7(32'hba85abac),
	.w8(32'hbbe02b70),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3813572e),
	.w1(32'h3a4efe68),
	.w2(32'hba40f9a7),
	.w3(32'hbb0658a1),
	.w4(32'hb9a89e33),
	.w5(32'hba823a4e),
	.w6(32'hba604c5c),
	.w7(32'h39aee996),
	.w8(32'hb9c56538),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f4a47),
	.w1(32'h3a1a042c),
	.w2(32'hbc2d8fcc),
	.w3(32'hbbf3df48),
	.w4(32'h3bb31980),
	.w5(32'hbbbd1d92),
	.w6(32'hbc16154a),
	.w7(32'h3a697dca),
	.w8(32'hbbe293d7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf5795),
	.w1(32'h3a06d139),
	.w2(32'hbbcd7ce5),
	.w3(32'hbb9825c6),
	.w4(32'h3b377c50),
	.w5(32'hbb634343),
	.w6(32'hbbc3a293),
	.w7(32'h3a89ca57),
	.w8(32'hbba9dac2),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4460),
	.w1(32'hba46aab3),
	.w2(32'hbbcc51cc),
	.w3(32'hbb2c6518),
	.w4(32'hba89127e),
	.w5(32'hbbddc4e8),
	.w6(32'hbb57020a),
	.w7(32'hbaeb5b33),
	.w8(32'hbbd48a6d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ed55dc),
	.w1(32'h38f98f18),
	.w2(32'h39ca1edc),
	.w3(32'hb9193cfb),
	.w4(32'h395a4307),
	.w5(32'h39fddd42),
	.w6(32'h387a2c10),
	.w7(32'h39c6bb79),
	.w8(32'h3a1bc5ed),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9507f0),
	.w1(32'hbaef1c7f),
	.w2(32'hbb37e95a),
	.w3(32'hbb4b6817),
	.w4(32'hba4f6f24),
	.w5(32'hbad06e2c),
	.w6(32'hbae2d3d7),
	.w7(32'hb9e3be68),
	.w8(32'hbafdb604),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8e0ed),
	.w1(32'h35d8858d),
	.w2(32'h38c9eae4),
	.w3(32'h38b0ead6),
	.w4(32'hb82f1311),
	.w5(32'h38929392),
	.w6(32'h391b76e4),
	.w7(32'h38295b16),
	.w8(32'h39272c8d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33f1ab),
	.w1(32'h38e4ed2a),
	.w2(32'hbb17c30f),
	.w3(32'hb8f6b4c5),
	.w4(32'h393d9ee3),
	.w5(32'hba5518fd),
	.w6(32'hbabd079c),
	.w7(32'hba9ba264),
	.w8(32'hbb2eb425),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91cd39),
	.w1(32'h39d0af15),
	.w2(32'hba15dbf9),
	.w3(32'hbade43c4),
	.w4(32'h38a3e5b2),
	.w5(32'hb949ee6c),
	.w6(32'hbaca49b9),
	.w7(32'h39944f06),
	.w8(32'hba4cb750),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae6a8a),
	.w1(32'hba3d912f),
	.w2(32'hbba14efc),
	.w3(32'hbbd2b8d7),
	.w4(32'h3a415b25),
	.w5(32'hbb006276),
	.w6(32'hbbe19919),
	.w7(32'hbabe39ad),
	.w8(32'hbb8b06a1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38896e08),
	.w1(32'hb69a3e1b),
	.w2(32'h382429e0),
	.w3(32'h382f61b6),
	.w4(32'hb7a622d1),
	.w5(32'h37bcdac7),
	.w6(32'h388e4707),
	.w7(32'h37cf0b19),
	.w8(32'h38887559),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ae50de),
	.w1(32'h3890245f),
	.w2(32'h38d66815),
	.w3(32'h379a4334),
	.w4(32'h37d96106),
	.w5(32'h388cd35c),
	.w6(32'h39118db7),
	.w7(32'h38f484b6),
	.w8(32'h38cd01eb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd5c08),
	.w1(32'h3a8f832f),
	.w2(32'h39bd52d4),
	.w3(32'hb98ce147),
	.w4(32'h3b0ad870),
	.w5(32'h3aac91f6),
	.w6(32'hbaa60f61),
	.w7(32'h3accb47c),
	.w8(32'h39a037e2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ab25),
	.w1(32'hba6b719f),
	.w2(32'hbba6d6ca),
	.w3(32'hbb3eace1),
	.w4(32'h39ca21a9),
	.w5(32'hbb42f9b8),
	.w6(32'hbb8a0735),
	.w7(32'hbb1bb3e6),
	.w8(32'hbba1c3ac),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c5c03),
	.w1(32'h38041d93),
	.w2(32'hbab18f1b),
	.w3(32'hbb1f79e2),
	.w4(32'hb8b98f49),
	.w5(32'hba9b5b07),
	.w6(32'h3a9b916d),
	.w7(32'h3b14d405),
	.w8(32'hba934c18),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33b7b4),
	.w1(32'h39259d8f),
	.w2(32'hba5fbc37),
	.w3(32'hba6562e2),
	.w4(32'h3754d56c),
	.w5(32'hba2a62d2),
	.w6(32'hbaa827e5),
	.w7(32'hb98c658f),
	.w8(32'hba6d8da0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88d3aa),
	.w1(32'hbb89c1a7),
	.w2(32'hbc8bd4ab),
	.w3(32'hbc117a44),
	.w4(32'h39b8bbbf),
	.w5(32'hbc62354a),
	.w6(32'hbb9dd208),
	.w7(32'h3a0f7a3b),
	.w8(32'hbbd1be0d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc414362),
	.w1(32'h3b116576),
	.w2(32'hbb8fe171),
	.w3(32'hbc218cd5),
	.w4(32'h3bd28f7e),
	.w5(32'h3b19fa8e),
	.w6(32'hbc1e14ef),
	.w7(32'h3bc3a0b5),
	.w8(32'hba8082b6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4829b7),
	.w1(32'hba064471),
	.w2(32'hba1e7f53),
	.w3(32'hb96f785e),
	.w4(32'hbac232c8),
	.w5(32'hbaaee0e4),
	.w6(32'h3a02391a),
	.w7(32'hba2b705f),
	.w8(32'hba854622),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37945bf5),
	.w1(32'hb78f8420),
	.w2(32'hb71d0018),
	.w3(32'hb88f81e2),
	.w4(32'hb86c79f5),
	.w5(32'hb8041e62),
	.w6(32'hb72ad2f0),
	.w7(32'h37ac3bb8),
	.w8(32'h37e87116),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38532ba0),
	.w1(32'h38b8ad85),
	.w2(32'h38c56719),
	.w3(32'h388c8d45),
	.w4(32'h37faaf79),
	.w5(32'h377b19d0),
	.w6(32'h3902e83f),
	.w7(32'h3804240f),
	.w8(32'h382cdcfd),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8e97d),
	.w1(32'h373220f5),
	.w2(32'h38a06ff0),
	.w3(32'h38ae928d),
	.w4(32'hb77cb349),
	.w5(32'h3865824c),
	.w6(32'h38ff8105),
	.w7(32'h382021b2),
	.w8(32'h38eaf295),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398162d0),
	.w1(32'hbafd14ee),
	.w2(32'hbb53d078),
	.w3(32'hb9a190c3),
	.w4(32'hbb18d706),
	.w5(32'hbb29f72b),
	.w6(32'h392f2bcb),
	.w7(32'hbb059f72),
	.w8(32'hbb64c52e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb64d2),
	.w1(32'hbaeaf7be),
	.w2(32'hbb0ef590),
	.w3(32'hbb86a752),
	.w4(32'h39ff1cc2),
	.w5(32'hbb1f136b),
	.w6(32'hbb94fc45),
	.w7(32'hbb1fb100),
	.w8(32'hbc076e39),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bf0a6),
	.w1(32'hba1c6b3a),
	.w2(32'hbb903474),
	.w3(32'hbb843c95),
	.w4(32'h3b9c8118),
	.w5(32'hba01b20c),
	.w6(32'hbbe89022),
	.w7(32'h3b0d652b),
	.w8(32'hbb45ad22),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57847a),
	.w1(32'h3abf0414),
	.w2(32'h3a176c9a),
	.w3(32'hb9bfa4a4),
	.w4(32'h3ad092f5),
	.w5(32'h3a10d810),
	.w6(32'hbad83e91),
	.w7(32'hba23cafe),
	.w8(32'hbb0002ea),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe12933),
	.w1(32'hbb983d86),
	.w2(32'hbc2e36ab),
	.w3(32'hbb7a3590),
	.w4(32'hba90c6eb),
	.w5(32'hbbf8a03c),
	.w6(32'hbbb0a66c),
	.w7(32'hbb455089),
	.w8(32'hbc0b8158),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb021fd2),
	.w1(32'hba39c12e),
	.w2(32'hbb041bd2),
	.w3(32'hbb0aec45),
	.w4(32'hbaaa2a03),
	.w5(32'hbb202d27),
	.w6(32'hbb13274a),
	.w7(32'hbaa34623),
	.w8(32'hbac9b5de),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934b46e),
	.w1(32'h386fe0eb),
	.w2(32'h393a3d9d),
	.w3(32'h391b5bde),
	.w4(32'h38284ab8),
	.w5(32'h3923c2d2),
	.w6(32'h395ec1e6),
	.w7(32'h38ed4794),
	.w8(32'h396e6adb),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8655b0),
	.w1(32'hba45047f),
	.w2(32'hba0359fe),
	.w3(32'hba271192),
	.w4(32'hb845b180),
	.w5(32'h3a1dd228),
	.w6(32'hba05bb52),
	.w7(32'h3987ee70),
	.w8(32'h3a8bbf86),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af32c4),
	.w1(32'h3892da8e),
	.w2(32'h39b71d5e),
	.w3(32'h399e4f47),
	.w4(32'h37a9139f),
	.w5(32'h399ad32e),
	.w6(32'h39f9ec30),
	.w7(32'h395de034),
	.w8(32'h39fe5d77),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb858025),
	.w1(32'h3a376ba2),
	.w2(32'hbb0f0e53),
	.w3(32'hbb0fcf72),
	.w4(32'h3b321e2b),
	.w5(32'hb9deab07),
	.w6(32'hbb894bb5),
	.w7(32'h38b90b83),
	.w8(32'hbba22a47),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb32eee),
	.w1(32'h3bd9eb9b),
	.w2(32'h389e2330),
	.w3(32'hbb50794d),
	.w4(32'h3c17ed99),
	.w5(32'h3b3b7972),
	.w6(32'hbc199dbb),
	.w7(32'h3b9aab70),
	.w8(32'hbb41a8a3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabdcd7),
	.w1(32'h39a3b695),
	.w2(32'hbb8992fc),
	.w3(32'hbb2f7d80),
	.w4(32'h3b476859),
	.w5(32'hbaece094),
	.w6(32'hbbb642d8),
	.w7(32'hb7f7bf46),
	.w8(32'hbbbd6a68),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904067d),
	.w1(32'h3acd0bfc),
	.w2(32'hb93398b3),
	.w3(32'hba027662),
	.w4(32'h3a619650),
	.w5(32'hba023974),
	.w6(32'hbae3f6fb),
	.w7(32'h39084bec),
	.w8(32'hba95f73e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4919f),
	.w1(32'h3acc5b31),
	.w2(32'hbb473fee),
	.w3(32'hbb2fcd0f),
	.w4(32'h3bac4423),
	.w5(32'h39879f0a),
	.w6(32'hbbcc4527),
	.w7(32'h3aa80989),
	.w8(32'hbbaaa8c8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb642528),
	.w1(32'h3811f05a),
	.w2(32'hbb38ff86),
	.w3(32'hbb3f7237),
	.w4(32'h3a0e2d28),
	.w5(32'hbad8d6ea),
	.w6(32'hbb4b181b),
	.w7(32'hba58e3b9),
	.w8(32'hbb160fdc),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc185ca3),
	.w1(32'h3acaf2f4),
	.w2(32'hbbb8193a),
	.w3(32'hbbfc699c),
	.w4(32'h3ba79565),
	.w5(32'hbb7dc35f),
	.w6(32'hbc01e996),
	.w7(32'h3aa1980a),
	.w8(32'hbbbdabb4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389aa327),
	.w1(32'hb74d03a1),
	.w2(32'h386db450),
	.w3(32'h388ad9fa),
	.w4(32'hb75bc07d),
	.w5(32'h38593bcc),
	.w6(32'h39131243),
	.w7(32'h38827f29),
	.w8(32'h3910fab3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914f9ff),
	.w1(32'h3904e5ba),
	.w2(32'h38ceaca4),
	.w3(32'hb8349eae),
	.w4(32'hb8d0c94f),
	.w5(32'hb94eb7ed),
	.w6(32'h37480864),
	.w7(32'h391c8ae1),
	.w8(32'h38a49bea),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcafe52),
	.w1(32'h3aa37dfb),
	.w2(32'hbb9d04ac),
	.w3(32'hbb933053),
	.w4(32'h3a104b2c),
	.w5(32'hbbb5ef44),
	.w6(32'hbbe6fe86),
	.w7(32'hba4faff3),
	.w8(32'hbbf54f3f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4556a),
	.w1(32'h3a9a2652),
	.w2(32'hbbc0dcb5),
	.w3(32'hbb821d09),
	.w4(32'h3a9207b4),
	.w5(32'hbc1520ec),
	.w6(32'hbbbcf637),
	.w7(32'hba6370e0),
	.w8(32'hbc11c6da),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb194d),
	.w1(32'h3a4c6fa0),
	.w2(32'hbb937b6e),
	.w3(32'hbb3defa3),
	.w4(32'h3b93fb20),
	.w5(32'hbaac32c9),
	.w6(32'hbbd50b52),
	.w7(32'h3a9de059),
	.w8(32'hbb97170d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72b702),
	.w1(32'hba8b50f8),
	.w2(32'hba8d695e),
	.w3(32'hbb9ca8d6),
	.w4(32'hbbb6ce1e),
	.w5(32'hbb26e7ef),
	.w6(32'h3b124f85),
	.w7(32'hba0b8b40),
	.w8(32'hba874d4b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb973b35f),
	.w1(32'hb981e6b8),
	.w2(32'hb90d7003),
	.w3(32'hb8ea13bb),
	.w4(32'hb949ce93),
	.w5(32'hb75d82aa),
	.w6(32'hb792f349),
	.w7(32'hb94357d6),
	.w8(32'h39010053),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8358e4),
	.w1(32'hb9b54f8e),
	.w2(32'h3956d55d),
	.w3(32'hba3c6232),
	.w4(32'hb9f64184),
	.w5(32'hb87da242),
	.w6(32'hba0a473e),
	.w7(32'hb965d031),
	.w8(32'h3930c590),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd4518),
	.w1(32'hbad5f87c),
	.w2(32'hbbe811bb),
	.w3(32'hbb49f151),
	.w4(32'hbbeb1b10),
	.w5(32'hbc1f7b08),
	.w6(32'h3ab9af79),
	.w7(32'hbb104f17),
	.w8(32'hbbd91aab),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc634c36),
	.w1(32'hbba9f658),
	.w2(32'hbc0ef23d),
	.w3(32'hbc1591b7),
	.w4(32'hbb3662ca),
	.w5(32'hbc1a5dd0),
	.w6(32'hbbe70663),
	.w7(32'hbb0ffb99),
	.w8(32'hbbe35ceb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e9430),
	.w1(32'hbb7e282f),
	.w2(32'hbb60c723),
	.w3(32'hbbd5d4a8),
	.w4(32'hbbbc13e1),
	.w5(32'hbb96da1e),
	.w6(32'hbb57ce46),
	.w7(32'hbb79f755),
	.w8(32'hbbae7770),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99cc26),
	.w1(32'h3be67751),
	.w2(32'h3ae42aad),
	.w3(32'hbb1c2f79),
	.w4(32'h3bcce336),
	.w5(32'h3abb4410),
	.w6(32'hbbae0e54),
	.w7(32'h3b697e21),
	.w8(32'hbae7d12b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f4110),
	.w1(32'h3b12a09d),
	.w2(32'hbb6ed893),
	.w3(32'hbb34bfca),
	.w4(32'h3bd3e281),
	.w5(32'h3a720c51),
	.w6(32'hbbb00c5d),
	.w7(32'h3b7cc620),
	.w8(32'hbb1956e3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b8bcd2),
	.w1(32'h381f066a),
	.w2(32'h38869508),
	.w3(32'h38a57f70),
	.w4(32'h380db2cd),
	.w5(32'h38662bbd),
	.w6(32'h38cb9eb4),
	.w7(32'h38808e72),
	.w8(32'h38b53838),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f1ae3a),
	.w1(32'h3858bd89),
	.w2(32'h38c002dc),
	.w3(32'h38e73398),
	.w4(32'h383a8ee4),
	.w5(32'h38b8f16f),
	.w6(32'h391b34c0),
	.w7(32'h38bc07d0),
	.w8(32'h390c1080),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6290f2),
	.w1(32'h39bc97e1),
	.w2(32'h3a062463),
	.w3(32'h37ccefd1),
	.w4(32'hba4578ad),
	.w5(32'hba2cd8ec),
	.w6(32'h38d3d943),
	.w7(32'hba31a030),
	.w8(32'hb90704d8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e25808),
	.w1(32'hb7fdeac7),
	.w2(32'h38757681),
	.w3(32'h38daa044),
	.w4(32'hb7f8f8a9),
	.w5(32'h3839aa61),
	.w6(32'h392d6012),
	.w7(32'h37b44854),
	.w8(32'h38f894a4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba6c5c),
	.w1(32'hbafe7935),
	.w2(32'hbb117929),
	.w3(32'hba5b95fd),
	.w4(32'hbafac177),
	.w5(32'hbb16a326),
	.w6(32'hba03fb40),
	.w7(32'hbaa2184d),
	.w8(32'hbadbe910),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc804b4),
	.w1(32'hbaf21490),
	.w2(32'hbbaf9e51),
	.w3(32'hbae52a77),
	.w4(32'h3a317cb7),
	.w5(32'hbb90675b),
	.w6(32'hbaeae578),
	.w7(32'hba1a7af2),
	.w8(32'hbbb8d229),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94fd82),
	.w1(32'hb6d4ce33),
	.w2(32'hbb20a05e),
	.w3(32'hbb835dea),
	.w4(32'h3a248e20),
	.w5(32'hbadfa826),
	.w6(32'hbb9e14ab),
	.w7(32'hbb0718d1),
	.w8(32'hbbae387f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6d479),
	.w1(32'h389b3e45),
	.w2(32'h38ea8bc2),
	.w3(32'h3909fbeb),
	.w4(32'h38de9123),
	.w5(32'h39193bcd),
	.w6(32'h391257bc),
	.w7(32'h392d7a82),
	.w8(32'h392cf525),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb889b22),
	.w1(32'hbb6154e9),
	.w2(32'hbc0bc47d),
	.w3(32'hbb9b2a1d),
	.w4(32'hbba2570a),
	.w5(32'hbc1a0a24),
	.w6(32'hb9e07dc9),
	.w7(32'hba91e7f3),
	.w8(32'hbc134e1e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62c017),
	.w1(32'hbac40004),
	.w2(32'hbb19d963),
	.w3(32'hbb1d268d),
	.w4(32'hbabfa4bc),
	.w5(32'hbb29705d),
	.w6(32'hbae723fe),
	.w7(32'hbac0c260),
	.w8(32'hbb164358),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37df521f),
	.w1(32'hb9454198),
	.w2(32'h397e8c88),
	.w3(32'hb9549df8),
	.w4(32'hb9b13265),
	.w5(32'h38dceaba),
	.w6(32'hb829a1d3),
	.w7(32'hb8a17384),
	.w8(32'hb8cb1f4c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf0ac6),
	.w1(32'hba9ef133),
	.w2(32'hbb453aa1),
	.w3(32'hbb07ad31),
	.w4(32'hbad30bd3),
	.w5(32'hbb3c2ac9),
	.w6(32'hbaa82405),
	.w7(32'hbadf23e8),
	.w8(32'hbb28ff4a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ed525),
	.w1(32'h391d9711),
	.w2(32'h395b2589),
	.w3(32'h3920771b),
	.w4(32'h390bc580),
	.w5(32'h3963d008),
	.w6(32'h390c7191),
	.w7(32'h38e51df6),
	.w8(32'h39530d4d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9768212),
	.w1(32'hb850a680),
	.w2(32'hb80c0221),
	.w3(32'hb87bebe3),
	.w4(32'h3986aa57),
	.w5(32'h394aed61),
	.w6(32'hba0abfcf),
	.w7(32'hb9c74f67),
	.w8(32'hba0c233c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b7964),
	.w1(32'h38fabfb4),
	.w2(32'h391720a0),
	.w3(32'h3912bf01),
	.w4(32'h38b29b17),
	.w5(32'h38d618af),
	.w6(32'h391a9888),
	.w7(32'h388e65a0),
	.w8(32'h38d3d9fa),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f77de0),
	.w1(32'h3893d70d),
	.w2(32'h38c6369c),
	.w3(32'h38a8ba82),
	.w4(32'h3811ea3f),
	.w5(32'h387339db),
	.w6(32'h38e8ae15),
	.w7(32'h38a4461a),
	.w8(32'h38c6c235),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13a499),
	.w1(32'h3b1687c3),
	.w2(32'h393c9eb0),
	.w3(32'hba7d13a9),
	.w4(32'h3af26959),
	.w5(32'hba42eaaf),
	.w6(32'hbb7c1ff1),
	.w7(32'h3a10751c),
	.w8(32'hba812847),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9928f),
	.w1(32'hbb1ceac9),
	.w2(32'hbc12ae46),
	.w3(32'hbb9d8485),
	.w4(32'hbacd0c5a),
	.w5(32'hbbe8b862),
	.w6(32'hbb9302ed),
	.w7(32'hbb34d349),
	.w8(32'hbbffcc9d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94fdc8),
	.w1(32'hbaa61a62),
	.w2(32'hbba372ee),
	.w3(32'hbadd704f),
	.w4(32'hba15add9),
	.w5(32'hbb92c00a),
	.w6(32'hba2dc8db),
	.w7(32'hb880b4f0),
	.w8(32'hbb4b6c5e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba338ec),
	.w1(32'hbb3edbd3),
	.w2(32'hbbc984af),
	.w3(32'hbbc12068),
	.w4(32'hbb431cf1),
	.w5(32'hbbac1b11),
	.w6(32'hbb8d00c8),
	.w7(32'hbb85d9dc),
	.w8(32'hbbb3f696),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39496ea5),
	.w1(32'h39a01bb2),
	.w2(32'h38d10482),
	.w3(32'h382339e1),
	.w4(32'h39987071),
	.w5(32'h3950f037),
	.w6(32'hb97734ad),
	.w7(32'h38309ca0),
	.w8(32'hb7018769),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6288e),
	.w1(32'hba006f05),
	.w2(32'hb92dddf4),
	.w3(32'hb942acab),
	.w4(32'hb9b6b823),
	.w5(32'h365ec426),
	.w6(32'hb8cf39ab),
	.w7(32'hb99dd418),
	.w8(32'hb888c89a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3820d861),
	.w1(32'hb7b2e07e),
	.w2(32'h38051a0a),
	.w3(32'h37b881bf),
	.w4(32'hb827dc76),
	.w5(32'h37a5f3c5),
	.w6(32'h384aa592),
	.w7(32'hb6e6d2da),
	.w8(32'h38668acc),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a97671),
	.w1(32'h38827340),
	.w2(32'h3874a578),
	.w3(32'h38b655de),
	.w4(32'hb5422496),
	.w5(32'h37546911),
	.w6(32'h38f74645),
	.w7(32'h377de1c7),
	.w8(32'h37819232),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc297b40),
	.w1(32'hbb84fbc6),
	.w2(32'hbbc94a36),
	.w3(32'hbbae71fd),
	.w4(32'hbae3a704),
	.w5(32'hbb4f5788),
	.w6(32'hbbaea745),
	.w7(32'hbaf75f18),
	.w8(32'hbb8e67a4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d4d0e9),
	.w1(32'hb875ce1f),
	.w2(32'h388fabcd),
	.w3(32'hb79cc508),
	.w4(32'hb8ea8191),
	.w5(32'hb7501ae5),
	.w6(32'h37d0887e),
	.w7(32'hb87a5352),
	.w8(32'h37f10524),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f82aa2),
	.w1(32'h3b10d848),
	.w2(32'hbaa0c7c6),
	.w3(32'hb81f9575),
	.w4(32'h3ae88cd6),
	.w5(32'hba75cf9d),
	.w6(32'hbae081db),
	.w7(32'h3a0c4281),
	.w8(32'hbaf8bab6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5c5be),
	.w1(32'h39462cb4),
	.w2(32'hba64c2f9),
	.w3(32'hbae532b4),
	.w4(32'h39915e41),
	.w5(32'hb9b33a8b),
	.w6(32'hbaa7330b),
	.w7(32'h3a3986d9),
	.w8(32'h39487f03),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388d9a57),
	.w1(32'h38042a8c),
	.w2(32'h37b96e08),
	.w3(32'h386ea250),
	.w4(32'h37ce6692),
	.w5(32'h37b78161),
	.w6(32'h38c9380f),
	.w7(32'h3843527b),
	.w8(32'h3821f3df),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf63ae),
	.w1(32'hba2e3595),
	.w2(32'hba365cd9),
	.w3(32'hba8a9e1e),
	.w4(32'h38ae39c2),
	.w5(32'hba388fbd),
	.w6(32'hba54ac2f),
	.w7(32'hba79676d),
	.w8(32'hbae48362),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f5ee6),
	.w1(32'hb94d998e),
	.w2(32'hb80fe8ce),
	.w3(32'h378a1e25),
	.w4(32'hb58af1c9),
	.w5(32'h391846f2),
	.w6(32'hb7b5223f),
	.w7(32'hb857dadd),
	.w8(32'hb87bb23b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfce7c3),
	.w1(32'hbb86ed74),
	.w2(32'hbc0fe7b0),
	.w3(32'hbbd5d4d2),
	.w4(32'hb9f64a06),
	.w5(32'hba82cd50),
	.w6(32'hbbeb8802),
	.w7(32'hbb53ee16),
	.w8(32'hbb7f6259),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a29988),
	.w1(32'hbb009207),
	.w2(32'h3af70f0c),
	.w3(32'h372f81d9),
	.w4(32'hba21d52f),
	.w5(32'h3b1ea002),
	.w6(32'hbaae6011),
	.w7(32'h39acccd8),
	.w8(32'hb91bd53a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50cbc9),
	.w1(32'h3c32e783),
	.w2(32'h3be76ac5),
	.w3(32'h3a33b011),
	.w4(32'h3ba97f73),
	.w5(32'h3b690ad3),
	.w6(32'hbc07e7d8),
	.w7(32'h3a821055),
	.w8(32'h3b06a479),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule