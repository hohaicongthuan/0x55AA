module layer_8_featuremap_165(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47f23c),
	.w1(32'h3c1cf32b),
	.w2(32'h3c5d3d68),
	.w3(32'h3ac3fc88),
	.w4(32'h398d1ed1),
	.w5(32'hb93a41de),
	.w6(32'h3c124ac9),
	.w7(32'hbbcfa5d1),
	.w8(32'hbc04e0d4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3781c6),
	.w1(32'hb9fe347e),
	.w2(32'hbba5bd32),
	.w3(32'hbab72a95),
	.w4(32'hbae90029),
	.w5(32'hbbbcdaaa),
	.w6(32'h3a1983e5),
	.w7(32'hbb5efc27),
	.w8(32'hba6e3860),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa11593),
	.w1(32'h3bd7bf6e),
	.w2(32'h3c649341),
	.w3(32'h3a2a2465),
	.w4(32'h3bb5f020),
	.w5(32'h3b95b484),
	.w6(32'h3c40bd88),
	.w7(32'h3c188a26),
	.w8(32'h3c535a2b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ce2f5),
	.w1(32'h3c15a499),
	.w2(32'h3bc53d1f),
	.w3(32'h3bbfe909),
	.w4(32'h3c2611c2),
	.w5(32'h3aac9a1a),
	.w6(32'h3bc8f11e),
	.w7(32'h3becae25),
	.w8(32'h3bb84bef),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b91ea4),
	.w1(32'h3bc8d6e3),
	.w2(32'h3acbd4ee),
	.w3(32'hbbe6f119),
	.w4(32'h3aaba7bd),
	.w5(32'h3af6cd39),
	.w6(32'h3b6edc08),
	.w7(32'h3a85eebf),
	.w8(32'h3b8a3cf5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1b22b),
	.w1(32'hbab9c809),
	.w2(32'hbcfaea96),
	.w3(32'h3b9ecff1),
	.w4(32'hbc224eea),
	.w5(32'hbc9cd976),
	.w6(32'h3b7e5741),
	.w7(32'hbc618e11),
	.w8(32'hbca57fb7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd054801),
	.w1(32'hbb1d335c),
	.w2(32'h3a03c70e),
	.w3(32'hbc85167c),
	.w4(32'hb9a2622a),
	.w5(32'h3ac7c3c4),
	.w6(32'hbbbfa4e7),
	.w7(32'hba85bccb),
	.w8(32'hba29ca66),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5aa18),
	.w1(32'hbc78bbbb),
	.w2(32'hbb01d984),
	.w3(32'hbb920c06),
	.w4(32'hbc372f94),
	.w5(32'hbb1d5e7b),
	.w6(32'h3b5a386a),
	.w7(32'hbbea4950),
	.w8(32'h3b457a0e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00e067),
	.w1(32'h3a015fac),
	.w2(32'h3a46487a),
	.w3(32'h3c29dc95),
	.w4(32'hbbab3312),
	.w5(32'h3a56d69f),
	.w6(32'hbc681195),
	.w7(32'hbb9c014c),
	.w8(32'hbb9e3135),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917ce5f),
	.w1(32'h3b41f562),
	.w2(32'h3a463899),
	.w3(32'h3b1dbd5f),
	.w4(32'hba77e956),
	.w5(32'hbbb421df),
	.w6(32'hb9c6a587),
	.w7(32'h3b898cb8),
	.w8(32'h3a9a8dec),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadfc17),
	.w1(32'hba7cc422),
	.w2(32'hbb953309),
	.w3(32'hbc361107),
	.w4(32'h3ab29ea9),
	.w5(32'hbb96ba7c),
	.w6(32'hbbbf72ce),
	.w7(32'hbca4d8b6),
	.w8(32'hbc4bdca3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8571ad),
	.w1(32'h3bf93c6b),
	.w2(32'h3c2c88b5),
	.w3(32'hbbc47603),
	.w4(32'h3ba07aa9),
	.w5(32'h3bd36f91),
	.w6(32'h3b91b091),
	.w7(32'h3b1783f8),
	.w8(32'h3b997f94),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c010bdc),
	.w1(32'hbc760820),
	.w2(32'hbc8f7d64),
	.w3(32'h3bd8c041),
	.w4(32'hbba00344),
	.w5(32'hbc8dee25),
	.w6(32'hbc4d9d22),
	.w7(32'hbc62109a),
	.w8(32'hbc1cf3a4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dceeb),
	.w1(32'h395c512c),
	.w2(32'hb9af1cb6),
	.w3(32'hbcbfab2a),
	.w4(32'hb90772de),
	.w5(32'h3afc16bf),
	.w6(32'hbc1434f7),
	.w7(32'hbb5940be),
	.w8(32'hbb837490),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12e9e9),
	.w1(32'hbbe8964f),
	.w2(32'h3aeeebe7),
	.w3(32'h3bb589ac),
	.w4(32'hbb64963c),
	.w5(32'h3b4bb85c),
	.w6(32'hbc38e085),
	.w7(32'hbaa75afb),
	.w8(32'hba9ad7a0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6cb4d),
	.w1(32'h3c3ac19c),
	.w2(32'h3bced58e),
	.w3(32'hb89f8f67),
	.w4(32'h3bf9f6ea),
	.w5(32'hbb09c869),
	.w6(32'h3ba5e9aa),
	.w7(32'hba42f999),
	.w8(32'hbbad11b0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc394d6),
	.w1(32'hbc23122a),
	.w2(32'hbcbdb46e),
	.w3(32'hbbcfdcca),
	.w4(32'hbc31e4c1),
	.w5(32'hbc8a6b74),
	.w6(32'hbc8723d6),
	.w7(32'hbc9e421d),
	.w8(32'hbc80daaa),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0ee23),
	.w1(32'h3ce5b649),
	.w2(32'h3cd9a8f0),
	.w3(32'hbca1c13d),
	.w4(32'h3c750507),
	.w5(32'h3c61952a),
	.w6(32'h3cc9438d),
	.w7(32'h3ccda9c6),
	.w8(32'h3c847348),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfd5005),
	.w1(32'hba0fa4d1),
	.w2(32'hbc3a8ab1),
	.w3(32'h3c2ccd12),
	.w4(32'hbb288149),
	.w5(32'hbc0d23cc),
	.w6(32'h3c42278b),
	.w7(32'hba206e65),
	.w8(32'h395d1733),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02d809),
	.w1(32'hbb57335d),
	.w2(32'h3b698588),
	.w3(32'hbc108d57),
	.w4(32'hbaed2e38),
	.w5(32'h3b05519a),
	.w6(32'hbbf00510),
	.w7(32'h3a77f71b),
	.w8(32'hbac59299),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390718e9),
	.w1(32'h3c3bd979),
	.w2(32'h3caed1ce),
	.w3(32'hbb254ab3),
	.w4(32'h3b90eefb),
	.w5(32'h3bf1f803),
	.w6(32'h3b166a3f),
	.w7(32'h3c84534c),
	.w8(32'h3ba318af),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5551bb),
	.w1(32'hbd2dce7e),
	.w2(32'hbd8257a5),
	.w3(32'h3c06255a),
	.w4(32'hbd10dbc2),
	.w5(32'hbd1f27b9),
	.w6(32'hbc4bd475),
	.w7(32'hbd419d1a),
	.w8(32'hbd02a117),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd259702),
	.w1(32'hbbc216b9),
	.w2(32'h3c07ef6e),
	.w3(32'hbc78dbde),
	.w4(32'hba20a08e),
	.w5(32'h3c5e028c),
	.w6(32'hbc4eac9f),
	.w7(32'hbc226e63),
	.w8(32'hbab3f67c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93be53),
	.w1(32'hbd1d18f4),
	.w2(32'hbd7080b4),
	.w3(32'h3ca3d907),
	.w4(32'hbcc1088d),
	.w5(32'hbd1653f7),
	.w6(32'hbc8ac266),
	.w7(32'hbd03e360),
	.w8(32'hbd12a68a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a68f0),
	.w1(32'hb9711d80),
	.w2(32'h3aec1674),
	.w3(32'hbccb1d86),
	.w4(32'hbb90b083),
	.w5(32'hbb78193b),
	.w6(32'h3b63944a),
	.w7(32'h3bcc8011),
	.w8(32'h3bae02dd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c246e),
	.w1(32'h3b8ee17a),
	.w2(32'h3c1897ee),
	.w3(32'hbbb3fb41),
	.w4(32'hbbd06614),
	.w5(32'hb92cdff1),
	.w6(32'hb96133ab),
	.w7(32'h3baf2ce8),
	.w8(32'h3c07f606),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58b797),
	.w1(32'h3c35edb4),
	.w2(32'h3bc508c7),
	.w3(32'hbb503332),
	.w4(32'h3a362b76),
	.w5(32'hb9075625),
	.w6(32'h3c485fa6),
	.w7(32'h3c3cc3cd),
	.w8(32'hbb9818b0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f8321),
	.w1(32'h3c54bc75),
	.w2(32'h3c491515),
	.w3(32'h3bf76b17),
	.w4(32'h3c242f00),
	.w5(32'h3b339a8d),
	.w6(32'h3b803472),
	.w7(32'h3b8d3d17),
	.w8(32'h3b6ac107),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23ccde),
	.w1(32'h39a4f296),
	.w2(32'h3c0f85de),
	.w3(32'h3a61ce89),
	.w4(32'hb8511a82),
	.w5(32'h3c1e922f),
	.w6(32'hbc1206c5),
	.w7(32'hbb21e41d),
	.w8(32'hbb591e9a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbadf08),
	.w1(32'hba1e3a3a),
	.w2(32'hbb0dea32),
	.w3(32'h3b4e5c78),
	.w4(32'h3b9c74f3),
	.w5(32'h3bd8d298),
	.w6(32'hb924bab5),
	.w7(32'h3a704fbe),
	.w8(32'hbbe89683),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fc46b),
	.w1(32'hbb34bdf0),
	.w2(32'h3c1da4f5),
	.w3(32'h3baa9307),
	.w4(32'h3ba6cb2e),
	.w5(32'hbb4603c4),
	.w6(32'h3b6544e6),
	.w7(32'h3c03ea99),
	.w8(32'h3bc219d3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b4ae8),
	.w1(32'hbc6249f1),
	.w2(32'hba921c39),
	.w3(32'hbb8e2a67),
	.w4(32'hbbb09248),
	.w5(32'hbaa37c42),
	.w6(32'hbba41aa9),
	.w7(32'hbbbff2ca),
	.w8(32'h3b837103),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c228582),
	.w1(32'h3c5d450d),
	.w2(32'h3c6821c9),
	.w3(32'h3c249e22),
	.w4(32'h3b8c8fca),
	.w5(32'h3b671671),
	.w6(32'h3b776b51),
	.w7(32'h3c611344),
	.w8(32'h3c8faecb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e8016),
	.w1(32'h3cbf4e27),
	.w2(32'h3d1d7e6a),
	.w3(32'h3b27b4d3),
	.w4(32'h3bf116a3),
	.w5(32'h3c6c57ff),
	.w6(32'h3c3cf5c7),
	.w7(32'h3ca954a3),
	.w8(32'hbb915583),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca73167),
	.w1(32'h3ab643bb),
	.w2(32'h3bc1aee0),
	.w3(32'h3b9597f4),
	.w4(32'hba5f2ed4),
	.w5(32'hba9a66c3),
	.w6(32'h3b45560b),
	.w7(32'h3b8e07b6),
	.w8(32'h3c172592),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b466479),
	.w1(32'h3cb93fd4),
	.w2(32'h3d184347),
	.w3(32'h3bc6329b),
	.w4(32'h3ca4b9ed),
	.w5(32'h3ca7beb3),
	.w6(32'h3cbeccf5),
	.w7(32'h3cb15731),
	.w8(32'h3c7bb36c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01abf1),
	.w1(32'hbbee2317),
	.w2(32'hbc08a018),
	.w3(32'h3c80449d),
	.w4(32'hbc0f986f),
	.w5(32'hbc027ca8),
	.w6(32'hbbfde792),
	.w7(32'hbbe9ae83),
	.w8(32'hbc10f17f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc040d82),
	.w1(32'hbbef8445),
	.w2(32'hba6f3f9d),
	.w3(32'hbba872a9),
	.w4(32'hbb4e8139),
	.w5(32'h3aabcd63),
	.w6(32'hbc3b2c5a),
	.w7(32'hbbbe06b1),
	.w8(32'hbb62f777),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b332e68),
	.w1(32'hbd3e1ff9),
	.w2(32'hbd9e3d9d),
	.w3(32'h3b65023a),
	.w4(32'hbc92aa9a),
	.w5(32'hbd1bc10b),
	.w6(32'hbd11f4d3),
	.w7(32'hbd3efe45),
	.w8(32'hbcdf3893),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd02756f),
	.w1(32'hbcdb6260),
	.w2(32'hbd53dec0),
	.w3(32'hbc8b269a),
	.w4(32'hbc9a7fc1),
	.w5(32'hbd19a996),
	.w6(32'hbcaa6ad0),
	.w7(32'hbced4171),
	.w8(32'hbcbab3d5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd269cc5),
	.w1(32'hbb205f3b),
	.w2(32'h3b6e2d11),
	.w3(32'hbccee504),
	.w4(32'h38e77765),
	.w5(32'h3bb44a22),
	.w6(32'hb7dfd643),
	.w7(32'h3bcbe5a7),
	.w8(32'h3a9c00fc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e34f5a),
	.w1(32'hba040c42),
	.w2(32'hbb0a1043),
	.w3(32'h3b88c9b2),
	.w4(32'h3b0c78e0),
	.w5(32'hbad9428e),
	.w6(32'hbbcd76c7),
	.w7(32'hb9b2169e),
	.w8(32'hba46cdc6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b1cdee),
	.w1(32'h3a299d8b),
	.w2(32'h3b3c7116),
	.w3(32'h3b3fe8a4),
	.w4(32'hbbbecefb),
	.w5(32'h3b269e90),
	.w6(32'hb8ccd07b),
	.w7(32'hb9f5c2e4),
	.w8(32'hbaba3aff),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0bd8b),
	.w1(32'h3a856f89),
	.w2(32'h3b7bb9b2),
	.w3(32'h3c22a629),
	.w4(32'h3c1d7b06),
	.w5(32'h3bb8e355),
	.w6(32'h3c1a9243),
	.w7(32'h3c0d5369),
	.w8(32'h3c267094),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fd53e),
	.w1(32'h3c92998e),
	.w2(32'h3c875573),
	.w3(32'h3c825840),
	.w4(32'h3c013513),
	.w5(32'h3bc40afe),
	.w6(32'hbaa63b17),
	.w7(32'h3c114241),
	.w8(32'hba02c3e8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b431d76),
	.w1(32'h3b1fb494),
	.w2(32'hbafff62b),
	.w3(32'h3b0124d5),
	.w4(32'h3b908fd3),
	.w5(32'hbb1f9095),
	.w6(32'hbb0f14b7),
	.w7(32'hbac1114e),
	.w8(32'hbaf4d33b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb505975),
	.w1(32'h3bcfac63),
	.w2(32'h3c15d8a9),
	.w3(32'hbaedc68b),
	.w4(32'hbb5eb0d8),
	.w5(32'h3ba0a61c),
	.w6(32'h3bc5a700),
	.w7(32'h3c65346c),
	.w8(32'h3bc13ca3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c275fc3),
	.w1(32'hbb69f8ef),
	.w2(32'hbce1e3ac),
	.w3(32'h3ace5b9f),
	.w4(32'h3b8457fc),
	.w5(32'hbbb30d34),
	.w6(32'h3b1384a4),
	.w7(32'hbc477df6),
	.w8(32'hbc09eb10),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd36fea),
	.w1(32'hbc18064f),
	.w2(32'hbbf1ab67),
	.w3(32'h39e638de),
	.w4(32'hbb8f8259),
	.w5(32'h3bad3572),
	.w6(32'h3b255fbc),
	.w7(32'h3bdd5b8f),
	.w8(32'h3ba0fdcc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6b440),
	.w1(32'h3c46b9fc),
	.w2(32'h3be9aae5),
	.w3(32'h3c5819ea),
	.w4(32'h3a6761a0),
	.w5(32'hb9977834),
	.w6(32'h3c011d5d),
	.w7(32'h3b59b60c),
	.w8(32'hba687a4e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01480b),
	.w1(32'h3b8f5fb8),
	.w2(32'h3b19d5ea),
	.w3(32'hbb6eba85),
	.w4(32'h3aa55367),
	.w5(32'h3bb942c4),
	.w6(32'h3ae472d2),
	.w7(32'h3bc9a06e),
	.w8(32'hb96fb7b2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10fd18),
	.w1(32'hbc7544e2),
	.w2(32'hbbf6aba6),
	.w3(32'h3b160206),
	.w4(32'hbba3993f),
	.w5(32'hbb91886e),
	.w6(32'hbbda0e53),
	.w7(32'hbb43856e),
	.w8(32'hbba9b8a8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8ee88),
	.w1(32'hbaea1901),
	.w2(32'hb9d92e93),
	.w3(32'hbaac4e6a),
	.w4(32'hb9abb52f),
	.w5(32'h3a9b3547),
	.w6(32'h39f4be40),
	.w7(32'hb9e9a4c1),
	.w8(32'h3a1d5912),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0f0d1),
	.w1(32'hbc7987fa),
	.w2(32'hbbd70033),
	.w3(32'h3bde506e),
	.w4(32'hbc04443e),
	.w5(32'hbbbe7909),
	.w6(32'h39f458b7),
	.w7(32'hba5ab132),
	.w8(32'h3bd84512),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee3ef7),
	.w1(32'h3c53bd02),
	.w2(32'h3bbc4e95),
	.w3(32'h3c1c3658),
	.w4(32'hbb295806),
	.w5(32'hbacc8331),
	.w6(32'h3c19f38f),
	.w7(32'h3bf6abb0),
	.w8(32'h3b9129ca),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3c18a),
	.w1(32'h3d1aab91),
	.w2(32'h3d6edd2c),
	.w3(32'h3b7dcd7e),
	.w4(32'h3c9fab1c),
	.w5(32'h3cee21d2),
	.w6(32'h3cb81a0e),
	.w7(32'h3d048228),
	.w8(32'h3c9e9cc3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08faa0),
	.w1(32'hbcaf245b),
	.w2(32'hbc2787dc),
	.w3(32'h3c7876c1),
	.w4(32'hbc2c4ef0),
	.w5(32'hbac7adfb),
	.w6(32'hbc6f9a07),
	.w7(32'hbc4c2223),
	.w8(32'hbc10db35),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77fdc7),
	.w1(32'hbb42db6c),
	.w2(32'hbb95574d),
	.w3(32'hbbee4fa8),
	.w4(32'hbb8af780),
	.w5(32'hbba0357c),
	.w6(32'hbbafc175),
	.w7(32'hbb2b1f44),
	.w8(32'hba33dc59),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c254c),
	.w1(32'hbb3d2842),
	.w2(32'hbb2312df),
	.w3(32'hbb498d8c),
	.w4(32'hbad928a6),
	.w5(32'hba193460),
	.w6(32'hb9e7ca51),
	.w7(32'hbb29ad2e),
	.w8(32'hba0082ac),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb395a58),
	.w1(32'hbd2db1de),
	.w2(32'hbd5e88f1),
	.w3(32'hb8b3c1cd),
	.w4(32'hbcdfe546),
	.w5(32'hbd046f3e),
	.w6(32'hbc807083),
	.w7(32'hbd27571b),
	.w8(32'hbcee2a06),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd16931a),
	.w1(32'hbb820b63),
	.w2(32'hbba94bad),
	.w3(32'hbc9854bd),
	.w4(32'hbb76288d),
	.w5(32'h3b73e8ca),
	.w6(32'h39d1169f),
	.w7(32'h3b6e47f6),
	.w8(32'hbbba6042),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc178d26),
	.w1(32'hbbaafa81),
	.w2(32'h3baa6907),
	.w3(32'h3b6e80a4),
	.w4(32'h3b802c6f),
	.w5(32'h3c23edb6),
	.w6(32'hbc30a58c),
	.w7(32'h3a2bf186),
	.w8(32'h3b4a2ff9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d8dae),
	.w1(32'h38d0c5ac),
	.w2(32'h3c3168cc),
	.w3(32'h3bcb5424),
	.w4(32'h3b952a81),
	.w5(32'h3bd1d79b),
	.w6(32'hbbaf9b69),
	.w7(32'h3aac29f6),
	.w8(32'h3bce5bf0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f7991),
	.w1(32'hbb961161),
	.w2(32'h3b095e82),
	.w3(32'h3bd41c4a),
	.w4(32'hbb42a1cb),
	.w5(32'h3ab8c156),
	.w6(32'hb983e03d),
	.w7(32'h3b8af3db),
	.w8(32'hb8800720),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3dfea),
	.w1(32'hbba1c9c1),
	.w2(32'hb93deeef),
	.w3(32'h3bcbac7b),
	.w4(32'h3b204932),
	.w5(32'hba1098ea),
	.w6(32'hbbbfd1a4),
	.w7(32'hba497fe4),
	.w8(32'h3b55f7d2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89004d),
	.w1(32'hbd059cd9),
	.w2(32'hbd821b61),
	.w3(32'h39f936e8),
	.w4(32'hbcc44f06),
	.w5(32'hbd229741),
	.w6(32'hbc3602c0),
	.w7(32'hbced58ba),
	.w8(32'hbcac9183),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd245b96),
	.w1(32'h3ce1a9c0),
	.w2(32'h3cd755b9),
	.w3(32'hbcd12b72),
	.w4(32'h3bbc017b),
	.w5(32'h3c895108),
	.w6(32'h3c3319b6),
	.w7(32'h3ca0a4cb),
	.w8(32'h3b5f4abe),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48f655),
	.w1(32'h3c28a69a),
	.w2(32'h3c3ba4a6),
	.w3(32'h3c9b076e),
	.w4(32'h3bb245df),
	.w5(32'h3c262a46),
	.w6(32'h3af43ea9),
	.w7(32'h3b3357f3),
	.w8(32'hbb834140),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d1d62),
	.w1(32'h3cb4062f),
	.w2(32'h3d086188),
	.w3(32'h3c2dd959),
	.w4(32'h3b90269c),
	.w5(32'h3c4169c0),
	.w6(32'h3c7d95b6),
	.w7(32'h3ca982be),
	.w8(32'h3c078148),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd703ea),
	.w1(32'hbc21361e),
	.w2(32'hb837dbde),
	.w3(32'h3c2e1842),
	.w4(32'h3b02546d),
	.w5(32'h3c1089ac),
	.w6(32'h3b874e2b),
	.w7(32'h3bd1dcf9),
	.w8(32'hbb270e18),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49595e),
	.w1(32'hbb7af379),
	.w2(32'h3bb70156),
	.w3(32'h3c73f52f),
	.w4(32'h3b847b66),
	.w5(32'h3c492647),
	.w6(32'hbc25f50b),
	.w7(32'h39f44c6a),
	.w8(32'h3b6f5962),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd235e),
	.w1(32'h3be9c00f),
	.w2(32'h3cdfb167),
	.w3(32'h3b9363bd),
	.w4(32'hba9d27a0),
	.w5(32'h3c28a767),
	.w6(32'h39c50fa5),
	.w7(32'h3c7cee85),
	.w8(32'h3c465ed7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc7ebf),
	.w1(32'h3cbd762c),
	.w2(32'h3d023981),
	.w3(32'h3c919cfc),
	.w4(32'h3be0c323),
	.w5(32'h3cb42508),
	.w6(32'h3c1a794b),
	.w7(32'h3c9c61bc),
	.w8(32'h3c5e845a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf53437),
	.w1(32'hbb40d8b3),
	.w2(32'h3c0ca2d4),
	.w3(32'h3cb17084),
	.w4(32'hba882687),
	.w5(32'h3b09cb5c),
	.w6(32'hbbaaf41e),
	.w7(32'h3aef41ef),
	.w8(32'hba9cba20),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca82c8),
	.w1(32'hbc1ac078),
	.w2(32'hbbb1b3cf),
	.w3(32'h3b245260),
	.w4(32'hbc09d56b),
	.w5(32'hbb4f11c4),
	.w6(32'hbc63764e),
	.w7(32'hbbd36859),
	.w8(32'hbb6707bf),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1aacbc),
	.w1(32'hbbd37119),
	.w2(32'hbcdf3909),
	.w3(32'h3a39a1df),
	.w4(32'hba5eb963),
	.w5(32'hbc1eb00b),
	.w6(32'hbb2c2718),
	.w7(32'hbcb39b10),
	.w8(32'hbb14e029),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64f092),
	.w1(32'hbb882b68),
	.w2(32'h3ad8007e),
	.w3(32'hbb03d3df),
	.w4(32'hb9cbc8c6),
	.w5(32'h3abb3812),
	.w6(32'hbb5c53f2),
	.w7(32'hbb5e9241),
	.w8(32'hbb2e3dc5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be67920),
	.w1(32'hbaf4f4b2),
	.w2(32'hbb45ac8a),
	.w3(32'h3c47c828),
	.w4(32'hba300860),
	.w5(32'hbb8599bd),
	.w6(32'hbab39671),
	.w7(32'hbb8498b6),
	.w8(32'hbb7dfcc8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf50b6c),
	.w1(32'h3bd6a82a),
	.w2(32'h3bac78ab),
	.w3(32'h3bea35d5),
	.w4(32'h3c1f4351),
	.w5(32'h3bb39ce3),
	.w6(32'h3b251a59),
	.w7(32'h3b9b60dc),
	.w8(32'hbb6b2d81),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb136fc),
	.w1(32'h3cf6b4de),
	.w2(32'h3d3ed64d),
	.w3(32'hbbd1bcf9),
	.w4(32'h3c63c060),
	.w5(32'h3ca938be),
	.w6(32'h3ca6ec90),
	.w7(32'h3d025b6d),
	.w8(32'h3c14f1b6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb6275f),
	.w1(32'h3983f199),
	.w2(32'h3c214e90),
	.w3(32'h3c9c7762),
	.w4(32'hbaa32ea9),
	.w5(32'h3ba9722d),
	.w6(32'h3b85dba1),
	.w7(32'h3c2367b8),
	.w8(32'h3c49a745),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beea1c7),
	.w1(32'h3bee5bac),
	.w2(32'h3c078f42),
	.w3(32'h3c17e9b3),
	.w4(32'h39907d70),
	.w5(32'hb9f63db3),
	.w6(32'hbb48486d),
	.w7(32'hb988a2f2),
	.w8(32'hba3394ec),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59abc6),
	.w1(32'hbb881598),
	.w2(32'hbc2fec2d),
	.w3(32'h3bb23aa4),
	.w4(32'h3bc57d76),
	.w5(32'h3afa1bd4),
	.w6(32'hbb17f668),
	.w7(32'hbc1a46a4),
	.w8(32'hbb9fd388),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99950c),
	.w1(32'hbc165758),
	.w2(32'hbcb14414),
	.w3(32'h3bae950c),
	.w4(32'hbc051a0c),
	.w5(32'hbbc6a657),
	.w6(32'hbb01c4e8),
	.w7(32'hbc4454dc),
	.w8(32'hbc1aa1e1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83372c),
	.w1(32'h3c15f988),
	.w2(32'h3c27b390),
	.w3(32'hbaec435e),
	.w4(32'h3a072251),
	.w5(32'h3b23d91e),
	.w6(32'h3c3bed9f),
	.w7(32'h3c68e655),
	.w8(32'h3c42a00a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfd7cd),
	.w1(32'h3b24f74b),
	.w2(32'h3bf46841),
	.w3(32'h3bb74fd4),
	.w4(32'h3c201b74),
	.w5(32'hba80c9b4),
	.w6(32'h3b9d060b),
	.w7(32'h3be44373),
	.w8(32'hbb84ec2f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32e365),
	.w1(32'hbba3eca4),
	.w2(32'hbbf3d7ed),
	.w3(32'hbb41ade5),
	.w4(32'hbbd8d54c),
	.w5(32'hbc608cf8),
	.w6(32'hbbbc3f7a),
	.w7(32'hbbd5a122),
	.w8(32'hbbf6157c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8c91),
	.w1(32'hbb6ad270),
	.w2(32'hbb17d6d7),
	.w3(32'hbc85d5a3),
	.w4(32'hbab3e859),
	.w5(32'h3b3ca74f),
	.w6(32'hbbbcd88c),
	.w7(32'hbba83651),
	.w8(32'hbb7f01e4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a1ce6),
	.w1(32'hbb6e9fc4),
	.w2(32'hbba71fe8),
	.w3(32'h3b25788b),
	.w4(32'hba7e0712),
	.w5(32'hbbd7b164),
	.w6(32'h3acfd959),
	.w7(32'h3b0456ae),
	.w8(32'h3b1d26f8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba55feb),
	.w1(32'h3c16dbed),
	.w2(32'h3c9f557c),
	.w3(32'hbb5c2936),
	.w4(32'h3c234b84),
	.w5(32'h3c336771),
	.w6(32'h3bb8466c),
	.w7(32'h3bed1c95),
	.w8(32'h3c48021f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9caa77),
	.w1(32'h3c9e45b2),
	.w2(32'h3d12b00d),
	.w3(32'h3cad5939),
	.w4(32'h3c578fc2),
	.w5(32'h3cc7eac6),
	.w6(32'h3c51c827),
	.w7(32'h3c885f98),
	.w8(32'h3c4b3e31),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2716a),
	.w1(32'h3c4aacc3),
	.w2(32'h3cdab7c8),
	.w3(32'h3c922bd2),
	.w4(32'h3b941a73),
	.w5(32'h3c93fe39),
	.w6(32'hbb794bcb),
	.w7(32'h3b96a97d),
	.w8(32'h3987050f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80225d),
	.w1(32'h3a689a76),
	.w2(32'hba8a5abe),
	.w3(32'h3c7dfb8b),
	.w4(32'h3b55eb48),
	.w5(32'hba9e0e13),
	.w6(32'h3abab5cd),
	.w7(32'h3942f566),
	.w8(32'h3b22c23b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb497432),
	.w1(32'hba9e9578),
	.w2(32'hbbfc8e1d),
	.w3(32'hbb89b0e3),
	.w4(32'hbb885433),
	.w5(32'hbbcb4401),
	.w6(32'hb9d08166),
	.w7(32'hbb8e61ee),
	.w8(32'hbafd52bf),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ff0ce),
	.w1(32'hbaefbb94),
	.w2(32'hbbbc51dc),
	.w3(32'hbb9b4a4a),
	.w4(32'hbb69e932),
	.w5(32'h3a0dd2cd),
	.w6(32'hb8b68a08),
	.w7(32'hbc11ef60),
	.w8(32'hbb82a76d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6734f9),
	.w1(32'h3b9af34c),
	.w2(32'h3c181cc2),
	.w3(32'hbaa57948),
	.w4(32'h3b1dfe7d),
	.w5(32'h3a8e5878),
	.w6(32'h3b1aee55),
	.w7(32'h3bd3dc8b),
	.w8(32'h3b91dc78),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc8616),
	.w1(32'hbca2b8e2),
	.w2(32'hbcf65b67),
	.w3(32'h3b14fcff),
	.w4(32'hbc831a07),
	.w5(32'hbc2879b3),
	.w6(32'hbc61d8c1),
	.w7(32'hbcacbe68),
	.w8(32'hbad7a8d9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc51330),
	.w1(32'hbcb1a5a9),
	.w2(32'hbd3e7222),
	.w3(32'h3beb4f0a),
	.w4(32'hbbcb01ce),
	.w5(32'hbcb0163b),
	.w6(32'hbc9f332c),
	.w7(32'hbcca3f20),
	.w8(32'hbbbb08a6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8bf02),
	.w1(32'hbd35aaf5),
	.w2(32'hbd791135),
	.w3(32'hbc9261e0),
	.w4(32'hbc5d4f09),
	.w5(32'hbd068670),
	.w6(32'hbd065777),
	.w7(32'hbd164ad7),
	.w8(32'hbc687266),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0018c0),
	.w1(32'hbafff9b4),
	.w2(32'hbb714685),
	.w3(32'hbca8502b),
	.w4(32'hbc66073e),
	.w5(32'hbc083987),
	.w6(32'h3bd0ad8c),
	.w7(32'h3b11883c),
	.w8(32'h3b1ddc5d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32120d),
	.w1(32'hbc413d5f),
	.w2(32'hbab25d5c),
	.w3(32'hbb835d5b),
	.w4(32'hbc33dd06),
	.w5(32'hbc38a12e),
	.w6(32'hbb25a77b),
	.w7(32'hba91332a),
	.w8(32'hbb6eea36),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe68628),
	.w1(32'h3c6e93d8),
	.w2(32'h3cc7d65f),
	.w3(32'hbb377b6b),
	.w4(32'h3895acb9),
	.w5(32'h3bee10fd),
	.w6(32'h3c16f3a5),
	.w7(32'h3c02be4c),
	.w8(32'h3c024851),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af93855),
	.w1(32'hbbea2478),
	.w2(32'hbbf5fcaa),
	.w3(32'hbc1a1952),
	.w4(32'hbbf551a4),
	.w5(32'hbbf95c9d),
	.w6(32'hbc4de477),
	.w7(32'hbc837643),
	.w8(32'hbc3b2711),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dae47),
	.w1(32'hbafcb809),
	.w2(32'hba47d3dc),
	.w3(32'hbc0c7c8d),
	.w4(32'hbbbd9835),
	.w5(32'hba85de99),
	.w6(32'hbbb562fa),
	.w7(32'hbb55c4ff),
	.w8(32'hbaea5d0d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8a831),
	.w1(32'hbca81ee2),
	.w2(32'hbbe7c938),
	.w3(32'h3b9328df),
	.w4(32'hbc2d5504),
	.w5(32'hbbbb0bb5),
	.w6(32'hbc2ec661),
	.w7(32'h3af1699f),
	.w8(32'hbc2284bb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390460b0),
	.w1(32'h3b300978),
	.w2(32'h3b21a8c3),
	.w3(32'hbc18e4c0),
	.w4(32'h3bead037),
	.w5(32'h3b541e18),
	.w6(32'hba95fb17),
	.w7(32'h399ebe1a),
	.w8(32'hbb3f8bab),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4d930),
	.w1(32'hbb470f29),
	.w2(32'h3b0432df),
	.w3(32'hbb4facc2),
	.w4(32'h3bbdf6bf),
	.w5(32'hbb771c72),
	.w6(32'hbae0152c),
	.w7(32'h3b822cfb),
	.w8(32'h3b2ccf9a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a2e9b),
	.w1(32'hba910382),
	.w2(32'h3b573548),
	.w3(32'h3a226c62),
	.w4(32'hbb5359f1),
	.w5(32'hbb48d830),
	.w6(32'h3c1b4b22),
	.w7(32'h3c9c950c),
	.w8(32'h3c304cca),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c929c),
	.w1(32'h3c1255d2),
	.w2(32'h3c77b96f),
	.w3(32'hbb8d39cc),
	.w4(32'h3c25e53c),
	.w5(32'h3c6d87a5),
	.w6(32'h3a902119),
	.w7(32'h3b155cf6),
	.w8(32'h3b843c42),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcabaaa),
	.w1(32'h3ad3b5cd),
	.w2(32'hbb131ca6),
	.w3(32'h3c2cd154),
	.w4(32'h3ad2a571),
	.w5(32'hba53c890),
	.w6(32'h3b5a5aee),
	.w7(32'hb8e8ef6f),
	.w8(32'h3aa90911),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcf80e),
	.w1(32'hbc146a0f),
	.w2(32'hbc2d114f),
	.w3(32'h3b4d7639),
	.w4(32'hbc76acdc),
	.w5(32'hbc09be9c),
	.w6(32'hbc7bc428),
	.w7(32'hbbd8fdc6),
	.w8(32'hbb69637c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72efd0),
	.w1(32'h3b012bdd),
	.w2(32'h3b78f54e),
	.w3(32'h3b1b36d1),
	.w4(32'h3b86e368),
	.w5(32'h3ab344cd),
	.w6(32'hbaf095c7),
	.w7(32'h3b192d63),
	.w8(32'h3b98e578),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d299a),
	.w1(32'hbc5c9368),
	.w2(32'hbcf63455),
	.w3(32'hbb0b7a79),
	.w4(32'h3a932cc4),
	.w5(32'hbc8a8d28),
	.w6(32'hbb61b9ba),
	.w7(32'hbca5cf94),
	.w8(32'hbbaecd75),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40a813),
	.w1(32'h3b512528),
	.w2(32'h3c2db515),
	.w3(32'hbc0ddea4),
	.w4(32'hbb5cd86c),
	.w5(32'h3bb7e8c1),
	.w6(32'h3ae99ff7),
	.w7(32'h3b4db119),
	.w8(32'h3aefae87),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60815f),
	.w1(32'hba6ba418),
	.w2(32'h3b88c20a),
	.w3(32'h3bf54d14),
	.w4(32'h3b485b0c),
	.w5(32'hbab83e24),
	.w6(32'h3b10735b),
	.w7(32'h3ab4812f),
	.w8(32'hbb39ebbb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a3772),
	.w1(32'hb9a449a8),
	.w2(32'h3a447e86),
	.w3(32'hbbddcf30),
	.w4(32'h3a2b812d),
	.w5(32'hb9fca6fd),
	.w6(32'h3b4679e0),
	.w7(32'h3afa464c),
	.w8(32'h3b06849a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b949d),
	.w1(32'h3b38694d),
	.w2(32'h3a2fe97e),
	.w3(32'h3ab7baea),
	.w4(32'h3c1aa68e),
	.w5(32'h3c1060a0),
	.w6(32'h3bb5b8d1),
	.w7(32'h3ba32c54),
	.w8(32'hbbbd0acd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc2f3b),
	.w1(32'h3a7f360b),
	.w2(32'hb9be6cce),
	.w3(32'h3a9088fc),
	.w4(32'hba4669d5),
	.w5(32'hbb0653ea),
	.w6(32'hbb41c746),
	.w7(32'hbb30f66f),
	.w8(32'hbb4d5e9f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f63e7),
	.w1(32'h3b93369e),
	.w2(32'hbb17a612),
	.w3(32'h3ad657d3),
	.w4(32'h3b4ca288),
	.w5(32'hbc5c296d),
	.w6(32'h3b77a1c7),
	.w7(32'h3be56e3b),
	.w8(32'hba835b36),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35addf),
	.w1(32'hbab2152b),
	.w2(32'h3bbd3fb0),
	.w3(32'hbbac7571),
	.w4(32'h3b2c9138),
	.w5(32'h3c553c25),
	.w6(32'hba59d8a2),
	.w7(32'h3b719b26),
	.w8(32'hb9f60421),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58bb39),
	.w1(32'h3d1963d3),
	.w2(32'h3d60bff9),
	.w3(32'h3c648d4b),
	.w4(32'h3c88159a),
	.w5(32'h3ce6f5f0),
	.w6(32'h3cca306a),
	.w7(32'h3d0911e4),
	.w8(32'h3b7a1a82),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01db5d),
	.w1(32'hb7afb747),
	.w2(32'h3c293a49),
	.w3(32'h3cb10a02),
	.w4(32'h3bc9ddb9),
	.w5(32'hb9953b41),
	.w6(32'h3bbf4184),
	.w7(32'h39a667fa),
	.w8(32'hbbedeb6a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5059ed),
	.w1(32'h3bd64713),
	.w2(32'h3adf7249),
	.w3(32'h3becdc5f),
	.w4(32'h3b17cf5c),
	.w5(32'h3960d8fd),
	.w6(32'h3b541ccb),
	.w7(32'h3b55b212),
	.w8(32'h3b7d1e27),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be6383),
	.w1(32'hbc56eb2e),
	.w2(32'hbd3568b5),
	.w3(32'h3a94c757),
	.w4(32'hbbd39fb6),
	.w5(32'hbcc7a0c1),
	.w6(32'hbba3ccaf),
	.w7(32'hbcb06b36),
	.w8(32'hbc01dbce),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabdbb1),
	.w1(32'hbc12741c),
	.w2(32'hbc8a86b6),
	.w3(32'hbc198559),
	.w4(32'hbc0d9c61),
	.w5(32'hbc041343),
	.w6(32'h3b6b747a),
	.w7(32'h3bc9a8c7),
	.w8(32'hbbc3d18d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5a7dc),
	.w1(32'hbc85d81d),
	.w2(32'hbd1a0c02),
	.w3(32'hbbfffe08),
	.w4(32'hbbaaac93),
	.w5(32'hbc8959fe),
	.w6(32'hbb81feaf),
	.w7(32'hbca3547b),
	.w8(32'hbc87d053),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0b561),
	.w1(32'h3b1eda9f),
	.w2(32'hbb789077),
	.w3(32'hbba80659),
	.w4(32'h39dfdfe9),
	.w5(32'hbb25d987),
	.w6(32'h3b5eec17),
	.w7(32'h3b336c7a),
	.w8(32'h3aa51984),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9376ad),
	.w1(32'hbc159a44),
	.w2(32'hbbfe4887),
	.w3(32'hbadc41c1),
	.w4(32'hbb445d75),
	.w5(32'hbbba7657),
	.w6(32'hbc982169),
	.w7(32'hbc82fe1e),
	.w8(32'hbc5c8d1f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule