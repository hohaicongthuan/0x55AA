module layer_10_featuremap_248(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06efd7),
	.w1(32'h3b562485),
	.w2(32'h3a67eb56),
	.w3(32'hbb9c1fb5),
	.w4(32'hba77a6e3),
	.w5(32'h3a37b364),
	.w6(32'hbae858f0),
	.w7(32'h3b88e382),
	.w8(32'hbae22ffe),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa647ee),
	.w1(32'hb9c9d7c6),
	.w2(32'h3bfb981a),
	.w3(32'h3b9d8f30),
	.w4(32'hb9ffb245),
	.w5(32'hbbc85a73),
	.w6(32'h3b6b3695),
	.w7(32'h3aa6f84f),
	.w8(32'hbb95e6b4),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae293a5),
	.w1(32'h3a485c3b),
	.w2(32'h3b1176fd),
	.w3(32'hbba74fc0),
	.w4(32'hbaeaa776),
	.w5(32'h3b2c6ee3),
	.w6(32'hbb5ee8c8),
	.w7(32'hb9c55905),
	.w8(32'h3a9747f5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92a0e0),
	.w1(32'h3b27c8db),
	.w2(32'h3b3ff078),
	.w3(32'hbaee528d),
	.w4(32'h3ac4d212),
	.w5(32'h3b4a6be5),
	.w6(32'h3a81d369),
	.w7(32'h3afe0e4a),
	.w8(32'hbc24241e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c030fcf),
	.w1(32'h3b959562),
	.w2(32'h3c038068),
	.w3(32'hba279527),
	.w4(32'h3bb44cf6),
	.w5(32'h3af97031),
	.w6(32'hbc32aca4),
	.w7(32'h3a6634e2),
	.w8(32'h3a9712f2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abddc37),
	.w1(32'hba46b5e2),
	.w2(32'hbadf3ff9),
	.w3(32'hb98e2659),
	.w4(32'hb97fa68d),
	.w5(32'h3c16fecc),
	.w6(32'hba99ca68),
	.w7(32'hba185e21),
	.w8(32'h3bb5c653),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8b327),
	.w1(32'hba2686e3),
	.w2(32'hb8aac7e5),
	.w3(32'h3b1644f9),
	.w4(32'hbadb25a6),
	.w5(32'hbb7e27db),
	.w6(32'hbba54c9a),
	.w7(32'hbab6a010),
	.w8(32'hbba5e606),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af507db),
	.w1(32'h3b3c6be8),
	.w2(32'h3b1a2a63),
	.w3(32'hbc21d20f),
	.w4(32'hbb44fc63),
	.w5(32'h3b6b4027),
	.w6(32'hbbacea31),
	.w7(32'h3ad44191),
	.w8(32'h3be71506),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8e629),
	.w1(32'h3b26b247),
	.w2(32'h3a6770c2),
	.w3(32'h3ad6f4d3),
	.w4(32'h3b1efc7d),
	.w5(32'h3b1d767d),
	.w6(32'h3b40eaec),
	.w7(32'h3b09e7e4),
	.w8(32'h3a2706d3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb520ec6),
	.w1(32'hba9e4583),
	.w2(32'hbc279b4d),
	.w3(32'hbb52142d),
	.w4(32'hbb18ccf2),
	.w5(32'hbbeab17a),
	.w6(32'hbba5c4f7),
	.w7(32'hbb067463),
	.w8(32'hbbff71ce),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4fd50),
	.w1(32'hba8c6ddc),
	.w2(32'hbb00b51b),
	.w3(32'hbbc8c38e),
	.w4(32'hbb53e95e),
	.w5(32'hbbad65d4),
	.w6(32'hbbe2cac3),
	.w7(32'hbaf1422c),
	.w8(32'hbb274e31),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be95d57),
	.w1(32'h3c4b12c0),
	.w2(32'h3bf38ecb),
	.w3(32'hbb363a26),
	.w4(32'h3b2897cf),
	.w5(32'hbc61d38c),
	.w6(32'hbb307c80),
	.w7(32'h3bfead8f),
	.w8(32'hbc2f2c67),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc343a1e),
	.w1(32'hbbf1cd50),
	.w2(32'hbc528a70),
	.w3(32'hbc4c9db1),
	.w4(32'hbbaae9eb),
	.w5(32'hbb89f001),
	.w6(32'hbb9bd6a4),
	.w7(32'hba89eca6),
	.w8(32'hbad92623),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08b247),
	.w1(32'h39040bcc),
	.w2(32'hbae99412),
	.w3(32'hba4c4f9f),
	.w4(32'hbb6a440e),
	.w5(32'hbb3d0f8b),
	.w6(32'h3b5c0c19),
	.w7(32'hb9d69413),
	.w8(32'hbaded607),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9808a0),
	.w1(32'h3bc2be9b),
	.w2(32'h3b0f8167),
	.w3(32'hbaff3b47),
	.w4(32'h3bbd9a1f),
	.w5(32'hbb8928c9),
	.w6(32'hbafdd691),
	.w7(32'h3b90b962),
	.w8(32'hb95fd653),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb743e54),
	.w1(32'hbb2310d0),
	.w2(32'hbb9e6456),
	.w3(32'hbc62ec26),
	.w4(32'hbba0b175),
	.w5(32'hbbd8c127),
	.w6(32'hbc0c5545),
	.w7(32'h3b67e351),
	.w8(32'hbb88ed33),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b032e38),
	.w1(32'h3c2ca3da),
	.w2(32'h3bdc80b0),
	.w3(32'hba7138c2),
	.w4(32'hbb5b8ae2),
	.w5(32'hbb356394),
	.w6(32'h3b81662b),
	.w7(32'h3a0fee55),
	.w8(32'hba437c64),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6d0c7),
	.w1(32'hbb2a38a7),
	.w2(32'hbb8b356b),
	.w3(32'hbac58e05),
	.w4(32'hbb984af2),
	.w5(32'hbbc1fb48),
	.w6(32'h3b47abe5),
	.w7(32'h3b0f7431),
	.w8(32'h3a190571),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6905cb),
	.w1(32'hbb6c452e),
	.w2(32'hbb2b9a68),
	.w3(32'hbb8b367f),
	.w4(32'hbb06dece),
	.w5(32'h3a62970b),
	.w6(32'hba95dc9c),
	.w7(32'h3add6d4c),
	.w8(32'h3abf7db5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b779d2d),
	.w1(32'h3b413177),
	.w2(32'hba3f2a0d),
	.w3(32'h3ae74e5b),
	.w4(32'hba507fae),
	.w5(32'hbb1f6cde),
	.w6(32'h3b1fbf14),
	.w7(32'hba14f266),
	.w8(32'h3b4b47aa),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e95809),
	.w1(32'h39091d19),
	.w2(32'h389d5e92),
	.w3(32'hbbb6a028),
	.w4(32'hb8051392),
	.w5(32'h3bddd3a4),
	.w6(32'hba0aaa8d),
	.w7(32'h3be65555),
	.w8(32'h3b1e3ec6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78193c),
	.w1(32'h3a9c908e),
	.w2(32'h3929e7c2),
	.w3(32'h3b8d3115),
	.w4(32'h3bcb8a6c),
	.w5(32'hbb56016d),
	.w6(32'hbb35cb31),
	.w7(32'h394b2767),
	.w8(32'hbb4c9c7c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba729dc),
	.w1(32'hba8c6a35),
	.w2(32'hbaafe11d),
	.w3(32'hbc2a3a95),
	.w4(32'hbb6baf80),
	.w5(32'hbbf744b7),
	.w6(32'hbc223aa6),
	.w7(32'hbafd651a),
	.w8(32'hbb74fe4d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17b786),
	.w1(32'hba9c631f),
	.w2(32'hbc40ecdf),
	.w3(32'hbc6b3100),
	.w4(32'hbc13f53d),
	.w5(32'hbb6b55c4),
	.w6(32'hbac663bd),
	.w7(32'h3b00fece),
	.w8(32'hbb6e2da5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3205e5),
	.w1(32'hbb5bfd47),
	.w2(32'hbb9ec6b1),
	.w3(32'h396c1cb4),
	.w4(32'hbac052d4),
	.w5(32'hbaa644ec),
	.w6(32'hbb92fcfd),
	.w7(32'hbba1e9cf),
	.w8(32'hbb37950b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b588504),
	.w1(32'h3b9bbed0),
	.w2(32'hba92617e),
	.w3(32'hbb56b472),
	.w4(32'h3a715b85),
	.w5(32'h3b8bce95),
	.w6(32'hbb6cad42),
	.w7(32'hb9307c9a),
	.w8(32'h3b9eee35),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9729f8),
	.w1(32'h3a6aee53),
	.w2(32'h3b3b12df),
	.w3(32'hbb1e7065),
	.w4(32'h3ab88758),
	.w5(32'h3b2dce92),
	.w6(32'hbaf9f552),
	.w7(32'h3b09741e),
	.w8(32'h3ba0c46b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd5fd6),
	.w1(32'h3a58e144),
	.w2(32'hbb85de27),
	.w3(32'h3a7ed4d9),
	.w4(32'hbb09d177),
	.w5(32'h3b8224cf),
	.w6(32'h3b634916),
	.w7(32'hbb019453),
	.w8(32'h3ad4146e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c8d73),
	.w1(32'hb9d30711),
	.w2(32'hbac4c134),
	.w3(32'h3b30602a),
	.w4(32'h3b193610),
	.w5(32'hbb68808c),
	.w6(32'h3a6e7796),
	.w7(32'h3b7fc1e6),
	.w8(32'hbb132d4b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba049020),
	.w1(32'h3a7a8d2c),
	.w2(32'hb96eb8e0),
	.w3(32'hbc12a1c0),
	.w4(32'hbb825930),
	.w5(32'hbb8c8fea),
	.w6(32'hbbc1633f),
	.w7(32'h3aa9056c),
	.w8(32'hbc045451),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb7e1),
	.w1(32'hbc08e958),
	.w2(32'hbc17a663),
	.w3(32'h3b094975),
	.w4(32'hbad73e81),
	.w5(32'hbbc305bf),
	.w6(32'hbbfd4f0e),
	.w7(32'hbc0e21f7),
	.w8(32'hba9602a1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7587da),
	.w1(32'h3bd87eb5),
	.w2(32'h3b8fa3e1),
	.w3(32'hbb22081d),
	.w4(32'hbb8ed7c8),
	.w5(32'h3ad2c11b),
	.w6(32'hbb623fac),
	.w7(32'hbb5c3f50),
	.w8(32'h3c0f4c95),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a66ce),
	.w1(32'hbad53baa),
	.w2(32'h39835e43),
	.w3(32'h3b09ee23),
	.w4(32'hbb0259a5),
	.w5(32'hbbbe9deb),
	.w6(32'hbb9b54ce),
	.w7(32'hbb5ba39e),
	.w8(32'hbb3a9e7a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb271c2f),
	.w1(32'hbb35fb7f),
	.w2(32'hbad090a7),
	.w3(32'h3a5a5556),
	.w4(32'hbb17f231),
	.w5(32'hba4e3387),
	.w6(32'h3a09cce0),
	.w7(32'h3ac92a50),
	.w8(32'hba3de827),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af06539),
	.w1(32'hbb02dce3),
	.w2(32'hb91c7d0d),
	.w3(32'hb953f2b1),
	.w4(32'h3957ab42),
	.w5(32'h3992bdbf),
	.w6(32'hbaf062b0),
	.w7(32'h3a8ce444),
	.w8(32'hbabbb415),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc86fc7),
	.w1(32'hbba26fe9),
	.w2(32'hbb801d2b),
	.w3(32'hba66d20f),
	.w4(32'hbb76f51e),
	.w5(32'hbaf941a0),
	.w6(32'h3b0ec6bb),
	.w7(32'h3aaf3f44),
	.w8(32'hba463fc8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6192be),
	.w1(32'hbbe7a022),
	.w2(32'hbc0d1acb),
	.w3(32'h39b06b39),
	.w4(32'h3aa0908e),
	.w5(32'h3b3392af),
	.w6(32'hbb8f1e76),
	.w7(32'h3b952189),
	.w8(32'h3bb34db0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb779668),
	.w1(32'hbc0e5e37),
	.w2(32'hbb018931),
	.w3(32'hbb4e1cfb),
	.w4(32'h3bc5f5ef),
	.w5(32'h3b8a1dba),
	.w6(32'hbbee3445),
	.w7(32'hba8a9e5c),
	.w8(32'hbc1dd491),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a49d3c),
	.w1(32'h3b235d70),
	.w2(32'hbb6fa927),
	.w3(32'h3c1f8349),
	.w4(32'h3b6ca4d4),
	.w5(32'h3b1778f6),
	.w6(32'hbb8ed7c9),
	.w7(32'hbc05c99d),
	.w8(32'hbac485e9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c0fce),
	.w1(32'hbb28f606),
	.w2(32'h3b62fb88),
	.w3(32'h3a4688c6),
	.w4(32'h3b575712),
	.w5(32'hbb622139),
	.w6(32'hbba7b8af),
	.w7(32'h3bb2e4fb),
	.w8(32'hbb0789d0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ec4cc),
	.w1(32'h3b2159d8),
	.w2(32'hb9b1bc76),
	.w3(32'hbb5063e8),
	.w4(32'h3a5fe08d),
	.w5(32'h3bbd1f92),
	.w6(32'h3aaafe45),
	.w7(32'h3b3fbbef),
	.w8(32'hba7ea611),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2fb4a),
	.w1(32'h3b5a87c1),
	.w2(32'hba2f9bc3),
	.w3(32'hb9234b51),
	.w4(32'h3ab612a6),
	.w5(32'hbb80ed53),
	.w6(32'hbc13e29e),
	.w7(32'hbb554167),
	.w8(32'hbab3659c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7b4cc),
	.w1(32'hbc350a25),
	.w2(32'hbbbad08a),
	.w3(32'hbc0abac6),
	.w4(32'hbb8da1ef),
	.w5(32'hbbaa1018),
	.w6(32'hbbc7c2db),
	.w7(32'hbaee1032),
	.w8(32'hbbc7a69b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50c6b9),
	.w1(32'h3abaf3d1),
	.w2(32'h3b63bcee),
	.w3(32'hbb035744),
	.w4(32'hb95247f1),
	.w5(32'hb756a101),
	.w6(32'h3b86ab11),
	.w7(32'h3bc7b63d),
	.w8(32'h39c8ed11),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba982656),
	.w1(32'h3a547900),
	.w2(32'hbba006cb),
	.w3(32'h3a8ef835),
	.w4(32'h3b50cd2b),
	.w5(32'hbad1db26),
	.w6(32'hbb96c935),
	.w7(32'h39849cd5),
	.w8(32'hbbb7d436),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae27f7f),
	.w1(32'hbb9184da),
	.w2(32'hbbcf50ec),
	.w3(32'h3ad87e07),
	.w4(32'hbb7b60e5),
	.w5(32'hbba95f4c),
	.w6(32'hbbe42935),
	.w7(32'hbb9f0ed5),
	.w8(32'hbbaa7422),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d02b7),
	.w1(32'h3a3acd0c),
	.w2(32'h3b32d220),
	.w3(32'hbb318013),
	.w4(32'h3a2d111f),
	.w5(32'h3b4d7999),
	.w6(32'hbbc78a8d),
	.w7(32'hbae7595a),
	.w8(32'h3aa2e392),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b2c67),
	.w1(32'hbaec1c45),
	.w2(32'hbb755d44),
	.w3(32'h3a8bbd36),
	.w4(32'h3b6a32fb),
	.w5(32'hbc062f72),
	.w6(32'h39dc6147),
	.w7(32'h3b55e4e8),
	.w8(32'hbb042079),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba60878),
	.w1(32'hbb3edbc2),
	.w2(32'hbbc61263),
	.w3(32'hbb462025),
	.w4(32'hba30d803),
	.w5(32'h3c4d654f),
	.w6(32'h3b7677b4),
	.w7(32'h3a5fafec),
	.w8(32'h3bc7d3cd),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f7a8),
	.w1(32'h3ac4cf3b),
	.w2(32'h3b420586),
	.w3(32'h3ab2113a),
	.w4(32'h3bdf9acf),
	.w5(32'h3ba343c6),
	.w6(32'hbc1da9b6),
	.w7(32'h3a041d4a),
	.w8(32'h3bdde6b6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b428949),
	.w1(32'hbbc75e77),
	.w2(32'hbb988d0f),
	.w3(32'hb9230a82),
	.w4(32'hbbc48dbf),
	.w5(32'hbb2fc8c3),
	.w6(32'h3b2ea5f6),
	.w7(32'hbbf00e47),
	.w8(32'h3aa80ee3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba685b57),
	.w1(32'hba3d38a7),
	.w2(32'h3b04585b),
	.w3(32'hbb0a177b),
	.w4(32'hbb21216a),
	.w5(32'hbb7f91b7),
	.w6(32'h3b4dcc21),
	.w7(32'hbaa55972),
	.w8(32'hbb5e0824),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f45a4),
	.w1(32'h39bc353a),
	.w2(32'hbb23c1a3),
	.w3(32'hbbd70532),
	.w4(32'hbbba5ce8),
	.w5(32'hbc06338d),
	.w6(32'hbb319dcd),
	.w7(32'hbb0f89b4),
	.w8(32'hbbc53b8f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba21f62),
	.w1(32'hbbede28e),
	.w2(32'hbb8b1e5c),
	.w3(32'hbc239e7e),
	.w4(32'h3b7b96d2),
	.w5(32'hbb8f2dd7),
	.w6(32'hbc474e21),
	.w7(32'h3c689531),
	.w8(32'hbb1153ea),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22c8f2),
	.w1(32'h3aff4d57),
	.w2(32'hbb1e3e3a),
	.w3(32'hba9d91f2),
	.w4(32'hbb1df639),
	.w5(32'hbadc33cc),
	.w6(32'h3b1c55e3),
	.w7(32'hb992351b),
	.w8(32'hbba64b02),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9531fb),
	.w1(32'hbb42ba21),
	.w2(32'hbb841d61),
	.w3(32'h391ee722),
	.w4(32'hbb2be0c4),
	.w5(32'hbaf7291f),
	.w6(32'hbacb82f1),
	.w7(32'hba98a368),
	.w8(32'hba85d9b2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac9b85),
	.w1(32'hba979ad4),
	.w2(32'hbb7ea537),
	.w3(32'hb9d0e72d),
	.w4(32'h3a9f36d3),
	.w5(32'hbb724cd3),
	.w6(32'h3b05c840),
	.w7(32'h3b086230),
	.w8(32'hbbbc60de),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff184c),
	.w1(32'hba0071a5),
	.w2(32'h3a80d33e),
	.w3(32'hbac6b7c2),
	.w4(32'h3a8f474d),
	.w5(32'h3c70c39b),
	.w6(32'hbb0721a4),
	.w7(32'h3bdde179),
	.w8(32'h3c19e284),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c273666),
	.w1(32'h3b822c30),
	.w2(32'h3b97dea9),
	.w3(32'h3a89372f),
	.w4(32'h3bf9670d),
	.w5(32'h3c3a2d26),
	.w6(32'hbc192215),
	.w7(32'h3a9f4723),
	.w8(32'h3b80a439),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b6bf9),
	.w1(32'hbc1fbd44),
	.w2(32'hbbfb0593),
	.w3(32'h3c602414),
	.w4(32'h3c2ca490),
	.w5(32'h3a27a8a5),
	.w6(32'h3a1938dc),
	.w7(32'hbbb717ac),
	.w8(32'hbb41c40f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea01bc),
	.w1(32'h3ac233a1),
	.w2(32'hbbacbf7e),
	.w3(32'h3b79f76f),
	.w4(32'h3b44cf75),
	.w5(32'hbb0257b5),
	.w6(32'hbb3e7722),
	.w7(32'hba8c9f52),
	.w8(32'hbbfb01ba),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42da83),
	.w1(32'h39c4251f),
	.w2(32'hbb81528d),
	.w3(32'hbbed2ef5),
	.w4(32'hbbf6ac45),
	.w5(32'hb9cf0a93),
	.w6(32'hbc1e75ac),
	.w7(32'hbc071fdd),
	.w8(32'hbb81c305),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b094a40),
	.w1(32'h39d63c2c),
	.w2(32'h3a63a096),
	.w3(32'h3a98f976),
	.w4(32'hb9f5fc1a),
	.w5(32'hbab1dc95),
	.w6(32'hbb220478),
	.w7(32'hbaf75322),
	.w8(32'hbb0dd60d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa08dae),
	.w1(32'hbaa1c652),
	.w2(32'h3a09fb60),
	.w3(32'hba87002d),
	.w4(32'h3b56eccf),
	.w5(32'h3b05dda3),
	.w6(32'h39a0db6c),
	.w7(32'h3bde4f1d),
	.w8(32'h3a449a2a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41291b),
	.w1(32'hbbc26bcc),
	.w2(32'hba6f58f1),
	.w3(32'hbb65d9dd),
	.w4(32'hba53b723),
	.w5(32'h3ad4d520),
	.w6(32'hbb62b159),
	.w7(32'h3b08de7a),
	.w8(32'hbb89370f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac66e09),
	.w1(32'h3b0a345b),
	.w2(32'hbb61c625),
	.w3(32'hba037e0d),
	.w4(32'h37fa171c),
	.w5(32'hbb913bd4),
	.w6(32'hba4982c5),
	.w7(32'hbac4b3c4),
	.w8(32'hbbe95315),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38888ea8),
	.w1(32'h3bdb00c7),
	.w2(32'h3a0f67dc),
	.w3(32'hbbca8583),
	.w4(32'hbb393d11),
	.w5(32'hbbbd9d24),
	.w6(32'hbb84e092),
	.w7(32'h39aa4381),
	.w8(32'hbb836f51),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa64b08),
	.w1(32'hbb1f09a8),
	.w2(32'hbb90e04a),
	.w3(32'hba9042b2),
	.w4(32'h3b29655b),
	.w5(32'hba509207),
	.w6(32'h3b63d503),
	.w7(32'h3b755891),
	.w8(32'h3b06fe32),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6cbe3),
	.w1(32'h3ac9a2ac),
	.w2(32'hbb82760a),
	.w3(32'hbb84243c),
	.w4(32'hbb901201),
	.w5(32'hbb1deea1),
	.w6(32'h39738ed5),
	.w7(32'hba2da26d),
	.w8(32'hba2fa25a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17944b),
	.w1(32'h38ddb0ef),
	.w2(32'hbb112ca4),
	.w3(32'h39cfaf52),
	.w4(32'h3b909283),
	.w5(32'h38a81e91),
	.w6(32'hbb228e05),
	.w7(32'h3b2c0ded),
	.w8(32'hbaad9fee),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b543c),
	.w1(32'hbb023c4b),
	.w2(32'h39c460ef),
	.w3(32'hbbaacf7b),
	.w4(32'h3a5787a7),
	.w5(32'hbbeeb9fc),
	.w6(32'hba828a47),
	.w7(32'h3ab7d91d),
	.w8(32'hbb3e6b1b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb117b7a),
	.w1(32'h3ba6f123),
	.w2(32'h3b8bc8e3),
	.w3(32'hbb8ccddd),
	.w4(32'hbb26d183),
	.w5(32'hba9a5245),
	.w6(32'hbabd151b),
	.w7(32'h3b220891),
	.w8(32'hb901f497),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dad04),
	.w1(32'h3a850500),
	.w2(32'hbb9e6b22),
	.w3(32'h395f93ba),
	.w4(32'hbabf8ab3),
	.w5(32'hbb0d330d),
	.w6(32'h3bafee82),
	.w7(32'hb9ca601f),
	.w8(32'hba942e95),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbababbd6),
	.w1(32'hbbc07b6a),
	.w2(32'hb61a0d34),
	.w3(32'h3b7f7992),
	.w4(32'h3b035a98),
	.w5(32'hbbcddfd2),
	.w6(32'h3aca7913),
	.w7(32'h3b9a9ea1),
	.w8(32'hbb9d97b3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac99e7a),
	.w1(32'h3b43c2f3),
	.w2(32'h3b8cfc88),
	.w3(32'hbb9ab3ad),
	.w4(32'hba4ddc7e),
	.w5(32'hbc28b8ce),
	.w6(32'hbb28fda2),
	.w7(32'h3bdba657),
	.w8(32'hbbbeecc9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc332370),
	.w1(32'hbbe0a30c),
	.w2(32'hbbf278c4),
	.w3(32'hbb2d132d),
	.w4(32'hbbb03574),
	.w5(32'h386b4140),
	.w6(32'h3b7c9539),
	.w7(32'hba838a8d),
	.w8(32'hba736b78),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77517c),
	.w1(32'hbb0e1f74),
	.w2(32'hbb61c6b8),
	.w3(32'hbb00c6fa),
	.w4(32'h399e3303),
	.w5(32'hbbdef6b6),
	.w6(32'hbb1a7e74),
	.w7(32'h3ac95225),
	.w8(32'hbb81f257),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39462333),
	.w1(32'h3b978099),
	.w2(32'h3b8594a7),
	.w3(32'hbba89cda),
	.w4(32'hbb7d79d0),
	.w5(32'hbb5238ee),
	.w6(32'hbbcf0dad),
	.w7(32'hbb0e4bdf),
	.w8(32'hbad60f7e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94c1bc),
	.w1(32'h3a042bec),
	.w2(32'hbb996133),
	.w3(32'hbba4b5d6),
	.w4(32'hbb4d05b6),
	.w5(32'hbae92747),
	.w6(32'hbb37d532),
	.w7(32'hba7b765a),
	.w8(32'hbaf22c01),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb777f7),
	.w1(32'h3b6993b0),
	.w2(32'hba19812b),
	.w3(32'h39e75a98),
	.w4(32'hba68e9ed),
	.w5(32'hbb2a3b67),
	.w6(32'h3af21f68),
	.w7(32'hb8dd5699),
	.w8(32'hbb2d2d16),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba430b28),
	.w1(32'h3a3aacd3),
	.w2(32'hbbd5f487),
	.w3(32'hbb93e37e),
	.w4(32'h3b86ba43),
	.w5(32'hbb988439),
	.w6(32'hbb7b290b),
	.w7(32'h3b6f8a07),
	.w8(32'hbb5f5a67),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fb41f),
	.w1(32'hbb05d0b5),
	.w2(32'hbb863b79),
	.w3(32'h39cf8176),
	.w4(32'hb845bc59),
	.w5(32'hbbc09adb),
	.w6(32'h389584da),
	.w7(32'h3acb2797),
	.w8(32'hbb7663b2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e65a1),
	.w1(32'hbbdd3149),
	.w2(32'hbb048363),
	.w3(32'hbbfa073f),
	.w4(32'hbbb1f383),
	.w5(32'hbaf63bd9),
	.w6(32'hbc06f358),
	.w7(32'hbb18f0b6),
	.w8(32'h3b7929f6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05c557),
	.w1(32'h3c2501ee),
	.w2(32'h3ba075a1),
	.w3(32'h3b1d78df),
	.w4(32'h3bb7293b),
	.w5(32'hbb0ead32),
	.w6(32'h3c436deb),
	.w7(32'h3c24f47e),
	.w8(32'hb9b9c8bc),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6a5ae),
	.w1(32'h3931250c),
	.w2(32'h3ae152ee),
	.w3(32'hbb2b023a),
	.w4(32'hba127910),
	.w5(32'hba9803d4),
	.w6(32'hbb1463cb),
	.w7(32'h3a9c2380),
	.w8(32'hbb93f34b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fd1d1),
	.w1(32'hba6a10bf),
	.w2(32'hbbde375e),
	.w3(32'h3ac7fb01),
	.w4(32'hbb35dddc),
	.w5(32'hba452cc1),
	.w6(32'hbb2d2d8a),
	.w7(32'hbbab38d8),
	.w8(32'h39d49264),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7d073),
	.w1(32'h3b96c4ac),
	.w2(32'h3be89e28),
	.w3(32'hbbe5443b),
	.w4(32'h3ad5d8a2),
	.w5(32'h3b904aca),
	.w6(32'hbc0eec43),
	.w7(32'h3b978a72),
	.w8(32'h3b1008df),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24fcb6),
	.w1(32'hb98d7ad0),
	.w2(32'hba824e59),
	.w3(32'h3b9d2e1c),
	.w4(32'h3b9040df),
	.w5(32'h3bdd71f2),
	.w6(32'h3b113ee6),
	.w7(32'hba523892),
	.w8(32'h3b7371b5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7582a),
	.w1(32'h3b4cf61a),
	.w2(32'h3b3f2a62),
	.w3(32'h3b3925cb),
	.w4(32'h3b36169f),
	.w5(32'hbc12dc97),
	.w6(32'hbb8da550),
	.w7(32'hb98f83f8),
	.w8(32'hba9621fa),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e68e6),
	.w1(32'hba99bc9c),
	.w2(32'hbbfc0399),
	.w3(32'hbc6b7dce),
	.w4(32'hbc0c3b6c),
	.w5(32'hbbb6a692),
	.w6(32'hbb3bc256),
	.w7(32'hbb9ce8c5),
	.w8(32'h3b5b45a5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b020b78),
	.w1(32'hbb2dcf63),
	.w2(32'hbad50912),
	.w3(32'hbb09b0c2),
	.w4(32'hbbd42f09),
	.w5(32'hbb331657),
	.w6(32'hb9a7a977),
	.w7(32'hbb565c23),
	.w8(32'hbb78092d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0b64b),
	.w1(32'h3b8d7d29),
	.w2(32'hbb587945),
	.w3(32'hbb4f02eb),
	.w4(32'hbb9e1e11),
	.w5(32'hbc12d0ec),
	.w6(32'h3a273ce6),
	.w7(32'hba51dea9),
	.w8(32'hbc0efe73),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76d659),
	.w1(32'h3c736ec3),
	.w2(32'h3c361c9f),
	.w3(32'hbbe9e84b),
	.w4(32'hbb01b69a),
	.w5(32'hbb515f04),
	.w6(32'hbbf302d7),
	.w7(32'hbbaffd46),
	.w8(32'hbb4d83b2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4d122),
	.w1(32'h3b9639ab),
	.w2(32'h3b3be1cc),
	.w3(32'h3b01fdc2),
	.w4(32'h3b36bca0),
	.w5(32'hbb92d039),
	.w6(32'h3b70068f),
	.w7(32'h3bc6e420),
	.w8(32'h3ade89f5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2e172),
	.w1(32'hb98a3f69),
	.w2(32'hbb1b1137),
	.w3(32'hbbd384bf),
	.w4(32'hbb006632),
	.w5(32'hbbc1849a),
	.w6(32'hbb5d041f),
	.w7(32'h38e4ba98),
	.w8(32'hbaa93816),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3baf8),
	.w1(32'hbb142c80),
	.w2(32'hbb1e25fd),
	.w3(32'hbb8c546b),
	.w4(32'hbacee6aa),
	.w5(32'h3b82a35c),
	.w6(32'hbbbfd389),
	.w7(32'hbb265871),
	.w8(32'h3b2932e8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a254a2c),
	.w1(32'hba36600f),
	.w2(32'hb93e71a3),
	.w3(32'h3ada31ad),
	.w4(32'hba15d52e),
	.w5(32'hbb1d6281),
	.w6(32'h3ac3b537),
	.w7(32'hba91b64e),
	.w8(32'h3a474bfb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec5712),
	.w1(32'h3abdfc97),
	.w2(32'hbc0d336a),
	.w3(32'hbaf5980e),
	.w4(32'hbb27d1b1),
	.w5(32'hba25234d),
	.w6(32'h3afb0b79),
	.w7(32'hbb6442f0),
	.w8(32'h391e0196),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af96cc8),
	.w1(32'hb9cbd1f1),
	.w2(32'h3b437a57),
	.w3(32'h3ba3c3d4),
	.w4(32'h3b60e8c8),
	.w5(32'hbb56ca05),
	.w6(32'hbc116729),
	.w7(32'hba4f9ac6),
	.w8(32'hb94e251a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb957029),
	.w1(32'hbaf20946),
	.w2(32'hbaecefcf),
	.w3(32'h3a83868a),
	.w4(32'hbb8dd101),
	.w5(32'hbbd8dba9),
	.w6(32'hbba053da),
	.w7(32'h3b870321),
	.w8(32'hb987622c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc694448),
	.w1(32'hbb475e96),
	.w2(32'hbb23a4c8),
	.w3(32'hbbc58af4),
	.w4(32'h3b57aa7a),
	.w5(32'hbb8e5db6),
	.w6(32'hbc4d7ead),
	.w7(32'hbbc71155),
	.w8(32'h3d024a2d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b848d58),
	.w1(32'h3c2a3ea7),
	.w2(32'hbc0622bc),
	.w3(32'h3c803e48),
	.w4(32'h3c70f29d),
	.w5(32'hbc27763d),
	.w6(32'h3d39532c),
	.w7(32'h3cb90382),
	.w8(32'hbbc33d6d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc061376),
	.w1(32'hbc5853b0),
	.w2(32'hbcac0616),
	.w3(32'h3bf83b9d),
	.w4(32'h3b6d7525),
	.w5(32'hbc092396),
	.w6(32'hbaeac034),
	.w7(32'h3aea66c7),
	.w8(32'hbb99634b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a432c80),
	.w1(32'h3bc1b2c2),
	.w2(32'hbafaaeb9),
	.w3(32'hbb919f7d),
	.w4(32'hbaad464c),
	.w5(32'h3a6970ce),
	.w6(32'h3b2587dc),
	.w7(32'h3b8f4ff6),
	.w8(32'h39d1aacf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd847e0),
	.w1(32'hbc14fa3d),
	.w2(32'hbc153b73),
	.w3(32'h3b6cbf33),
	.w4(32'h3b8fd22f),
	.w5(32'h3bbfc164),
	.w6(32'hbc18a251),
	.w7(32'hbc2de29d),
	.w8(32'h3b2f902f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24d01a),
	.w1(32'hbae5aa6a),
	.w2(32'hbb137566),
	.w3(32'h3baae9d6),
	.w4(32'h3be49f7e),
	.w5(32'hbc1a0c75),
	.w6(32'hba69ea78),
	.w7(32'hba0da23b),
	.w8(32'h3af9b910),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb040485),
	.w1(32'h3b54183e),
	.w2(32'h3a91cfb8),
	.w3(32'hbb984d5c),
	.w4(32'hbb18c70a),
	.w5(32'hbbd0b570),
	.w6(32'h3c0ea6d0),
	.w7(32'h3c215802),
	.w8(32'hbaabc000),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a7562),
	.w1(32'hbb59bb93),
	.w2(32'hb93f2c22),
	.w3(32'hbb85e184),
	.w4(32'hbad962b6),
	.w5(32'h3b1b0b8a),
	.w6(32'hbb512ed1),
	.w7(32'hbaaa9947),
	.w8(32'h3a6d8eef),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd51dbd),
	.w1(32'hbbaee45b),
	.w2(32'hbb1be1e5),
	.w3(32'h3b092ca9),
	.w4(32'h3bb517b9),
	.w5(32'hbb9186cb),
	.w6(32'hbc269bd4),
	.w7(32'h3a46a80b),
	.w8(32'hbb2b2a18),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac944a3),
	.w1(32'hba009702),
	.w2(32'hba9fe9ef),
	.w3(32'hbac90b14),
	.w4(32'hba3c56e4),
	.w5(32'hb90d72a0),
	.w6(32'hbbf9dc28),
	.w7(32'hbb9381dd),
	.w8(32'h3ae04cd0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03c6d2),
	.w1(32'hbb6c56ed),
	.w2(32'h3a9f88f5),
	.w3(32'hbac14b8f),
	.w4(32'hba5b4642),
	.w5(32'hbc83062c),
	.w6(32'h3a28e0be),
	.w7(32'h3a18856b),
	.w8(32'hbc8d7034),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88482b),
	.w1(32'hbc859643),
	.w2(32'hbc0e0488),
	.w3(32'hbce09571),
	.w4(32'hbc780d44),
	.w5(32'hbb2f6641),
	.w6(32'hbc5052ee),
	.w7(32'hbc89111d),
	.w8(32'h3a386535),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c017d7d),
	.w1(32'h3a63ef19),
	.w2(32'h3ba7804d),
	.w3(32'h3a92e285),
	.w4(32'h3b00df92),
	.w5(32'hbc9c165e),
	.w6(32'hbbca4b9e),
	.w7(32'h3b5d647c),
	.w8(32'h3c4578e7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb520b),
	.w1(32'h3c3825da),
	.w2(32'hbbfdf1b3),
	.w3(32'hbc8b9f31),
	.w4(32'hbc915b3b),
	.w5(32'h39cc5d76),
	.w6(32'hbbb4adba),
	.w7(32'h3a97c450),
	.w8(32'h3b202be0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5ef31),
	.w1(32'h3beadcc9),
	.w2(32'h3ad8d863),
	.w3(32'hbb89ca89),
	.w4(32'h3b34a8a6),
	.w5(32'hbc6872c4),
	.w6(32'h3a080d41),
	.w7(32'hbac99459),
	.w8(32'hbb8bf220),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb830f61),
	.w1(32'hbc221e8d),
	.w2(32'hbc403667),
	.w3(32'hbc4fb246),
	.w4(32'hbc0fbf30),
	.w5(32'h38fe15a9),
	.w6(32'h3c524165),
	.w7(32'hbc8769dc),
	.w8(32'hbb2dd551),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9ef9e),
	.w1(32'hbaab33e7),
	.w2(32'hba356568),
	.w3(32'hbad5c519),
	.w4(32'hba914ba0),
	.w5(32'hb913855b),
	.w6(32'hbbc04750),
	.w7(32'hbba26fa2),
	.w8(32'hbb5830be),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e8c1f),
	.w1(32'hbac45fc6),
	.w2(32'h3a96c55a),
	.w3(32'h3b1c7b92),
	.w4(32'hbbc194fe),
	.w5(32'h3c159ae4),
	.w6(32'h3b8a504e),
	.w7(32'h3adb297a),
	.w8(32'h3c1ee1b2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2d09d),
	.w1(32'h3b3d1548),
	.w2(32'h3b68e51b),
	.w3(32'h3c16709a),
	.w4(32'h3abc1c89),
	.w5(32'hbaaa8483),
	.w6(32'h3aaef488),
	.w7(32'h3b898cbf),
	.w8(32'h3aa6a930),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25bbb4),
	.w1(32'hbbdc1ff7),
	.w2(32'hbbe38e54),
	.w3(32'hbb9201ad),
	.w4(32'hbc016725),
	.w5(32'h3c7abe19),
	.w6(32'hbb9c2e0c),
	.w7(32'hbbac0106),
	.w8(32'hbcb53cf1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb235b41),
	.w1(32'hbc6a4c96),
	.w2(32'h3aeb1976),
	.w3(32'h3b7d83c3),
	.w4(32'h3cacddc3),
	.w5(32'hbb886b38),
	.w6(32'hbbfac3ce),
	.w7(32'hbca72afb),
	.w8(32'hbb9947d1),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e68d3),
	.w1(32'hbb4cda7f),
	.w2(32'hbb00af82),
	.w3(32'hbb10f1e8),
	.w4(32'hbbda1f6a),
	.w5(32'h3b98f0ab),
	.w6(32'h3982aae9),
	.w7(32'hb91f3d83),
	.w8(32'hbb3dd86c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85aa3d),
	.w1(32'hbb804ee0),
	.w2(32'hbb2d2714),
	.w3(32'h3ba3a760),
	.w4(32'h3b5d2a98),
	.w5(32'hbb874ed9),
	.w6(32'h3adb9e33),
	.w7(32'hbba97d01),
	.w8(32'h399a2b87),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9072d9),
	.w1(32'hba8841d0),
	.w2(32'h3b9016d2),
	.w3(32'hbb35f904),
	.w4(32'hbb5218f3),
	.w5(32'hbbebde72),
	.w6(32'h3b991716),
	.w7(32'h3c04d969),
	.w8(32'h3b8d1fa1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c065edc),
	.w1(32'h39b2fc91),
	.w2(32'h3b2bf83d),
	.w3(32'hbbff4dbe),
	.w4(32'hbbccfa50),
	.w5(32'h3cc8870c),
	.w6(32'h3c2a426f),
	.w7(32'h3b4d9ef2),
	.w8(32'h3d28160b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ad0e7),
	.w1(32'h3ce210e8),
	.w2(32'h3ca257aa),
	.w3(32'h3ccaca17),
	.w4(32'h3b1a6f11),
	.w5(32'hbbe6d6c9),
	.w6(32'h3cb534b2),
	.w7(32'h3c03e3ab),
	.w8(32'h392da1a3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad02098),
	.w1(32'hbbc9949d),
	.w2(32'hbb62cfd0),
	.w3(32'hbb83c287),
	.w4(32'hbb30e33d),
	.w5(32'hbba13914),
	.w6(32'h3b98a22c),
	.w7(32'h3b098ab9),
	.w8(32'h3bd466ca),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10192e),
	.w1(32'h3c6c4763),
	.w2(32'hbb384dd7),
	.w3(32'hbc00d55d),
	.w4(32'hbb8beffc),
	.w5(32'hbc39260e),
	.w6(32'hbb5d328d),
	.w7(32'hbc071c46),
	.w8(32'hbb9f1e23),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d66fd),
	.w1(32'hbb010c44),
	.w2(32'hbbfaaea6),
	.w3(32'hbbab873b),
	.w4(32'hbbaea4f3),
	.w5(32'hbaf67596),
	.w6(32'hbbd2e0cc),
	.w7(32'hbb9f2353),
	.w8(32'h39bee735),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231bec),
	.w1(32'hbaaf4dcb),
	.w2(32'h3ac52493),
	.w3(32'hba4ea09c),
	.w4(32'h3b31cdd5),
	.w5(32'hbc04b5d5),
	.w6(32'hbb5b8b74),
	.w7(32'h3a6fa4e9),
	.w8(32'h3c396861),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04b87c),
	.w1(32'h3c1b6b4e),
	.w2(32'h3a5fe1a5),
	.w3(32'hbbc02b9e),
	.w4(32'hbc2dddf6),
	.w5(32'h39e38b26),
	.w6(32'h3cf164da),
	.w7(32'h3bb2481f),
	.w8(32'h3af09c47),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b988bf),
	.w1(32'h3a339d6f),
	.w2(32'hba38fda1),
	.w3(32'hbb400c81),
	.w4(32'h39586f68),
	.w5(32'hbb977340),
	.w6(32'h3af41d61),
	.w7(32'h3b3e851b),
	.w8(32'h3b836d0a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03d15e),
	.w1(32'hbc979ada),
	.w2(32'hbc1b920e),
	.w3(32'h39e4e6aa),
	.w4(32'hbb0164d4),
	.w5(32'hbbb31fac),
	.w6(32'h3c53b0be),
	.w7(32'h3b82f4c4),
	.w8(32'h3b23423e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb5b78),
	.w1(32'hbb0b7186),
	.w2(32'hbb4298fb),
	.w3(32'hbb228587),
	.w4(32'hbb0f3c84),
	.w5(32'hbb9b6b91),
	.w6(32'h3b4db5a5),
	.w7(32'h3aaa1f79),
	.w8(32'h3b7eb4bf),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb247bf3),
	.w1(32'hbb305ed3),
	.w2(32'hbba3b815),
	.w3(32'hbb3cfe10),
	.w4(32'hbb9cf264),
	.w5(32'hbc4a1967),
	.w6(32'h3b3a7bd9),
	.w7(32'h3ae1c7c7),
	.w8(32'hbc177a12),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cea6d),
	.w1(32'h391cced9),
	.w2(32'hbbb08472),
	.w3(32'hbc2796dd),
	.w4(32'hbb800aec),
	.w5(32'h3a1dd847),
	.w6(32'hbc181eda),
	.w7(32'hbb5ee6ce),
	.w8(32'h3b251c69),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59d4c5),
	.w1(32'hb983fc93),
	.w2(32'h389d7963),
	.w3(32'hba882fd0),
	.w4(32'hb9afa843),
	.w5(32'hbbb0526b),
	.w6(32'hbba69b9b),
	.w7(32'hbb3711cb),
	.w8(32'hba1498cc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8554d7),
	.w1(32'hbad5b9bd),
	.w2(32'hbb30bffe),
	.w3(32'hba7794fd),
	.w4(32'hba67067d),
	.w5(32'hbb28ce9d),
	.w6(32'h3b5bd251),
	.w7(32'h3b1e7645),
	.w8(32'h3b9a1a73),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dc9b5),
	.w1(32'hba99c84d),
	.w2(32'hb8814443),
	.w3(32'h3bc98b16),
	.w4(32'h3b8d315b),
	.w5(32'h3b280f58),
	.w6(32'h3bfa6a15),
	.w7(32'h3b911ae2),
	.w8(32'hbbb4a6b5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da5ba9),
	.w1(32'hba82aeea),
	.w2(32'h3b86e6bd),
	.w3(32'hbb28cd12),
	.w4(32'h3b65afa0),
	.w5(32'h3a20c8ea),
	.w6(32'hbb059015),
	.w7(32'hbad755ab),
	.w8(32'hbc766400),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5afe14),
	.w1(32'h3b466172),
	.w2(32'hba8a3a11),
	.w3(32'h3985b2ca),
	.w4(32'hb988771c),
	.w5(32'h3c84b0df),
	.w6(32'hbc3906b8),
	.w7(32'hbc405b8c),
	.w8(32'hbc00bba4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba04234),
	.w1(32'h3c584b4a),
	.w2(32'h3cafba38),
	.w3(32'h3c16b1de),
	.w4(32'hba87cba0),
	.w5(32'h3bcbdcca),
	.w6(32'h3b3f0c7e),
	.w7(32'hbb21cd57),
	.w8(32'h3b458f40),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5af903),
	.w1(32'h3a9212dd),
	.w2(32'h3b8e9183),
	.w3(32'h3b0d21c9),
	.w4(32'h3ae59fba),
	.w5(32'hbc1a4a4e),
	.w6(32'h3b342b5e),
	.w7(32'h3b82bb79),
	.w8(32'hbb79f402),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a7fda),
	.w1(32'hbb819069),
	.w2(32'hbb86bcdf),
	.w3(32'hbc3ce5cd),
	.w4(32'hbbed165d),
	.w5(32'hbb62a361),
	.w6(32'hbbeb4067),
	.w7(32'hbbfe1765),
	.w8(32'h3a7598f8),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaa54c),
	.w1(32'hba9ee2d6),
	.w2(32'h3ac7d1b1),
	.w3(32'hbb773588),
	.w4(32'h3b822ea7),
	.w5(32'hbb597be8),
	.w6(32'hbb12219b),
	.w7(32'hba90be7e),
	.w8(32'h3a1bd786),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b429),
	.w1(32'hbbb91734),
	.w2(32'hbbec3f62),
	.w3(32'hbb63b7fe),
	.w4(32'hba8c162d),
	.w5(32'h3b4b6a52),
	.w6(32'hba9d5eb7),
	.w7(32'hbb757cf7),
	.w8(32'hbb8a5bc4),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa291ed),
	.w1(32'h3b44aaac),
	.w2(32'h3b72451c),
	.w3(32'h3b062e44),
	.w4(32'hbab93e7e),
	.w5(32'hbc15d01a),
	.w6(32'hbbd56940),
	.w7(32'hb92d6f80),
	.w8(32'hbc31d59b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0d32f),
	.w1(32'hbc3e1a56),
	.w2(32'hbc609338),
	.w3(32'hbc276f28),
	.w4(32'hbc77ac87),
	.w5(32'hbbe76de3),
	.w6(32'hbbe83cd6),
	.w7(32'hbb6e1c66),
	.w8(32'hbb368713),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa85580),
	.w1(32'hb90a9e3b),
	.w2(32'h3abb9fd2),
	.w3(32'hbbc1433b),
	.w4(32'hbb26bcfd),
	.w5(32'hbb0c9e2e),
	.w6(32'h3ae35a19),
	.w7(32'h3b1bfc57),
	.w8(32'hbb2358a0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b2616),
	.w1(32'h3b17d03c),
	.w2(32'h399e3023),
	.w3(32'hbb81f7ab),
	.w4(32'hbaa69cce),
	.w5(32'hbcb1cf9f),
	.w6(32'hbbee51f0),
	.w7(32'h3ac42ed3),
	.w8(32'hbbba01ee),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad3f91),
	.w1(32'h3cc1c967),
	.w2(32'h3c53743d),
	.w3(32'hbc365d21),
	.w4(32'hbc3a9a3f),
	.w5(32'hbc21253f),
	.w6(32'h3b6d765a),
	.w7(32'h3c9b478e),
	.w8(32'h3bd2e24d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74ed80),
	.w1(32'hbb7c5fb4),
	.w2(32'hbb9fd6f0),
	.w3(32'hbb75edce),
	.w4(32'hbc422ed5),
	.w5(32'h3b916b60),
	.w6(32'h3b114b20),
	.w7(32'hbc027343),
	.w8(32'h3b5e3997),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeaccd),
	.w1(32'hbb45830a),
	.w2(32'hbc19197a),
	.w3(32'h3c68fd85),
	.w4(32'h3bfa687f),
	.w5(32'hbb0c4c21),
	.w6(32'h3d0ddb97),
	.w7(32'h3bc7136f),
	.w8(32'hbb236f24),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66700b),
	.w1(32'hbb99d0be),
	.w2(32'hbb82a4fd),
	.w3(32'hbbd74d3e),
	.w4(32'hbb352cf1),
	.w5(32'hbb92162f),
	.w6(32'hbb745d6f),
	.w7(32'hbbdb746a),
	.w8(32'hbbd8ff64),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1d1b3),
	.w1(32'hbb139a9f),
	.w2(32'h3b0190d1),
	.w3(32'hbb09d546),
	.w4(32'h3a0eb0bb),
	.w5(32'h39abc839),
	.w6(32'hbb57bd30),
	.w7(32'h3b4527b6),
	.w8(32'h3a5bd439),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae967eb),
	.w1(32'hb9082d27),
	.w2(32'h3a52d22c),
	.w3(32'h3a7d670f),
	.w4(32'hbaccff84),
	.w5(32'h3ce00853),
	.w6(32'hbbe17811),
	.w7(32'hbb7f7735),
	.w8(32'h3cae7261),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac52ce7),
	.w1(32'h3a93df2c),
	.w2(32'h3c8124ce),
	.w3(32'h3cedf813),
	.w4(32'h3bc3e897),
	.w5(32'hbc1833a1),
	.w6(32'h3ccf2867),
	.w7(32'h3cd6eff7),
	.w8(32'hbc25de4d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b01f2),
	.w1(32'hbb8ee9f9),
	.w2(32'hbaba8eb1),
	.w3(32'hbbfcafe9),
	.w4(32'hbbc6e66c),
	.w5(32'h3b240b29),
	.w6(32'hba2f4c38),
	.w7(32'h3a884e08),
	.w8(32'hb98bf4a4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4da8d1),
	.w1(32'h3b5ace1b),
	.w2(32'h3aa5847b),
	.w3(32'h3ba468ea),
	.w4(32'hbc077747),
	.w5(32'h3b4b5958),
	.w6(32'hbbe76dc2),
	.w7(32'hbbd71916),
	.w8(32'h3c18a8a9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3eda3),
	.w1(32'h3c67a1a4),
	.w2(32'h3c2e22f6),
	.w3(32'hbb0177ed),
	.w4(32'h3b913291),
	.w5(32'h3b3c07ca),
	.w6(32'h3c28cd44),
	.w7(32'hbb0057d8),
	.w8(32'h3b935e8f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c93c5),
	.w1(32'hbaa872a6),
	.w2(32'hbbb32ca4),
	.w3(32'h3b2fc42d),
	.w4(32'h3be92588),
	.w5(32'hbb7bbe12),
	.w6(32'hbc07e9ce),
	.w7(32'hbc0e07fa),
	.w8(32'hbae1e8dd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37da41),
	.w1(32'hbc0c87c8),
	.w2(32'hb9e5a2a3),
	.w3(32'hbbdcf6ff),
	.w4(32'hbbd4d3b7),
	.w5(32'hbc44d032),
	.w6(32'hb9935df1),
	.w7(32'hbb5dd0c7),
	.w8(32'hbc98abfe),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee4b2d),
	.w1(32'hbc84eefa),
	.w2(32'hbb219f47),
	.w3(32'hbc3b7b01),
	.w4(32'hbc279951),
	.w5(32'hbc2f165a),
	.w6(32'hbbe50d28),
	.w7(32'hbc123253),
	.w8(32'h3b48f22e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd1098),
	.w1(32'h3c60bdfe),
	.w2(32'hb7bd4397),
	.w3(32'hbb52da33),
	.w4(32'h3bae147d),
	.w5(32'h3b2193df),
	.w6(32'h3c78b32c),
	.w7(32'h3bda8877),
	.w8(32'hbb9941d0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd77426),
	.w1(32'h3b9bdb08),
	.w2(32'h3c24f700),
	.w3(32'h3bfdfed6),
	.w4(32'hbaa48417),
	.w5(32'hbbac133d),
	.w6(32'hbb52dc36),
	.w7(32'hbbaddba0),
	.w8(32'hbb2f5cb5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e53d98),
	.w1(32'hbbb37dea),
	.w2(32'hbb830c97),
	.w3(32'hbaeb9687),
	.w4(32'hbab59de1),
	.w5(32'hbad1c561),
	.w6(32'hbb319e40),
	.w7(32'hbafa9188),
	.w8(32'hbb4c57e0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc5f4d),
	.w1(32'hbb69f4aa),
	.w2(32'hbb222c15),
	.w3(32'h3bbf129f),
	.w4(32'h3badd471),
	.w5(32'hbad79d2b),
	.w6(32'h3bb5e16c),
	.w7(32'h3bc4938e),
	.w8(32'hbba24e2d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba060587),
	.w1(32'h3b09399a),
	.w2(32'h3b2b1533),
	.w3(32'hbbcd78ae),
	.w4(32'hba8fa540),
	.w5(32'hbbf1b097),
	.w6(32'hbc840852),
	.w7(32'h3b74f889),
	.w8(32'hbc1b1244),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c7789),
	.w1(32'hbb985ca4),
	.w2(32'h3ba92e49),
	.w3(32'hbbd10cf4),
	.w4(32'hb9d35eb0),
	.w5(32'hbc6ff89b),
	.w6(32'hbc3502d3),
	.w7(32'hba1a626e),
	.w8(32'hbc3e97a1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18c0f7),
	.w1(32'hbc128ac9),
	.w2(32'hbc2a0f2f),
	.w3(32'hbc17393b),
	.w4(32'hbb45c99d),
	.w5(32'hbb4f8cd7),
	.w6(32'hbb1a73e6),
	.w7(32'hbbf40b10),
	.w8(32'h3b55b83f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a3e0c),
	.w1(32'h3ad4d3a0),
	.w2(32'hbacc865f),
	.w3(32'hbbdc4db9),
	.w4(32'hbbb2b378),
	.w5(32'h3a168bd6),
	.w6(32'h3b3fa49e),
	.w7(32'h3c0cea9b),
	.w8(32'h3b86df1f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88b652),
	.w1(32'hbbcd9dfe),
	.w2(32'h3b9635ed),
	.w3(32'h3ac19319),
	.w4(32'h3b0d06fb),
	.w5(32'h3a07dbbe),
	.w6(32'h39d43c12),
	.w7(32'h3bc4759f),
	.w8(32'hbbf7a008),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b78d0),
	.w1(32'hbb2f8fab),
	.w2(32'hbbd8f9c2),
	.w3(32'h3b50afb7),
	.w4(32'h3be54006),
	.w5(32'hbc22cd6b),
	.w6(32'h3a27de82),
	.w7(32'h386d403c),
	.w8(32'hbbdae6a5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc02667),
	.w1(32'hbb1b5663),
	.w2(32'hbbd6392e),
	.w3(32'hbb2fb02f),
	.w4(32'hbb832533),
	.w5(32'h3aa8b44d),
	.w6(32'hbacd4db4),
	.w7(32'hbbc971ae),
	.w8(32'h3a993081),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace413b),
	.w1(32'hbaeb5f15),
	.w2(32'hbba404f7),
	.w3(32'hbb31a6d7),
	.w4(32'h3a0dd8d3),
	.w5(32'hb9347d0f),
	.w6(32'h3a8491b9),
	.w7(32'hbb285209),
	.w8(32'h3aa5b82f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e1279),
	.w1(32'h3ba82b18),
	.w2(32'h3bc724f2),
	.w3(32'h39cb036f),
	.w4(32'h3b9c8dbe),
	.w5(32'hba02ee7a),
	.w6(32'hbba7bb1c),
	.w7(32'h3a2d974e),
	.w8(32'hb9d43ce5),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b980dd0),
	.w1(32'h3b0b54f0),
	.w2(32'hba87ec4f),
	.w3(32'hba68d557),
	.w4(32'hbaf28226),
	.w5(32'hbbef1c55),
	.w6(32'h3ad17c3e),
	.w7(32'h3a2a760d),
	.w8(32'hbb4d2a4b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fad7d),
	.w1(32'hb9c292d1),
	.w2(32'h3ae880cc),
	.w3(32'hbbc80d66),
	.w4(32'hbb48a57b),
	.w5(32'hb9a0d543),
	.w6(32'hbbdbad78),
	.w7(32'hba96cf7a),
	.w8(32'h3aede4af),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8090b0),
	.w1(32'hbba95dec),
	.w2(32'h3c4ebb12),
	.w3(32'hbcaad490),
	.w4(32'hbc38c0c8),
	.w5(32'hbb4b243a),
	.w6(32'h39c6cb0c),
	.w7(32'hbbbae66c),
	.w8(32'h3b8aade3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba271cc),
	.w1(32'hbbe60cd2),
	.w2(32'hbb22c8eb),
	.w3(32'hba2d6c13),
	.w4(32'hbb21f625),
	.w5(32'h3bda0554),
	.w6(32'h3b9e9898),
	.w7(32'h3bbdf30d),
	.w8(32'hbcb2f5f8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4db5ac),
	.w1(32'hbc63871b),
	.w2(32'h3c28c58e),
	.w3(32'hbc5fae5d),
	.w4(32'hbb3d938e),
	.w5(32'hba82a033),
	.w6(32'hbccedf38),
	.w7(32'hbcb8e3cd),
	.w8(32'hbb02febb),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae89965),
	.w1(32'hbb2e027b),
	.w2(32'h3b073f99),
	.w3(32'hbbc3f7df),
	.w4(32'hbb968caa),
	.w5(32'hbbe0708d),
	.w6(32'hbbfbeea6),
	.w7(32'hbafae1ca),
	.w8(32'hbc694e75),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a949771),
	.w1(32'hbaf8182b),
	.w2(32'hbbdfe914),
	.w3(32'hbbeed148),
	.w4(32'hbbaa4959),
	.w5(32'hbb50de17),
	.w6(32'hbbc075a0),
	.w7(32'hbc18c687),
	.w8(32'hbbcfcddd),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb635870),
	.w1(32'hbc79f935),
	.w2(32'hbbe017d7),
	.w3(32'hba8704a9),
	.w4(32'hbba2a4b2),
	.w5(32'hbb79e488),
	.w6(32'h3bc673c0),
	.w7(32'h3b818227),
	.w8(32'hbc1b8ba8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb928bfd),
	.w1(32'hbbba09dc),
	.w2(32'h3a3eb10c),
	.w3(32'hbbcdc060),
	.w4(32'hbbaf0e05),
	.w5(32'hbb34162a),
	.w6(32'hbbff86bb),
	.w7(32'h3ad65d52),
	.w8(32'hbc160409),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d86ab),
	.w1(32'hbc1afc22),
	.w2(32'hba0912ae),
	.w3(32'hb982a5fe),
	.w4(32'hbaf1147b),
	.w5(32'hbbe5bdce),
	.w6(32'hbbdfd6a0),
	.w7(32'h3be177ad),
	.w8(32'h3adbd374),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44d41c),
	.w1(32'hbb04af1b),
	.w2(32'hba0e1bff),
	.w3(32'hbbecc452),
	.w4(32'hbb85ca42),
	.w5(32'h3a890d7b),
	.w6(32'hbbc1b093),
	.w7(32'hbb8c28bf),
	.w8(32'hbaece383),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec616f),
	.w1(32'hbb781030),
	.w2(32'hbbb03e5a),
	.w3(32'hbb27b2d2),
	.w4(32'hbb91caff),
	.w5(32'hbb8f0ce1),
	.w6(32'hbb04c925),
	.w7(32'hbb781145),
	.w8(32'hbb74b79b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc1273),
	.w1(32'hbbf7b375),
	.w2(32'hbae0d5ed),
	.w3(32'h3ae1e1d6),
	.w4(32'h3b057ba9),
	.w5(32'hbba256df),
	.w6(32'hb994791d),
	.w7(32'h3ad63fd2),
	.w8(32'hbb350f56),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc2dec),
	.w1(32'hbb3ca361),
	.w2(32'hbb13cc8e),
	.w3(32'hbc3c47b2),
	.w4(32'hbc1f4dc4),
	.w5(32'h3b93a197),
	.w6(32'hb9239e7f),
	.w7(32'hbb9d3985),
	.w8(32'hbcf08ec9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79423d),
	.w1(32'h3b1ccee9),
	.w2(32'h3ca81b5f),
	.w3(32'hba8e7ae6),
	.w4(32'h3bc45080),
	.w5(32'hbc80f535),
	.w6(32'hbc3754e1),
	.w7(32'hbcc145cf),
	.w8(32'hbc864a4c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc488e57),
	.w1(32'hbc8eb771),
	.w2(32'h3861994d),
	.w3(32'hbca1f6ba),
	.w4(32'hbc8715c5),
	.w5(32'hba049dec),
	.w6(32'hbc3a9485),
	.w7(32'h3b00d163),
	.w8(32'hbc7f2754),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90a167),
	.w1(32'hbc22faff),
	.w2(32'hbc17b4ad),
	.w3(32'hbbee780f),
	.w4(32'h3880368b),
	.w5(32'h3a224cc6),
	.w6(32'hbc8f2980),
	.w7(32'hbc95bfd1),
	.w8(32'hbc1c27fe),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53cb85),
	.w1(32'hba92d02a),
	.w2(32'h3c030ae0),
	.w3(32'h3b1062a2),
	.w4(32'h3a4c28c7),
	.w5(32'hbbaf6bf2),
	.w6(32'h3c0d84d1),
	.w7(32'hbc0d0193),
	.w8(32'hbb1e0ad3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab661b),
	.w1(32'hbb13e4b3),
	.w2(32'hbb468414),
	.w3(32'hba2bb6ba),
	.w4(32'h3aae2cb9),
	.w5(32'h3bab164e),
	.w6(32'h3bb1c8b1),
	.w7(32'h3b767f57),
	.w8(32'h3b44ac61),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a46b7),
	.w1(32'hbb1d0ce2),
	.w2(32'h3acf0f33),
	.w3(32'hbb623d77),
	.w4(32'h3b92e38c),
	.w5(32'hb9ea7e94),
	.w6(32'hbc098210),
	.w7(32'h3b09c433),
	.w8(32'h3b8f1475),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f20b7),
	.w1(32'hbc6d697b),
	.w2(32'hbc544d39),
	.w3(32'h3c418bb1),
	.w4(32'h3c0fa450),
	.w5(32'h3bea3d4c),
	.w6(32'hba188ee7),
	.w7(32'hbbecff90),
	.w8(32'hba7285bd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b151d6c),
	.w1(32'h3b113729),
	.w2(32'hbb1f4330),
	.w3(32'h3a9b6c39),
	.w4(32'h3bb86e93),
	.w5(32'hbbb2964e),
	.w6(32'hbc899cd6),
	.w7(32'h3b214d10),
	.w8(32'hbb7fe262),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b292c01),
	.w1(32'h3bd1d45e),
	.w2(32'h3be311a2),
	.w3(32'hbb98a1d5),
	.w4(32'hbba84469),
	.w5(32'hbb32c056),
	.w6(32'hbb87d178),
	.w7(32'h3ba9f4de),
	.w8(32'hbbfa21e7),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904d107),
	.w1(32'h3b91e670),
	.w2(32'hbb245b8b),
	.w3(32'hbbf59682),
	.w4(32'h3ae9acf9),
	.w5(32'hbb8beb15),
	.w6(32'h39b4d46a),
	.w7(32'hbb329c10),
	.w8(32'h3ba625ac),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cdf9c),
	.w1(32'hbae85cda),
	.w2(32'hbb1f8c60),
	.w3(32'hbc0cf010),
	.w4(32'hbb696f32),
	.w5(32'hbb0fd8c7),
	.w6(32'h3b2ae0c0),
	.w7(32'hbb041085),
	.w8(32'hbbd4dc22),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44176a),
	.w1(32'h3a0f68c3),
	.w2(32'h3bba8745),
	.w3(32'hbbe19285),
	.w4(32'hbb6d5bb1),
	.w5(32'hbb0f67d0),
	.w6(32'hba12dd9a),
	.w7(32'hba83113e),
	.w8(32'hbb1a2e85),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabebdbe),
	.w1(32'hbb34355b),
	.w2(32'h3a710932),
	.w3(32'hb916f4f1),
	.w4(32'hbab7959b),
	.w5(32'h3a8971a7),
	.w6(32'hba6b284a),
	.w7(32'h3ac1e610),
	.w8(32'h3b5bff02),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e99b3),
	.w1(32'h3b5d27c4),
	.w2(32'h395db47a),
	.w3(32'hb99286a7),
	.w4(32'h3a964a41),
	.w5(32'hbc88d439),
	.w6(32'h3b978f07),
	.w7(32'h3b97676a),
	.w8(32'h3aa0e6c8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f5aea),
	.w1(32'hbc51e982),
	.w2(32'hbcab6a8a),
	.w3(32'hbb759161),
	.w4(32'hbbcfe2d3),
	.w5(32'hbb538d80),
	.w6(32'h3ba51f95),
	.w7(32'hbb22d6ae),
	.w8(32'h3bb4ad8d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a264cde),
	.w1(32'h3b85c7f9),
	.w2(32'h3bd1f8b6),
	.w3(32'h3a0f599a),
	.w4(32'hb86244be),
	.w5(32'h3b5647aa),
	.w6(32'h3bbd883a),
	.w7(32'h3bd6e922),
	.w8(32'hb8940aae),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b004948),
	.w1(32'h38af7bf1),
	.w2(32'hbb9d8974),
	.w3(32'hbb73457b),
	.w4(32'h3b655c75),
	.w5(32'hbb9b4138),
	.w6(32'hbbe386a4),
	.w7(32'h3b16fa4e),
	.w8(32'h3aefbf49),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e6aa8),
	.w1(32'hba2aa012),
	.w2(32'h3a9d462b),
	.w3(32'hbabfea5c),
	.w4(32'hba9bc4ad),
	.w5(32'hbb86ff1f),
	.w6(32'h3b4964c0),
	.w7(32'h3b8a53e0),
	.w8(32'hbb3b74d1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b287e66),
	.w1(32'h3bdbda01),
	.w2(32'hbb3e4702),
	.w3(32'hbbb95562),
	.w4(32'hbb82d57a),
	.w5(32'hbb8c2a22),
	.w6(32'hbc35771e),
	.w7(32'hbb2c7be6),
	.w8(32'hbb1bd808),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40190d),
	.w1(32'hba287722),
	.w2(32'hbb70677d),
	.w3(32'hbb26b182),
	.w4(32'hbaab3ae4),
	.w5(32'h3b49a453),
	.w6(32'h3a70ea7d),
	.w7(32'hba8da27c),
	.w8(32'h3cbb5370),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c118a57),
	.w1(32'h3c347c11),
	.w2(32'hbc1493a9),
	.w3(32'h3d2bad65),
	.w4(32'h3cfb4da3),
	.w5(32'h3b16c83e),
	.w6(32'h3cf114d7),
	.w7(32'h3c22c47a),
	.w8(32'h3a6fc72d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe988d),
	.w1(32'hbb14a5a4),
	.w2(32'hbb3135f4),
	.w3(32'hba7cc485),
	.w4(32'h3aa3df13),
	.w5(32'hbb5f10c8),
	.w6(32'h3b136ec0),
	.w7(32'h3b806fd6),
	.w8(32'h3c0aebcd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f22f8),
	.w1(32'h3d0dcf1c),
	.w2(32'h3ca58f2e),
	.w3(32'h3bf80f2d),
	.w4(32'h3bd0a3ad),
	.w5(32'hbc2d7489),
	.w6(32'h3bbd9166),
	.w7(32'h3d033edf),
	.w8(32'h3aa58039),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab710f2),
	.w1(32'hbbb97728),
	.w2(32'hbbc0289a),
	.w3(32'h3b659879),
	.w4(32'hbbd02fa8),
	.w5(32'hbbc8ac71),
	.w6(32'h3c3eba0d),
	.w7(32'hba4cc893),
	.w8(32'hba6ce251),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf53a2c),
	.w1(32'hba510fe7),
	.w2(32'hbc1be962),
	.w3(32'hbb66bb54),
	.w4(32'hba1e162a),
	.w5(32'hbc0afdb1),
	.w6(32'h3b93e1bc),
	.w7(32'hbbb0969c),
	.w8(32'h3c889c83),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0d220),
	.w1(32'hbc3fff91),
	.w2(32'hbc725407),
	.w3(32'h3bf4dff4),
	.w4(32'hbb6c0c3e),
	.w5(32'hbb001780),
	.w6(32'h3cba7f10),
	.w7(32'h3c298d60),
	.w8(32'h3b51aaee),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ceadc),
	.w1(32'hbb3c7b2c),
	.w2(32'h3a9b8692),
	.w3(32'hbb021135),
	.w4(32'hbb0fb707),
	.w5(32'hbbf0306c),
	.w6(32'hbb0f7799),
	.w7(32'hbacd9688),
	.w8(32'h3b7c3b2c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371a7338),
	.w1(32'h3bba5ce8),
	.w2(32'h3a2a2570),
	.w3(32'hbbe60161),
	.w4(32'hbb141aea),
	.w5(32'h3b0e1567),
	.w6(32'h3b708dee),
	.w7(32'h3ad074f1),
	.w8(32'h3b9f4ec4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb474bc4),
	.w1(32'hbaec3930),
	.w2(32'hba43c219),
	.w3(32'hbb87b4dc),
	.w4(32'hbb647d2d),
	.w5(32'h3b02c9cc),
	.w6(32'h3b8ef3a5),
	.w7(32'hbb21df32),
	.w8(32'h385ff517),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3f5ab),
	.w1(32'hbc29b13c),
	.w2(32'hbbaf2ecb),
	.w3(32'hbb045505),
	.w4(32'hbc051ea8),
	.w5(32'hbb280204),
	.w6(32'h3b9b7b50),
	.w7(32'h3bb4a8cf),
	.w8(32'h3c09d425),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38fd98),
	.w1(32'h39a537f2),
	.w2(32'h3a27b480),
	.w3(32'hbba1e71d),
	.w4(32'hbadbab46),
	.w5(32'h3bd0178c),
	.w6(32'h3c2b87d0),
	.w7(32'hbb9e3a3e),
	.w8(32'h3b27b86a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01b156),
	.w1(32'hbb9ee8b5),
	.w2(32'hbacf880e),
	.w3(32'h3b0191d9),
	.w4(32'hba74689b),
	.w5(32'hbbc85705),
	.w6(32'h3bab7e52),
	.w7(32'h3b8f75ae),
	.w8(32'hbb087de0),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb628c),
	.w1(32'h3a38133f),
	.w2(32'hbb040020),
	.w3(32'hbb3d94ad),
	.w4(32'hbb092887),
	.w5(32'h3b823961),
	.w6(32'h3a1f5634),
	.w7(32'hb98f79dd),
	.w8(32'h3c411ab3),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6701f0),
	.w1(32'h3b854b6a),
	.w2(32'h3bc02235),
	.w3(32'hbb7eb50f),
	.w4(32'hbb55cdcd),
	.w5(32'h3b614de5),
	.w6(32'h3c675e44),
	.w7(32'h3c26d526),
	.w8(32'hb9971d12),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d5a70),
	.w1(32'h3b844506),
	.w2(32'h3b6cb2fd),
	.w3(32'hbb8808cf),
	.w4(32'hbb0bcbdc),
	.w5(32'h3c128577),
	.w6(32'hbbd35548),
	.w7(32'h3b97dead),
	.w8(32'h3a439f1c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57b87e),
	.w1(32'h3b42975f),
	.w2(32'hbaae13ba),
	.w3(32'h3b8df3f1),
	.w4(32'hbbba80c6),
	.w5(32'h3bbc06c4),
	.w6(32'hbbe97216),
	.w7(32'hbc13c201),
	.w8(32'h3b7d8344),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8476ee),
	.w1(32'h3b4be724),
	.w2(32'h3af74a67),
	.w3(32'h3ba81ae7),
	.w4(32'h3b86eda0),
	.w5(32'hbbbdf093),
	.w6(32'h3c394dc2),
	.w7(32'h3bb65cec),
	.w8(32'hbc427534),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c140f),
	.w1(32'hbbd1d206),
	.w2(32'hbc2f540b),
	.w3(32'hbc2dc49e),
	.w4(32'hbc51f5ad),
	.w5(32'hbc360976),
	.w6(32'hbc5e4e7c),
	.w7(32'hbbe81452),
	.w8(32'hbb97d4fd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5563),
	.w1(32'hbb76950f),
	.w2(32'hbb88038f),
	.w3(32'hbbfeeac4),
	.w4(32'hbbdb3bdc),
	.w5(32'hbc0ca825),
	.w6(32'hbbc3400c),
	.w7(32'hbb8d0e61),
	.w8(32'hbc2f4375),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b4ac9),
	.w1(32'h39a64214),
	.w2(32'hbad131d0),
	.w3(32'hbb8d823c),
	.w4(32'hbb6cfe6a),
	.w5(32'h392d322b),
	.w6(32'hbc277a5b),
	.w7(32'hbb9e5930),
	.w8(32'h39887cf6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a55195),
	.w1(32'hbb507398),
	.w2(32'hbb5e7797),
	.w3(32'hbb2553d5),
	.w4(32'h39b326d8),
	.w5(32'hbb788c7b),
	.w6(32'hb9cd704b),
	.w7(32'h3b172f1d),
	.w8(32'hbc631f8c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc534ea6),
	.w1(32'hbc8eedd3),
	.w2(32'hbc131b00),
	.w3(32'hbbed04dd),
	.w4(32'hbb1a4e54),
	.w5(32'hbb3cc9b6),
	.w6(32'hbc980292),
	.w7(32'hbc4af768),
	.w8(32'h3c25efd2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7a60f),
	.w1(32'h3b9ba1f6),
	.w2(32'h3b561c3e),
	.w3(32'hbba7ff26),
	.w4(32'hba6032d4),
	.w5(32'hbbac0269),
	.w6(32'h3c0f0e53),
	.w7(32'h3bc03c05),
	.w8(32'hbaf7e296),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa15196),
	.w1(32'h3a6e02d2),
	.w2(32'hbafb7c45),
	.w3(32'h3a0461ef),
	.w4(32'hba930523),
	.w5(32'hbb50a319),
	.w6(32'hbb5fa182),
	.w7(32'h3a31046f),
	.w8(32'hbba58ffb),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35b708),
	.w1(32'hbc245918),
	.w2(32'hba99ca35),
	.w3(32'hbb810590),
	.w4(32'h3b4e171f),
	.w5(32'hbb57932c),
	.w6(32'hbbceb9ee),
	.w7(32'hbba53e54),
	.w8(32'hbb15b01f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395957e9),
	.w1(32'h3b2722d0),
	.w2(32'hbb90a04a),
	.w3(32'hbae63db4),
	.w4(32'hbb89c7fd),
	.w5(32'h3bdf06ab),
	.w6(32'hb98dcd68),
	.w7(32'hbb589015),
	.w8(32'h3bb8ffc0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7f65),
	.w1(32'h3bd23653),
	.w2(32'h3c04318b),
	.w3(32'h3bbc17e0),
	.w4(32'h3c0660de),
	.w5(32'h3b8ac7ed),
	.w6(32'h3c659840),
	.w7(32'h3c2ae968),
	.w8(32'h3bbc33a4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3f390),
	.w1(32'h3b5b88a4),
	.w2(32'hb9b8d55a),
	.w3(32'h3ba98708),
	.w4(32'hbb5c74d4),
	.w5(32'hbbac5b8f),
	.w6(32'h3bc36225),
	.w7(32'hbb0a10ec),
	.w8(32'hbb171d6c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2247a9),
	.w1(32'h3b65a911),
	.w2(32'h3a631c36),
	.w3(32'hbb887b16),
	.w4(32'hb95e66f7),
	.w5(32'h3b46d95e),
	.w6(32'h3b91f667),
	.w7(32'h3ac12f26),
	.w8(32'hbad9d07b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa484c),
	.w1(32'hbb013cd7),
	.w2(32'hbbc6f4d0),
	.w3(32'hbb8057a9),
	.w4(32'hbb95b503),
	.w5(32'h3b871bec),
	.w6(32'hbb0a0d40),
	.w7(32'h39b3135d),
	.w8(32'h3bdd15b7),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be836e3),
	.w1(32'h3c30fc10),
	.w2(32'h3c0ec862),
	.w3(32'h3c0f62dc),
	.w4(32'h3ba0abc0),
	.w5(32'hbae98bed),
	.w6(32'h3c29b379),
	.w7(32'h3c2e756b),
	.w8(32'h3b2d4cc9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1234a),
	.w1(32'h3a5c2171),
	.w2(32'hbbb75af6),
	.w3(32'h3b803f8f),
	.w4(32'h3b71b66e),
	.w5(32'h3ad25c52),
	.w6(32'hbb0a1ec7),
	.w7(32'hba17d3c1),
	.w8(32'hbc0e1b04),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe52e8c),
	.w1(32'hbbc4133f),
	.w2(32'hba2e78b4),
	.w3(32'hba90a9ce),
	.w4(32'h39fad34e),
	.w5(32'h39a87917),
	.w6(32'hbb9b02c7),
	.w7(32'h3af450b0),
	.w8(32'hbb663b7d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973ea0),
	.w1(32'hbb771ba6),
	.w2(32'hbb9630e0),
	.w3(32'hbb5f9f09),
	.w4(32'hbb7324f6),
	.w5(32'h3b1c1fa3),
	.w6(32'hbb90d9b8),
	.w7(32'hbb035e5d),
	.w8(32'h3b35cdd5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba3236),
	.w1(32'h3be2916b),
	.w2(32'h3ba5b9ea),
	.w3(32'h3befebfc),
	.w4(32'h3bbdefea),
	.w5(32'hbc263426),
	.w6(32'h3c05c1a0),
	.w7(32'h3b9dbd5b),
	.w8(32'hbb823b14),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefb180),
	.w1(32'hbbc347b9),
	.w2(32'hbc2c64ff),
	.w3(32'hbc8bfde4),
	.w4(32'hbc28cb91),
	.w5(32'h3b40c447),
	.w6(32'hbc081ef2),
	.w7(32'hbc31b26d),
	.w8(32'h3b8b5f04),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11e866),
	.w1(32'h3b84fdec),
	.w2(32'h38e1d7e0),
	.w3(32'h3b07f388),
	.w4(32'h3b52d714),
	.w5(32'h3a0abb25),
	.w6(32'h3bae2bc3),
	.w7(32'h3bba44f1),
	.w8(32'hbbf7b1c1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca678a),
	.w1(32'h3b19d9f4),
	.w2(32'h3b156f9d),
	.w3(32'h3b94b47e),
	.w4(32'h3af8097d),
	.w5(32'hbab810cd),
	.w6(32'h3c897d6c),
	.w7(32'hbb7f2dd6),
	.w8(32'hbb9c0b09),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed154),
	.w1(32'hbc09270e),
	.w2(32'hbb9353ca),
	.w3(32'hbbfc49a5),
	.w4(32'hbbf48ffc),
	.w5(32'h3bcaaa70),
	.w6(32'hbba54dcc),
	.w7(32'hbb3174d6),
	.w8(32'h3bd416bc),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9abb7d),
	.w1(32'h3ba5d659),
	.w2(32'h3bd27fef),
	.w3(32'h3b7deb90),
	.w4(32'h3b57b63d),
	.w5(32'h3b83758e),
	.w6(32'h3be178b6),
	.w7(32'h3b928185),
	.w8(32'h3b6b5936),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b475e72),
	.w1(32'h3b55c1d2),
	.w2(32'hbb170daa),
	.w3(32'h3bec01c0),
	.w4(32'h3b0e359b),
	.w5(32'h3af660d3),
	.w6(32'hbaf2bff3),
	.w7(32'hbafdbf6e),
	.w8(32'h3a90b104),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05d349),
	.w1(32'h3bbcc74e),
	.w2(32'h3c0e45e2),
	.w3(32'h3b29d438),
	.w4(32'h39b54803),
	.w5(32'h387ce51e),
	.w6(32'hbb0b051d),
	.w7(32'h3b070c95),
	.w8(32'h3aa2a44b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acca10e),
	.w1(32'h3a2188c5),
	.w2(32'h3af7ea29),
	.w3(32'h397c210b),
	.w4(32'hba1314fe),
	.w5(32'hba5244c6),
	.w6(32'h3931da74),
	.w7(32'h3ad3ef08),
	.w8(32'hbb97cb5e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f244f),
	.w1(32'hbb8ccc3d),
	.w2(32'hbb17fa7a),
	.w3(32'h3b02a8b8),
	.w4(32'h3aeab1a1),
	.w5(32'h3b908127),
	.w6(32'hbbe165eb),
	.w7(32'hba1da044),
	.w8(32'h3b1c6e6c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b292f67),
	.w1(32'h3bda1c98),
	.w2(32'h3c06f3ec),
	.w3(32'h3b4e624e),
	.w4(32'h3ac8e13d),
	.w5(32'h3a7ff5d7),
	.w6(32'h3b74d7a1),
	.w7(32'hb9a9f796),
	.w8(32'hba65e2b1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c2327),
	.w1(32'hbbe757ab),
	.w2(32'hbbf7b4ed),
	.w3(32'hbb4e383d),
	.w4(32'h3a2cf9b4),
	.w5(32'h3b82b656),
	.w6(32'hbbad5f1f),
	.w7(32'h3ace1a23),
	.w8(32'h3c24900f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule