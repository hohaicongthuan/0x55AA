module layer_8_featuremap_252(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf2a61b),
	.w1(32'hbb5d704b),
	.w2(32'hbbd87bb6),
	.w3(32'h3c5b0b9b),
	.w4(32'hbaf156a9),
	.w5(32'hbaf773f8),
	.w6(32'hba702afa),
	.w7(32'hbb80f962),
	.w8(32'hbbc12a1c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0385d9),
	.w1(32'h3b826de0),
	.w2(32'hbbf4368e),
	.w3(32'h3bbdb144),
	.w4(32'h3bd26ad1),
	.w5(32'hbafb46ea),
	.w6(32'h3c20d8f5),
	.w7(32'h3b9d4c55),
	.w8(32'h3c06166f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc8c14),
	.w1(32'h3bf7c62e),
	.w2(32'h3bb80a02),
	.w3(32'h3a6977da),
	.w4(32'h3b22086e),
	.w5(32'h3bad653d),
	.w6(32'h3b87e029),
	.w7(32'h3bd8d850),
	.w8(32'h3bb4a536),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04b5f3),
	.w1(32'h3b9fab80),
	.w2(32'h3b8252ce),
	.w3(32'h3b99af28),
	.w4(32'h3c39a809),
	.w5(32'h3c6446a7),
	.w6(32'hbafd3191),
	.w7(32'h3b78f173),
	.w8(32'hba2c5a54),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4198af),
	.w1(32'hbac6b947),
	.w2(32'hbca3edf7),
	.w3(32'h3c815070),
	.w4(32'hba2a6b2c),
	.w5(32'hbc9123b6),
	.w6(32'h3bc72cdd),
	.w7(32'hbae409fe),
	.w8(32'hbb88fe01),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce144b4),
	.w1(32'h3b53c202),
	.w2(32'hbc80a356),
	.w3(32'hbcb74b4c),
	.w4(32'hbb63c007),
	.w5(32'hbc0b211c),
	.w6(32'h3b4b9778),
	.w7(32'hbb82f268),
	.w8(32'hbc4bd9e7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44213b),
	.w1(32'hbba8ac39),
	.w2(32'h3bad4fc7),
	.w3(32'hbbfe0f6d),
	.w4(32'hbbebeefa),
	.w5(32'h3b8f0429),
	.w6(32'hbc23903a),
	.w7(32'hbae6efda),
	.w8(32'h38e10fe7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc66fce),
	.w1(32'h3b59bd41),
	.w2(32'hbbdd3527),
	.w3(32'h3b9596c9),
	.w4(32'hbaadadfd),
	.w5(32'h3a14a4f7),
	.w6(32'h3b0e9418),
	.w7(32'hbb34a339),
	.w8(32'hbc1aeb0a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aef86),
	.w1(32'hbc5484a8),
	.w2(32'hbd0db1ef),
	.w3(32'h390db2ff),
	.w4(32'hbc659c20),
	.w5(32'hbd047083),
	.w6(32'hbbf6d595),
	.w7(32'hbc89c786),
	.w8(32'hbc34c478),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1302df),
	.w1(32'hb98f48c5),
	.w2(32'hbaec99c1),
	.w3(32'hbd067b24),
	.w4(32'hbb060327),
	.w5(32'hbc479b61),
	.w6(32'hbbd2e3f5),
	.w7(32'hbbff8e08),
	.w8(32'h3c280ddb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c271318),
	.w1(32'h3c11f619),
	.w2(32'h3bceeb5f),
	.w3(32'hbbff1458),
	.w4(32'h3b87c921),
	.w5(32'hbac82790),
	.w6(32'h3bcd6bc8),
	.w7(32'h3bd9b9aa),
	.w8(32'h3c014631),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab76845),
	.w1(32'h3a940cd5),
	.w2(32'h3c0c5530),
	.w3(32'h3bdc87a5),
	.w4(32'h3a9e7b28),
	.w5(32'h3c674412),
	.w6(32'hb9599588),
	.w7(32'h3a766bf7),
	.w8(32'h3c83c6cb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d018b01),
	.w1(32'hbb4d7066),
	.w2(32'hbb93d82c),
	.w3(32'h3d273929),
	.w4(32'hbbb35be9),
	.w5(32'hbc1e7b6b),
	.w6(32'hbbdd7a45),
	.w7(32'hbc05d254),
	.w8(32'hbbba6a40),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb945e75),
	.w1(32'h3b97424c),
	.w2(32'h3bf5c601),
	.w3(32'hbbf62da5),
	.w4(32'h3993d7b2),
	.w5(32'hbac88e0d),
	.w6(32'h3aa7d4e8),
	.w7(32'h3b77278d),
	.w8(32'hba0b5a6e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3dcb8),
	.w1(32'hbc327784),
	.w2(32'hbc7059f5),
	.w3(32'h3ae821fa),
	.w4(32'hbc3e88be),
	.w5(32'hbc6641ff),
	.w6(32'hbc6b24ef),
	.w7(32'hbc91496b),
	.w8(32'hbca13d8a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91cbe0),
	.w1(32'hbb465e92),
	.w2(32'hbbc53807),
	.w3(32'hbca960de),
	.w4(32'hbbb0f917),
	.w5(32'hbc4237e3),
	.w6(32'hbb7948a6),
	.w7(32'hbc0c3375),
	.w8(32'h3b8ee625),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fc50a),
	.w1(32'h3ac22001),
	.w2(32'hbbe338f4),
	.w3(32'hb7d983e3),
	.w4(32'hbc073cbe),
	.w5(32'hbb4c66ca),
	.w6(32'hbbcad69a),
	.w7(32'hbb566c63),
	.w8(32'hbb1ca33e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0475f7),
	.w1(32'h3c02145b),
	.w2(32'h3baf66cb),
	.w3(32'h3bf9111a),
	.w4(32'h3c282f3e),
	.w5(32'h3b15e819),
	.w6(32'h3bc817c4),
	.w7(32'h3b004218),
	.w8(32'h3a48ace8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f6f60),
	.w1(32'hbc7b22a7),
	.w2(32'hbcceb8be),
	.w3(32'h3ab6181e),
	.w4(32'hbc836942),
	.w5(32'hbcb763ff),
	.w6(32'hbc37411b),
	.w7(32'hbc692fed),
	.w8(32'hbc5eda75),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8669b1),
	.w1(32'hbc632e65),
	.w2(32'h3b108f22),
	.w3(32'hbc1ae18b),
	.w4(32'hbc7b4a09),
	.w5(32'hbb5ae5ac),
	.w6(32'hbc9be399),
	.w7(32'hbc3d6797),
	.w8(32'hbc27d4ac),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93f167),
	.w1(32'h3bce0819),
	.w2(32'h3ba97848),
	.w3(32'hbb09b1be),
	.w4(32'h3aa448cb),
	.w5(32'h3bcc4201),
	.w6(32'h3be2e0b6),
	.w7(32'hbb09056b),
	.w8(32'h3b3f6192),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b360002),
	.w1(32'h3b9c58fe),
	.w2(32'h3a179545),
	.w3(32'h3b83fe9f),
	.w4(32'h3b9102c3),
	.w5(32'hba812747),
	.w6(32'h3c11983c),
	.w7(32'h3a79037f),
	.w8(32'hbbb8651a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91f556),
	.w1(32'hbab7b657),
	.w2(32'hbc37d86c),
	.w3(32'h3b07d7c0),
	.w4(32'hbb1eb964),
	.w5(32'hbc205b06),
	.w6(32'h393f764f),
	.w7(32'hbb9bb155),
	.w8(32'hbc1918a5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d1970),
	.w1(32'h3bf678c9),
	.w2(32'h3aaa2f30),
	.w3(32'hbb40eeae),
	.w4(32'hbb407611),
	.w5(32'hbb2797a1),
	.w6(32'h3bac3b0c),
	.w7(32'hbb0534cd),
	.w8(32'hbb8dc779),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e26ae),
	.w1(32'hbc5511bb),
	.w2(32'hbb9c14ae),
	.w3(32'h3a8c1ff8),
	.w4(32'hbc484ffd),
	.w5(32'hbbee59ec),
	.w6(32'hbbb0ccef),
	.w7(32'h39e9d647),
	.w8(32'hba66edba),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc47052),
	.w1(32'h3b71412f),
	.w2(32'h3ba3882a),
	.w3(32'h3b893759),
	.w4(32'hbb44efe2),
	.w5(32'h3bdeb262),
	.w6(32'h3baa23b3),
	.w7(32'h3c1f74ca),
	.w8(32'h3bbffc5c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13a5d6),
	.w1(32'hbba1d5e4),
	.w2(32'hbbb88c4e),
	.w3(32'h3b5d2bbd),
	.w4(32'hbc098dfa),
	.w5(32'hbbb2c6ac),
	.w6(32'h3bac4940),
	.w7(32'h3b3ce84c),
	.w8(32'h3af5be9f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b6b1c),
	.w1(32'h3a89a9f3),
	.w2(32'h3b20942e),
	.w3(32'hbbdf878f),
	.w4(32'hbc15fca3),
	.w5(32'h39b6d569),
	.w6(32'hb9b871c8),
	.w7(32'hbb1299ad),
	.w8(32'hbb167c63),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ec025),
	.w1(32'h399cd3fe),
	.w2(32'hbc0f501b),
	.w3(32'hba38f448),
	.w4(32'hbb3cf231),
	.w5(32'hbbe33346),
	.w6(32'h3c0ad1f8),
	.w7(32'hbc300c3e),
	.w8(32'hb91185ac),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ccc27),
	.w1(32'hbb64749b),
	.w2(32'hbc0b684b),
	.w3(32'h3c67f72c),
	.w4(32'hbc27ad4e),
	.w5(32'hbc0e265f),
	.w6(32'hbbba01a0),
	.w7(32'hbbb2222b),
	.w8(32'hba89c95a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70eeecd),
	.w1(32'hba92eaff),
	.w2(32'h3c1d4211),
	.w3(32'h3abc2a73),
	.w4(32'hbb4fc7d9),
	.w5(32'h3bcfbe10),
	.w6(32'h3a5f982a),
	.w7(32'h3bb26487),
	.w8(32'h3c135880),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98c458),
	.w1(32'h3c31e825),
	.w2(32'h3b885fc7),
	.w3(32'h3c897d70),
	.w4(32'h3c1e8bcf),
	.w5(32'h3aeddc15),
	.w6(32'h3c50413b),
	.w7(32'h3bd9c5d2),
	.w8(32'h3b313def),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2390be),
	.w1(32'hbad3f735),
	.w2(32'hbb0a90b9),
	.w3(32'h3c0deec4),
	.w4(32'h3a571950),
	.w5(32'hba80c8fc),
	.w6(32'hba4ba0f9),
	.w7(32'hbb40b5e6),
	.w8(32'hbaecccbb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3dd26e),
	.w1(32'h390a4644),
	.w2(32'h3b4c9ed7),
	.w3(32'h3b6f8761),
	.w4(32'h3b2c5ab8),
	.w5(32'h3bc45fc2),
	.w6(32'hbb199f4c),
	.w7(32'h3bfb2e1a),
	.w8(32'h389284ca),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814c2c),
	.w1(32'h3ac6ef28),
	.w2(32'h3ba6bf24),
	.w3(32'hbaba181e),
	.w4(32'hbac1d841),
	.w5(32'h3c2ca829),
	.w6(32'hbb92fc5d),
	.w7(32'h3b43a1c9),
	.w8(32'h39feae3e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb655b03),
	.w1(32'hbaa3313e),
	.w2(32'h3b242472),
	.w3(32'h3c3d6ef0),
	.w4(32'h3af1da50),
	.w5(32'h3b5be73f),
	.w6(32'hbb878894),
	.w7(32'hbb0fcec7),
	.w8(32'hbbc0d5c0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399af2cb),
	.w1(32'h3c4edddc),
	.w2(32'h3bccdbe1),
	.w3(32'h3a8215ef),
	.w4(32'h3c9b6c1f),
	.w5(32'h3c93266f),
	.w6(32'h3c013251),
	.w7(32'hbb449390),
	.w8(32'hbc33fa1a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba3e88),
	.w1(32'h3bbc2ffb),
	.w2(32'hbc5d6b09),
	.w3(32'h3c0a4683),
	.w4(32'h3c1fcf5b),
	.w5(32'hbb8c501d),
	.w6(32'h3bdfdda8),
	.w7(32'hbacd150e),
	.w8(32'h3b808f56),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ea52f),
	.w1(32'h3ba422e4),
	.w2(32'h3a534027),
	.w3(32'hbb864ea1),
	.w4(32'h3a72017c),
	.w5(32'hbb48c760),
	.w6(32'h3b094e9e),
	.w7(32'hbbaa4a64),
	.w8(32'hba986b93),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0c2ac),
	.w1(32'h3976616a),
	.w2(32'h3b1319eb),
	.w3(32'hbb07a573),
	.w4(32'h3a992dbd),
	.w5(32'hba8e2c1f),
	.w6(32'h3a9df20f),
	.w7(32'h3a73afdf),
	.w8(32'h3a75961b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a588efc),
	.w1(32'h3bc7f117),
	.w2(32'h3c766406),
	.w3(32'h3bb0a107),
	.w4(32'h3bf28c6d),
	.w5(32'h3c9aaf20),
	.w6(32'h3c0493b0),
	.w7(32'h3c67d9b7),
	.w8(32'h3ca96a1d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb388c4),
	.w1(32'h3cbd0902),
	.w2(32'h3c725fed),
	.w3(32'h3cb9c3ac),
	.w4(32'h3cd94903),
	.w5(32'h3c96c5ec),
	.w6(32'h3c95315f),
	.w7(32'h3c4b9e1b),
	.w8(32'h3c32c934),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b27cc),
	.w1(32'hbc6dbc10),
	.w2(32'h3b181d56),
	.w3(32'h3c7406f8),
	.w4(32'hbc32ecdc),
	.w5(32'h3aaa2647),
	.w6(32'hbc8788fa),
	.w7(32'hbbd73f52),
	.w8(32'h3ba09dd6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6122b3),
	.w1(32'h3a100ec7),
	.w2(32'hbb8190d9),
	.w3(32'h3c1d6e2e),
	.w4(32'h3c198d9b),
	.w5(32'h3b70a7d5),
	.w6(32'h3a198b69),
	.w7(32'hbb99c07a),
	.w8(32'hbc072d00),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba176771),
	.w1(32'h3b875da8),
	.w2(32'hbba52a4a),
	.w3(32'hbb4e4499),
	.w4(32'hbb87416d),
	.w5(32'hbbefa9b6),
	.w6(32'hba97d398),
	.w7(32'hbbf308b1),
	.w8(32'hbb3b1007),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8c791),
	.w1(32'h3b353130),
	.w2(32'h3ca74aab),
	.w3(32'hbba154ac),
	.w4(32'h3a80cb15),
	.w5(32'h3c96f364),
	.w6(32'hbba703ec),
	.w7(32'h3bdf530c),
	.w8(32'h3c18107c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8a4ec),
	.w1(32'hbc149a3b),
	.w2(32'hba767ae1),
	.w3(32'h3c972e40),
	.w4(32'hbc447cd2),
	.w5(32'h3ab0b22a),
	.w6(32'hbbe615b1),
	.w7(32'hbb8c08d1),
	.w8(32'h3b6bcc6d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932a16),
	.w1(32'h3b6d0c8a),
	.w2(32'hb8e66f5c),
	.w3(32'h3b8fed23),
	.w4(32'hbb0f83f8),
	.w5(32'h3b664d39),
	.w6(32'h3b946ffc),
	.w7(32'h3b078705),
	.w8(32'hbad2a590),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad15b20),
	.w1(32'h3b64c812),
	.w2(32'h3a70cc69),
	.w3(32'h3c0f943a),
	.w4(32'hbb4d036e),
	.w5(32'hbba2c212),
	.w6(32'h3b9fc8c2),
	.w7(32'hba8da46b),
	.w8(32'hbbdc7130),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf42b0e),
	.w1(32'hbb81cffe),
	.w2(32'hbae6f044),
	.w3(32'h3a0f0c50),
	.w4(32'hbaaf79af),
	.w5(32'hbbace24c),
	.w6(32'hb9c2bab1),
	.w7(32'hbbc7fdac),
	.w8(32'hbc085ddf),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccb45a),
	.w1(32'hbc3a09ac),
	.w2(32'hbba6ad1f),
	.w3(32'hbc2a730e),
	.w4(32'hbb0f7c8f),
	.w5(32'h3b4de291),
	.w6(32'hbb2e0026),
	.w7(32'hba2f1499),
	.w8(32'hbb2ce569),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94bac8),
	.w1(32'hbc64c60c),
	.w2(32'hbcb1882c),
	.w3(32'hbbc4c6c9),
	.w4(32'hbc9879ea),
	.w5(32'hbca9d982),
	.w6(32'hbc09bf31),
	.w7(32'hbc867a9f),
	.w8(32'hbc511ad4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4ffe9),
	.w1(32'hb78b5c92),
	.w2(32'hbcd5993e),
	.w3(32'hbc580c31),
	.w4(32'hb98cfc57),
	.w5(32'hbcaac55c),
	.w6(32'h3bc43f50),
	.w7(32'hbbd705a1),
	.w8(32'hbc12ae70),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06db74),
	.w1(32'hbbf27b2f),
	.w2(32'hbc994b8a),
	.w3(32'hbcdf2366),
	.w4(32'hbc23cfeb),
	.w5(32'hbbfcef38),
	.w6(32'hbb3e0f53),
	.w7(32'hbc8bc7df),
	.w8(32'hbb9be560),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2dc14),
	.w1(32'h3b8c6703),
	.w2(32'h3c0fd110),
	.w3(32'h3b25d971),
	.w4(32'hbb685115),
	.w5(32'h3bf7ef58),
	.w6(32'h3b79edf7),
	.w7(32'h3ba90153),
	.w8(32'h3c0dbb42),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20fa06),
	.w1(32'h3bd8bcf6),
	.w2(32'h3b5ee3e0),
	.w3(32'h3c10f0bc),
	.w4(32'hba7c4454),
	.w5(32'hbb32ab9e),
	.w6(32'h3b113719),
	.w7(32'h3bae2d9a),
	.w8(32'hb954ed35),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af709bc),
	.w1(32'hbbc5d8b9),
	.w2(32'h3a117718),
	.w3(32'hbb871056),
	.w4(32'hbc2a2d0e),
	.w5(32'h3baa74d1),
	.w6(32'hbc029c1e),
	.w7(32'hbba4c702),
	.w8(32'hbc364056),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c948f),
	.w1(32'h3c47c8b7),
	.w2(32'h3bebbec3),
	.w3(32'h3a3ccaee),
	.w4(32'h3c504622),
	.w5(32'h3c375558),
	.w6(32'h3bbfb345),
	.w7(32'hbb95b951),
	.w8(32'hbc3a5dc8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcd561),
	.w1(32'hbb608e9f),
	.w2(32'h3bf279c6),
	.w3(32'h39e283c9),
	.w4(32'hbb5d69c3),
	.w5(32'h3c1e8659),
	.w6(32'hbb06bd4e),
	.w7(32'h3b7c9914),
	.w8(32'h3c4651b0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ea3fc),
	.w1(32'h3c007f39),
	.w2(32'h3bc6278d),
	.w3(32'h3c862f69),
	.w4(32'h3b717cdf),
	.w5(32'h3c1c17fc),
	.w6(32'hbaa44489),
	.w7(32'h3bb1f63d),
	.w8(32'h3af1ad28),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af232a9),
	.w1(32'hbba0ae70),
	.w2(32'hbbf3e0ab),
	.w3(32'h3af4aa00),
	.w4(32'hbba5938b),
	.w5(32'hbba18c51),
	.w6(32'h3be223e6),
	.w7(32'h3b96c68a),
	.w8(32'hbb1762f0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52e959),
	.w1(32'hbaa4bf47),
	.w2(32'hbc5f8919),
	.w3(32'hbc085da1),
	.w4(32'hbaee1419),
	.w5(32'h3c03cf69),
	.w6(32'hbc5a65ba),
	.w7(32'hbcb64d2e),
	.w8(32'hbd1ce257),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0caf6),
	.w1(32'h3c832cd1),
	.w2(32'h3bb5101b),
	.w3(32'h3ca4f697),
	.w4(32'h3c52c3d5),
	.w5(32'h3b9c229f),
	.w6(32'h3c564327),
	.w7(32'h3bbe2400),
	.w8(32'hbb02979a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bb03d),
	.w1(32'hbc8a2693),
	.w2(32'hbb089948),
	.w3(32'hba9ad040),
	.w4(32'hbc1ff0f5),
	.w5(32'h3c0801e4),
	.w6(32'hbc40b558),
	.w7(32'h3af9bd4a),
	.w8(32'h3c4290d3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c540558),
	.w1(32'hbb87c1d3),
	.w2(32'h3bb75841),
	.w3(32'h3cb4ac75),
	.w4(32'h3ae3408a),
	.w5(32'h3c4f3981),
	.w6(32'hbbc5ea5f),
	.w7(32'h3b2ac589),
	.w8(32'h3c592bab),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae2a0e),
	.w1(32'h3afccd3d),
	.w2(32'h3c64b675),
	.w3(32'h3ccf0a5f),
	.w4(32'h3919ef10),
	.w5(32'h3c653b3e),
	.w6(32'hba22dbca),
	.w7(32'h3b231429),
	.w8(32'h3bcb999e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c125d59),
	.w1(32'hbbf99b42),
	.w2(32'hbc69f5dc),
	.w3(32'h3bdf7db3),
	.w4(32'hba900598),
	.w5(32'hbb8e0d32),
	.w6(32'hbb9b2c10),
	.w7(32'hbbbbc149),
	.w8(32'h3bb70f47),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc2bea),
	.w1(32'h3aed8baf),
	.w2(32'h3a01adcf),
	.w3(32'h3b9e7709),
	.w4(32'h3a1dab6a),
	.w5(32'hbae2ff5a),
	.w6(32'h3ba351b0),
	.w7(32'h3bd7c043),
	.w8(32'h3a5e12bf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fb554),
	.w1(32'h3b1da1b4),
	.w2(32'hba71d5df),
	.w3(32'hbb13ccba),
	.w4(32'h3b3f5aa5),
	.w5(32'hbb5ab6aa),
	.w6(32'hbbb6fe73),
	.w7(32'h3b038e2d),
	.w8(32'hbb2ed9f8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b452f7a),
	.w1(32'h3bf12adf),
	.w2(32'h3b7906bd),
	.w3(32'hbab17529),
	.w4(32'hbaf74243),
	.w5(32'h3b061347),
	.w6(32'hba1fcc99),
	.w7(32'h3c0bda48),
	.w8(32'h3c2b94ad),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3803ff),
	.w1(32'hbd4053bf),
	.w2(32'hbd2e39f5),
	.w3(32'h3bee46a4),
	.w4(32'hbd40fd09),
	.w5(32'hbd26a03c),
	.w6(32'hbd1ad474),
	.w7(32'hbcbe07a8),
	.w8(32'h3bfcbc2d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0866d),
	.w1(32'h3b0d5cfb),
	.w2(32'h3a488d66),
	.w3(32'hbc164e4c),
	.w4(32'hbb2e9322),
	.w5(32'h3b01b3a2),
	.w6(32'hb81a63a4),
	.w7(32'hba8cd8e7),
	.w8(32'h3b5b6e93),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14a91f),
	.w1(32'hb9cef717),
	.w2(32'h3ad27399),
	.w3(32'h3bddd287),
	.w4(32'h3b47f367),
	.w5(32'h3ac04955),
	.w6(32'h3b4b1156),
	.w7(32'h3b9cfdf6),
	.w8(32'h3b30d2fe),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb5649),
	.w1(32'h3a595800),
	.w2(32'h3b6918de),
	.w3(32'h3aad8fc2),
	.w4(32'hb9c76a8a),
	.w5(32'hbc053115),
	.w6(32'hbad7382a),
	.w7(32'hb90c93fa),
	.w8(32'h3b856ae5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed930b),
	.w1(32'hbc475025),
	.w2(32'hbce59c93),
	.w3(32'h3a801463),
	.w4(32'hbcb2d1ec),
	.w5(32'hbd006822),
	.w6(32'hbc0c3209),
	.w7(32'hbc7b0332),
	.w8(32'hbca6f1af),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd843a9),
	.w1(32'h3a86eefe),
	.w2(32'hbb4b0dc0),
	.w3(32'hbc4e0c66),
	.w4(32'h3af82f8f),
	.w5(32'hbae75eeb),
	.w6(32'hbb237250),
	.w7(32'hbb3a25d3),
	.w8(32'hbbffa3f6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5d173),
	.w1(32'h390788d3),
	.w2(32'h3be8c3f7),
	.w3(32'hbbf2c974),
	.w4(32'hb9470188),
	.w5(32'h3ba7c7f9),
	.w6(32'hbb46747d),
	.w7(32'h3a9b240c),
	.w8(32'h3b846d1e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9a42),
	.w1(32'h3c41faa5),
	.w2(32'h3ca9d7f6),
	.w3(32'h3c1f6e68),
	.w4(32'h3c44b9a0),
	.w5(32'h3ca5f7e4),
	.w6(32'h3beed2a9),
	.w7(32'h3c0af239),
	.w8(32'hba938fd2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9802029),
	.w1(32'hbc227a4b),
	.w2(32'hbb9d07af),
	.w3(32'h3b4d2b40),
	.w4(32'hbbe1fac6),
	.w5(32'hbc28391b),
	.w6(32'hbb99abe5),
	.w7(32'hbbcec99a),
	.w8(32'h3ad51b94),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd15ba9),
	.w1(32'h3c1ab3a5),
	.w2(32'h3be59a9c),
	.w3(32'hbb6e8814),
	.w4(32'h3b206001),
	.w5(32'h3b136408),
	.w6(32'h3b338542),
	.w7(32'h3beeeb7e),
	.w8(32'h3bdb80a7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a933),
	.w1(32'h3b70cda4),
	.w2(32'h3c1ff4eb),
	.w3(32'h3a2581e5),
	.w4(32'h389a0ce3),
	.w5(32'h3b34ef45),
	.w6(32'h3baa48dc),
	.w7(32'h3c114ba0),
	.w8(32'h3b295fcf),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5857a1),
	.w1(32'h3b508978),
	.w2(32'h3bad112a),
	.w3(32'h3c142978),
	.w4(32'h3adcc8f1),
	.w5(32'hbb25458f),
	.w6(32'h3acb9f82),
	.w7(32'h3aed5c6c),
	.w8(32'h3a377f71),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b07a1),
	.w1(32'h39246ae4),
	.w2(32'hbb4b160a),
	.w3(32'hbbdce842),
	.w4(32'h3ae00581),
	.w5(32'h39d1c9f5),
	.w6(32'hba4e4f91),
	.w7(32'h3b2b3a08),
	.w8(32'h3b801581),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b763b),
	.w1(32'h3c0a38f2),
	.w2(32'h3b12226b),
	.w3(32'hb96702fb),
	.w4(32'h3b743b81),
	.w5(32'h3c2ee3d5),
	.w6(32'h3b2e2766),
	.w7(32'h3c2da6d7),
	.w8(32'h3bc6a627),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ea2a8),
	.w1(32'h3bc57a12),
	.w2(32'h3bdae653),
	.w3(32'h3bac7c23),
	.w4(32'hb92725b3),
	.w5(32'h3a0948fb),
	.w6(32'h3c0a2486),
	.w7(32'h3c6cd735),
	.w8(32'h3c162213),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0423f3),
	.w1(32'hbb59c70a),
	.w2(32'hbb325fc5),
	.w3(32'hb9ee62e4),
	.w4(32'h3ae72381),
	.w5(32'h3b58f28d),
	.w6(32'h3be6fb4b),
	.w7(32'h3be1862b),
	.w8(32'h3b2e9e83),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2df840),
	.w1(32'hbb120099),
	.w2(32'h3bad48c6),
	.w3(32'h3b2d2a07),
	.w4(32'hbc309ff5),
	.w5(32'hbc45589c),
	.w6(32'h3c0b6118),
	.w7(32'h3c7fc8ff),
	.w8(32'h3ca0b0a2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21e43a),
	.w1(32'h3bb674cc),
	.w2(32'h3c4fc609),
	.w3(32'hbca3a77b),
	.w4(32'h3bcf5be5),
	.w5(32'h3c28751a),
	.w6(32'h3b98237a),
	.w7(32'h3c145652),
	.w8(32'h3c286bd6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac6242),
	.w1(32'hbb9c30e5),
	.w2(32'h3b629df9),
	.w3(32'h3cc7ec7d),
	.w4(32'hbc6be93e),
	.w5(32'hbb3c51a2),
	.w6(32'h3c12db5b),
	.w7(32'h3c82bbb5),
	.w8(32'h3ca44e22),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c30e2),
	.w1(32'h3ba5b80e),
	.w2(32'h3bddebd5),
	.w3(32'hb98e7906),
	.w4(32'hbbba9eb3),
	.w5(32'hbb1b610b),
	.w6(32'h3aa96a3e),
	.w7(32'h3ae239f6),
	.w8(32'h3b2e482e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a547f56),
	.w1(32'hbb869041),
	.w2(32'hbbe353ef),
	.w3(32'h3bf85409),
	.w4(32'hba088ff8),
	.w5(32'h3b5727ba),
	.w6(32'h38de377c),
	.w7(32'hbbb6f29f),
	.w8(32'hbadbdf42),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92680f),
	.w1(32'hbbd8bbe9),
	.w2(32'h397d7a73),
	.w3(32'h3b1f0dfe),
	.w4(32'hbb70977a),
	.w5(32'h3b90e508),
	.w6(32'hbad0552a),
	.w7(32'h3ae80e3d),
	.w8(32'h3b7416c0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4878be),
	.w1(32'hbb2d2f8c),
	.w2(32'hbb1bfbe0),
	.w3(32'h3b6d5e1a),
	.w4(32'hbb4690c4),
	.w5(32'hba967ff2),
	.w6(32'hbba69c60),
	.w7(32'hbb5c86df),
	.w8(32'h3b8a7368),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb836c9),
	.w1(32'h38f63868),
	.w2(32'hbad3f37f),
	.w3(32'h3bc591ba),
	.w4(32'h3b3f610f),
	.w5(32'h3afa5194),
	.w6(32'h3ba72663),
	.w7(32'h3afca7b1),
	.w8(32'h3b98036b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1080f5),
	.w1(32'h3c44b1ea),
	.w2(32'h3c3d5b94),
	.w3(32'h3bc15d5e),
	.w4(32'h3c91d249),
	.w5(32'h3c3942dc),
	.w6(32'h3c3f0786),
	.w7(32'h3c578d08),
	.w8(32'h3c1f8664),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02629c),
	.w1(32'h3cc445a5),
	.w2(32'h3cae09d2),
	.w3(32'h3c863791),
	.w4(32'h3c4c7c08),
	.w5(32'h3bd84ba5),
	.w6(32'h3cc0250c),
	.w7(32'h3c9fdb4c),
	.w8(32'h3c1efe29),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be958ae),
	.w1(32'h3c0c38c4),
	.w2(32'h3c011c4d),
	.w3(32'hbb54d828),
	.w4(32'h3be8dc10),
	.w5(32'h3b871af8),
	.w6(32'hba323d3c),
	.w7(32'h3a8548d4),
	.w8(32'h3b0e55b5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0dbc4),
	.w1(32'h3aeffb37),
	.w2(32'h38cab6f2),
	.w3(32'h39998c2f),
	.w4(32'h3ac507e3),
	.w5(32'hba170cb6),
	.w6(32'hba20aef1),
	.w7(32'h3c0aa041),
	.w8(32'h3bddccde),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52f2e6),
	.w1(32'hbc11d7a9),
	.w2(32'hbc0bc092),
	.w3(32'hbb9c37b3),
	.w4(32'h3b0c4c20),
	.w5(32'hbc43f02a),
	.w6(32'hbaba83c8),
	.w7(32'hbc07ca18),
	.w8(32'hbb0b4515),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a5a70),
	.w1(32'hbc29adfb),
	.w2(32'h3bf2155e),
	.w3(32'hbc0eb6d7),
	.w4(32'hbc1d6d66),
	.w5(32'hbba3b5e9),
	.w6(32'hba624b96),
	.w7(32'hb98075b1),
	.w8(32'h3b053d46),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae174d6),
	.w1(32'h3b87671c),
	.w2(32'h3b18ac1b),
	.w3(32'hbbd2caf3),
	.w4(32'h3c2ec434),
	.w5(32'h3c1da939),
	.w6(32'h3bc749fa),
	.w7(32'h3bd2ae43),
	.w8(32'h3bb6627c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff22f3),
	.w1(32'hbb7215aa),
	.w2(32'hbbc6819f),
	.w3(32'hbb983a98),
	.w4(32'hba05eab4),
	.w5(32'hbbb0eca5),
	.w6(32'hbbb33ef4),
	.w7(32'hbc1a690b),
	.w8(32'hbbfd99ef),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6734f),
	.w1(32'h3ba13f9e),
	.w2(32'hbb45d94a),
	.w3(32'hbb9f98b1),
	.w4(32'hbaa1c162),
	.w5(32'hbc3d668f),
	.w6(32'h3b40b182),
	.w7(32'h3a916781),
	.w8(32'hbb8ab73e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb448dc5),
	.w1(32'hbb8885f3),
	.w2(32'h3b93396e),
	.w3(32'hbbcbd07c),
	.w4(32'hbbaedb88),
	.w5(32'h3a9bbbbd),
	.w6(32'hbae1ec1f),
	.w7(32'hba0c559c),
	.w8(32'h3b4807e0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b075f36),
	.w1(32'hbad6a6cf),
	.w2(32'h3b9e3755),
	.w3(32'hbaccebf7),
	.w4(32'hbaed483d),
	.w5(32'h3ade6878),
	.w6(32'h3b0367ad),
	.w7(32'h3b24ded2),
	.w8(32'hbb8392b6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf94d5),
	.w1(32'hbb0bbb72),
	.w2(32'h3aaa1dbd),
	.w3(32'hbbdf7076),
	.w4(32'hbbbcc78c),
	.w5(32'hbab7bea8),
	.w6(32'hbbbf8184),
	.w7(32'hbba48fe6),
	.w8(32'hbc0c91d9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eaf36),
	.w1(32'hbb09daec),
	.w2(32'h3c2c63c3),
	.w3(32'hbc218fa3),
	.w4(32'hbbf8da18),
	.w5(32'hbbde3267),
	.w6(32'h3b9846c3),
	.w7(32'h3c57920d),
	.w8(32'h3c8f3d6a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86935b),
	.w1(32'hbb6d3ee9),
	.w2(32'h3b2c66e4),
	.w3(32'hbc195521),
	.w4(32'h3998c587),
	.w5(32'h3c3e4600),
	.w6(32'hbb7dbccd),
	.w7(32'hbc205f88),
	.w8(32'hbc20457a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36deeba3),
	.w1(32'h3a5b3418),
	.w2(32'h3c083f5e),
	.w3(32'h3c38ec58),
	.w4(32'h3bc2d3c6),
	.w5(32'h3c41dfc7),
	.w6(32'h3b9a784c),
	.w7(32'h3bb18395),
	.w8(32'h3b90aac2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0b29c),
	.w1(32'h3c5009f0),
	.w2(32'h3a6bd213),
	.w3(32'h3ba02394),
	.w4(32'h3c6e6f3d),
	.w5(32'h3b39f398),
	.w6(32'h3c882425),
	.w7(32'h3c169144),
	.w8(32'h3bdc0bb0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73235c),
	.w1(32'hbb34f877),
	.w2(32'hbba1098f),
	.w3(32'hb9162093),
	.w4(32'h3a3b152f),
	.w5(32'hbacacf9f),
	.w6(32'hbb714eb7),
	.w7(32'h3b63f62e),
	.w8(32'hba94b59e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b1f3a),
	.w1(32'h3bb5148f),
	.w2(32'h3cebf74a),
	.w3(32'hba53acc9),
	.w4(32'h3c1d05f0),
	.w5(32'h3d052ae4),
	.w6(32'h3b04afba),
	.w7(32'h3c8b1558),
	.w8(32'h3cded70a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3b77a8),
	.w1(32'hbb670c47),
	.w2(32'hbc207cf7),
	.w3(32'h3d48e4f1),
	.w4(32'hbbb6ac15),
	.w5(32'hbbdfde01),
	.w6(32'hbaeaeec4),
	.w7(32'hbb6ea848),
	.w8(32'hbc056f57),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf1244),
	.w1(32'h3bcf093b),
	.w2(32'h3bf014d7),
	.w3(32'hbc02f56b),
	.w4(32'h3a8b15ec),
	.w5(32'h3c19b8e1),
	.w6(32'h3b82471e),
	.w7(32'h3a909e7a),
	.w8(32'hb910bcad),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfab56c),
	.w1(32'hbc4518ea),
	.w2(32'hbb9a891a),
	.w3(32'h3c2cf7ca),
	.w4(32'hbc3dca05),
	.w5(32'hbb675e89),
	.w6(32'hbbf5b003),
	.w7(32'hbb2474d9),
	.w8(32'h3b9fa636),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ce18b),
	.w1(32'h3c17aafb),
	.w2(32'hba73ccc9),
	.w3(32'hb9956dfc),
	.w4(32'h3c49dd85),
	.w5(32'h3b4a58e0),
	.w6(32'h3c4ea0f9),
	.w7(32'h3bde9ba9),
	.w8(32'h3bd98374),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba731672),
	.w1(32'hbbf77110),
	.w2(32'hbc2f5f4c),
	.w3(32'h3b667a2b),
	.w4(32'hbb503302),
	.w5(32'hbc59e24e),
	.w6(32'hbb742bfa),
	.w7(32'hbbded1a3),
	.w8(32'hbc1a812f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e1713),
	.w1(32'hbc438671),
	.w2(32'hbbddb6fa),
	.w3(32'hbcdbd75a),
	.w4(32'hbb628266),
	.w5(32'hbc29c396),
	.w6(32'hbc0f3cee),
	.w7(32'hbb1a9686),
	.w8(32'hba3a4a86),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe809dc),
	.w1(32'h3a52a70c),
	.w2(32'hb9607ebc),
	.w3(32'hbc33770f),
	.w4(32'h3c110d04),
	.w5(32'hba0daf8f),
	.w6(32'h3ac6a15d),
	.w7(32'h3b9e680a),
	.w8(32'hbb0e153b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caf36a),
	.w1(32'h3b431c89),
	.w2(32'hbc5efa84),
	.w3(32'h3b12b474),
	.w4(32'h36610181),
	.w5(32'hbc90d672),
	.w6(32'h3c2644a8),
	.w7(32'hba3c3fba),
	.w8(32'hbba4a2cf),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51dea7),
	.w1(32'h3b51af26),
	.w2(32'h3ab7e9bc),
	.w3(32'hbc7fa159),
	.w4(32'h3c0dbac5),
	.w5(32'h3b033ae3),
	.w6(32'h3b99a9c0),
	.w7(32'h398cea1b),
	.w8(32'hb95b0951),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c99cd),
	.w1(32'hbc474b2b),
	.w2(32'hbbb90e76),
	.w3(32'hbbd91c0e),
	.w4(32'hbbc7962a),
	.w5(32'hbbc5b5dc),
	.w6(32'hbc36ca2a),
	.w7(32'hbbdacbe6),
	.w8(32'h398a63a4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef549d),
	.w1(32'hbcac0b78),
	.w2(32'hbc8fc0bf),
	.w3(32'h3c0295e1),
	.w4(32'hbc66b5cd),
	.w5(32'hbc3c93be),
	.w6(32'hbc6d246f),
	.w7(32'hbc3d9d2a),
	.w8(32'hbb2788a3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00be6d),
	.w1(32'hbb2b427a),
	.w2(32'hbbad33f0),
	.w3(32'hbade0871),
	.w4(32'h3bba059b),
	.w5(32'hbbb4a1da),
	.w6(32'hba8100f2),
	.w7(32'hbb41295d),
	.w8(32'hbb8d6944),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc131aa8),
	.w1(32'h3be810fd),
	.w2(32'h39a6143d),
	.w3(32'hbc454f76),
	.w4(32'h3bbb5704),
	.w5(32'h3be6fc08),
	.w6(32'h3b9ae225),
	.w7(32'h3a76ad5a),
	.w8(32'hbaa3d072),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf73faa),
	.w1(32'h3ab917af),
	.w2(32'hbb38548f),
	.w3(32'h3ba4fce7),
	.w4(32'h3ba84ec0),
	.w5(32'hba9c7aba),
	.w6(32'h3a16d760),
	.w7(32'hba6d3a7e),
	.w8(32'hbbe531a0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb674e2f),
	.w1(32'hbae99a7a),
	.w2(32'h3a0dda84),
	.w3(32'hbb0ed280),
	.w4(32'h39a0184c),
	.w5(32'hba4da50e),
	.w6(32'h39a7d17a),
	.w7(32'hbaadc193),
	.w8(32'h3a85cc4e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3c924),
	.w1(32'hbc027a1d),
	.w2(32'h3ac2814d),
	.w3(32'h399d598c),
	.w4(32'hbc527c2b),
	.w5(32'hbb54ff23),
	.w6(32'hbade40ba),
	.w7(32'hbb164f65),
	.w8(32'hbbb083b2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule