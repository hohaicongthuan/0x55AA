module layer_8_featuremap_68(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c2040),
	.w1(32'hbb9bdd1c),
	.w2(32'h3bfdb84d),
	.w3(32'hbc2f4e4d),
	.w4(32'hbc1a73a8),
	.w5(32'hbb10d639),
	.w6(32'hbb0b9f0f),
	.w7(32'hbbc79900),
	.w8(32'hbbf6596e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb8931),
	.w1(32'h3bc62780),
	.w2(32'h3b86a9dd),
	.w3(32'h3c074e50),
	.w4(32'h3b805d14),
	.w5(32'hb8867686),
	.w6(32'h3ba6c521),
	.w7(32'h3add6d42),
	.w8(32'hba9e2382),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44520e),
	.w1(32'hbb7b92c2),
	.w2(32'hbb11b8a9),
	.w3(32'hba39b718),
	.w4(32'hbb339780),
	.w5(32'hbb4dd27a),
	.w6(32'hbadd7061),
	.w7(32'hbb31c860),
	.w8(32'hbbca4f3a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08c553),
	.w1(32'hbb9443d9),
	.w2(32'hba95ddda),
	.w3(32'h3864330d),
	.w4(32'h3b29af40),
	.w5(32'h3b185485),
	.w6(32'hb907f4d2),
	.w7(32'hbba9e860),
	.w8(32'h3a88e3b8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeafa9),
	.w1(32'h3b5e0f4a),
	.w2(32'h3b0df0dd),
	.w3(32'h3b389a8d),
	.w4(32'hbacccea0),
	.w5(32'hbb36ed26),
	.w6(32'h3b6ef5d4),
	.w7(32'hbaaf9716),
	.w8(32'h38dfc6a6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd38518),
	.w1(32'h3bba8e27),
	.w2(32'h3abd923e),
	.w3(32'h3b9232e7),
	.w4(32'h39843dea),
	.w5(32'h3a97a7a3),
	.w6(32'hbb1b70d3),
	.w7(32'hba931d7c),
	.w8(32'h3bc16729),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a104d84),
	.w1(32'h3a70af04),
	.w2(32'h3a2f8c95),
	.w3(32'h39a53854),
	.w4(32'h3a3b53e1),
	.w5(32'h3a359e96),
	.w6(32'h3a3f7675),
	.w7(32'h39767736),
	.w8(32'hb9295ecc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dde99),
	.w1(32'h3b1ae107),
	.w2(32'h3bb80c91),
	.w3(32'hbba43911),
	.w4(32'hbb16ded9),
	.w5(32'h3a8fc083),
	.w6(32'hbb3de954),
	.w7(32'hbbe6174f),
	.w8(32'hbbc3b297),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cc77c),
	.w1(32'hb80eb61b),
	.w2(32'h37551e01),
	.w3(32'h39c37c08),
	.w4(32'hbb8c85de),
	.w5(32'hbbdaa94c),
	.w6(32'hba1ba695),
	.w7(32'hbb88b32e),
	.w8(32'hbbe6ccc4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf44f1),
	.w1(32'h3b879bea),
	.w2(32'h3c32b884),
	.w3(32'h3b082b79),
	.w4(32'hbb3ba2e2),
	.w5(32'hba39e0db),
	.w6(32'hbb6bcd16),
	.w7(32'hbb43e3b8),
	.w8(32'hbbc8ed5e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8f949),
	.w1(32'hbb2db59c),
	.w2(32'h3b3af4d4),
	.w3(32'hbc2bb97b),
	.w4(32'hbbca2eb8),
	.w5(32'h3a49e23f),
	.w6(32'h3a3caa33),
	.w7(32'hbbd34065),
	.w8(32'hbbaddbb9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f7680),
	.w1(32'hb96882a4),
	.w2(32'h3bd18b81),
	.w3(32'hb854f888),
	.w4(32'hbb74c19c),
	.w5(32'h3af16e20),
	.w6(32'h3b3ad95c),
	.w7(32'hbbd733f2),
	.w8(32'hbc2189a7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b806693),
	.w1(32'h3b4da81b),
	.w2(32'h3b4ee27c),
	.w3(32'h3b3b31ec),
	.w4(32'hba6b3979),
	.w5(32'hbb5441eb),
	.w6(32'h3a9100f5),
	.w7(32'hb793751a),
	.w8(32'h3b072bf6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31a23b),
	.w1(32'h3ac60b88),
	.w2(32'h3a7bb798),
	.w3(32'h3b413272),
	.w4(32'h3ad8610a),
	.w5(32'h39a74d9e),
	.w6(32'h3adbd2db),
	.w7(32'h3a959fcf),
	.w8(32'hb9d9ce37),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbf374),
	.w1(32'h3ac0e2e0),
	.w2(32'h3a843797),
	.w3(32'h3ac629fa),
	.w4(32'h3aaebc36),
	.w5(32'h3a1ef9ed),
	.w6(32'h3a8d9338),
	.w7(32'h3a6126ff),
	.w8(32'hba17900c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070b06),
	.w1(32'hbab73d48),
	.w2(32'hbac9ce50),
	.w3(32'hbab9edf4),
	.w4(32'hba82c4fe),
	.w5(32'hba746c30),
	.w6(32'hbaa49f03),
	.w7(32'hba7c8200),
	.w8(32'hbaa6b360),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84fe31),
	.w1(32'hbbb2caef),
	.w2(32'hbbad169e),
	.w3(32'hbb867828),
	.w4(32'hbba9ba40),
	.w5(32'hbb7a179a),
	.w6(32'hbb3f66a6),
	.w7(32'hbae60e2a),
	.w8(32'h3a1728ff),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a9e89),
	.w1(32'h3b42a315),
	.w2(32'h3c13867e),
	.w3(32'h3a0d3730),
	.w4(32'hbb2028b9),
	.w5(32'hbb107553),
	.w6(32'h3b81e686),
	.w7(32'hbae71805),
	.w8(32'hbbed1c48),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8d3f8),
	.w1(32'hbbe35ce4),
	.w2(32'h3d2f86c1),
	.w3(32'hbca072af),
	.w4(32'h3c300917),
	.w5(32'h3d341efd),
	.w6(32'h3c691f8c),
	.w7(32'hbc74c525),
	.w8(32'hbc3983bd),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5e4c1),
	.w1(32'h3bb9d16e),
	.w2(32'h3c65c718),
	.w3(32'hbb8f4daa),
	.w4(32'hbc3c820e),
	.w5(32'hbb5208b9),
	.w6(32'h3aa169b1),
	.w7(32'h3b5fd6b5),
	.w8(32'h3c1bb40a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed09aa),
	.w1(32'hb97d2849),
	.w2(32'hbb71fe42),
	.w3(32'hbb0036f7),
	.w4(32'hbc01afbd),
	.w5(32'hbbad8f0d),
	.w6(32'hb9d520a1),
	.w7(32'hb98b222b),
	.w8(32'hbb206e2a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c074469),
	.w1(32'h3b86a8b5),
	.w2(32'hba13cb58),
	.w3(32'h3c12eb30),
	.w4(32'h3b58f88d),
	.w5(32'hbae57744),
	.w6(32'h3b9c847e),
	.w7(32'hbad28de7),
	.w8(32'hbbb9cc6c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85fa3c),
	.w1(32'hbc355d5f),
	.w2(32'h3c696d22),
	.w3(32'hbd1893cb),
	.w4(32'hbcae7638),
	.w5(32'h3ba91cf2),
	.w6(32'h3964af9e),
	.w7(32'hbc2fa537),
	.w8(32'hbc9ad900),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83e4e3),
	.w1(32'h3b7043d7),
	.w2(32'h3b3fb378),
	.w3(32'h38e0ba9d),
	.w4(32'hbb76045c),
	.w5(32'hbba6c81f),
	.w6(32'hbb85968c),
	.w7(32'hba914590),
	.w8(32'hba89c279),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7fd37),
	.w1(32'hbb44ca4f),
	.w2(32'hbb995669),
	.w3(32'hbbc22871),
	.w4(32'hbb904250),
	.w5(32'hbb7dd3f1),
	.w6(32'hbc0a64c9),
	.w7(32'hbb35c047),
	.w8(32'hbba1921c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb385611),
	.w1(32'hbb2c4678),
	.w2(32'h3c22936b),
	.w3(32'hbbcea630),
	.w4(32'hbb855345),
	.w5(32'h3c2befaa),
	.w6(32'h3b8d6981),
	.w7(32'hbb7e56c1),
	.w8(32'hbb912ca5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a20cf),
	.w1(32'hba89dbd9),
	.w2(32'h39163cd1),
	.w3(32'h3a353ba7),
	.w4(32'hba394851),
	.w5(32'h3855ed35),
	.w6(32'h3a9f517a),
	.w7(32'h3aa7ee65),
	.w8(32'h3a8ccea7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8ab5b),
	.w1(32'hbceb8c77),
	.w2(32'h3d010ba1),
	.w3(32'hbd9e7452),
	.w4(32'hbcb9702e),
	.w5(32'h3e0d8f3d),
	.w6(32'h3dcefb25),
	.w7(32'h3d7ee7e4),
	.w8(32'h3ce6fd23),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e1830),
	.w1(32'hbad341be),
	.w2(32'h3bf1be00),
	.w3(32'hbb2ae121),
	.w4(32'hbb64a97d),
	.w5(32'h3b1e4c9a),
	.w6(32'h3b47ac26),
	.w7(32'h3ad94cb5),
	.w8(32'h39703a96),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f11b2d),
	.w1(32'h3a18f166),
	.w2(32'hba0506e7),
	.w3(32'hba118ec5),
	.w4(32'hbac6b833),
	.w5(32'hbb3309f9),
	.w6(32'hba8d2798),
	.w7(32'hbb0cf9f8),
	.w8(32'hbb024d68),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb50711),
	.w1(32'h3b40a71d),
	.w2(32'h3ba6813d),
	.w3(32'h3c01de15),
	.w4(32'h3be31065),
	.w5(32'h3befccfa),
	.w6(32'h3bc17120),
	.w7(32'h3c00d59a),
	.w8(32'h3bc67f47),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bc0b4),
	.w1(32'h3a4b0a46),
	.w2(32'hb83c15dc),
	.w3(32'hba767838),
	.w4(32'hbb2b4274),
	.w5(32'hbab4c7ca),
	.w6(32'h3a2669ec),
	.w7(32'h3ae1a913),
	.w8(32'h3b710ea9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392383f0),
	.w1(32'hbb24edca),
	.w2(32'hbae6b92d),
	.w3(32'h3ab15bcc),
	.w4(32'hbabb4dbe),
	.w5(32'hbb20c462),
	.w6(32'h3aa8bce3),
	.w7(32'h3aabb1a9),
	.w8(32'h3aa5f66f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ccb219),
	.w1(32'hbb1c5d0e),
	.w2(32'hba70dc46),
	.w3(32'h37c366d2),
	.w4(32'hba929bd0),
	.w5(32'hba88d4ff),
	.w6(32'h3afa0723),
	.w7(32'h3b095b80),
	.w8(32'h3b3163ec),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5329ad),
	.w1(32'h3c4a259f),
	.w2(32'h3c184819),
	.w3(32'h3c32793e),
	.w4(32'h3bb7f9b9),
	.w5(32'h3a18b03a),
	.w6(32'h3b75f943),
	.w7(32'h3b947f69),
	.w8(32'h3b2899e5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa249f2),
	.w1(32'hbac291d9),
	.w2(32'h3c5280a1),
	.w3(32'h3ad5037d),
	.w4(32'h3bad2a1f),
	.w5(32'h3c81191d),
	.w6(32'h3c5be968),
	.w7(32'h3bfe0459),
	.w8(32'h3b0d370d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39b799),
	.w1(32'hbb4ef4cd),
	.w2(32'hbb10b22b),
	.w3(32'hbae3d727),
	.w4(32'hbb4c382d),
	.w5(32'hbb2ec810),
	.w6(32'hbace6532),
	.w7(32'hba4fd028),
	.w8(32'hba2d5a07),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf1b86),
	.w1(32'h3b4f1b48),
	.w2(32'h392eb2e6),
	.w3(32'h3b9f48ff),
	.w4(32'h3b07434b),
	.w5(32'hbaf09bcd),
	.w6(32'h3b92f72c),
	.w7(32'h3ac02b9f),
	.w8(32'h3a085aef),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b223470),
	.w1(32'h3b1a80f7),
	.w2(32'h3abb5f94),
	.w3(32'h3b278a44),
	.w4(32'h3b06499c),
	.w5(32'h3a628ee8),
	.w6(32'h3ad87585),
	.w7(32'h3ab0028b),
	.w8(32'h3926a0a1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4dbbe7),
	.w1(32'hba810c5f),
	.w2(32'hba594649),
	.w3(32'hbaf94078),
	.w4(32'hba5b45b1),
	.w5(32'h39e52d6e),
	.w6(32'hbb222472),
	.w7(32'hba927f4c),
	.w8(32'hb9d00c2a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc700f49),
	.w1(32'hbbd776e3),
	.w2(32'h3c82f709),
	.w3(32'hbb8e903c),
	.w4(32'hbbc5adfd),
	.w5(32'h3ba7dc37),
	.w6(32'h3c16aa18),
	.w7(32'hbbe73310),
	.w8(32'hbc0215e9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb457af1),
	.w1(32'h384f2aec),
	.w2(32'h3bc614fc),
	.w3(32'hbadafb6e),
	.w4(32'h3a7909fe),
	.w5(32'h3ba81280),
	.w6(32'h3aecbc7c),
	.w7(32'hbac75395),
	.w8(32'h3b143cd8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a970526),
	.w1(32'hb848dfb4),
	.w2(32'hbab1dc07),
	.w3(32'h39dbc857),
	.w4(32'h39d6b1c7),
	.w5(32'hba2fcaf5),
	.w6(32'hb7e7d1c6),
	.w7(32'hba9cf5fe),
	.w8(32'hbaa996f1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba98358),
	.w1(32'hbbdc55e6),
	.w2(32'hba90deb1),
	.w3(32'hbc07afc0),
	.w4(32'hbba81c50),
	.w5(32'h3b07535c),
	.w6(32'h398c5a7a),
	.w7(32'hbb74121c),
	.w8(32'hbad9590f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7affc),
	.w1(32'hb9af515a),
	.w2(32'h3c391db2),
	.w3(32'hbc05009a),
	.w4(32'h3b1b513c),
	.w5(32'h3c707113),
	.w6(32'h3bc7a35d),
	.w7(32'hbba2a0ba),
	.w8(32'hbb3810c7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad66fc5),
	.w1(32'h3bc1cd55),
	.w2(32'h3c51797d),
	.w3(32'h3ae7aeeb),
	.w4(32'h3beb1ce5),
	.w5(32'h3c488285),
	.w6(32'h3ba36521),
	.w7(32'h3af45894),
	.w8(32'h3ad3b5d5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dcf8d),
	.w1(32'hbab84d3a),
	.w2(32'hba8af45a),
	.w3(32'hbb069b5a),
	.w4(32'hbab6626d),
	.w5(32'hbaaf6d72),
	.w6(32'hba50c5a3),
	.w7(32'hbac53dcf),
	.w8(32'h3ad91dfb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49eace),
	.w1(32'hbbbfc840),
	.w2(32'h3be17e10),
	.w3(32'hbc6bd9a7),
	.w4(32'hbb8e9461),
	.w5(32'h3c03d2cd),
	.w6(32'h3b60a14e),
	.w7(32'hbbae080f),
	.w8(32'hbc1a4873),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015841),
	.w1(32'hba826e8a),
	.w2(32'h39f9c75c),
	.w3(32'hbacab084),
	.w4(32'hbb0f1d62),
	.w5(32'hba71b79c),
	.w6(32'hb90b58a9),
	.w7(32'hbb230171),
	.w8(32'h3a50ec52),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9ea0b),
	.w1(32'hbb48a915),
	.w2(32'h3be6cdf9),
	.w3(32'h3ba3c5a2),
	.w4(32'h3b2b5a30),
	.w5(32'h3c1a1485),
	.w6(32'h3c03c517),
	.w7(32'hbb9c5eef),
	.w8(32'hbb59316f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a7370),
	.w1(32'h3c68e97b),
	.w2(32'h3c151b23),
	.w3(32'h3c369e46),
	.w4(32'h3c14f218),
	.w5(32'h3af7db64),
	.w6(32'h3ba1d4d3),
	.w7(32'h3b5441f3),
	.w8(32'h3acfe680),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5c0ce),
	.w1(32'h3a72397e),
	.w2(32'h3cdc84f0),
	.w3(32'hbc7f3a25),
	.w4(32'h3c29ec88),
	.w5(32'h3d148191),
	.w6(32'h3b892d94),
	.w7(32'hbbe831ad),
	.w8(32'h3c3ced8e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa43454),
	.w1(32'hb9f79c63),
	.w2(32'h3b9fe8a3),
	.w3(32'hbbd16a1e),
	.w4(32'hbb82875d),
	.w5(32'h3a8f9641),
	.w6(32'hbab58c44),
	.w7(32'hbad6bc3f),
	.w8(32'hbb449f5b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee66a),
	.w1(32'hb8b7d541),
	.w2(32'h3c4c8e37),
	.w3(32'hbb973609),
	.w4(32'hbc18118e),
	.w5(32'hbc0c6863),
	.w6(32'hbba67a80),
	.w7(32'hbbd158cb),
	.w8(32'hbc17dd6d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b35137),
	.w1(32'h39cc11e1),
	.w2(32'h39eee7c9),
	.w3(32'hb7af1abb),
	.w4(32'h38c158f8),
	.w5(32'hb9e42d91),
	.w6(32'hb9ee4710),
	.w7(32'h39381d34),
	.w8(32'hba810293),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bf247),
	.w1(32'h3bc50c41),
	.w2(32'h3cc7385c),
	.w3(32'hbc09f713),
	.w4(32'hbb8a743d),
	.w5(32'h3ca31d19),
	.w6(32'h3c15aa32),
	.w7(32'hb8b56ae4),
	.w8(32'hbc8389cc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b703612),
	.w1(32'h3c032be4),
	.w2(32'h3c02b24a),
	.w3(32'hbab899c5),
	.w4(32'hbb8e3bf6),
	.w5(32'hbbd2ee3c),
	.w6(32'hbb9c47c9),
	.w7(32'hbb5d6a59),
	.w8(32'hbb88b759),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc32b3e),
	.w1(32'hbb2df006),
	.w2(32'h3b1c9a2c),
	.w3(32'hbb944a59),
	.w4(32'h3b80dd53),
	.w5(32'h3bdf2f14),
	.w6(32'h3b027508),
	.w7(32'hbbb70396),
	.w8(32'hba47047b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015a2f),
	.w1(32'hbbb0ed6f),
	.w2(32'hbb650212),
	.w3(32'hbc066905),
	.w4(32'hbb750762),
	.w5(32'h3b8310ba),
	.w6(32'h3ac13815),
	.w7(32'hb9ec3041),
	.w8(32'h398f3c9c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04b44e),
	.w1(32'h3b2fc0f2),
	.w2(32'h3b240920),
	.w3(32'hbad0cc32),
	.w4(32'hb8a782ab),
	.w5(32'h39efd175),
	.w6(32'h3b942813),
	.w7(32'h3b04c181),
	.w8(32'h3b1895d2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eb545),
	.w1(32'hbb183cfb),
	.w2(32'hbb626ecf),
	.w3(32'hbbb24cad),
	.w4(32'hbb861d1d),
	.w5(32'hbb86ebd0),
	.w6(32'hbaf676f7),
	.w7(32'hbb2a1465),
	.w8(32'hbaa51ebd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa239f0),
	.w1(32'h3b16eaae),
	.w2(32'h3abe5ba8),
	.w3(32'h39921fbf),
	.w4(32'h3a8bd51a),
	.w5(32'h3b21b1ba),
	.w6(32'hb99e0403),
	.w7(32'h38b073b3),
	.w8(32'h3a26fe24),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18326e),
	.w1(32'h3c380fe8),
	.w2(32'h3cd22cb2),
	.w3(32'h3a406f72),
	.w4(32'hb8579780),
	.w5(32'h3c165a0c),
	.w6(32'h3b98fee6),
	.w7(32'hba294bee),
	.w8(32'hbb6fb834),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20dd85),
	.w1(32'h3b1e7bbf),
	.w2(32'h3b67da33),
	.w3(32'h3a3bace8),
	.w4(32'h3b085b12),
	.w5(32'h3b603642),
	.w6(32'hb9566b9d),
	.w7(32'hba1e5555),
	.w8(32'h3a8d89bb),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ae3b0),
	.w1(32'hb84b38cb),
	.w2(32'h3a02072a),
	.w3(32'h3952355d),
	.w4(32'hba507358),
	.w5(32'h39f5b6c6),
	.w6(32'h3a8fddbe),
	.w7(32'hb95711ce),
	.w8(32'h3a1e6430),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bba87),
	.w1(32'hbb159392),
	.w2(32'h3ae8871a),
	.w3(32'hbb73c721),
	.w4(32'hbabe04f7),
	.w5(32'h3b0f6f17),
	.w6(32'h3b099eb5),
	.w7(32'hbac57631),
	.w8(32'hbae7610f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3612352e),
	.w1(32'hbb24dfed),
	.w2(32'hbb33acf1),
	.w3(32'hbb793941),
	.w4(32'hbb997cb7),
	.w5(32'hbb47b542),
	.w6(32'hbb1297e3),
	.w7(32'hbb8a054a),
	.w8(32'hbb3613ef),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c882b0),
	.w1(32'h3b8fdd2a),
	.w2(32'h3c3a8d75),
	.w3(32'h3b652759),
	.w4(32'h3bd6c837),
	.w5(32'h3bf9c599),
	.w6(32'h3ba30912),
	.w7(32'h3b078d65),
	.w8(32'hbb81909c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58373e),
	.w1(32'h39fcb2f7),
	.w2(32'h3a9b2f3e),
	.w3(32'h3ab371b6),
	.w4(32'h3aa5e012),
	.w5(32'h3ad1d3eb),
	.w6(32'h3ae5e692),
	.w7(32'h3b0ff7ac),
	.w8(32'h3b75815d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87cd22),
	.w1(32'hbce8a4b9),
	.w2(32'hbc272069),
	.w3(32'hbd0728fa),
	.w4(32'hbc87fcdc),
	.w5(32'h3c6f8ca2),
	.w6(32'h3c40b868),
	.w7(32'hbb952d55),
	.w8(32'hbc665a2c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c09b3),
	.w1(32'h3a40a547),
	.w2(32'hb79569b5),
	.w3(32'h3a6a0005),
	.w4(32'h3a895c07),
	.w5(32'h3a4fa88f),
	.w6(32'h3a7485d6),
	.w7(32'h3a0eae5f),
	.w8(32'h3b0239dd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98da61),
	.w1(32'h3b8a88db),
	.w2(32'h3b9e9bbc),
	.w3(32'hbb231fe3),
	.w4(32'hbb10b3a8),
	.w5(32'hbae89a7d),
	.w6(32'h3abdcdbd),
	.w7(32'h3a77ebef),
	.w8(32'h3b36baa1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a8a65),
	.w1(32'h3a1000a7),
	.w2(32'hb98d4d76),
	.w3(32'h3a5b6f24),
	.w4(32'h3aad3838),
	.w5(32'h3a38e261),
	.w6(32'h3b0512e1),
	.w7(32'h3ab9abde),
	.w8(32'h3a3acf31),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c244f),
	.w1(32'h3b2d0392),
	.w2(32'h3b967840),
	.w3(32'hbab057d7),
	.w4(32'hbbac9759),
	.w5(32'hbb791c42),
	.w6(32'h3bd106d5),
	.w7(32'h3b4e88fb),
	.w8(32'hbb95ab71),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e928c),
	.w1(32'h3aefc835),
	.w2(32'h3ab33666),
	.w3(32'h3b280012),
	.w4(32'h3ad20b5a),
	.w5(32'h3ad301c3),
	.w6(32'h3b18a03c),
	.w7(32'h3af3fe46),
	.w8(32'hba1947ce),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd9f89),
	.w1(32'h3b4b5cbd),
	.w2(32'h3b66cb5b),
	.w3(32'hbb8dbc74),
	.w4(32'hbbb2892f),
	.w5(32'hbadfcaeb),
	.w6(32'h3a069ee9),
	.w7(32'hbaa0d709),
	.w8(32'h3b25d349),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a408553),
	.w1(32'h3a2f8df5),
	.w2(32'hb99deb38),
	.w3(32'h3a876386),
	.w4(32'h3a4412d3),
	.w5(32'h39bcef97),
	.w6(32'h3a78f8d7),
	.w7(32'h392121b6),
	.w8(32'h3b195ee9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd2a54),
	.w1(32'hbbe17cc0),
	.w2(32'h3be39117),
	.w3(32'hbc1f6d62),
	.w4(32'hbb104fd0),
	.w5(32'h3c3315ec),
	.w6(32'h3c0261b4),
	.w7(32'h38fb234a),
	.w8(32'hbbcbaf31),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a1b26),
	.w1(32'h3bd0e4c9),
	.w2(32'h3c8e837b),
	.w3(32'hbb34bc9a),
	.w4(32'h3b21e473),
	.w5(32'h3c1e4ef2),
	.w6(32'hb984d226),
	.w7(32'h3b8a8b1b),
	.w8(32'h3a370808),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53627d),
	.w1(32'hbb1acac6),
	.w2(32'hbb04d7a3),
	.w3(32'hbb8d0ba2),
	.w4(32'hbb3170aa),
	.w5(32'hbae56014),
	.w6(32'hbb437d6e),
	.w7(32'hbb2f39c0),
	.w8(32'hba0e104a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba232120),
	.w1(32'h3a3459fa),
	.w2(32'h38eaf8a2),
	.w3(32'hba3d524e),
	.w4(32'hba96ae9a),
	.w5(32'hb9fb2ccb),
	.w6(32'h3abdd78d),
	.w7(32'h3a88ad16),
	.w8(32'h3ac3bace),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b99f8),
	.w1(32'h3b024f28),
	.w2(32'hbb709e50),
	.w3(32'hbbd6c7e1),
	.w4(32'hbc075c9b),
	.w5(32'hbb8b4d82),
	.w6(32'hbbad631a),
	.w7(32'hbb84ffac),
	.w8(32'h3b2b7229),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec433),
	.w1(32'hb90b740a),
	.w2(32'h3bd95f85),
	.w3(32'hbbd1e39b),
	.w4(32'hbb958292),
	.w5(32'h3b6d9025),
	.w6(32'h3be790c2),
	.w7(32'hbb3725c5),
	.w8(32'hbc162f98),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79d8b6),
	.w1(32'h3c30e9b3),
	.w2(32'h3d04aadf),
	.w3(32'h3cb2b1d0),
	.w4(32'h3cc7fcd7),
	.w5(32'h3b66ecac),
	.w6(32'h3c256bc6),
	.w7(32'hbb508ec1),
	.w8(32'h3bdc2a0e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8821ee),
	.w1(32'hbc164ebb),
	.w2(32'h3c177cf6),
	.w3(32'hbcb0796d),
	.w4(32'hbbb4faf2),
	.w5(32'h3c099252),
	.w6(32'h3be35e8d),
	.w7(32'hbc1f75b0),
	.w8(32'hbc6d9364),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf75c6a),
	.w1(32'h3c26d381),
	.w2(32'h3bd19c40),
	.w3(32'hbaf455c3),
	.w4(32'hbb1bacec),
	.w5(32'h3b206b0c),
	.w6(32'hbaf6a43f),
	.w7(32'hbb8ce4e9),
	.w8(32'h3b74eb9c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac47c8d),
	.w1(32'hba966bc2),
	.w2(32'hbac8ad03),
	.w3(32'hba66fa78),
	.w4(32'hb9606e74),
	.w5(32'hba911388),
	.w6(32'hbad7c808),
	.w7(32'hbaea0a9c),
	.w8(32'h39bccac3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41d0a6),
	.w1(32'h3a41ac0b),
	.w2(32'hba1eae17),
	.w3(32'hb9385b24),
	.w4(32'hb8e70f38),
	.w5(32'hba1479f0),
	.w6(32'h3a3f2e5e),
	.w7(32'h3941a94b),
	.w8(32'h3acddc7a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa5538),
	.w1(32'h3a9cf660),
	.w2(32'h3aa16698),
	.w3(32'h3a83257e),
	.w4(32'h3ab9974b),
	.w5(32'h3a18957d),
	.w6(32'h3aaf8008),
	.w7(32'h3a9f13b2),
	.w8(32'hbb30c7e3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ddfa8),
	.w1(32'h3b3910a3),
	.w2(32'h3a53eef3),
	.w3(32'hbac3ecbb),
	.w4(32'hba8c5fa9),
	.w5(32'hbadbcd7e),
	.w6(32'h3ab56d84),
	.w7(32'h39e82ac9),
	.w8(32'h3a21f112),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d3d03),
	.w1(32'h3ba471b8),
	.w2(32'h3b477b09),
	.w3(32'hbaa78204),
	.w4(32'hbaf66464),
	.w5(32'hbaf483b9),
	.w6(32'hbb42d71c),
	.w7(32'hba44b3f6),
	.w8(32'h3a7faa4a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d1d99),
	.w1(32'h3a41f60c),
	.w2(32'h3a49311f),
	.w3(32'hb9832a51),
	.w4(32'h3ac66b80),
	.w5(32'h3a88b047),
	.w6(32'h397a3bf5),
	.w7(32'h398bd143),
	.w8(32'hbb012da5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9ca3d),
	.w1(32'h3a61cda6),
	.w2(32'h39bddb53),
	.w3(32'hbbbde285),
	.w4(32'hbb722013),
	.w5(32'hbb6b7796),
	.w6(32'h3a908ecf),
	.w7(32'h3b4c71fd),
	.w8(32'h3bbc2389),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68ec90),
	.w1(32'h3a9f4ca4),
	.w2(32'h3b9e42f1),
	.w3(32'hb9fcd9d7),
	.w4(32'hbb2352f2),
	.w5(32'h3a92f87f),
	.w6(32'h3b3bd60f),
	.w7(32'hba08883d),
	.w8(32'hbbae6383),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b956d60),
	.w1(32'h3c181de4),
	.w2(32'h3c0fa594),
	.w3(32'h3bdf36f1),
	.w4(32'h3b9cc2fc),
	.w5(32'h3a455cec),
	.w6(32'hbb312536),
	.w7(32'hbb8ca29a),
	.w8(32'hbb11179c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90929f6),
	.w1(32'h3a787d53),
	.w2(32'h3c46b052),
	.w3(32'hbb85724e),
	.w4(32'h3ad8a0d9),
	.w5(32'h3ba30c43),
	.w6(32'h3708084c),
	.w7(32'h38c499f2),
	.w8(32'h3b28567b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae3679),
	.w1(32'h3c3e9b70),
	.w2(32'h3c8c4d30),
	.w3(32'h3aecc2fd),
	.w4(32'h3adf9084),
	.w5(32'h3b9fa8d7),
	.w6(32'h3ba206e0),
	.w7(32'hba512fda),
	.w8(32'h3b910312),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8de97b),
	.w1(32'hb80f94bc),
	.w2(32'hb99088f2),
	.w3(32'hbae18472),
	.w4(32'hb9b8e0af),
	.w5(32'hbaa2eec4),
	.w6(32'hbad2a69f),
	.w7(32'hba3becd6),
	.w8(32'h3b048898),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71e8da),
	.w1(32'h3a8fd117),
	.w2(32'h3ad31931),
	.w3(32'h3ab76822),
	.w4(32'h3a90e7de),
	.w5(32'h3b2a59fd),
	.w6(32'h3aca76d8),
	.w7(32'h3b13ca0b),
	.w8(32'hb89ae2e0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16fd74),
	.w1(32'h39617bed),
	.w2(32'hba5efc5d),
	.w3(32'hb9bdd165),
	.w4(32'hb8979c28),
	.w5(32'hb9ab885a),
	.w6(32'h393dbd06),
	.w7(32'hb99521b7),
	.w8(32'hb9a654b2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f2832c),
	.w1(32'hba2213e7),
	.w2(32'hb996f263),
	.w3(32'hba311230),
	.w4(32'h37d93451),
	.w5(32'hb970eb17),
	.w6(32'hb97f76b5),
	.w7(32'h3937bda8),
	.w8(32'h3af2a989),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b675304),
	.w1(32'h3a5310b9),
	.w2(32'hbb0aceff),
	.w3(32'h3b13efd4),
	.w4(32'hbae5ace4),
	.w5(32'hbb91701c),
	.w6(32'h3a923d50),
	.w7(32'hbb1dd591),
	.w8(32'hbb42365a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47d048),
	.w1(32'h3b380185),
	.w2(32'h3b1c7570),
	.w3(32'hbabd9ba5),
	.w4(32'h3a795db4),
	.w5(32'h3b31a00e),
	.w6(32'hba015194),
	.w7(32'h3ad97458),
	.w8(32'hb682a4a7),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74d64a),
	.w1(32'h3b44fa8e),
	.w2(32'hbb0fc306),
	.w3(32'hbb8c37fa),
	.w4(32'hbb9200e6),
	.w5(32'hbbfa0ba8),
	.w6(32'hbb845644),
	.w7(32'hba9ab2e5),
	.w8(32'h3a3aa4d4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368a90e7),
	.w1(32'hba303655),
	.w2(32'hbacaf5e8),
	.w3(32'hba60a587),
	.w4(32'hbadf5284),
	.w5(32'hbb4a7ba3),
	.w6(32'hbb4a5e5f),
	.w7(32'hbb3428b7),
	.w8(32'hbb1803b9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc155646),
	.w1(32'hbc3e2642),
	.w2(32'hbb0f5409),
	.w3(32'hbc893517),
	.w4(32'hbc132ddf),
	.w5(32'h3bc9ae75),
	.w6(32'h3bd92de8),
	.w7(32'hbb0d48a1),
	.w8(32'hba4bee8c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3e163),
	.w1(32'hba8c037b),
	.w2(32'hb984e588),
	.w3(32'h3baff2c5),
	.w4(32'hbb377c0f),
	.w5(32'hba542661),
	.w6(32'h3b800a62),
	.w7(32'h399a9139),
	.w8(32'hba615249),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b274c7f),
	.w1(32'hba132b50),
	.w2(32'hbab275ec),
	.w3(32'hb876d5e4),
	.w4(32'hbb8e386c),
	.w5(32'hbbd4fd1b),
	.w6(32'hba16af74),
	.w7(32'hbaf72e84),
	.w8(32'hbad64626),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6f31e),
	.w1(32'h3aa6565a),
	.w2(32'h3ab1f0cf),
	.w3(32'h3a86759e),
	.w4(32'h37c50502),
	.w5(32'hb9ae973f),
	.w6(32'h39e2f6cd),
	.w7(32'h3a6efc50),
	.w8(32'h3a7153a3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd717a),
	.w1(32'h3a2fc295),
	.w2(32'hba46fd98),
	.w3(32'hbb68cef4),
	.w4(32'hbb9f53b1),
	.w5(32'hbbf44439),
	.w6(32'hbb7d60b4),
	.w7(32'hbb39ef93),
	.w8(32'hbaccd2f1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90ed9b),
	.w1(32'h3ac31e9c),
	.w2(32'h3a8c28a6),
	.w3(32'h3b8d8cd4),
	.w4(32'hbae84c63),
	.w5(32'hbb93f28f),
	.w6(32'h3aab64d5),
	.w7(32'hbb51b1ec),
	.w8(32'hbad1e37c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8332f7),
	.w1(32'h3995d256),
	.w2(32'h3b8cf649),
	.w3(32'hba0013a4),
	.w4(32'h3ab5393d),
	.w5(32'h3bac0f5f),
	.w6(32'h3ba5a507),
	.w7(32'hbaca0e16),
	.w8(32'hbb0d6a6b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e89f5),
	.w1(32'hbb7e4f2b),
	.w2(32'hbbe0fdca),
	.w3(32'hbb445d14),
	.w4(32'hbb97f4ab),
	.w5(32'hbbaadcbb),
	.w6(32'hbb9ae8ef),
	.w7(32'hbbb2c5b1),
	.w8(32'hbbc68212),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a14f5),
	.w1(32'hba57e839),
	.w2(32'hba75c9ec),
	.w3(32'hba7a2cfc),
	.w4(32'hba8ca2a5),
	.w5(32'hbabbab2a),
	.w6(32'hbad09c66),
	.w7(32'hba99385e),
	.w8(32'hba79bc39),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e91ea),
	.w1(32'hbad8e172),
	.w2(32'h3a44dcf8),
	.w3(32'h3a55de9b),
	.w4(32'h3a55fec5),
	.w5(32'h3968b9b5),
	.w6(32'hbabe821b),
	.w7(32'hba65777a),
	.w8(32'h38e7da48),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4045d8),
	.w1(32'hbb47acf7),
	.w2(32'hbb8c545c),
	.w3(32'hbb5e3f7f),
	.w4(32'hbb66457d),
	.w5(32'hbba3f5b9),
	.w6(32'hbb133e8d),
	.w7(32'hbb29a474),
	.w8(32'h39e35a12),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b3426),
	.w1(32'h3a7dde8c),
	.w2(32'h3b2414e9),
	.w3(32'hba81af90),
	.w4(32'hbb731302),
	.w5(32'hba785acd),
	.w6(32'h3b3483a0),
	.w7(32'h3b1ecb1e),
	.w8(32'hbb7328e5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c930c),
	.w1(32'hbc0f2e9b),
	.w2(32'hbb3bc57c),
	.w3(32'hbc820bb5),
	.w4(32'hbc38fa9e),
	.w5(32'hba754930),
	.w6(32'hba86bab0),
	.w7(32'hbc01fd19),
	.w8(32'hbb375b18),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10254f),
	.w1(32'h3a47639d),
	.w2(32'hba9c4de0),
	.w3(32'h3a734ab7),
	.w4(32'h3b0fa32e),
	.w5(32'hb9d407d8),
	.w6(32'h3ad596da),
	.w7(32'hba3e81f1),
	.w8(32'hbb0f465a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d87b3),
	.w1(32'hbb6d0b98),
	.w2(32'hb9fac7a2),
	.w3(32'hbb257b45),
	.w4(32'hbb27d8ac),
	.w5(32'hbad4d525),
	.w6(32'hbb75d53a),
	.w7(32'hbad580f7),
	.w8(32'hbbc86532),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19eae5),
	.w1(32'h3c45279c),
	.w2(32'h3c23cb1e),
	.w3(32'hbbbc4230),
	.w4(32'hbc4f9f2f),
	.w5(32'hbc703d29),
	.w6(32'hbc32dc5c),
	.w7(32'hb9fed0fa),
	.w8(32'h3bb9c913),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b85422),
	.w1(32'hba2bd19a),
	.w2(32'h3b915223),
	.w3(32'h3ae09f7b),
	.w4(32'h3bccce98),
	.w5(32'h3bd9c44f),
	.w6(32'h3ba33553),
	.w7(32'h3b3e9fb8),
	.w8(32'h3bef0ac6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad91c46),
	.w1(32'h3993fcee),
	.w2(32'h3a9f9693),
	.w3(32'h3b2375e4),
	.w4(32'h3a531214),
	.w5(32'h3aacb163),
	.w6(32'h3ae9557b),
	.w7(32'h3b1c95b9),
	.w8(32'h3b6f8538),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32030f),
	.w1(32'h3bbc375e),
	.w2(32'h3bb02928),
	.w3(32'h39932264),
	.w4(32'h3b7d4834),
	.w5(32'h3bb374bc),
	.w6(32'h38c5bb5c),
	.w7(32'h3b12ac57),
	.w8(32'h3b8d878d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bae116),
	.w1(32'hbb633abc),
	.w2(32'hbb9e4183),
	.w3(32'h3aa162d0),
	.w4(32'hbb018c0a),
	.w5(32'hbb6bd7a7),
	.w6(32'h3aae9cfd),
	.w7(32'hba8da96f),
	.w8(32'hbb532901),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b574292),
	.w1(32'hbb651c9e),
	.w2(32'hb9ae2c2c),
	.w3(32'h3a98c43c),
	.w4(32'hbb3633e6),
	.w5(32'hba3db5f1),
	.w6(32'h3b515e18),
	.w7(32'hbac62628),
	.w8(32'h39df1de2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30a32a),
	.w1(32'h3b206c8e),
	.w2(32'h3bc02dff),
	.w3(32'hba0ae025),
	.w4(32'hbb15756e),
	.w5(32'h3a1caf3f),
	.w6(32'hbac0dd48),
	.w7(32'h3a978e73),
	.w8(32'h3a7760b3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac22e2e),
	.w1(32'hbbf22343),
	.w2(32'h3b6870ca),
	.w3(32'hbbd11588),
	.w4(32'hbb5164ea),
	.w5(32'h3bd07833),
	.w6(32'h38ff7899),
	.w7(32'h3b31dc10),
	.w8(32'h3abc472e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule