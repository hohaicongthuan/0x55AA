module layer_8_featuremap_157(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3d2bc),
	.w1(32'hbaf6936c),
	.w2(32'h3be491d0),
	.w3(32'h3c589564),
	.w4(32'h3c44deeb),
	.w5(32'h3b95c885),
	.w6(32'hbc109491),
	.w7(32'h3bf606bb),
	.w8(32'hbc941123),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b827e6a),
	.w1(32'h3c04a425),
	.w2(32'hbb96c0a5),
	.w3(32'hbb744e37),
	.w4(32'hbacfafb4),
	.w5(32'h3c0f6af1),
	.w6(32'hbbac1205),
	.w7(32'hba99b07f),
	.w8(32'hbc50fcf5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00f2c9),
	.w1(32'h3b3c7f12),
	.w2(32'hbb950f52),
	.w3(32'hba3bf2cb),
	.w4(32'hbab891bb),
	.w5(32'h3b9b54de),
	.w6(32'hbb8b2771),
	.w7(32'h3ac45e4f),
	.w8(32'h3b101c36),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43eb53),
	.w1(32'h3b5e6197),
	.w2(32'hbbe143a2),
	.w3(32'h3bd9dcf2),
	.w4(32'h3a2ef054),
	.w5(32'hbc0fa30a),
	.w6(32'hbc41869e),
	.w7(32'hba3d680b),
	.w8(32'h3cadbd0f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca065b),
	.w1(32'hbc08d92a),
	.w2(32'hbb8d55bb),
	.w3(32'hbc91390a),
	.w4(32'h3c893c1e),
	.w5(32'hbc2192d8),
	.w6(32'h3c01b4b9),
	.w7(32'hbcb8fea4),
	.w8(32'h3ce2fb10),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16997d),
	.w1(32'hbc680f1a),
	.w2(32'h3bca0b99),
	.w3(32'hbcb9cd82),
	.w4(32'h3c3719ec),
	.w5(32'hbc865042),
	.w6(32'h3aa2f667),
	.w7(32'hbc8fcc45),
	.w8(32'h3d1e8427),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc575071),
	.w1(32'hbc8458d7),
	.w2(32'hbc88b137),
	.w3(32'h3a93faf0),
	.w4(32'hbb192308),
	.w5(32'hbb21b0e7),
	.w6(32'h3c130463),
	.w7(32'hbc4e4df0),
	.w8(32'h3cd2a10e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dfdaa),
	.w1(32'h3b9bc51f),
	.w2(32'h3aea90cc),
	.w3(32'hbcaddd66),
	.w4(32'h3b073e2f),
	.w5(32'h3bc8a51f),
	.w6(32'hbc9194af),
	.w7(32'hbb57aa06),
	.w8(32'h3c88b39d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38dcd8),
	.w1(32'h3bd1d914),
	.w2(32'hbb894b47),
	.w3(32'h3c5fe8dc),
	.w4(32'hbc7bb79d),
	.w5(32'hbc8fc7de),
	.w6(32'hbc2df9ce),
	.w7(32'hbc2f08aa),
	.w8(32'h3bfb803e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45cc5d),
	.w1(32'hbc17260c),
	.w2(32'hbb9bd519),
	.w3(32'hbbad09a1),
	.w4(32'hbb026b91),
	.w5(32'hbbb0095e),
	.w6(32'h3ae3a889),
	.w7(32'h3a964427),
	.w8(32'h3ca5aa73),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14bed5),
	.w1(32'h3c0a6f31),
	.w2(32'hbc62e931),
	.w3(32'h3ae3775a),
	.w4(32'hbc132c38),
	.w5(32'h3b70544b),
	.w6(32'hbc57908c),
	.w7(32'h3ba6d5f5),
	.w8(32'hbc4f4a0f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc502c40),
	.w1(32'hbac9321d),
	.w2(32'hbc1332af),
	.w3(32'h3c68f6a5),
	.w4(32'hbb300926),
	.w5(32'hbb80d4d4),
	.w6(32'hbc124a39),
	.w7(32'hbc1d36ec),
	.w8(32'hbb951dcc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd38701),
	.w1(32'h3c477949),
	.w2(32'hbeb1b856),
	.w3(32'hb9911c25),
	.w4(32'h3eaa1a42),
	.w5(32'h3f96c953),
	.w6(32'hbc0c6678),
	.w7(32'hbf1aa07a),
	.w8(32'hbf1e417d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf3b2d46),
	.w1(32'h3ee73a5a),
	.w2(32'hbed11dee),
	.w3(32'hbed5830d),
	.w4(32'h3e963a6e),
	.w5(32'hbf68898e),
	.w6(32'h3fb52132),
	.w7(32'h3fb6f2d4),
	.w8(32'hbf89f25a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbfb900f9),
	.w1(32'hbf311557),
	.w2(32'hbf3f883e),
	.w3(32'hbf350d3d),
	.w4(32'h3f73d6b4),
	.w5(32'hbe8395dd),
	.w6(32'hbee00fba),
	.w7(32'h3fc586c0),
	.w8(32'hbe2c73b4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fae04e9),
	.w1(32'h3e2cf42f),
	.w2(32'h3eafea55),
	.w3(32'hbf35ca86),
	.w4(32'h3e5d78ea),
	.w5(32'h3f05ec25),
	.w6(32'h3faf743d),
	.w7(32'hbf344d6c),
	.w8(32'hbe6f96d5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf15b209),
	.w1(32'hbfd1bc9b),
	.w2(32'hbfb4d19f),
	.w3(32'hbf815504),
	.w4(32'h3f79df23),
	.w5(32'hbdd490df),
	.w6(32'h3e9ca5aa),
	.w7(32'hbf8da50d),
	.w8(32'h3f1aa09b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fce01ed),
	.w1(32'h3f1115ca),
	.w2(32'h3e0a4073),
	.w3(32'hbc43fb3e),
	.w4(32'hbea22a8b),
	.w5(32'hbeeeed01),
	.w6(32'hbe76d97c),
	.w7(32'h3f0ee60e),
	.w8(32'hbf3ffd10),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e9897e6),
	.w1(32'h3f13efe4),
	.w2(32'hbe95a861),
	.w3(32'h3fa006f7),
	.w4(32'h3e9c7314),
	.w5(32'hbf9b8e1e),
	.w6(32'h3e62ac3b),
	.w7(32'h3d02298f),
	.w8(32'hbf27ceb3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf5d09c8),
	.w1(32'hbf63cbc3),
	.w2(32'hbdcb24da),
	.w3(32'h3fa34f45),
	.w4(32'h3f0fac30),
	.w5(32'h3dd060a2),
	.w6(32'hbe1cc704),
	.w7(32'hbf097dc0),
	.w8(32'hbf77959b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fac2123),
	.w1(32'h3ea42727),
	.w2(32'h3f687099),
	.w3(32'hbf539ed4),
	.w4(32'h3d570f28),
	.w5(32'h3fa99d5d),
	.w6(32'hbf1f493c),
	.w7(32'h3e83ae27),
	.w8(32'hbf2b0e8e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3faa9671),
	.w1(32'hbf35b6c5),
	.w2(32'hbf293085),
	.w3(32'hbdab85be),
	.w4(32'h3e9012c4),
	.w5(32'h3e5fb64f),
	.w6(32'hbf0cf3f8),
	.w7(32'hbecc4b2c),
	.w8(32'hbf164f97),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf48f07a),
	.w1(32'h3e53db9c),
	.w2(32'hbe99e0b8),
	.w3(32'h3ed0a03e),
	.w4(32'hbf02dc7e),
	.w5(32'hbf47f993),
	.w6(32'hbea43b3c),
	.w7(32'h3f8ef9dd),
	.w8(32'hbec4dc43),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1d01d4),
	.w1(32'h3eaf4728),
	.w2(32'hbdcf95ea),
	.w3(32'h3ee3abfe),
	.w4(32'hbe801b94),
	.w5(32'h3e97ea91),
	.w6(32'h3f920725),
	.w7(32'hbeb21992),
	.w8(32'h3f0b5b8b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8f1609),
	.w1(32'h3d832f9c),
	.w2(32'h3ea5400c),
	.w3(32'h3effecb4),
	.w4(32'h3e1cd234),
	.w5(32'hbf818832),
	.w6(32'hbdfd6d51),
	.w7(32'hbf4d0f10),
	.w8(32'hbf317dcc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fdc078d),
	.w1(32'h3dacee9e),
	.w2(32'h3f76e34d),
	.w3(32'hbe30cccd),
	.w4(32'hbf4d836e),
	.w5(32'hbf1fb361),
	.w6(32'h3ef73678),
	.w7(32'hbf29db3e),
	.w8(32'h3f73f255),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf686316),
	.w1(32'hbf3f66d2),
	.w2(32'hbf7d0091),
	.w3(32'h3f1200ca),
	.w4(32'h3ef18f85),
	.w5(32'h3e2b1f4a),
	.w6(32'h3f1708d3),
	.w7(32'hbded489d),
	.w8(32'h3f99d9e3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f05a103),
	.w1(32'hbf066339),
	.w2(32'h3f9ee565),
	.w3(32'hbf1495d7),
	.w4(32'h3e9b97fc),
	.w5(32'h3f29c2ef),
	.w6(32'h3f6ad415),
	.w7(32'h3ea3238d),
	.w8(32'h3f45377f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbef9099e),
	.w1(32'hbede62d2),
	.w2(32'hbf23d5f7),
	.w3(32'hbec4c946),
	.w4(32'h3e2727cb),
	.w5(32'h3f632a42),
	.w6(32'hbea1df45),
	.w7(32'hbf72aefe),
	.w8(32'hbf86a649),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf2e8256),
	.w1(32'h3eaeb8d6),
	.w2(32'hbeef04e9),
	.w3(32'h3e08ac25),
	.w4(32'hbe0d4b18),
	.w5(32'hbec6ee24),
	.w6(32'hbf8f2f0e),
	.w7(32'hbf64d23d),
	.w8(32'hbf85f50a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf4ace11),
	.w1(32'hbebd96ac),
	.w2(32'hbef70ef8),
	.w3(32'h3f9f37c2),
	.w4(32'hbf5c4f69),
	.w5(32'hbebf9463),
	.w6(32'hbf5ec03b),
	.w7(32'h3f05573a),
	.w8(32'hbeffb13e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e931831),
	.w1(32'hbf329b5a),
	.w2(32'hbe846113),
	.w3(32'hbeeb3b16),
	.w4(32'h3f0c4131),
	.w5(32'h3f9a31f7),
	.w6(32'hbee16dfb),
	.w7(32'h3ff6ef1d),
	.w8(32'h3d5f0340),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeef0660),
	.w1(32'hbf1154a9),
	.w2(32'hbf511030),
	.w3(32'hbf7b4032),
	.w4(32'hbf7c84a5),
	.w5(32'hbbfe9433),
	.w6(32'hbfe3361a),
	.w7(32'h3e0cf5e1),
	.w8(32'hbf82b022),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ed90a26),
	.w1(32'h3ea877ea),
	.w2(32'h3f27840c),
	.w3(32'hbf6e28b2),
	.w4(32'h3edf388e),
	.w5(32'hbf66b0c0),
	.w6(32'h3f47d214),
	.w7(32'h3e6d67e2),
	.w8(32'hbf07c1b1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf831baa),
	.w1(32'hbdf8db90),
	.w2(32'hbf31ccef),
	.w3(32'hbf128d51),
	.w4(32'h3e69e414),
	.w5(32'hbea1ac8d),
	.w6(32'h3f82c7e4),
	.w7(32'hbf2884a2),
	.w8(32'h3f43ef84),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3eba8182),
	.w1(32'hbe7898ca),
	.w2(32'hbf34cdc4),
	.w3(32'hbe5a9192),
	.w4(32'hbdc4bb67),
	.w5(32'hbf170970),
	.w6(32'h3d00afcc),
	.w7(32'h3ebf1f5b),
	.w8(32'hbf35b812),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf4c50cf),
	.w1(32'hbf575c11),
	.w2(32'hbf829e7c),
	.w3(32'hbf1d6089),
	.w4(32'hbf930baf),
	.w5(32'h3eea3f0b),
	.w6(32'hbf96085a),
	.w7(32'h3ec3a16d),
	.w8(32'h3f66b6ca),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f52b3b8),
	.w1(32'hbf306a4d),
	.w2(32'hbf15ee17),
	.w3(32'hbe7488f0),
	.w4(32'hbf432275),
	.w5(32'hbe347900),
	.w6(32'hbebe9733),
	.w7(32'h3f14e2b8),
	.w8(32'hbe923399),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf02e1a3),
	.w1(32'h3ef442a1),
	.w2(32'h3ec89253),
	.w3(32'hbf551a8f),
	.w4(32'hbe894106),
	.w5(32'h3e1a5b68),
	.w6(32'hbf30c6cd),
	.w7(32'h3ef79aeb),
	.w8(32'hbfbef5f9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec982b1),
	.w1(32'h3dc6424e),
	.w2(32'h3e8cbc68),
	.w3(32'hbdf4cc9a),
	.w4(32'h3e6a03ea),
	.w5(32'hbf61e6ce),
	.w6(32'hbf70399f),
	.w7(32'h3f967408),
	.w8(32'h3f33158c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e7ef56f),
	.w1(32'hbf1bf5af),
	.w2(32'hbe9fb9f8),
	.w3(32'hbf3e88c0),
	.w4(32'hbe9f7e92),
	.w5(32'hbf0a8d64),
	.w6(32'h3f8193fc),
	.w7(32'hbf2a383f),
	.w8(32'h3f9e2fbc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ec221d6),
	.w1(32'h3f188324),
	.w2(32'h3f8e47e3),
	.w3(32'h3f8fda1b),
	.w4(32'h3fa873e3),
	.w5(32'h3f1ce79c),
	.w6(32'h3f8b6186),
	.w7(32'h3f33ebb3),
	.w8(32'h3f93ece7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2613c1),
	.w1(32'h3f562570),
	.w2(32'h3f042f01),
	.w3(32'h3f1577be),
	.w4(32'h3fcbeff8),
	.w5(32'h3f1085da),
	.w6(32'h3fc5def7),
	.w7(32'h3fb14d48),
	.w8(32'h3f209ef2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f951eaf),
	.w1(32'h3f6e1f5c),
	.w2(32'h3f5fc7c8),
	.w3(32'h3f92c5c4),
	.w4(32'h3f4f7297),
	.w5(32'h3f812979),
	.w6(32'h3faac45c),
	.w7(32'h3f8a1d3f),
	.w8(32'h3f59ec43),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fa91272),
	.w1(32'h3e8aa567),
	.w2(32'h3f82e804),
	.w3(32'h3fa21f8b),
	.w4(32'h3f8d0391),
	.w5(32'h3f8784c2),
	.w6(32'h3f67eb4f),
	.w7(32'h3fcddb4e),
	.w8(32'h3f8f27f3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fba4f3c),
	.w1(32'h3f6e5600),
	.w2(32'h3f181767),
	.w3(32'h3fbab245),
	.w4(32'h3f8fc5e2),
	.w5(32'h3fafb62d),
	.w6(32'h3f953231),
	.w7(32'h3f8ace82),
	.w8(32'h3f1d4f30),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fa86c7d),
	.w1(32'h3f82e041),
	.w2(32'h3f8421ff),
	.w3(32'h3f995827),
	.w4(32'h3f6b0599),
	.w5(32'h3eb9cd9b),
	.w6(32'h3f8518f7),
	.w7(32'h3f97e634),
	.w8(32'h3f4a8d6f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f9f17ad),
	.w1(32'h3f8eb0ed),
	.w2(32'h3fa49646),
	.w3(32'h3f1fdebe),
	.w4(32'h3ef58985),
	.w5(32'h3fbd9541),
	.w6(32'h3fa6a084),
	.w7(32'h3fa779a3),
	.w8(32'h3f383dd9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f413faa),
	.w1(32'h3fbead3e),
	.w2(32'h3f009b8b),
	.w3(32'h3e817579),
	.w4(32'h3f3ad24f),
	.w5(32'h3f936e64),
	.w6(32'h3f2059d8),
	.w7(32'h3f8d64ba),
	.w8(32'h3f79b6c8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f30d739),
	.w1(32'h3fa92d4f),
	.w2(32'h3fb1369d),
	.w3(32'h3f693e9d),
	.w4(32'h3f4687d3),
	.w5(32'h3fa2b048),
	.w6(32'h3f9050d3),
	.w7(32'h3f4ab99c),
	.w8(32'h3f6ee620),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fab5ba4),
	.w1(32'h3f284ede),
	.w2(32'h3ebd6a0a),
	.w3(32'h3f47beae),
	.w4(32'h3f2e8927),
	.w5(32'h3f906dea),
	.w6(32'h3f013598),
	.w7(32'h3f28873b),
	.w8(32'h3f848331),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f29bff0),
	.w1(32'h3f933872),
	.w2(32'h3f8521ab),
	.w3(32'h3f674b59),
	.w4(32'h3f87c88b),
	.w5(32'h3f48a52c),
	.w6(32'h3f8f5cbc),
	.w7(32'hba394756),
	.w8(32'h3fa98cee),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d71854a),
	.w1(32'h3f4f1421),
	.w2(32'h3f76ff0a),
	.w3(32'h3f98ee34),
	.w4(32'h3f63ba89),
	.w5(32'h3fb5a275),
	.w6(32'h3f139b4e),
	.w7(32'h3fa245cd),
	.w8(32'h3f1d7d5c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f314986),
	.w1(32'h3f9d49fa),
	.w2(32'h3edaf959),
	.w3(32'h3f2cf6f8),
	.w4(32'h3f1b4a80),
	.w5(32'h3f5b04a9),
	.w6(32'h3faf5755),
	.w7(32'h3eef495d),
	.w8(32'h3f67020d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f9e8b9c),
	.w1(32'h3f815246),
	.w2(32'h3f5ddd7e),
	.w3(32'h3f2756c0),
	.w4(32'h3dee49c7),
	.w5(32'h3f82d50a),
	.w6(32'hb79da856),
	.w7(32'h3f578b1e),
	.w8(32'h3f34f348),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ef7d75e),
	.w1(32'h3f56b699),
	.w2(32'h3f4076be),
	.w3(32'h3f9445a1),
	.w4(32'h3f8356ef),
	.w5(32'h3f7ae35f),
	.w6(32'h3f7d12f1),
	.w7(32'h3f25cc34),
	.w8(32'h3faeff89),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f555288),
	.w1(32'h3f841c16),
	.w2(32'h3f920a6d),
	.w3(32'h3f825016),
	.w4(32'h3f2c0cac),
	.w5(32'h3f8bbbb9),
	.w6(32'h3ed3df6a),
	.w7(32'h3f8c87d5),
	.w8(32'h3f62d716),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fbc6434),
	.w1(32'h3fb30da5),
	.w2(32'h3f9d315f),
	.w3(32'h3f58cc69),
	.w4(32'h3fa4cd4d),
	.w5(32'h3f17448e),
	.w6(32'h3fa07de8),
	.w7(32'h3e2769fa),
	.w8(32'h3f9f6ba5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f6c5382),
	.w1(32'h3fb882d0),
	.w2(32'h3facb2f6),
	.w3(32'h3f2579d1),
	.w4(32'h3f9d5ac9),
	.w5(32'h3f1eb43f),
	.w6(32'h3f3ad4fc),
	.w7(32'h3f195174),
	.w8(32'h3fa42733),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f0ff1fa),
	.w1(32'h3fa68eb0),
	.w2(32'h3f17d57e),
	.w3(32'h388289c9),
	.w4(32'h3edd3ed8),
	.w5(32'h3f912154),
	.w6(32'h3f7ec211),
	.w7(32'h3f1d2a29),
	.w8(32'h3f8e901a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3ce1d8),
	.w1(32'h3f459e0f),
	.w2(32'h3f9c3e20),
	.w3(32'h3f0be4e6),
	.w4(32'h3e228935),
	.w5(32'h3f8e7069),
	.w6(32'h3f8fd09d),
	.w7(32'h3fa847bc),
	.w8(32'h3fbe455b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f592168),
	.w1(32'h3fb6a972),
	.w2(32'h3f0cbf27),
	.w3(32'h3fac35be),
	.w4(32'h3fb7f3bd),
	.w5(32'h3f00502a),
	.w6(32'h3f91edc1),
	.w7(32'h3fa7000d),
	.w8(32'h3f617da3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3fa277e1),
	.w1(32'h3f7f90d5),
	.w2(32'h3f8215b7),
	.w3(32'h3f6c49db),
	.w4(32'h3fa3a005),
	.w5(32'h3f5d7e90),
	.w6(32'h3f8a2f6e),
	.w7(32'h3f566b20),
	.w8(32'h3f16ca17),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f865368),
	.w1(32'h3f7ed43d),
	.w2(32'h3f4eec22),
	.w3(32'h3f93a69c),
	.w4(32'h3f3897ff),
	.w5(32'h3e9041e0),
	.w6(32'h3f3344e9),
	.w7(32'h3f701287),
	.w8(32'h3e49559a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f8f7c68),
	.w1(32'h3f909965),
	.w2(32'h3f9fb7a0),
	.w3(32'h3f3ac1e4),
	.w4(32'h3f0e437d),
	.w5(32'h3f7862f6),
	.w6(32'h3da3099e),
	.w7(32'h3f88ed0d),
	.w8(32'h3f4d12b1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cee661a),
	.w1(32'h3f505c1c),
	.w2(32'h3f36530d),
	.w3(32'h3f8aac1a),
	.w4(32'h3f635482),
	.w5(32'h3fa22aeb),
	.w6(32'h3f1d7768),
	.w7(32'h3f969a0d),
	.w8(32'h3f9e964d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f9b786e),
	.w1(32'h3f9be571),
	.w2(32'h3f6b39e3),
	.w3(32'h3f89902e),
	.w4(32'h3f92b955),
	.w5(32'h3f8cef7c),
	.w6(32'h3f56f784),
	.w7(32'h3f8dd75a),
	.w8(32'h3f73d24d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f8546e7),
	.w1(32'h3f50761c),
	.w2(32'h3f970d7b),
	.w3(32'h3fbc3fe6),
	.w4(32'h3f534434),
	.w5(32'h3f8507e8),
	.w6(32'h3f820ca6),
	.w7(32'h3fa0408b),
	.w8(32'h3e64dd14),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f890c26),
	.w1(32'h3f638deb),
	.w2(32'h3f9ba2f9),
	.w3(32'h3f9a75ef),
	.w4(32'h3f496709),
	.w5(32'h3f9e1b98),
	.w6(32'h3f652c55),
	.w7(32'h3f9e9080),
	.w8(32'h3fa119b2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3efa98af),
	.w1(32'h3d81fd34),
	.w2(32'hbc8878f8),
	.w3(32'h3f8a0c6a),
	.w4(32'h3ead1e4f),
	.w5(32'h3f391005),
	.w6(32'h3f870130),
	.w7(32'hbebd55f7),
	.w8(32'h3e2223ed),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e406851),
	.w1(32'h3dd50953),
	.w2(32'hbe70ea62),
	.w3(32'hbe8a8042),
	.w4(32'h3fd091e8),
	.w5(32'hbf6ee165),
	.w6(32'hbfc1682b),
	.w7(32'h3e3a6187),
	.w8(32'hbe08b63f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbfa3afd6),
	.w1(32'hbf349a11),
	.w2(32'hbee6ae3c),
	.w3(32'h3ea9b896),
	.w4(32'hbe4a4a27),
	.w5(32'hbf449c73),
	.w6(32'hbf519546),
	.w7(32'hbe8fd940),
	.w8(32'h3f89b318),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe4f7b04),
	.w1(32'hbf0abc57),
	.w2(32'h3e425b38),
	.w3(32'hbfb2b0c2),
	.w4(32'hbf797703),
	.w5(32'h3ecba1b9),
	.w6(32'h3df80539),
	.w7(32'h3f6142d0),
	.w8(32'hbe940d16),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdaf959c),
	.w1(32'h3f0c55e4),
	.w2(32'h3d1c2ab9),
	.w3(32'h3e18d524),
	.w4(32'hbddc6898),
	.w5(32'h3ee3a092),
	.w6(32'hbf8064c2),
	.w7(32'hbe950e82),
	.w8(32'hbee9732e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e3fb841),
	.w1(32'hbe8871df),
	.w2(32'h3e9e1cb7),
	.w3(32'hbe950665),
	.w4(32'hbf906d6c),
	.w5(32'hbc90e519),
	.w6(32'hbeecc84c),
	.w7(32'hbf215ed0),
	.w8(32'hbf5a8515),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec9c518),
	.w1(32'h3e4c0ad9),
	.w2(32'hbdf86527),
	.w3(32'hbf40b3aa),
	.w4(32'hbda5f96f),
	.w5(32'hbf110ad7),
	.w6(32'h3f87afc1),
	.w7(32'h3e2b485f),
	.w8(32'hbe5a7906),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdde8fb8),
	.w1(32'hc06b4a28),
	.w2(32'hbe90b681),
	.w3(32'hbf4cd01c),
	.w4(32'h3e4e1a8c),
	.w5(32'hbdfdbd5c),
	.w6(32'hbf25fc4d),
	.w7(32'hbd4a9c06),
	.w8(32'h3f43ebcb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe95c1f9),
	.w1(32'hbef61cd3),
	.w2(32'hbf647fb6),
	.w3(32'h3d92cc8e),
	.w4(32'h3f181e65),
	.w5(32'hbe13b1fb),
	.w6(32'hbe1150bb),
	.w7(32'h3eb9924b),
	.w8(32'hbe57c207),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbea19d42),
	.w1(32'h3ec7ed2c),
	.w2(32'hbea63850),
	.w3(32'hbfbb2323),
	.w4(32'hbfda6c0d),
	.w5(32'h3dc7e554),
	.w6(32'hbf6ac899),
	.w7(32'h3e986086),
	.w8(32'hbee6125c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e9dc1eb),
	.w1(32'hbf542a49),
	.w2(32'hbd6ddbd4),
	.w3(32'hbef8492f),
	.w4(32'h40470011),
	.w5(32'h3e4090da),
	.w6(32'hbe41e50d),
	.w7(32'h3f15d179),
	.w8(32'hbf104583),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ab2aa),
	.w1(32'hbf295f7d),
	.w2(32'h3f884193),
	.w3(32'h3eb03b5d),
	.w4(32'hbdef4fc3),
	.w5(32'hbf9b2591),
	.w6(32'hbeee5545),
	.w7(32'hbf0f45b6),
	.w8(32'h3eaf4777),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbfcf9f9d),
	.w1(32'hbf2f6d11),
	.w2(32'hbe79f4db),
	.w3(32'h3f0db8fb),
	.w4(32'hbde0d23e),
	.w5(32'hbf16ec99),
	.w6(32'hbfc1ca80),
	.w7(32'h3d9b8692),
	.w8(32'hbfa541ea),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe3b59db),
	.w1(32'hbec02804),
	.w2(32'h38ad44af),
	.w3(32'hbfe94d7a),
	.w4(32'h3e19d747),
	.w5(32'h3f05be77),
	.w6(32'h3ce772b7),
	.w7(32'h3eb981db),
	.w8(32'h3c54995f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe925dd6),
	.w1(32'h3fc980d6),
	.w2(32'hba2505ba),
	.w3(32'hbeeea4e9),
	.w4(32'hbd3d5c4d),
	.w5(32'h3d4c1744),
	.w6(32'hbf03d48a),
	.w7(32'hbe73ce4b),
	.w8(32'hbf9b6fbd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf22c970),
	.w1(32'h3ef3fdb8),
	.w2(32'hbec297ac),
	.w3(32'h3f7ea04c),
	.w4(32'hbe0a5bd8),
	.w5(32'hbf3a5a09),
	.w6(32'hbf8e29d3),
	.w7(32'h3f04c6b0),
	.w8(32'hbfbbbc7d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbfc7dd40),
	.w1(32'hc03580f1),
	.w2(32'hbe9180cb),
	.w3(32'hbe224865),
	.w4(32'hbdfc9361),
	.w5(32'h3f939084),
	.w6(32'hbe7cdbb6),
	.w7(32'h3ec3c74a),
	.w8(32'hbf80e4b2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbee6428f),
	.w1(32'hbe6f3481),
	.w2(32'h3e67f15d),
	.w3(32'h3ebfff1a),
	.w4(32'hbcd89ee0),
	.w5(32'hbda96f1e),
	.w6(32'h3f7f3bd3),
	.w7(32'h3d3735d5),
	.w8(32'hbe707236),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f732759),
	.w1(32'hbe920cb6),
	.w2(32'h3c81be41),
	.w3(32'hbe8bc7b9),
	.w4(32'h3f2855e0),
	.w5(32'hbe0da462),
	.w6(32'h3ec9687a),
	.w7(32'h36fb29b4),
	.w8(32'hbe595626),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e193585),
	.w1(32'hbf22f3ed),
	.w2(32'h3e0dd769),
	.w3(32'hbf40d0bc),
	.w4(32'hbef32367),
	.w5(32'hbfca849c),
	.w6(32'h3f3dcbff),
	.w7(32'hbdb87597),
	.w8(32'hbd394fc7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf0667cd),
	.w1(32'hbf3159dd),
	.w2(32'hbfe5c5fb),
	.w3(32'hc0097c95),
	.w4(32'h3e93ee27),
	.w5(32'hbd944612),
	.w6(32'hbd95642e),
	.w7(32'h3e556d3e),
	.w8(32'hbf8cf831),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeac8697),
	.w1(32'hbe3a266c),
	.w2(32'h3eff6095),
	.w3(32'hbf825dc0),
	.w4(32'h3ea45a1c),
	.w5(32'h3b97fb63),
	.w6(32'h3f8c56a8),
	.w7(32'hbd894662),
	.w8(32'hbebb5fe3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdc273a6),
	.w1(32'hbf96ee8b),
	.w2(32'h3e3d7129),
	.w3(32'hbe278ab2),
	.w4(32'hbe93ddad),
	.w5(32'h3f0d4dcd),
	.w6(32'h3deec30c),
	.w7(32'hbe9c0a2a),
	.w8(32'hbfba3d13),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf2dd4b8),
	.w1(32'h3ea01dfb),
	.w2(32'hbd104ff0),
	.w3(32'h3fa72fc9),
	.w4(32'hbfb74485),
	.w5(32'hbe9c67a9),
	.w6(32'h3e4ef80e),
	.w7(32'h3dfeeb5b),
	.w8(32'h3ebe2c58),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe30234e),
	.w1(32'hbe8c4029),
	.w2(32'h3f5d45e9),
	.w3(32'h3c5460db),
	.w4(32'hbe2b4e25),
	.w5(32'h3ec470cc),
	.w6(32'hbe94cca6),
	.w7(32'hbdf90866),
	.w8(32'hc0222792),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1bab05),
	.w1(32'h3f0cb67c),
	.w2(32'hbdbc6cb8),
	.w3(32'h3eb412c9),
	.w4(32'hbf506536),
	.w5(32'hbeff7e2f),
	.w6(32'hbf08fca2),
	.w7(32'h3cd8013d),
	.w8(32'hbedbd0f6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe2f0931),
	.w1(32'hbe489a86),
	.w2(32'hbecc9cf2),
	.w3(32'h3ee9116d),
	.w4(32'hbe98fdfe),
	.w5(32'h3e081b2b),
	.w6(32'hbe9474f8),
	.w7(32'hbfd5f15b),
	.w8(32'hbe7f4e03),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbebd98a1),
	.w1(32'h3f62f7fd),
	.w2(32'hbf7d2895),
	.w3(32'hbf50e8ba),
	.w4(32'h3e2ca965),
	.w5(32'hbf062ceb),
	.w6(32'hbef0fe09),
	.w7(32'hbfd71839),
	.w8(32'h3dce6d52),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe87ade2),
	.w1(32'hbfbbdc0d),
	.w2(32'hbf0a7888),
	.w3(32'h3ebb9df0),
	.w4(32'h3e5aac41),
	.w5(32'h3f0bbfb5),
	.w6(32'hbf68159c),
	.w7(32'hbea2758f),
	.w8(32'h3d2fa69f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e9b74bf),
	.w1(32'h3e8ac7d5),
	.w2(32'h3f90e751),
	.w3(32'h3f3dfe79),
	.w4(32'h3e237279),
	.w5(32'h3f80de62),
	.w6(32'h3e0608b6),
	.w7(32'h3f832bcf),
	.w8(32'h3f120b41),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e0753e5),
	.w1(32'h3e9983b8),
	.w2(32'h3d89f413),
	.w3(32'h3eb1b9a4),
	.w4(32'h3ed37e60),
	.w5(32'h3f12df38),
	.w6(32'h3dbf5e83),
	.w7(32'h3ddffcac),
	.w8(32'h3f57c84f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e7bf864),
	.w1(32'h40102366),
	.w2(32'h3f11aa36),
	.w3(32'h3ef1001e),
	.w4(32'h3e3560f2),
	.w5(32'h3e9e14f7),
	.w6(32'h3e8d2384),
	.w7(32'h3f01e5bc),
	.w8(32'h3edbd90f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2b18ef),
	.w1(32'h3e5b19d0),
	.w2(32'h3db3c8f2),
	.w3(32'h3eebbc54),
	.w4(32'h3ee5b1f5),
	.w5(32'h3ed8a5cf),
	.w6(32'h3d6a1256),
	.w7(32'h3eba2725),
	.w8(32'h3e5cfb2f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ecc9cee),
	.w1(32'h3f476fc2),
	.w2(32'h3fa051bc),
	.w3(32'h3ec7a28a),
	.w4(32'h3eb01a61),
	.w5(32'h3e215ef4),
	.w6(32'h3efe7847),
	.w7(32'h3e22d7fb),
	.w8(32'h3fa8d2c8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f43836c),
	.w1(32'h3ea63f75),
	.w2(32'h3e275fa8),
	.w3(32'h3e8f4736),
	.w4(32'h3f333f49),
	.w5(32'h3eab9398),
	.w6(32'h3e6e8368),
	.w7(32'h3ea889ce),
	.w8(32'h3f0f51ac),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3de7a5ba),
	.w1(32'h3d173cde),
	.w2(32'h3e91dbd4),
	.w3(32'h3e376ce5),
	.w4(32'h3f119d08),
	.w5(32'h3f660496),
	.w6(32'h3e40cdd0),
	.w7(32'h3ef1537f),
	.w8(32'h3e1e6a79),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3db9489a),
	.w1(32'h3f0b9107),
	.w2(32'h3ec3d97c),
	.w3(32'h3e592353),
	.w4(32'h3e4fc21f),
	.w5(32'h3ea478a1),
	.w6(32'h3ee25eea),
	.w7(32'h3db9cbc5),
	.w8(32'h3f351b23),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3eb0f449),
	.w1(32'h3f54205a),
	.w2(32'h3e7ea085),
	.w3(32'h3f8e4715),
	.w4(32'h3f2e002a),
	.w5(32'h3f2059a5),
	.w6(32'h3ea66182),
	.w7(32'h3f212333),
	.w8(32'h3f10c6d4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dfa4d05),
	.w1(32'h3d942f74),
	.w2(32'h3f164374),
	.w3(32'h3e71e3e5),
	.w4(32'h3e6a8bb3),
	.w5(32'h3e8c9063),
	.w6(32'h3df47bb4),
	.w7(32'h3dc6662c),
	.w8(32'h3f396e1c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ebcbd71),
	.w1(32'h3e65377c),
	.w2(32'h3e87c252),
	.w3(32'h3e94e2ab),
	.w4(32'h39cc3d07),
	.w5(32'h3f2dfca6),
	.w6(32'h3f0d7a64),
	.w7(32'h3ea7a066),
	.w8(32'h3b162e88),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ef990d2),
	.w1(32'h3e832c92),
	.w2(32'h3fd28939),
	.w3(32'h3f01904f),
	.w4(32'h400b4d28),
	.w5(32'h3e3de5e5),
	.w6(32'h3ee180bc),
	.w7(32'h3e9eae74),
	.w8(32'h3da72d12),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f6c84c5),
	.w1(32'h3f2d0034),
	.w2(32'h3e781836),
	.w3(32'h3e8ad37a),
	.w4(32'h3de18fb2),
	.w5(32'h3e3cadb0),
	.w6(32'h3ea01beb),
	.w7(32'h3eee5522),
	.w8(32'h3e58d9d6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e545fdc),
	.w1(32'h3b8aa8e6),
	.w2(32'h3e596a6a),
	.w3(32'h38adcc6f),
	.w4(32'h3ec49c0b),
	.w5(32'h3ec4fd7b),
	.w6(32'h3eac3683),
	.w7(32'h3eeb97db),
	.w8(32'h3de53bcf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e4f67fe),
	.w1(32'h3ec900b7),
	.w2(32'h3e683747),
	.w3(32'h3ec69d64),
	.w4(32'h3de4a4c5),
	.w5(32'h3f4c705d),
	.w6(32'h3eb7207c),
	.w7(32'h3f226726),
	.w8(32'h3e894b28),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e99724e),
	.w1(32'h3e116e11),
	.w2(32'h3e794909),
	.w3(32'h3ef121cf),
	.w4(32'h3eb07278),
	.w5(32'h3f1eb2de),
	.w6(32'h3f0b3e3a),
	.w7(32'h3f011b10),
	.w8(32'h3ea6de78),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e006a1b),
	.w1(32'h3ebec948),
	.w2(32'h3f1fe011),
	.w3(32'h3f8a6620),
	.w4(32'h3d93e28d),
	.w5(32'h3edfffa2),
	.w6(32'h3e652b8d),
	.w7(32'h3e45c231),
	.w8(32'h3e0f6550),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dbeff8b),
	.w1(32'h3e5d76f0),
	.w2(32'h3dfbb46b),
	.w3(32'h3e04f737),
	.w4(32'h3e92c981),
	.w5(32'h3e5758d0),
	.w6(32'h3e767cce),
	.w7(32'h3e7e496b),
	.w8(32'h3f38c3d4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38950edd),
	.w1(32'h3eb2fc74),
	.w2(32'h3e677600),
	.w3(32'h3ea098c1),
	.w4(32'h3dcb04c8),
	.w5(32'h3f083dd7),
	.w6(32'h3f0e9307),
	.w7(32'h3e58b630),
	.w8(32'h3efcfbca),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e445fd1),
	.w1(32'h3c8fd50f),
	.w2(32'h3e5c01a9),
	.w3(32'h3ee5c857),
	.w4(32'h3e52320c),
	.w5(32'h3f11b590),
	.w6(32'h3f150f30),
	.w7(32'h3e50b8f2),
	.w8(32'h3f9c01a7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e80e2cc),
	.w1(32'h3f9ecb1b),
	.w2(32'h3e4b73ec),
	.w3(32'h3f05cdf1),
	.w4(32'h3e686d10),
	.w5(32'h3eb77815),
	.w6(32'h3e916830),
	.w7(32'h3ed61d07),
	.w8(32'h3f0bca39),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ec0aa35),
	.w1(32'h3e358cdc),
	.w2(32'h3e81498e),
	.w3(32'h3e45201b),
	.w4(32'h3e49a77a),
	.w5(32'h3f210ad4),
	.w6(32'h3ea58b58),
	.w7(32'h3ee5c5c9),
	.w8(32'h3e559125),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e394153),
	.w1(32'h3f4deded),
	.w2(32'h3d13c29e),
	.w3(32'h3e339f0c),
	.w4(32'h3ea3ace9),
	.w5(32'h3d6346c8),
	.w6(32'h3e9fcc40),
	.w7(32'h3f053b98),
	.w8(32'h3ef318ac),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dfbc9ed),
	.w1(32'h3d994d1c),
	.w2(32'h3e6ff5a8),
	.w3(32'h3bc8dd4e),
	.w4(32'h3e4cd583),
	.w5(32'h3d845520),
	.w6(32'h3e5f266c),
	.w7(32'h3e2f2527),
	.w8(32'h3c37bcbf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e2e2b93),
	.w1(32'h3f3caf64),
	.w2(32'h3e8c2aa8),
	.w3(32'h3e6062cf),
	.w4(32'h3f0d09eb),
	.w5(32'h3e9af10b),
	.w6(32'h3e139fbf),
	.w7(32'h3e497945),
	.w8(32'h3f19bfaa),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e7194ef),
	.w1(32'h3eaeeb16),
	.w2(32'h3f229dd8),
	.w3(32'h3eb4d442),
	.w4(32'h3e38b361),
	.w5(32'h3e5c1b21),
	.w6(32'h3ef82baa),
	.w7(32'h3e248153),
	.w8(32'h3ed02c5b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f9a6f16),
	.w1(32'h3e29dffd),
	.w2(32'h3ec1f2f8),
	.w3(32'h3ec742ca),
	.w4(32'h3f233d1a),
	.w5(32'h3e3bced5),
	.w6(32'h3dd7b17d),
	.w7(32'h3ef84cdd),
	.w8(32'h3f1feca1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f4c9741),
	.w1(32'h3e83abd6),
	.w2(32'h3e8db581),
	.w3(32'h3e047871),
	.w4(32'h3e68de1d),
	.w5(32'h3effa122),
	.w6(32'h3f22d5fe),
	.w7(32'h3f662008),
	.w8(32'h3d92217f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e89f500),
	.w1(32'hba98f84e),
	.w2(32'hba845032),
	.w3(32'h3e8c7317),
	.w4(32'h398d612a),
	.w5(32'hba51cae2),
	.w6(32'h3a25f798),
	.w7(32'h3afd96b5),
	.w8(32'h3ac53d59),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380b5cbe),
	.w1(32'h3c4ead0a),
	.w2(32'h3c669cef),
	.w3(32'h3a2d78a0),
	.w4(32'h3c1dc578),
	.w5(32'hbbaebe9d),
	.w6(32'hbb53e337),
	.w7(32'h3ac15309),
	.w8(32'hbbbd1093),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule