module layer_10_featuremap_493(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb530b40),
	.w1(32'hba26f5b1),
	.w2(32'h3abf8e32),
	.w3(32'hbb625bed),
	.w4(32'hbab8fc77),
	.w5(32'h3b762c59),
	.w6(32'hb8eaad3c),
	.w7(32'hbb6a4c51),
	.w8(32'h37720a5b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba568d34),
	.w1(32'hbac68c9f),
	.w2(32'hbb14fccc),
	.w3(32'hb9cf2aea),
	.w4(32'hbb170dfe),
	.w5(32'h3bda887e),
	.w6(32'hbaaaeebc),
	.w7(32'hbbcda9e4),
	.w8(32'h3b9028cd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad504a8),
	.w1(32'h3bff7eed),
	.w2(32'hbc82b240),
	.w3(32'h3c38e082),
	.w4(32'h3af026ac),
	.w5(32'h3d1d6ddd),
	.w6(32'h3bd479d4),
	.w7(32'hbc9cb23c),
	.w8(32'h3cd04146),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84c2d3),
	.w1(32'h392f0410),
	.w2(32'hbb84bfad),
	.w3(32'hbb954a21),
	.w4(32'hbb9315ec),
	.w5(32'hbc7adabe),
	.w6(32'hbadf9bfe),
	.w7(32'hbb6932de),
	.w8(32'hbc57c187),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55abd6),
	.w1(32'hbbe467b8),
	.w2(32'hbae1bd6f),
	.w3(32'hbbc63bbd),
	.w4(32'hbb9f4b73),
	.w5(32'h38ccf4b4),
	.w6(32'hbba7f76f),
	.w7(32'hbb669353),
	.w8(32'hbb0aa67c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f7fc1),
	.w1(32'hbadc6c54),
	.w2(32'h3ab2ac52),
	.w3(32'h39fc9a4f),
	.w4(32'h3ae1a31f),
	.w5(32'hbbd045a3),
	.w6(32'h3ab23cd5),
	.w7(32'h3b59d359),
	.w8(32'hbb7f35fd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea5bb3),
	.w1(32'hbbf2b42b),
	.w2(32'hbc9e5cfb),
	.w3(32'h3b804bd0),
	.w4(32'h3bcea83d),
	.w5(32'h3c87c979),
	.w6(32'hbbda2744),
	.w7(32'h39372166),
	.w8(32'h3c0fdf51),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca10cc2),
	.w1(32'h3c5ac893),
	.w2(32'h3d07fe04),
	.w3(32'hbc39efa3),
	.w4(32'h3cb1c01d),
	.w5(32'h3d318215),
	.w6(32'hbbfb6d59),
	.w7(32'h3c5f7685),
	.w8(32'h3cd6fb94),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04e0c3),
	.w1(32'hbb8faab8),
	.w2(32'hbc93c8a1),
	.w3(32'h3cc10b41),
	.w4(32'hbb8b9290),
	.w5(32'hbc99d952),
	.w6(32'h3c8317b2),
	.w7(32'hb9c2ef3d),
	.w8(32'hbcad8b6c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5197ad),
	.w1(32'h3b8cd6ca),
	.w2(32'h3bbeff65),
	.w3(32'h3bf467ed),
	.w4(32'h3bed2a1c),
	.w5(32'hba234588),
	.w6(32'hbc99930f),
	.w7(32'h3ba6153c),
	.w8(32'hba1f9b49),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b994c4b),
	.w1(32'hbab51f28),
	.w2(32'hbadd9682),
	.w3(32'hbb35fb20),
	.w4(32'h3b7350bd),
	.w5(32'h3c014e29),
	.w6(32'h3c283f92),
	.w7(32'h3b6665c7),
	.w8(32'h3bdeac43),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74e530),
	.w1(32'hbb7bf0d8),
	.w2(32'h3ae40948),
	.w3(32'h3b391548),
	.w4(32'hbb94ce19),
	.w5(32'hbb85d1c8),
	.w6(32'h3ad9b0d5),
	.w7(32'hb9d487f1),
	.w8(32'hbb2f98b2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0036ca),
	.w1(32'hbb9a602e),
	.w2(32'hbc031a8f),
	.w3(32'h380fbaf9),
	.w4(32'hbb66c4af),
	.w5(32'hba733382),
	.w6(32'h3b07004d),
	.w7(32'hbb92da45),
	.w8(32'h3a7ed479),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc790306),
	.w1(32'hbc85ccd0),
	.w2(32'hbc7821c0),
	.w3(32'hbc12ca8e),
	.w4(32'hbc40c6f4),
	.w5(32'hbbec0e88),
	.w6(32'h3bfa40dd),
	.w7(32'hbc0c3255),
	.w8(32'hbc6829c2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49e90c),
	.w1(32'h3ba249ea),
	.w2(32'h3b90ac17),
	.w3(32'hbc595fc2),
	.w4(32'h3b93c22e),
	.w5(32'h3c8b9ae3),
	.w6(32'hbc4c513a),
	.w7(32'hbb3e9146),
	.w8(32'h3bdf617c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaecd4),
	.w1(32'h39ef804f),
	.w2(32'hbbd2243b),
	.w3(32'hb850d3f7),
	.w4(32'hb9cc5a03),
	.w5(32'h3b833527),
	.w6(32'hbb2cd018),
	.w7(32'h3addd9fe),
	.w8(32'h3c031c7c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc258f3d),
	.w1(32'h3b99efa9),
	.w2(32'h3ba88506),
	.w3(32'hbc0632c4),
	.w4(32'hbb534c5e),
	.w5(32'hbc12c91c),
	.w6(32'h3a4ed7b4),
	.w7(32'hbb3bdfa1),
	.w8(32'hbb9cc91a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8879b86),
	.w1(32'h3c26edb5),
	.w2(32'h3b6253cd),
	.w3(32'h3a724da0),
	.w4(32'h3c07fe2e),
	.w5(32'h3bc493d5),
	.w6(32'hbc118333),
	.w7(32'hbb45c572),
	.w8(32'h3ae07f9d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97b8f7),
	.w1(32'hbb2471ea),
	.w2(32'hbc096417),
	.w3(32'hbbbd6459),
	.w4(32'hbc19b694),
	.w5(32'hbc8608cb),
	.w6(32'hbbdda684),
	.w7(32'hb9d95943),
	.w8(32'hbc261c6a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96af0d),
	.w1(32'h3aa78a27),
	.w2(32'h3c0457bf),
	.w3(32'hbaae13f7),
	.w4(32'h3bd84410),
	.w5(32'h3c89904e),
	.w6(32'hbbb4e37b),
	.w7(32'hbb29a22c),
	.w8(32'hbb139168),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb53c48),
	.w1(32'hb70f220b),
	.w2(32'hb98c22e0),
	.w3(32'h3bee8c65),
	.w4(32'hbb73ff3a),
	.w5(32'hbb50b087),
	.w6(32'h3a880dbf),
	.w7(32'hba55e2e7),
	.w8(32'hbb1754be),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c54d4),
	.w1(32'hbaea8324),
	.w2(32'h3b5e64ee),
	.w3(32'h3a732b24),
	.w4(32'hbad070bb),
	.w5(32'h3b3fd45d),
	.w6(32'hbaeb0612),
	.w7(32'h3b184804),
	.w8(32'h3c15ac28),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdf1c7),
	.w1(32'h3b81597a),
	.w2(32'h3bedf0dd),
	.w3(32'hbb4ca4bc),
	.w4(32'h3aaa188f),
	.w5(32'h3aead7e9),
	.w6(32'hbc208ec5),
	.w7(32'h3ae92f18),
	.w8(32'h3ba047ce),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c8d37),
	.w1(32'hbb83ac81),
	.w2(32'hbb3a32c1),
	.w3(32'h3c2c4866),
	.w4(32'h3beb89a9),
	.w5(32'h37199428),
	.w6(32'h3bde1eb2),
	.w7(32'h3bb4fbfa),
	.w8(32'h3b722554),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa83941),
	.w1(32'hbbee19b6),
	.w2(32'hbb174364),
	.w3(32'h3bbc4428),
	.w4(32'hbb9e7b31),
	.w5(32'h3b565c23),
	.w6(32'h3bba1ba6),
	.w7(32'hbbf31e41),
	.w8(32'hbc3c7789),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97e546),
	.w1(32'h3be223b4),
	.w2(32'h3bb57f9f),
	.w3(32'h3a6e8be3),
	.w4(32'h3b2d9bfb),
	.w5(32'hbbe816b0),
	.w6(32'hbb9c106b),
	.w7(32'hba830a29),
	.w8(32'h3b6fc3aa),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80065c),
	.w1(32'hbacffe4c),
	.w2(32'h3ae32502),
	.w3(32'h3b3562fc),
	.w4(32'hbb1fe84b),
	.w5(32'hbb70e2ec),
	.w6(32'hbaa0b71a),
	.w7(32'h3af2f9cd),
	.w8(32'hbc11a305),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba077f0),
	.w1(32'h3c26075a),
	.w2(32'h3b6e362f),
	.w3(32'h3b873ff7),
	.w4(32'h3c09620e),
	.w5(32'h3b01602d),
	.w6(32'hbc53cb9d),
	.w7(32'h3c0161af),
	.w8(32'h3bf7cd06),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e0dc3),
	.w1(32'hbbac4212),
	.w2(32'h3b842c29),
	.w3(32'h3ab1ab67),
	.w4(32'h3c5fab42),
	.w5(32'h3bb0a6b0),
	.w6(32'hbb05702f),
	.w7(32'h3c18f753),
	.w8(32'hbb32388b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f30cc),
	.w1(32'h3bf4f039),
	.w2(32'h3bac105d),
	.w3(32'h3bf5c35d),
	.w4(32'h3bee7d08),
	.w5(32'hbb0a71a9),
	.w6(32'h3b1ecc52),
	.w7(32'h3b9a23ee),
	.w8(32'h3aa74e76),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab80f9c),
	.w1(32'hbc33bd4a),
	.w2(32'hbbea687f),
	.w3(32'h3b6132c6),
	.w4(32'h3b67bf0a),
	.w5(32'hbbfef412),
	.w6(32'hbba78038),
	.w7(32'hbb097417),
	.w8(32'h3b8da4b0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19c4dc),
	.w1(32'h3be34210),
	.w2(32'h3a862a63),
	.w3(32'hbbf4d588),
	.w4(32'h3c850333),
	.w5(32'h3d1ca4fa),
	.w6(32'hbaf3bcf7),
	.w7(32'hbc551b92),
	.w8(32'h3c3c6966),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74c5bf),
	.w1(32'h3ab98879),
	.w2(32'hba2c7c92),
	.w3(32'hbabcb51b),
	.w4(32'h3b046de4),
	.w5(32'h3ca007f1),
	.w6(32'h3c77711b),
	.w7(32'hba0512a1),
	.w8(32'h3a661eda),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adab4eb),
	.w1(32'h3b6a93e6),
	.w2(32'hbbb31a3f),
	.w3(32'hba3632ac),
	.w4(32'hbb264f53),
	.w5(32'hbbaacb07),
	.w6(32'h39e0cd11),
	.w7(32'h3c1fe2a6),
	.w8(32'h3c123405),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57e339),
	.w1(32'hbc80becd),
	.w2(32'hbc70eebd),
	.w3(32'hbc017c72),
	.w4(32'hbd079507),
	.w5(32'hbd3f1d21),
	.w6(32'h3c335276),
	.w7(32'hbc8c024e),
	.w8(32'hbce563c4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2a5fd),
	.w1(32'h3b1ae317),
	.w2(32'h3b1bb6d4),
	.w3(32'hbd3ab18c),
	.w4(32'hbc082365),
	.w5(32'hbb439105),
	.w6(32'hbccfacd0),
	.w7(32'hbbac0850),
	.w8(32'h3ae3dfaf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaade24),
	.w1(32'hbc82594d),
	.w2(32'hbc48f7ba),
	.w3(32'hbb153041),
	.w4(32'hbc1b6dc4),
	.w5(32'hbb91ac65),
	.w6(32'hbb97dc28),
	.w7(32'hbb0f41f2),
	.w8(32'hbc822556),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87787f),
	.w1(32'hbc4d6135),
	.w2(32'hbc1f48f2),
	.w3(32'h3b969738),
	.w4(32'hbb207bad),
	.w5(32'h3c862804),
	.w6(32'h3af67302),
	.w7(32'hbc3dcad4),
	.w8(32'h38a4d373),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c2374),
	.w1(32'hbc10ac2a),
	.w2(32'hbc6dde3c),
	.w3(32'hbb707e47),
	.w4(32'hbc577d20),
	.w5(32'hbc4f0666),
	.w6(32'h3be9711e),
	.w7(32'h3b19239e),
	.w8(32'hbb534b8c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e974f),
	.w1(32'hbc1bc553),
	.w2(32'h3b2410b0),
	.w3(32'hbc0e7be2),
	.w4(32'h3a701bc5),
	.w5(32'h3c0a385a),
	.w6(32'hbabd7173),
	.w7(32'hba8be258),
	.w8(32'hbb1e5f6e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba864695),
	.w1(32'hbc5731ac),
	.w2(32'h3d0a5e82),
	.w3(32'h3ae27d31),
	.w4(32'hbc814cac),
	.w5(32'h3ba9aee3),
	.w6(32'h398a119b),
	.w7(32'hbcf34423),
	.w8(32'hbcfbeb20),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be71b98),
	.w1(32'hbb66a5a7),
	.w2(32'hbb5d34ef),
	.w3(32'h3c06cc94),
	.w4(32'hbc100ae4),
	.w5(32'hbbf682f7),
	.w6(32'hbaa2bb0b),
	.w7(32'hbc065971),
	.w8(32'hbbc1bd81),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30cae8),
	.w1(32'hbaf6ef68),
	.w2(32'hbad181c9),
	.w3(32'hbba747b9),
	.w4(32'h3bac8ce6),
	.w5(32'hbbeb4a24),
	.w6(32'hbaf25862),
	.w7(32'hbba742d5),
	.w8(32'hbbe6cc2c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc553447),
	.w1(32'h3baf732d),
	.w2(32'h3c007d14),
	.w3(32'hbc4755d8),
	.w4(32'h3b9bf26a),
	.w5(32'hbb2b5ae1),
	.w6(32'hbb7089ab),
	.w7(32'hba843ee1),
	.w8(32'hbb931050),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd046d5),
	.w1(32'hbb5e1a48),
	.w2(32'hbbacbad2),
	.w3(32'h3af8e818),
	.w4(32'hb9efbafd),
	.w5(32'hbbb530e9),
	.w6(32'h39d21e28),
	.w7(32'h3bff64f9),
	.w8(32'hbb9490b4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7000c),
	.w1(32'h3b8c9037),
	.w2(32'h39bcfe40),
	.w3(32'h3b771685),
	.w4(32'hbae9e57e),
	.w5(32'h3b8bb6b4),
	.w6(32'h3abb158c),
	.w7(32'hbb2b4c78),
	.w8(32'h3b253f71),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf413d0),
	.w1(32'hbbe1f0a8),
	.w2(32'hbbb625fe),
	.w3(32'hbc250d29),
	.w4(32'hbc1a2de9),
	.w5(32'hbbeb6a2b),
	.w6(32'hba1ae423),
	.w7(32'hba990f51),
	.w8(32'hbbad6edc),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd7ad6),
	.w1(32'h3b3e30a0),
	.w2(32'h3aa92715),
	.w3(32'hbc708a7e),
	.w4(32'hbbd7dfe4),
	.w5(32'h3a96f2d8),
	.w6(32'hbb375c03),
	.w7(32'hbb6254b2),
	.w8(32'hbb664696),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ebf59),
	.w1(32'hbc1ecbf8),
	.w2(32'hbc54042b),
	.w3(32'h3a491f2b),
	.w4(32'hbc498f74),
	.w5(32'hbd0cf11d),
	.w6(32'hbaeae845),
	.w7(32'hbb9c6efa),
	.w8(32'hbcaa17a3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d2dca),
	.w1(32'h3c4be91f),
	.w2(32'h3c752a79),
	.w3(32'hbc3136c1),
	.w4(32'h3c42bec6),
	.w5(32'h3c7acf78),
	.w6(32'hbc9b44f3),
	.w7(32'hbb97a72e),
	.w8(32'h3b5822e4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac80085),
	.w1(32'hba9ab822),
	.w2(32'h38b9ee38),
	.w3(32'h3c62e3e3),
	.w4(32'hb8eacf6d),
	.w5(32'hbbfa402c),
	.w6(32'h3c514ce5),
	.w7(32'hbb12d4af),
	.w8(32'hbb40dc91),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b808665),
	.w1(32'h3b909be1),
	.w2(32'hbb195860),
	.w3(32'h3b938a2c),
	.w4(32'hbb47a3f4),
	.w5(32'h3ad386ac),
	.w6(32'hb9cde567),
	.w7(32'h3c1a2fd4),
	.w8(32'hb9ca46a4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bddc46),
	.w1(32'h3ad0bbe3),
	.w2(32'h3c09475a),
	.w3(32'hbb1c6ee7),
	.w4(32'h3c3d9496),
	.w5(32'h3c22f3a0),
	.w6(32'hbc41e84a),
	.w7(32'h3b8ef1d9),
	.w8(32'h3c23027c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38d0f9),
	.w1(32'hbb812142),
	.w2(32'h3b1bb9e9),
	.w3(32'h3bcaf4ea),
	.w4(32'h3c01663b),
	.w5(32'h3c6f6f84),
	.w6(32'h3baf4c2f),
	.w7(32'h3b1df8ef),
	.w8(32'h39a88c6a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bee31),
	.w1(32'hbbf3dacf),
	.w2(32'hbb38fb4d),
	.w3(32'h3c126329),
	.w4(32'h3b6360bc),
	.w5(32'h3c0e45cb),
	.w6(32'h3b405ded),
	.w7(32'hba26dda6),
	.w8(32'h3c04cf5c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58e385),
	.w1(32'hbc2ff785),
	.w2(32'hbc11171c),
	.w3(32'hbc242846),
	.w4(32'h3a779aa2),
	.w5(32'h3c4529cc),
	.w6(32'hbb2b17b1),
	.w7(32'h3be30b44),
	.w8(32'hba35bc8b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1252a8),
	.w1(32'hbb2b352c),
	.w2(32'hbb6b6cbf),
	.w3(32'h3af3a5ad),
	.w4(32'hb82338da),
	.w5(32'hbaa79b4d),
	.w6(32'hbac9daa9),
	.w7(32'h3b534388),
	.w8(32'h396f972e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa41b72),
	.w1(32'hba10b22d),
	.w2(32'hbb032afb),
	.w3(32'h3b71458a),
	.w4(32'h3b4b743e),
	.w5(32'h3b939a01),
	.w6(32'hba724b7e),
	.w7(32'hbacb2a71),
	.w8(32'h3c77bfb4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a1f22),
	.w1(32'hbbb42666),
	.w2(32'hbba55ab1),
	.w3(32'hbb810a57),
	.w4(32'hba835b6f),
	.w5(32'hbc49325e),
	.w6(32'h3b5ac276),
	.w7(32'hb98c1373),
	.w8(32'hbc1a07ab),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb78f5),
	.w1(32'hbb236277),
	.w2(32'hbb09ae7b),
	.w3(32'h3b912fcf),
	.w4(32'hbc3ef0cd),
	.w5(32'hba82ef3f),
	.w6(32'h39ba8a54),
	.w7(32'h3b408441),
	.w8(32'hbc2cda94),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78e11b),
	.w1(32'hbb0f78e3),
	.w2(32'h3ab02cec),
	.w3(32'hbc4b74b9),
	.w4(32'hba4aee4c),
	.w5(32'hbadeb13e),
	.w6(32'hbbd94c5a),
	.w7(32'h395f281d),
	.w8(32'h3b8d8251),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba282ded),
	.w1(32'h3b8818c9),
	.w2(32'hbb17a0a7),
	.w3(32'h3ac808de),
	.w4(32'h3c22605a),
	.w5(32'h3b8bb093),
	.w6(32'hba363a13),
	.w7(32'h3b263b54),
	.w8(32'hba8f8b29),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d001),
	.w1(32'hbaabf288),
	.w2(32'h3bc6dc56),
	.w3(32'hbb1d1b5a),
	.w4(32'h3a83a216),
	.w5(32'h3bc89dc8),
	.w6(32'hbb3613f4),
	.w7(32'hbc783f6e),
	.w8(32'hbbf3a46f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a1557),
	.w1(32'h3a8d9ebc),
	.w2(32'hbb5b15e7),
	.w3(32'hbac92a53),
	.w4(32'h3ad38cbe),
	.w5(32'hbb7898bf),
	.w6(32'hbb5b202a),
	.w7(32'h3b2ec818),
	.w8(32'hb950251f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4605c7),
	.w1(32'h3bc2cec1),
	.w2(32'h3c743c07),
	.w3(32'hbb29bb6e),
	.w4(32'hba711e86),
	.w5(32'h3a67b474),
	.w6(32'h3bc3ec61),
	.w7(32'h3a0d88d1),
	.w8(32'hbb383f7e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2601cd),
	.w1(32'hbbe7e0df),
	.w2(32'hbc34f463),
	.w3(32'h3b6ff904),
	.w4(32'hbb44feb3),
	.w5(32'hbc18181f),
	.w6(32'h3b08323a),
	.w7(32'h3b9126e8),
	.w8(32'hbb3ab459),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30963e),
	.w1(32'hbaaed904),
	.w2(32'hbab2faaa),
	.w3(32'hbc2baf64),
	.w4(32'h3c1b25c1),
	.w5(32'h3c6ab74e),
	.w6(32'hbc00eeb0),
	.w7(32'h3b55abb3),
	.w8(32'h3b34a74d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b0c59),
	.w1(32'h3c100677),
	.w2(32'h3b4516bd),
	.w3(32'h3be53fb2),
	.w4(32'h3b320922),
	.w5(32'h3b6ed376),
	.w6(32'h3bfca379),
	.w7(32'hbbc51208),
	.w8(32'hbc205b39),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dc3e6),
	.w1(32'h3ac74c1a),
	.w2(32'h3bd28aeb),
	.w3(32'hbbb1af7f),
	.w4(32'hbc137f1e),
	.w5(32'hbb5eef84),
	.w6(32'hbbc6d115),
	.w7(32'hbbc71ae1),
	.w8(32'h3b00c613),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26391e),
	.w1(32'hba8c755b),
	.w2(32'hba08aaaf),
	.w3(32'hba613a18),
	.w4(32'hbba892f7),
	.w5(32'hbc1c475c),
	.w6(32'hbaf82488),
	.w7(32'hbba750ee),
	.w8(32'hbbee1215),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbc461),
	.w1(32'hbb0d292d),
	.w2(32'h38a415ac),
	.w3(32'hbc078c7a),
	.w4(32'hb828b055),
	.w5(32'hbc1643ac),
	.w6(32'hbbfeb5f7),
	.w7(32'h3a8f2963),
	.w8(32'h3a9b9c58),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a4d09),
	.w1(32'hbbdadfb4),
	.w2(32'h3ac7442a),
	.w3(32'hbb4ab4c0),
	.w4(32'hbc00d210),
	.w5(32'hbc6f6208),
	.w6(32'h3a5b4c4f),
	.w7(32'hba3c545a),
	.w8(32'hbba26df7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9c454),
	.w1(32'h3bb21680),
	.w2(32'hbb1e63e4),
	.w3(32'h3a1236db),
	.w4(32'h3aaae44a),
	.w5(32'h3ba078e5),
	.w6(32'h3b3cc95a),
	.w7(32'h3aab1017),
	.w8(32'hbab849ff),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc938e1),
	.w1(32'h3b17bb7b),
	.w2(32'hbb05e031),
	.w3(32'hb9ec5644),
	.w4(32'hbb45bf4a),
	.w5(32'h3b3e65e1),
	.w6(32'hb8994b6c),
	.w7(32'h3b83efa2),
	.w8(32'h3b5f880d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fbc66),
	.w1(32'h3b5a1c21),
	.w2(32'hb8fe5f8e),
	.w3(32'hbb1bdccb),
	.w4(32'hbb1ff576),
	.w5(32'h3baee2f6),
	.w6(32'h38a16f3c),
	.w7(32'hbba39e09),
	.w8(32'hbb8fd990),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2972e7),
	.w1(32'h3b141529),
	.w2(32'h3bcac1ce),
	.w3(32'h3b1aa489),
	.w4(32'h3b6b4a9a),
	.w5(32'h3c12f6a4),
	.w6(32'h3b7e3aed),
	.w7(32'hbb61cb4c),
	.w8(32'hb9f8a948),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4f0cd),
	.w1(32'hbb8675b7),
	.w2(32'hbba88d13),
	.w3(32'h3bb5c38b),
	.w4(32'hbaa75f13),
	.w5(32'h3b562c2f),
	.w6(32'h39cd03ad),
	.w7(32'h3a89f8b4),
	.w8(32'hba11072a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f6f0),
	.w1(32'h3a6dad45),
	.w2(32'hbc1ecf26),
	.w3(32'hbbad522e),
	.w4(32'hbc23dec2),
	.w5(32'h3cb8bc7c),
	.w6(32'hbbe40848),
	.w7(32'hbba8f331),
	.w8(32'hbbc564d8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57a3a9),
	.w1(32'h3b107920),
	.w2(32'h3abe832f),
	.w3(32'hbbacefdf),
	.w4(32'hbb2d9bbe),
	.w5(32'h3c4e9cef),
	.w6(32'h3ae1e75d),
	.w7(32'hbbc51034),
	.w8(32'h398851c9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc003fcc),
	.w1(32'hbc29b2c5),
	.w2(32'hbc81367c),
	.w3(32'h3add88fc),
	.w4(32'hbc090d47),
	.w5(32'hbc48c0da),
	.w6(32'h39ddc9bc),
	.w7(32'h3b814b26),
	.w8(32'hbae065b0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb95c96),
	.w1(32'h3bfddeae),
	.w2(32'h3c05ff91),
	.w3(32'hbc0874bc),
	.w4(32'h3bd26aa8),
	.w5(32'h3beb911d),
	.w6(32'hbb349c7d),
	.w7(32'h3b6aa71b),
	.w8(32'h3b5b6d35),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02bccd),
	.w1(32'hbb03a706),
	.w2(32'hba36638f),
	.w3(32'h3c3c9bab),
	.w4(32'hb98a108d),
	.w5(32'hbb8df76e),
	.w6(32'h3b91a9fa),
	.w7(32'h3b51c704),
	.w8(32'h3b54603a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0811c),
	.w1(32'hba98cc6d),
	.w2(32'hbae89233),
	.w3(32'hbb175d01),
	.w4(32'h3bd007ca),
	.w5(32'hbb3c73b0),
	.w6(32'hbb8e3905),
	.w7(32'h3c10dcf4),
	.w8(32'hb9d2f2f2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81be10),
	.w1(32'hb7b45ed2),
	.w2(32'hbb07317b),
	.w3(32'hb9fab620),
	.w4(32'hbabc1d77),
	.w5(32'hbb815a5b),
	.w6(32'h3a8354cd),
	.w7(32'hbbbaba15),
	.w8(32'h3b2652cf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922cc1),
	.w1(32'hbb6b62c5),
	.w2(32'h3b6f135b),
	.w3(32'h3b0eaaf7),
	.w4(32'hbaa99d55),
	.w5(32'hbb991c92),
	.w6(32'hba634098),
	.w7(32'hbb2585ee),
	.w8(32'h3bb5de01),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01da3b),
	.w1(32'hbadb1782),
	.w2(32'hbae3b14d),
	.w3(32'h3b9dc0eb),
	.w4(32'hbb5871f9),
	.w5(32'hbc2e209f),
	.w6(32'hb91883a9),
	.w7(32'hbbee4979),
	.w8(32'hbc03b2a0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae87e),
	.w1(32'h3baa69e7),
	.w2(32'hbc610e16),
	.w3(32'hbb49e495),
	.w4(32'hba07b5ad),
	.w5(32'h3d1cd635),
	.w6(32'h3aa3e3fe),
	.w7(32'hbc2657f5),
	.w8(32'h3a38c798),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2defa3),
	.w1(32'h395a3187),
	.w2(32'hbbd20b80),
	.w3(32'hbb8fe0e5),
	.w4(32'hbb532529),
	.w5(32'h3c89fa35),
	.w6(32'h3c2422c3),
	.w7(32'hbbb9d781),
	.w8(32'h3bcb8c5c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd18bdd),
	.w1(32'hbb268d06),
	.w2(32'h394cc3d4),
	.w3(32'hbae048fb),
	.w4(32'hbaf1d7f0),
	.w5(32'hbb45ee74),
	.w6(32'h3c1cb7cb),
	.w7(32'h3a2d9621),
	.w8(32'hbb60c766),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a894ef6),
	.w1(32'h3bb999ed),
	.w2(32'hbb28ce9a),
	.w3(32'hba8f70bc),
	.w4(32'h3b47c6bd),
	.w5(32'h3c4d5dc3),
	.w6(32'hbc177d43),
	.w7(32'h3a21bca0),
	.w8(32'h3c0864fb),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a7212),
	.w1(32'hbb9ebc5b),
	.w2(32'hbc000500),
	.w3(32'h3a501f23),
	.w4(32'hbb891465),
	.w5(32'hbbd490e4),
	.w6(32'h3aab8826),
	.w7(32'hbb5996eb),
	.w8(32'hbbb699bb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21771d),
	.w1(32'hbbd5280d),
	.w2(32'hbb5a06a2),
	.w3(32'hbc88d11c),
	.w4(32'hbc098b68),
	.w5(32'hbb8b4d72),
	.w6(32'hbc6e672f),
	.w7(32'hbc67294b),
	.w8(32'hbc3171ce),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acad907),
	.w1(32'hbc352da7),
	.w2(32'h3b4524d7),
	.w3(32'h3b902da7),
	.w4(32'hbb40a807),
	.w5(32'hbc6db767),
	.w6(32'hbbb1f566),
	.w7(32'h3a6b8e86),
	.w8(32'hbc1f8eea),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cf24a),
	.w1(32'hb9dc5c82),
	.w2(32'h3b150bf4),
	.w3(32'hbad75c93),
	.w4(32'hba11323b),
	.w5(32'h3b54a391),
	.w6(32'hbc42dc32),
	.w7(32'hbacd9f2e),
	.w8(32'hbaaef17b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25b58d),
	.w1(32'h3b094df2),
	.w2(32'hb912a50e),
	.w3(32'h3bb8c25a),
	.w4(32'hbc2b8145),
	.w5(32'hbb8ae9cc),
	.w6(32'h387b3518),
	.w7(32'h3ac886b1),
	.w8(32'hbb8ab252),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a871b83),
	.w1(32'hb8b0542e),
	.w2(32'hbbc599e5),
	.w3(32'hbaea7550),
	.w4(32'hbb6a9556),
	.w5(32'hbc4af06b),
	.w6(32'h3a10ba43),
	.w7(32'h3b481d66),
	.w8(32'hb8f35bb0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cea1d0),
	.w1(32'hbc070e09),
	.w2(32'hbb036cf9),
	.w3(32'hbc025768),
	.w4(32'hbc73b73b),
	.w5(32'hbc88f772),
	.w6(32'hbc1c4068),
	.w7(32'hbbd5b200),
	.w8(32'hbbb920df),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73f514),
	.w1(32'h3b574079),
	.w2(32'h3b1e3057),
	.w3(32'hbbadb599),
	.w4(32'h3b62f005),
	.w5(32'h3c10ca47),
	.w6(32'hbb845555),
	.w7(32'hbb4340f3),
	.w8(32'h3b8e9e8f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb771eef),
	.w1(32'hbbb522f9),
	.w2(32'h3b16305a),
	.w3(32'hbb3db08a),
	.w4(32'hbb993301),
	.w5(32'h39c9aba6),
	.w6(32'hba08f6d4),
	.w7(32'hba9a6e40),
	.w8(32'hba8a37f7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f50c5),
	.w1(32'hbbd0581f),
	.w2(32'hbb8513e1),
	.w3(32'hbbdafc5b),
	.w4(32'hbc07a40e),
	.w5(32'hbba08451),
	.w6(32'hbc1644ab),
	.w7(32'hbc39452a),
	.w8(32'hbc358a39),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe09119),
	.w1(32'h3b95e5a2),
	.w2(32'h3ad0404a),
	.w3(32'h3b03ae4d),
	.w4(32'hbb5644cb),
	.w5(32'h3adf65fe),
	.w6(32'hbbe25c2c),
	.w7(32'h3ac90a90),
	.w8(32'h3a4c64c0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac200a2),
	.w1(32'hbb07569d),
	.w2(32'h3bf6564b),
	.w3(32'hbb713bc0),
	.w4(32'hbb8624dc),
	.w5(32'hbb40c4de),
	.w6(32'h3aae188a),
	.w7(32'hba024e6c),
	.w8(32'h374e5663),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea0334),
	.w1(32'hbb829119),
	.w2(32'hbc17a90a),
	.w3(32'h3b86abb9),
	.w4(32'h38b7b32d),
	.w5(32'hbc33fe6e),
	.w6(32'hbc00d08b),
	.w7(32'hbbc401eb),
	.w8(32'hbc106f93),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd313ca),
	.w1(32'h3994d059),
	.w2(32'hbbcf4e2c),
	.w3(32'hbc297654),
	.w4(32'h3c32dd87),
	.w5(32'h3be1501c),
	.w6(32'hbb9f60c0),
	.w7(32'hba3f25d6),
	.w8(32'h3c600820),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ab266),
	.w1(32'hb9f633af),
	.w2(32'h3bfcc906),
	.w3(32'hbb86c26e),
	.w4(32'h3b9f1c5c),
	.w5(32'hbb45e7dd),
	.w6(32'hbb1a7b64),
	.w7(32'h3ba22301),
	.w8(32'hbabf4cb9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c404566),
	.w1(32'hbbcbe661),
	.w2(32'hbb892e69),
	.w3(32'h3bb066cc),
	.w4(32'hbbdd6f9e),
	.w5(32'hbb9ed3b3),
	.w6(32'hbac19242),
	.w7(32'hbacdba86),
	.w8(32'hbbe02f9b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f8ee5),
	.w1(32'h3a8ef2bc),
	.w2(32'hbb9f4a6d),
	.w3(32'hbba8f3ed),
	.w4(32'h3ba21096),
	.w5(32'h3aef7cdf),
	.w6(32'hbacf5d56),
	.w7(32'h38fb05e2),
	.w8(32'h3b0000e3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b481cde),
	.w1(32'hb9111648),
	.w2(32'h3c034d4a),
	.w3(32'hba55ed63),
	.w4(32'hbb0b9258),
	.w5(32'hba8a19c7),
	.w6(32'h3a1f34e1),
	.w7(32'h3b0ab441),
	.w8(32'hbb8f916b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8aa5),
	.w1(32'hbc3731a4),
	.w2(32'hbb74a296),
	.w3(32'h3a6f7d7f),
	.w4(32'hba7fd1ca),
	.w5(32'hbc27e64b),
	.w6(32'hbb3fc9d9),
	.w7(32'h3b9d9276),
	.w8(32'hbb5b5438),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd4f58),
	.w1(32'hb9fb7488),
	.w2(32'h3a8dd494),
	.w3(32'hbbbca8fa),
	.w4(32'h3be7bc4f),
	.w5(32'h3b785fe0),
	.w6(32'hbc0fea40),
	.w7(32'h3b8e6c58),
	.w8(32'h3bdc1051),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb1395),
	.w1(32'hbb66fdda),
	.w2(32'hbb734c6c),
	.w3(32'h3a28916e),
	.w4(32'h390d6276),
	.w5(32'hbc147c9c),
	.w6(32'h3aa865a7),
	.w7(32'hba7995b0),
	.w8(32'hba706845),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f8cb),
	.w1(32'h3ae56a64),
	.w2(32'h3b40cdba),
	.w3(32'h3bc737b4),
	.w4(32'hbaf63faa),
	.w5(32'hbb31fad0),
	.w6(32'h39facc24),
	.w7(32'h3b37fef2),
	.w8(32'hb999e045),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a180),
	.w1(32'h3b473933),
	.w2(32'hbaf5b491),
	.w3(32'hbb1387af),
	.w4(32'hbbdd06bd),
	.w5(32'hbc392028),
	.w6(32'hbb5a69df),
	.w7(32'h3b17569b),
	.w8(32'hb856fbb2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac54f64),
	.w1(32'hbb237f51),
	.w2(32'h3b20e94e),
	.w3(32'hbbe5a7ca),
	.w4(32'h3977be7e),
	.w5(32'hbb8679f0),
	.w6(32'hbc0bcb01),
	.w7(32'hba7b10d5),
	.w8(32'hbbda4d1d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a178a),
	.w1(32'hbb3b6c96),
	.w2(32'hbbdc84d0),
	.w3(32'hbb6bc24a),
	.w4(32'hbb37c00a),
	.w5(32'hbb31abc6),
	.w6(32'hbc15820c),
	.w7(32'hbbaa3dce),
	.w8(32'hb8099c1c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61884c),
	.w1(32'hb91fecf8),
	.w2(32'h3b64da6c),
	.w3(32'hbbaf6144),
	.w4(32'h392706d3),
	.w5(32'hba182485),
	.w6(32'h3b97290c),
	.w7(32'h3a540094),
	.w8(32'h3a8b0233),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a8ea7),
	.w1(32'h3a0794ff),
	.w2(32'hbb37a21a),
	.w3(32'hbb7369b4),
	.w4(32'h3a6f33fa),
	.w5(32'hbad3ee19),
	.w6(32'hba29d067),
	.w7(32'h3b8d01ad),
	.w8(32'h3bdd2093),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2c906),
	.w1(32'hbc2a26be),
	.w2(32'hbade2ff8),
	.w3(32'hbbe6e093),
	.w4(32'hba1e49ac),
	.w5(32'hbc0344ca),
	.w6(32'hbbbcd609),
	.w7(32'h3c55711c),
	.w8(32'hbb97f583),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f2bb),
	.w1(32'hbb008d94),
	.w2(32'hbb99d238),
	.w3(32'h3b75d527),
	.w4(32'hbc22b4c4),
	.w5(32'h3aab32bc),
	.w6(32'hbb61342e),
	.w7(32'hbaecf4b1),
	.w8(32'hbb936d0b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63fe75),
	.w1(32'h3b92d3bd),
	.w2(32'h3bad440d),
	.w3(32'h38194768),
	.w4(32'hbacea684),
	.w5(32'h3b8266c4),
	.w6(32'hba7aafdd),
	.w7(32'hbbb9cc07),
	.w8(32'hbc30f4bd),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0930e7),
	.w1(32'hbb9245f6),
	.w2(32'hbc130d2f),
	.w3(32'hbb81cc0a),
	.w4(32'hbba07c31),
	.w5(32'hbb5a72b0),
	.w6(32'hbba006c1),
	.w7(32'hbb9d92d6),
	.w8(32'h39bf0bb7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b778a),
	.w1(32'hbc11cdb6),
	.w2(32'h3ba5bd64),
	.w3(32'hbb8029d3),
	.w4(32'hbade0834),
	.w5(32'hbb69e82d),
	.w6(32'hbbca8141),
	.w7(32'h39811f33),
	.w8(32'hb9944cbe),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd73f97),
	.w1(32'hba65769c),
	.w2(32'hbb8be2c2),
	.w3(32'h39b8e225),
	.w4(32'hbbc73e8d),
	.w5(32'hbc1f51dd),
	.w6(32'hbb0dd44c),
	.w7(32'h3ac49d44),
	.w8(32'h3a8bd136),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e5336),
	.w1(32'hbc6e3a89),
	.w2(32'h3a9279b7),
	.w3(32'hbb5501e3),
	.w4(32'hbc101318),
	.w5(32'hbca925a0),
	.w6(32'hbb8106d9),
	.w7(32'h3b85fe9a),
	.w8(32'h395919e7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06c0c8),
	.w1(32'hbc2202c7),
	.w2(32'h3c34691a),
	.w3(32'h3b544b49),
	.w4(32'h3b3e9b2b),
	.w5(32'hbbef08e2),
	.w6(32'hbc4d9ee6),
	.w7(32'h3c039ea2),
	.w8(32'h3b4544ed),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee1750),
	.w1(32'hbabda6cc),
	.w2(32'hbb956bfe),
	.w3(32'h3be80709),
	.w4(32'hba9a2587),
	.w5(32'hbca7b920),
	.w6(32'hbb014e3c),
	.w7(32'hbb1c42c4),
	.w8(32'hbbfe2187),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb512249),
	.w1(32'hbc099753),
	.w2(32'hbbcd7a69),
	.w3(32'hbc0ede55),
	.w4(32'hbc31ffa1),
	.w5(32'hbc611375),
	.w6(32'hbbcd127b),
	.w7(32'hbc48e4f2),
	.w8(32'hbc2b1570),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03a1af),
	.w1(32'h3b3e6ed7),
	.w2(32'h3bf62f02),
	.w3(32'hbc3c149f),
	.w4(32'hba9b759c),
	.w5(32'hbabbde8d),
	.w6(32'hbc60ce4e),
	.w7(32'hbbc6f741),
	.w8(32'h3b3b0e7c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac566ce),
	.w1(32'hbb26836a),
	.w2(32'h3a8eb4d0),
	.w3(32'h3aeb1323),
	.w4(32'hbbb06ab6),
	.w5(32'h3c428877),
	.w6(32'hbbad4a1f),
	.w7(32'hbb87a1c5),
	.w8(32'hba7db95d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eee50),
	.w1(32'h3b6fd0d9),
	.w2(32'hbb182e11),
	.w3(32'hba85d295),
	.w4(32'hba2fb160),
	.w5(32'h3c4def5b),
	.w6(32'hba496ace),
	.w7(32'hbacbf6ee),
	.w8(32'h3b36bb8f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e05de),
	.w1(32'hbaa5028d),
	.w2(32'hbb78c6f2),
	.w3(32'h3a7487e2),
	.w4(32'h3ad286ce),
	.w5(32'h3be0b53e),
	.w6(32'h3c1606ce),
	.w7(32'hbb89eb5e),
	.w8(32'h3b599d83),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce007),
	.w1(32'hbb1d58ba),
	.w2(32'hba954d8a),
	.w3(32'hbba6cb35),
	.w4(32'hb994bd1f),
	.w5(32'hbb89e4cd),
	.w6(32'hbacc34b3),
	.w7(32'hbaa96df0),
	.w8(32'hbc4ee54c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2de799),
	.w1(32'hbbca635f),
	.w2(32'hbae43a7f),
	.w3(32'h3be58d7b),
	.w4(32'hba1f82b3),
	.w5(32'hbaef89ec),
	.w6(32'hba821b19),
	.w7(32'h3b1fcfde),
	.w8(32'h3bb8e5b5),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42770b),
	.w1(32'h3b3c46b8),
	.w2(32'h3b3cdeca),
	.w3(32'hbb8e4bc0),
	.w4(32'hba1a6260),
	.w5(32'hba8abf24),
	.w6(32'hbb0c5d67),
	.w7(32'h3c0e19ac),
	.w8(32'hbb31d0d8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb530a83),
	.w1(32'h3a23fe2a),
	.w2(32'hbb080f7d),
	.w3(32'h3b0ef9aa),
	.w4(32'hbb8a7ab0),
	.w5(32'h3bd1abb5),
	.w6(32'hbb30b2fd),
	.w7(32'hbbb04154),
	.w8(32'hbb43a716),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cede7),
	.w1(32'h3bb24f1a),
	.w2(32'h3af12182),
	.w3(32'h3b260664),
	.w4(32'hbaadb586),
	.w5(32'h3bc70b34),
	.w6(32'h3b2d6067),
	.w7(32'h3b6c54a5),
	.w8(32'hbbafb2d9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb6d23),
	.w1(32'h3acdce38),
	.w2(32'hbb80f5c3),
	.w3(32'hba363833),
	.w4(32'h3b5e9492),
	.w5(32'hba874951),
	.w6(32'hbbcb0bc6),
	.w7(32'h3bc94f29),
	.w8(32'hba8260ac),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bfe93),
	.w1(32'hba110318),
	.w2(32'h38edacfc),
	.w3(32'hbb930730),
	.w4(32'h3ac162c9),
	.w5(32'hbb5d560b),
	.w6(32'hbb937d54),
	.w7(32'h3bf2d84d),
	.w8(32'h39fc7bab),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2defe),
	.w1(32'hba42d2da),
	.w2(32'hbb0b7e41),
	.w3(32'h3b5282c9),
	.w4(32'hba9a4ea1),
	.w5(32'hbb19556f),
	.w6(32'h3a622da4),
	.w7(32'h3b816daa),
	.w8(32'h3c189806),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0878b9),
	.w1(32'hbc23b676),
	.w2(32'hbbb8b09c),
	.w3(32'hbae4cc62),
	.w4(32'hbba398f1),
	.w5(32'hbbddf388),
	.w6(32'h3bbb95ba),
	.w7(32'hbabdadee),
	.w8(32'hbb08a8db),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d390f),
	.w1(32'h3b108a66),
	.w2(32'hbc1886a5),
	.w3(32'hbaf6e75b),
	.w4(32'h3b142204),
	.w5(32'hbbd5edce),
	.w6(32'hbb496857),
	.w7(32'h3ae876f1),
	.w8(32'hbbe446e9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab301bc),
	.w1(32'hba93a719),
	.w2(32'hbbd19334),
	.w3(32'hbc0d00e5),
	.w4(32'h3c0065a0),
	.w5(32'hbb82c509),
	.w6(32'hbb874acf),
	.w7(32'hbb654d43),
	.w8(32'h3b0abaa8),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bda7a),
	.w1(32'h39181a87),
	.w2(32'h3bde246e),
	.w3(32'h3b231deb),
	.w4(32'h3b7c1da8),
	.w5(32'h3a75a65b),
	.w6(32'hbb526971),
	.w7(32'h3babcbd9),
	.w8(32'h3ba2f188),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75988a),
	.w1(32'h3b5594fd),
	.w2(32'h3ae1b71d),
	.w3(32'h3b4bc2ff),
	.w4(32'h3c10cc42),
	.w5(32'hbb23aa54),
	.w6(32'hbb7aab15),
	.w7(32'h3b8bfd87),
	.w8(32'h3b596821),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0a949),
	.w1(32'h3aa7f72b),
	.w2(32'hba2c8215),
	.w3(32'h3b2c5fb2),
	.w4(32'hbab9ba0f),
	.w5(32'h3ac84231),
	.w6(32'h386a14d8),
	.w7(32'h3b895c49),
	.w8(32'h3a66fc97),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98121d0),
	.w1(32'hbb27dccf),
	.w2(32'hbba04f03),
	.w3(32'h3a00cb3a),
	.w4(32'hba9e753f),
	.w5(32'h3b2d58d2),
	.w6(32'hbb16a3cc),
	.w7(32'hbb3c703d),
	.w8(32'hbafa7cf5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb2bd5),
	.w1(32'hbb9d4561),
	.w2(32'hba8ab9ba),
	.w3(32'hbb699bed),
	.w4(32'hbb81e389),
	.w5(32'hbc085193),
	.w6(32'hbc175592),
	.w7(32'h3aeaf9fc),
	.w8(32'h3b3e151e),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b278764),
	.w1(32'hbb1cfd2a),
	.w2(32'hbab59a19),
	.w3(32'hba9c5a0a),
	.w4(32'h3a4b3b13),
	.w5(32'hbc4b60cd),
	.w6(32'hbb270805),
	.w7(32'h3b41cd13),
	.w8(32'hbb53951c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecf15d),
	.w1(32'hbbfe31dd),
	.w2(32'hbba6f598),
	.w3(32'hbb15f146),
	.w4(32'hbb71d179),
	.w5(32'hbc1eae94),
	.w6(32'hbabd85c6),
	.w7(32'h39f5a102),
	.w8(32'hba995f9a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b62f8),
	.w1(32'hbb2260fb),
	.w2(32'hbbd15665),
	.w3(32'hba9afa93),
	.w4(32'hbb324d3f),
	.w5(32'hbc109d27),
	.w6(32'hbaf115d6),
	.w7(32'hbbc82406),
	.w8(32'hbb329979),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae5b5),
	.w1(32'hbb06ead9),
	.w2(32'h3b599502),
	.w3(32'hbb48eab9),
	.w4(32'h3a417753),
	.w5(32'hbbe684e5),
	.w6(32'hba95def8),
	.w7(32'hb9d7cecd),
	.w8(32'h3bf5d7e9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a6031),
	.w1(32'hbb45ddf1),
	.w2(32'hbaf6b305),
	.w3(32'hbb7c1183),
	.w4(32'h3b715d27),
	.w5(32'h3b09ce3f),
	.w6(32'hbbf52b16),
	.w7(32'h3b691497),
	.w8(32'h3b86378c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb027f7f),
	.w1(32'h3c40da29),
	.w2(32'hbbe7d924),
	.w3(32'h3b02ef51),
	.w4(32'h3c4efa67),
	.w5(32'hbbbcf9ed),
	.w6(32'hb9def005),
	.w7(32'hbb5e17fb),
	.w8(32'h3bc2692f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b476a73),
	.w1(32'hba9136a1),
	.w2(32'hbafa8437),
	.w3(32'hbb9caea5),
	.w4(32'hbc0307b4),
	.w5(32'hbc19eb8c),
	.w6(32'hbaefdeaf),
	.w7(32'h3ab8a5e9),
	.w8(32'hbb4920ed),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b977024),
	.w1(32'hbad37ea8),
	.w2(32'h3aaf2e06),
	.w3(32'h3ac7c65f),
	.w4(32'hbb91991d),
	.w5(32'hbb6670f9),
	.w6(32'hbb31600c),
	.w7(32'hbba370a7),
	.w8(32'hbb7c6d77),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba44862),
	.w1(32'h397a7166),
	.w2(32'h398b2ab4),
	.w3(32'h3bc4bc20),
	.w4(32'hbb745e28),
	.w5(32'hbc1ada7c),
	.w6(32'h39caff74),
	.w7(32'hbab8b32d),
	.w8(32'hbba95946),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabea6b2),
	.w1(32'hbb2ea0bb),
	.w2(32'h3b4f42c4),
	.w3(32'h38c952a1),
	.w4(32'h3be7c152),
	.w5(32'hba270cf8),
	.w6(32'hbaf3781a),
	.w7(32'hba883038),
	.w8(32'h3b695520),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95d970),
	.w1(32'hbc193ab4),
	.w2(32'hbb45b0c2),
	.w3(32'hbac40d26),
	.w4(32'hbbaf976b),
	.w5(32'hbc0b57ae),
	.w6(32'h3b1b79e8),
	.w7(32'h3b1f4d38),
	.w8(32'hbb347d9c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae269ab),
	.w1(32'hbbe251ea),
	.w2(32'hb71e12fd),
	.w3(32'hbbb4d240),
	.w4(32'hba91b749),
	.w5(32'hbb4256e4),
	.w6(32'hbc021b18),
	.w7(32'h3b13a641),
	.w8(32'h3aa5ae9f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b770f),
	.w1(32'h3aa62586),
	.w2(32'h3b0e1f79),
	.w3(32'hba94bab1),
	.w4(32'hba9a5a30),
	.w5(32'h3c69228a),
	.w6(32'h39d0e0e3),
	.w7(32'hbaabcc6f),
	.w8(32'hbbe95ee7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8fb31),
	.w1(32'h3bc7b8b3),
	.w2(32'hbb465773),
	.w3(32'hbb0406bc),
	.w4(32'h3b4ccdf7),
	.w5(32'h3c93605a),
	.w6(32'hbb8b12e0),
	.w7(32'hbaa5fc2c),
	.w8(32'h3b579559),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed3f6e),
	.w1(32'h3b100dfb),
	.w2(32'hba62d969),
	.w3(32'hbb173d49),
	.w4(32'hbc027a7d),
	.w5(32'hbc14e01e),
	.w6(32'h3bc27e29),
	.w7(32'hba9c8ad2),
	.w8(32'hbb72c870),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba210430),
	.w1(32'hbb24c7e5),
	.w2(32'hbbc367c0),
	.w3(32'hbb6bf7d5),
	.w4(32'h3c123aef),
	.w5(32'hbc18aef4),
	.w6(32'hbb97470c),
	.w7(32'h3c8309c7),
	.w8(32'hba812031),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe699f),
	.w1(32'h3b25e9d1),
	.w2(32'hbb32244d),
	.w3(32'hbbd8d9d1),
	.w4(32'h3b5ff75f),
	.w5(32'h3ba7ea9b),
	.w6(32'hbc083607),
	.w7(32'hbaf703ee),
	.w8(32'hbb894031),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8671d6),
	.w1(32'h3c140e91),
	.w2(32'h3aab43a2),
	.w3(32'h3b0e2e25),
	.w4(32'h39a8f0a6),
	.w5(32'h3c7f9f3d),
	.w6(32'h3ac8d5f8),
	.w7(32'hbb422614),
	.w8(32'h3bb5eb1e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb79506),
	.w1(32'h39f23b5b),
	.w2(32'hbb42801c),
	.w3(32'h3bd3df2b),
	.w4(32'hbb1c7387),
	.w5(32'h3cfd62fe),
	.w6(32'h3c805634),
	.w7(32'hbbf7b297),
	.w8(32'h3a7c0143),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb569f87),
	.w1(32'h36b58c8d),
	.w2(32'h39d2f0ca),
	.w3(32'h3ba55f92),
	.w4(32'h3b33ba56),
	.w5(32'h3b39171e),
	.w6(32'h3c47d712),
	.w7(32'h3bd5274f),
	.w8(32'h3ba106b3),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2027c2),
	.w1(32'h3bdcb172),
	.w2(32'hba34df1e),
	.w3(32'h3b421cfc),
	.w4(32'hbb6ef75d),
	.w5(32'h3cac9443),
	.w6(32'h3b2c0c8b),
	.w7(32'hbc348f39),
	.w8(32'hbb056f53),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47b6cb),
	.w1(32'hbbd69ab1),
	.w2(32'hb9dbb2ec),
	.w3(32'h3ac93de9),
	.w4(32'h3a0bffae),
	.w5(32'hbb05364c),
	.w6(32'h3bbb418a),
	.w7(32'h39f591ca),
	.w8(32'h39db8898),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb12d08),
	.w1(32'hbae8c000),
	.w2(32'h3bc0d87f),
	.w3(32'h39148df0),
	.w4(32'hbb922afa),
	.w5(32'hbb311880),
	.w6(32'hbbddb8ef),
	.w7(32'hbb468bd7),
	.w8(32'hbaa608d5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d9bc7),
	.w1(32'h3a23b8ce),
	.w2(32'hbbe11f24),
	.w3(32'h3aca424c),
	.w4(32'hba9ae444),
	.w5(32'hbb1bc074),
	.w6(32'hbb965401),
	.w7(32'hbbb4ed6e),
	.w8(32'hbc3faa35),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8113eb),
	.w1(32'h3b0afb7b),
	.w2(32'h3b89f0fe),
	.w3(32'hbb578cbb),
	.w4(32'hbb52c168),
	.w5(32'h3c012740),
	.w6(32'hbb92a222),
	.w7(32'hbbea00df),
	.w8(32'hbb6a7017),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de3040),
	.w1(32'h389bedcc),
	.w2(32'hbb8e9957),
	.w3(32'h3bacbce6),
	.w4(32'h38cc1a04),
	.w5(32'hbc352058),
	.w6(32'h39868745),
	.w7(32'h3b9c2baf),
	.w8(32'h3b67fac7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4288e),
	.w1(32'h3b9b2847),
	.w2(32'h3b89c174),
	.w3(32'hbb0ea5ff),
	.w4(32'h3b8c6634),
	.w5(32'hba86b9b6),
	.w6(32'hbb5a0d8e),
	.w7(32'h3b57c77d),
	.w8(32'h3ba72561),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a063284),
	.w1(32'hb910f504),
	.w2(32'hba327473),
	.w3(32'h3beb829c),
	.w4(32'h3b1687bf),
	.w5(32'hbb66dea1),
	.w6(32'h3b4e0437),
	.w7(32'hbb167e42),
	.w8(32'h3b2f7449),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ac619),
	.w1(32'h3addde85),
	.w2(32'h3b252ca4),
	.w3(32'hbb883d46),
	.w4(32'hbb4af3f5),
	.w5(32'hbb21e81f),
	.w6(32'h3bc9347b),
	.w7(32'hbb512bef),
	.w8(32'hbbfea0f4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934a2f),
	.w1(32'hbc1f0620),
	.w2(32'hbaaa0557),
	.w3(32'h3af41d44),
	.w4(32'h3b6bd8b9),
	.w5(32'hbc19abc6),
	.w6(32'hb9b75d58),
	.w7(32'h3c4aa933),
	.w8(32'h3c0960d2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b944aee),
	.w1(32'hbaeb37d1),
	.w2(32'h3b3386c9),
	.w3(32'hbaab79e3),
	.w4(32'hbb6792f4),
	.w5(32'h3a176559),
	.w6(32'hbbbc277c),
	.w7(32'hbbccbeb5),
	.w8(32'hbc15f3af),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea46ba),
	.w1(32'hbb1463af),
	.w2(32'hbb8dc9dd),
	.w3(32'h3b349551),
	.w4(32'h3a1e3232),
	.w5(32'hbc26037b),
	.w6(32'hbb301784),
	.w7(32'h3c352119),
	.w8(32'h3afa43df),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a996b4b),
	.w1(32'hba97e86e),
	.w2(32'h3b174df2),
	.w3(32'hbbc81905),
	.w4(32'h3b0c2161),
	.w5(32'h3b996d63),
	.w6(32'hbb93460d),
	.w7(32'h3be4706a),
	.w8(32'h3c27c5a7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a204c),
	.w1(32'h3baec89b),
	.w2(32'h3b04a952),
	.w3(32'hbb30a249),
	.w4(32'hbbc1423d),
	.w5(32'hbad2e8a1),
	.w6(32'h3b350bf6),
	.w7(32'hbb59e0a8),
	.w8(32'h38dea505),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba56cb5),
	.w1(32'h3b5f214b),
	.w2(32'hbbfa322b),
	.w3(32'hbba42f25),
	.w4(32'hba585607),
	.w5(32'h3c7e5145),
	.w6(32'hb7de6e76),
	.w7(32'hbbd9ccdf),
	.w8(32'h3a8f0a98),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc436107),
	.w1(32'h3bc1782c),
	.w2(32'hbb51f1aa),
	.w3(32'hbbd7114d),
	.w4(32'h3bd4ed7a),
	.w5(32'h3cb1f3d8),
	.w6(32'h3ae4499b),
	.w7(32'hba28e51f),
	.w8(32'hbacc0fe4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38336192),
	.w1(32'h3b761980),
	.w2(32'hbc1da3ee),
	.w3(32'hbbaf4da4),
	.w4(32'h3b4db996),
	.w5(32'h3d01517b),
	.w6(32'h3c049d4c),
	.w7(32'hbb9d063d),
	.w8(32'h3b178fa5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc442f30),
	.w1(32'hbb6202b2),
	.w2(32'hbaad7022),
	.w3(32'hbb5f4e3b),
	.w4(32'hbad1b034),
	.w5(32'hba8845ac),
	.w6(32'hb95345f1),
	.w7(32'h3a40d3eb),
	.w8(32'h3a9aae8f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22a2ba),
	.w1(32'hba97e339),
	.w2(32'h3a86a959),
	.w3(32'hbb77efaf),
	.w4(32'hbc216fb7),
	.w5(32'h3a3368fe),
	.w6(32'hbbacffec),
	.w7(32'hbbf8702a),
	.w8(32'hbbbbb9f7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24a020),
	.w1(32'h3b300fe3),
	.w2(32'hbac42d8a),
	.w3(32'h3aba369b),
	.w4(32'h3a2fbdfb),
	.w5(32'h3aecabd4),
	.w6(32'h3a5fa49f),
	.w7(32'hba9fb632),
	.w8(32'hbb1a7802),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd13852),
	.w1(32'h3c26ed02),
	.w2(32'hbc5a1a18),
	.w3(32'hbbdf1a75),
	.w4(32'h3ba88588),
	.w5(32'h3c131427),
	.w6(32'hba1936dc),
	.w7(32'h39c35b8a),
	.w8(32'h3b353d09),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaede376),
	.w1(32'hbb251bdb),
	.w2(32'hbc31db2d),
	.w3(32'hbbe180f1),
	.w4(32'hbb977775),
	.w5(32'hbc2a08b1),
	.w6(32'h3c511e6f),
	.w7(32'hba6b5b27),
	.w8(32'hbbafc676),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8880a),
	.w1(32'hbbaf7145),
	.w2(32'hbae14553),
	.w3(32'hbb92c35a),
	.w4(32'hbb97d46e),
	.w5(32'hbb4ac1fd),
	.w6(32'hbb9964b4),
	.w7(32'hbb33797f),
	.w8(32'hbbbf34ff),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2313b),
	.w1(32'h3b2f14c7),
	.w2(32'hbba0cdb0),
	.w3(32'hbb9879bf),
	.w4(32'h3a373d75),
	.w5(32'h3bcf87a1),
	.w6(32'hbc500230),
	.w7(32'hbb6f36d1),
	.w8(32'hbb16257b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a31a9),
	.w1(32'hbb184037),
	.w2(32'hbb989a30),
	.w3(32'h3b061e5c),
	.w4(32'h3a849b78),
	.w5(32'h3943cc87),
	.w6(32'h3b8c1fc7),
	.w7(32'h3baa52f1),
	.w8(32'h3bc5aa20),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4411f5),
	.w1(32'h3c0476ec),
	.w2(32'h3b59d569),
	.w3(32'hbafa713c),
	.w4(32'h3bb2a612),
	.w5(32'h3bf573c1),
	.w6(32'h3b21044a),
	.w7(32'h3afc99e6),
	.w8(32'h3b5a2a6e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a339c),
	.w1(32'hbbbd7331),
	.w2(32'h3b8163af),
	.w3(32'h3bc95659),
	.w4(32'hbb839c9e),
	.w5(32'hbc1412a8),
	.w6(32'h3b11cf1f),
	.w7(32'h3b2f7350),
	.w8(32'hbb6a3ce3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddb5e5),
	.w1(32'hbbbe6755),
	.w2(32'h3ac1495d),
	.w3(32'h3ba7fe8a),
	.w4(32'hba5d83e1),
	.w5(32'hbbbd8d48),
	.w6(32'hbbf09751),
	.w7(32'h3bc0fe7d),
	.w8(32'h3985b56c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd94652),
	.w1(32'hbbdc9b8f),
	.w2(32'h3bc07341),
	.w3(32'hbbdb1463),
	.w4(32'hbc1fc9b1),
	.w5(32'hbb9d55b4),
	.w6(32'h3b0fd472),
	.w7(32'h3b621b73),
	.w8(32'hbc07d557),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac73a19),
	.w1(32'hbc1d2401),
	.w2(32'hbbd4c846),
	.w3(32'h3ad4204b),
	.w4(32'hbc1ba594),
	.w5(32'hbad13df3),
	.w6(32'hbbe96fd0),
	.w7(32'hbc52bf01),
	.w8(32'hbba5dad1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9ea78),
	.w1(32'hba1ace19),
	.w2(32'hba5c6d0b),
	.w3(32'h3a4e1709),
	.w4(32'h397c38ee),
	.w5(32'hba179b32),
	.w6(32'h39ff07f1),
	.w7(32'hbb659b5d),
	.w8(32'hbaf1c0af),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83dd40),
	.w1(32'hbac89fa9),
	.w2(32'hbab7e92e),
	.w3(32'hbb0082a2),
	.w4(32'hba1f6976),
	.w5(32'h39f34ea0),
	.w6(32'hbb0545dc),
	.w7(32'hbb2e3384),
	.w8(32'hbb5ae098),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa76af2),
	.w1(32'h3b1d57a5),
	.w2(32'h39c9742b),
	.w3(32'h3a22afc9),
	.w4(32'hbac47373),
	.w5(32'hb9b833f6),
	.w6(32'h399be5c3),
	.w7(32'hbb07f908),
	.w8(32'hba39b9e3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c3c49),
	.w1(32'hb9669da4),
	.w2(32'h39d7aecb),
	.w3(32'hba5932ef),
	.w4(32'h3baaa80d),
	.w5(32'h3ac89594),
	.w6(32'hbb0156be),
	.w7(32'h3b7b993d),
	.w8(32'hb8f96df2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d07ef1),
	.w1(32'hb9ae5dbf),
	.w2(32'h3a02acdc),
	.w3(32'hbb120595),
	.w4(32'h37f698cf),
	.w5(32'hb8edbffe),
	.w6(32'h39a8e634),
	.w7(32'hba422ea1),
	.w8(32'hba921b6f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80353b),
	.w1(32'hbaa6b845),
	.w2(32'hba4791f4),
	.w3(32'hbaa0cd10),
	.w4(32'hb9ddfc03),
	.w5(32'h3ac49732),
	.w6(32'hbb1bb6a7),
	.w7(32'hbb17821d),
	.w8(32'hbb57477e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4b703ae),
	.w1(32'h39f1d59d),
	.w2(32'h387d7c75),
	.w3(32'hba509ecf),
	.w4(32'hb949797e),
	.w5(32'hbac0de4a),
	.w6(32'hbb03d495),
	.w7(32'h391a50ff),
	.w8(32'hb9bac84e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10bf1e),
	.w1(32'hba4c7dba),
	.w2(32'hbb103b5d),
	.w3(32'h3a31454e),
	.w4(32'hbac51ad3),
	.w5(32'hbb080a43),
	.w6(32'hb9d6b6db),
	.w7(32'hbb38c12b),
	.w8(32'hbb4d64ef),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bb20c),
	.w1(32'hba8fef42),
	.w2(32'hba334c4a),
	.w3(32'hbb03e516),
	.w4(32'hba8207b0),
	.w5(32'hbb482db1),
	.w6(32'hbb62f0d9),
	.w7(32'hb9d99099),
	.w8(32'hba6c38c9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bea31),
	.w1(32'h3b4230e2),
	.w2(32'hba95f631),
	.w3(32'h39219477),
	.w4(32'h3af77acb),
	.w5(32'h3960be56),
	.w6(32'hbaf781d0),
	.w7(32'h3a902667),
	.w8(32'hbb000917),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbe908),
	.w1(32'h39c947c3),
	.w2(32'h39ed5d01),
	.w3(32'h3ab4c8c4),
	.w4(32'h39ee0f77),
	.w5(32'h37f1ef1f),
	.w6(32'hb97c07d7),
	.w7(32'hbb41f6fd),
	.w8(32'hb953124f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa272ee),
	.w1(32'h3b857aa0),
	.w2(32'h3bb4b616),
	.w3(32'hbb39765a),
	.w4(32'h3b82dde8),
	.w5(32'h3b882dbe),
	.w6(32'hbb9ac98e),
	.w7(32'h3b9331ae),
	.w8(32'h3b5788ba),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82d64e),
	.w1(32'h3932f489),
	.w2(32'h3a0a468c),
	.w3(32'h3bba7ab7),
	.w4(32'hb98f5571),
	.w5(32'hba108d6b),
	.w6(32'h3b8c94a9),
	.w7(32'h38e70a95),
	.w8(32'hb9eac729),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1993e2),
	.w1(32'h3a3e21c1),
	.w2(32'h399306a8),
	.w3(32'hb90e0e65),
	.w4(32'h3a228058),
	.w5(32'hb98fcbc8),
	.w6(32'h3a12d87d),
	.w7(32'h3a0b5b02),
	.w8(32'h395e045d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a572c5a),
	.w1(32'h3aa0a757),
	.w2(32'h3ae81fe9),
	.w3(32'hba77a00c),
	.w4(32'h39c6d04e),
	.w5(32'h3b2116ef),
	.w6(32'hbb57a051),
	.w7(32'hb8b751ea),
	.w8(32'hba94a84d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1c732),
	.w1(32'h3983212f),
	.w2(32'h3a5607c3),
	.w3(32'hbb7bb326),
	.w4(32'h3aa20324),
	.w5(32'hbad203ca),
	.w6(32'hbb44ca06),
	.w7(32'h3aa31c52),
	.w8(32'h39c92a7d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ceae5),
	.w1(32'hba7f976d),
	.w2(32'hbb9d3779),
	.w3(32'hba3d83c8),
	.w4(32'hbb0f356e),
	.w5(32'hbb8201c7),
	.w6(32'hba6690af),
	.w7(32'hbb242a98),
	.w8(32'hbb5c46f7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07961e),
	.w1(32'hbb587dd7),
	.w2(32'hbb000b6a),
	.w3(32'hbb87a0f7),
	.w4(32'h3a2d6e85),
	.w5(32'hba8cc14a),
	.w6(32'hbac4eb7a),
	.w7(32'hba65a291),
	.w8(32'hb96202e6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6d59c),
	.w1(32'h39ef3174),
	.w2(32'h3a9c26c7),
	.w3(32'hba5f749c),
	.w4(32'hbb0ae67d),
	.w5(32'hba439dfb),
	.w6(32'hbb081ecc),
	.w7(32'hba8b2343),
	.w8(32'hba040ab4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb777776d),
	.w1(32'h39949f3d),
	.w2(32'hba009428),
	.w3(32'hbb54728c),
	.w4(32'hb9614f97),
	.w5(32'h3a6b1c7c),
	.w6(32'hbb114330),
	.w7(32'hba06239d),
	.w8(32'hb839452d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a3ff1),
	.w1(32'hbafb91a4),
	.w2(32'h3b4550c2),
	.w3(32'hbb407fe1),
	.w4(32'hbb439da4),
	.w5(32'hbb1fe5f2),
	.w6(32'hbb9964a5),
	.w7(32'hbb93c263),
	.w8(32'hbbacd644),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6717e2),
	.w1(32'h39f2c2fd),
	.w2(32'h3b06203a),
	.w3(32'hbb40aca4),
	.w4(32'h39d2287a),
	.w5(32'h399ef2b6),
	.w6(32'hbbbd628f),
	.w7(32'hbaa7f8be),
	.w8(32'hba2e14ee),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833a04),
	.w1(32'hbb8f916b),
	.w2(32'h3a6d28e8),
	.w3(32'hbb6255f8),
	.w4(32'h3ad28d85),
	.w5(32'h3b979432),
	.w6(32'hbbd821f8),
	.w7(32'hbb4d9931),
	.w8(32'hba408c0d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10c438),
	.w1(32'h3b0f6df9),
	.w2(32'h3b2aee10),
	.w3(32'h3a888387),
	.w4(32'h3a518949),
	.w5(32'hba91f0b4),
	.w6(32'h3ad6d987),
	.w7(32'h3a815f13),
	.w8(32'h394e3559),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf7d52),
	.w1(32'h3acdac9e),
	.w2(32'h3998bd5b),
	.w3(32'h3a2d43cf),
	.w4(32'h3aab41ba),
	.w5(32'hbae1bf7b),
	.w6(32'h3a0549c0),
	.w7(32'h3af94ae5),
	.w8(32'h39aff948),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85c046),
	.w1(32'hba1cfc8f),
	.w2(32'hba8ebfd5),
	.w3(32'h3a76b132),
	.w4(32'h3b57b771),
	.w5(32'h3b6bbd17),
	.w6(32'h3b4b3880),
	.w7(32'hbb1cdf7f),
	.w8(32'hba8f4644),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba860fd9),
	.w1(32'hb9957d05),
	.w2(32'hba828abe),
	.w3(32'hb9b69ec3),
	.w4(32'hba352348),
	.w5(32'h396c075c),
	.w6(32'hba2a41e5),
	.w7(32'hbb52c038),
	.w8(32'hb92a05a5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba845ccc),
	.w1(32'hb8082680),
	.w2(32'hbabf6cb0),
	.w3(32'h3a248854),
	.w4(32'h39d68fc7),
	.w5(32'h398649c6),
	.w6(32'h3ab4cb96),
	.w7(32'hba465964),
	.w8(32'hba6567df),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb294dfd),
	.w1(32'h3975913b),
	.w2(32'hba8e6fe8),
	.w3(32'h392a6659),
	.w4(32'hbb3aeb22),
	.w5(32'hbaa50986),
	.w6(32'h3a015202),
	.w7(32'hbb178750),
	.w8(32'h395a60d3),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba081c46),
	.w1(32'hbab086b9),
	.w2(32'hba5dae36),
	.w3(32'h3b1a1c2a),
	.w4(32'hbb212fe9),
	.w5(32'hbb443b16),
	.w6(32'hb9dd769c),
	.w7(32'hbb649987),
	.w8(32'hbb2c84ed),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb452811),
	.w1(32'h3a7aa622),
	.w2(32'h3b45d0eb),
	.w3(32'hbb4b0955),
	.w4(32'h3a5bff78),
	.w5(32'h3aefd288),
	.w6(32'hbbb8b865),
	.w7(32'hbac4f8cd),
	.w8(32'hb9947bcb),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a808f90),
	.w1(32'h39c2d71f),
	.w2(32'h38566825),
	.w3(32'h3af9f0e6),
	.w4(32'hba2022ef),
	.w5(32'hba72a5a2),
	.w6(32'h36934ba8),
	.w7(32'hba415490),
	.w8(32'hbaab2162),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ede9f),
	.w1(32'hbaf0ec35),
	.w2(32'hb9b4cfb2),
	.w3(32'hbacb4317),
	.w4(32'hbaa44704),
	.w5(32'hbb397d65),
	.w6(32'hba9244d8),
	.w7(32'hbaa1d3aa),
	.w8(32'hbb5284a3),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4e043),
	.w1(32'hbb0d211e),
	.w2(32'h3af5b2be),
	.w3(32'hbb3e75b6),
	.w4(32'hbb3c15fb),
	.w5(32'h3b402979),
	.w6(32'hbbb80f80),
	.w7(32'hbb661d4a),
	.w8(32'hba95da7d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb022c76),
	.w1(32'h38f0e0b5),
	.w2(32'hba79a980),
	.w3(32'hba9ce0c4),
	.w4(32'hb9f6fbea),
	.w5(32'hbb6dbda9),
	.w6(32'hbb724023),
	.w7(32'hba47bb19),
	.w8(32'hbb73db94),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02d8f9),
	.w1(32'hbaba4bb5),
	.w2(32'h36fec7c6),
	.w3(32'hbae1203b),
	.w4(32'hb9665a23),
	.w5(32'hba6ac052),
	.w6(32'hbb463979),
	.w7(32'hba231284),
	.w8(32'hba326f4e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33bfab),
	.w1(32'hba0ec5e9),
	.w2(32'hb812439a),
	.w3(32'hbb0c9dba),
	.w4(32'h3884725b),
	.w5(32'h38a9a3a8),
	.w6(32'hbb840add),
	.w7(32'hba4dcbdb),
	.w8(32'h3a772e0d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f98064),
	.w1(32'hb93a8f47),
	.w2(32'h3a981941),
	.w3(32'h3a6611a1),
	.w4(32'h3a192538),
	.w5(32'h3a9824f1),
	.w6(32'h3a9e209f),
	.w7(32'h3abd5a9a),
	.w8(32'h3a4a81f6),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb136c),
	.w1(32'hbaed7e96),
	.w2(32'hba8476d4),
	.w3(32'h39827e8a),
	.w4(32'hb98d37d4),
	.w5(32'h3a25a17f),
	.w6(32'h3aa23a9a),
	.w7(32'hba2816a5),
	.w8(32'h3a440499),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3851d6f3),
	.w1(32'hb688f2d5),
	.w2(32'h3b126265),
	.w3(32'hba3cb786),
	.w4(32'hba6246dc),
	.w5(32'h38717f74),
	.w6(32'h38d2dc56),
	.w7(32'hba39ba9d),
	.w8(32'hb70326cc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380beb85),
	.w1(32'hbb861257),
	.w2(32'hba8f34e7),
	.w3(32'hb995a58d),
	.w4(32'hbb680d87),
	.w5(32'hbb56df35),
	.w6(32'hbacea443),
	.w7(32'hbadddea3),
	.w8(32'hbaa09970),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03e86b),
	.w1(32'hba254053),
	.w2(32'hb81d19d3),
	.w3(32'hbaa0ba3e),
	.w4(32'hbb0b4e93),
	.w5(32'hb8381cad),
	.w6(32'hbb3dd2c3),
	.w7(32'hba4ae6c3),
	.w8(32'hbabc29ca),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bebcf),
	.w1(32'hbace8742),
	.w2(32'hbb1542d5),
	.w3(32'hbaadaf90),
	.w4(32'h3afbdd09),
	.w5(32'hbae26e2b),
	.w6(32'hbb3a9812),
	.w7(32'h39ff28ed),
	.w8(32'hba9c8a52),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ae0e8),
	.w1(32'hb9c3b0f8),
	.w2(32'h3a541bb6),
	.w3(32'hba08d8fe),
	.w4(32'h3b0cba34),
	.w5(32'h3b43fb78),
	.w6(32'hbab8ecf9),
	.w7(32'hba272117),
	.w8(32'h3a1900bb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59572c),
	.w1(32'hb9a5a360),
	.w2(32'h3b163c22),
	.w3(32'h3a719e35),
	.w4(32'h3b59c062),
	.w5(32'h3b84e69f),
	.w6(32'hbacfe33b),
	.w7(32'hba792ef7),
	.w8(32'h3a3e152a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39439dbc),
	.w1(32'hbacd9c93),
	.w2(32'hbade361b),
	.w3(32'h3aef481f),
	.w4(32'hb9cfca7d),
	.w5(32'hba2830ad),
	.w6(32'h39c7247d),
	.w7(32'hbb136a09),
	.w8(32'hbb01bd2a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c337d6),
	.w1(32'hb9591612),
	.w2(32'hba810073),
	.w3(32'h37d1fb11),
	.w4(32'hba61d9f3),
	.w5(32'h391856df),
	.w6(32'hbb2f0ac2),
	.w7(32'hba6fa4a1),
	.w8(32'h3a30722a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93dc970),
	.w1(32'hba937682),
	.w2(32'hb849bd22),
	.w3(32'hb9283644),
	.w4(32'hb972215f),
	.w5(32'h394e70a9),
	.w6(32'h3999e411),
	.w7(32'hba72adf0),
	.w8(32'hbb135841),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de6546),
	.w1(32'h3af3c172),
	.w2(32'h3b875613),
	.w3(32'h39893068),
	.w4(32'h3b07ec61),
	.w5(32'h3a441b3b),
	.w6(32'hb9ef961a),
	.w7(32'h3ac01b39),
	.w8(32'h3b536a22),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf4b62),
	.w1(32'hb928517e),
	.w2(32'h3ab2c007),
	.w3(32'hbac5bdb3),
	.w4(32'hb97f357e),
	.w5(32'h3a84af14),
	.w6(32'hb8fd0e54),
	.w7(32'hb9afe80d),
	.w8(32'h3a86e7f2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5dec84),
	.w1(32'hbaafdf44),
	.w2(32'hbaf8e1e4),
	.w3(32'hbae11062),
	.w4(32'hb96d45ab),
	.w5(32'hba0fa05e),
	.w6(32'hbb0ab76d),
	.w7(32'hbabc725f),
	.w8(32'hba854b64),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6c1b3),
	.w1(32'h39c1f23a),
	.w2(32'h399d752b),
	.w3(32'hba60aad0),
	.w4(32'h3b1118c1),
	.w5(32'h3b083508),
	.w6(32'hba74ed7d),
	.w7(32'h3a2e8983),
	.w8(32'hb9418fa8),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb007eac),
	.w1(32'h3b1322c5),
	.w2(32'h3a8414f4),
	.w3(32'hbafa93f9),
	.w4(32'hba8c5492),
	.w5(32'h3abbb19e),
	.w6(32'hba348364),
	.w7(32'h39915462),
	.w8(32'h3ab40024),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b3602),
	.w1(32'h38c0d4eb),
	.w2(32'h39ef6423),
	.w3(32'h3afe0705),
	.w4(32'hb8c18b43),
	.w5(32'h3981f12b),
	.w6(32'hba96f749),
	.w7(32'hba555ec0),
	.w8(32'hbaba0c2a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d5f1d),
	.w1(32'h38041042),
	.w2(32'h3aa9d13b),
	.w3(32'hbaa81a38),
	.w4(32'h3b238497),
	.w5(32'h3a3ca6ba),
	.w6(32'hbaa6fc14),
	.w7(32'h3a9319a4),
	.w8(32'hb9ead273),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a202c74),
	.w1(32'hb8f45dc2),
	.w2(32'h3b52517b),
	.w3(32'h3b48ca7c),
	.w4(32'hbad5358e),
	.w5(32'hbab06d1c),
	.w6(32'h3b39581b),
	.w7(32'hba9c3ed8),
	.w8(32'hba241ea6),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a031c),
	.w1(32'hb9a0372c),
	.w2(32'hbb4f1eac),
	.w3(32'hbb92df80),
	.w4(32'h3b0ee1d7),
	.w5(32'h3a884876),
	.w6(32'hbb9bf34f),
	.w7(32'h38f65be5),
	.w8(32'h3aced2b8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aa629),
	.w1(32'hba895e64),
	.w2(32'hbac3d5c2),
	.w3(32'hb94c1e0d),
	.w4(32'hb9eed72c),
	.w5(32'hbb6b668e),
	.w6(32'hba8ad4fb),
	.w7(32'hba3ac83e),
	.w8(32'hbb1d80ab),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b5d89),
	.w1(32'hb94af458),
	.w2(32'hb84a0384),
	.w3(32'h38ede01f),
	.w4(32'hbb1f1d85),
	.w5(32'hbaabc429),
	.w6(32'hbad7998f),
	.w7(32'hbaf98078),
	.w8(32'hba86ef25),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule