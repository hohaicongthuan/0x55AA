module layer_8_featuremap_22(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987b789),
	.w1(32'h3c251d0b),
	.w2(32'hbbf456cb),
	.w3(32'h3c1944dd),
	.w4(32'hbb41142a),
	.w5(32'hbcc60161),
	.w6(32'h3cc091e2),
	.w7(32'h3b89b6fd),
	.w8(32'hbc8db6aa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27b8e2),
	.w1(32'hbb8df0da),
	.w2(32'hbbbebd13),
	.w3(32'hbac602b8),
	.w4(32'hbba68087),
	.w5(32'h3ac04959),
	.w6(32'h3b618b95),
	.w7(32'h3bbc0d4b),
	.w8(32'h3c5affc8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f5bc4),
	.w1(32'hbb08e860),
	.w2(32'h3aa53221),
	.w3(32'hbc229bd9),
	.w4(32'hbb730093),
	.w5(32'h3be1932c),
	.w6(32'hbb46951d),
	.w7(32'h3bbecbee),
	.w8(32'h3c0c270e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bd9b7),
	.w1(32'h3c785e54),
	.w2(32'hbc9c8db5),
	.w3(32'h3cbef60d),
	.w4(32'h3c5091fc),
	.w5(32'h3c4463d4),
	.w6(32'h3bede605),
	.w7(32'h3adb3a46),
	.w8(32'hbc1c866c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6cfc5),
	.w1(32'hbc4074b1),
	.w2(32'hbb87a571),
	.w3(32'hbca35780),
	.w4(32'hbbd79e5a),
	.w5(32'h3b38aee7),
	.w6(32'hbc0c6e3c),
	.w7(32'h3b3bd840),
	.w8(32'h3d2f9f38),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7268d6),
	.w1(32'h3b817751),
	.w2(32'hbce1d261),
	.w3(32'hbb922d3c),
	.w4(32'hbccc8d1d),
	.w5(32'h3abbb0f6),
	.w6(32'hbc29492a),
	.w7(32'hbc1bb72e),
	.w8(32'h3d0607a4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb191106),
	.w1(32'hbad081d5),
	.w2(32'hbb790b37),
	.w3(32'h39feb978),
	.w4(32'h399c9289),
	.w5(32'hb863f8f7),
	.w6(32'hb9d10d70),
	.w7(32'h3aecc90d),
	.w8(32'hbc6b1297),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcff03c2),
	.w1(32'hbc3418e3),
	.w2(32'hbbb841eb),
	.w3(32'hbc95cb83),
	.w4(32'hbc35a6df),
	.w5(32'hbb9fbbb7),
	.w6(32'hbc036ca8),
	.w7(32'hbb462a7c),
	.w8(32'hbc0f2419),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8c869),
	.w1(32'hbc90ff72),
	.w2(32'hbc1d683c),
	.w3(32'hbc68cdd0),
	.w4(32'hbc47998f),
	.w5(32'h3b43ed77),
	.w6(32'hbad52751),
	.w7(32'h3c00fb03),
	.w8(32'hbb404311),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04425d),
	.w1(32'hbcdc987e),
	.w2(32'h3bd4208a),
	.w3(32'h3c666577),
	.w4(32'hbafcee05),
	.w5(32'hbcf4c5e0),
	.w6(32'h3c827f28),
	.w7(32'h3c7a3032),
	.w8(32'hbc695bba),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88baf4),
	.w1(32'h3a834b1b),
	.w2(32'hbc536c23),
	.w3(32'h3bb5af2c),
	.w4(32'hbb82f60c),
	.w5(32'hbc951d5c),
	.w6(32'h3cbc8cfd),
	.w7(32'h3b3e7510),
	.w8(32'hbcb82f4b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c085d96),
	.w1(32'hbaea84ec),
	.w2(32'h3a1df079),
	.w3(32'h3c6d0514),
	.w4(32'hbc2b5a0a),
	.w5(32'hbbd73611),
	.w6(32'h3ab1e84e),
	.w7(32'hbbd851ca),
	.w8(32'hbc53db4f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28f11c),
	.w1(32'hbbcb2c7c),
	.w2(32'h3ab65a4d),
	.w3(32'hbb735d48),
	.w4(32'h3a4dc16c),
	.w5(32'h3c3f628a),
	.w6(32'hbbafc12b),
	.w7(32'h3c151110),
	.w8(32'h3d82323e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6163ee),
	.w1(32'hbb944044),
	.w2(32'hbd669e32),
	.w3(32'h3c83466d),
	.w4(32'hbd05abf4),
	.w5(32'hbd5a4ca2),
	.w6(32'h3a9e90ac),
	.w7(32'hbcde44bd),
	.w8(32'h3ca556eb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdd38e1),
	.w1(32'h3a575006),
	.w2(32'hbce34c17),
	.w3(32'h3bf7e9ad),
	.w4(32'hbc20f5ef),
	.w5(32'hbcd0d6b3),
	.w6(32'h3baa57f6),
	.w7(32'hbc3bea2c),
	.w8(32'hbabe6bce),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb389a88),
	.w1(32'hbb4af43c),
	.w2(32'hba90cdaf),
	.w3(32'hbb3630d3),
	.w4(32'hbb250988),
	.w5(32'h3b33b7c9),
	.w6(32'hb9b12c26),
	.w7(32'h3b06b665),
	.w8(32'hbb997ae1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9495b1),
	.w1(32'h3b769b13),
	.w2(32'hbc0b049d),
	.w3(32'h3c0fe2db),
	.w4(32'h3b57057d),
	.w5(32'hbca46f3e),
	.w6(32'h3c07d9dc),
	.w7(32'h3c2b68ad),
	.w8(32'hbbefcd3f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbda9de),
	.w1(32'hbbedcbec),
	.w2(32'h3ae1dcf4),
	.w3(32'h3b316988),
	.w4(32'hbb5387e6),
	.w5(32'h3a9d2b00),
	.w6(32'hbb88da6f),
	.w7(32'h3bca25f8),
	.w8(32'hbc79fba4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3b5f09),
	.w1(32'h3c593bf7),
	.w2(32'hbc476490),
	.w3(32'h3caad93b),
	.w4(32'hbd1622f4),
	.w5(32'hbd948931),
	.w6(32'h3d60be19),
	.w7(32'hbd0ad64f),
	.w8(32'hbdc28512),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c18cd),
	.w1(32'hbb1d464b),
	.w2(32'hbc6fb048),
	.w3(32'hbccf78e6),
	.w4(32'hbd2b7612),
	.w5(32'hbabad32f),
	.w6(32'h3c24cbfd),
	.w7(32'hbcb1cbdd),
	.w8(32'hbc9f32a1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd15f10e),
	.w1(32'hbbc9aac1),
	.w2(32'h3d049950),
	.w3(32'hbcac6105),
	.w4(32'h3c86e12f),
	.w5(32'h3d08e7a3),
	.w6(32'hbc77c9b6),
	.w7(32'h3c8937a4),
	.w8(32'hbcaac526),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f6306),
	.w1(32'hbb2cdb79),
	.w2(32'h3ac90824),
	.w3(32'hbc4f4313),
	.w4(32'h39836467),
	.w5(32'h3c51d059),
	.w6(32'hbb9ddaff),
	.w7(32'h3be8db34),
	.w8(32'hbba2543c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd58b085),
	.w1(32'hbb872b15),
	.w2(32'h3d4300b8),
	.w3(32'h3b90da70),
	.w4(32'hbc25f6c8),
	.w5(32'hbc997e45),
	.w6(32'h3d0a8e7e),
	.w7(32'h3c23c77e),
	.w8(32'hbd8d8c74),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc921272),
	.w1(32'hbbf3ef7d),
	.w2(32'h3ba52b6c),
	.w3(32'hbcce6163),
	.w4(32'hbc44034e),
	.w5(32'h3c72b5d8),
	.w6(32'hbc4f7b41),
	.w7(32'h3c8d29c4),
	.w8(32'h3bda69fd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd211bf),
	.w1(32'hbc3779df),
	.w2(32'h3ca7d3ce),
	.w3(32'hbbba1724),
	.w4(32'hbb867cb0),
	.w5(32'h3c94a39d),
	.w6(32'hbc9286b7),
	.w7(32'h3b89b055),
	.w8(32'hbcbe2cd0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc689030),
	.w1(32'h3c48d5e4),
	.w2(32'h3d992908),
	.w3(32'h3cad3bf4),
	.w4(32'h3c8a96fb),
	.w5(32'h3d15ac2c),
	.w6(32'h3c8668d8),
	.w7(32'h3cfe7de7),
	.w8(32'hbcadcfbd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a8d39),
	.w1(32'h3b4eb9d9),
	.w2(32'h3d214a25),
	.w3(32'h3b35bd6a),
	.w4(32'h3c1bdb90),
	.w5(32'h3ce70142),
	.w6(32'hbbf2b3f5),
	.w7(32'h3c730187),
	.w8(32'hbcfb0bbc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdfa2170),
	.w1(32'hbdc1a5e4),
	.w2(32'h3eb0b2f3),
	.w3(32'h3d155af5),
	.w4(32'h3da6ece4),
	.w5(32'h3baff76d),
	.w6(32'h3dfefa49),
	.w7(32'h3dcb5f1d),
	.w8(32'hbdf44952),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c07db),
	.w1(32'hbb911cdf),
	.w2(32'h3cc6de3c),
	.w3(32'h3c4b7e0b),
	.w4(32'hbc6ba365),
	.w5(32'h3ba30fb6),
	.w6(32'hbaee4a8a),
	.w7(32'h3bf2f933),
	.w8(32'hbbece72e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b53a8b),
	.w1(32'h397d8373),
	.w2(32'hbbb8b4ca),
	.w3(32'h3a1f46fc),
	.w4(32'h3ae01a67),
	.w5(32'h39a5fe4f),
	.w6(32'h3b7fbb51),
	.w7(32'h3b274b9d),
	.w8(32'h3c860713),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2089dd),
	.w1(32'h3b2401a9),
	.w2(32'hbc9e1bca),
	.w3(32'hbbfa7c88),
	.w4(32'h3c9ba817),
	.w5(32'h3ceea0d2),
	.w6(32'h3cb24b8d),
	.w7(32'hbc452960),
	.w8(32'hbd9c8166),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8d24c5),
	.w1(32'hbb5f7dcd),
	.w2(32'h3d6104d2),
	.w3(32'hbce80da3),
	.w4(32'h3cd9c655),
	.w5(32'h3d8699a4),
	.w6(32'hbcb7f95e),
	.w7(32'h3c9f3f0d),
	.w8(32'h3c0e8fc6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb66773),
	.w1(32'hbc32ee1c),
	.w2(32'hbce0871e),
	.w3(32'hbbf8ca78),
	.w4(32'hbbd0d716),
	.w5(32'hb8d002b7),
	.w6(32'hbb9b7f9b),
	.w7(32'h3b8b1a72),
	.w8(32'h3a41953d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f12e0),
	.w1(32'hbb2b9f49),
	.w2(32'h3bcfb076),
	.w3(32'hbb268772),
	.w4(32'h3b056ef2),
	.w5(32'h3bb0837e),
	.w6(32'h3c1a18e4),
	.w7(32'hbbf03f90),
	.w8(32'h3d22851f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4d9d2d),
	.w1(32'hbcaa5eef),
	.w2(32'hbd7df6fc),
	.w3(32'h3a8e33f4),
	.w4(32'hbd4446a3),
	.w5(32'hbd55e2fc),
	.w6(32'hbc0dbb14),
	.w7(32'hbce5f735),
	.w8(32'h3bae05ea),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca645ed),
	.w1(32'hbc1b4f51),
	.w2(32'h3ae69457),
	.w3(32'h3c2602e0),
	.w4(32'hbb8cf912),
	.w5(32'hbc500598),
	.w6(32'h3c5b6d72),
	.w7(32'h3b6b6680),
	.w8(32'hbd6e2933),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd05df17),
	.w1(32'hbacc59ed),
	.w2(32'h3ccc7609),
	.w3(32'hbc265c40),
	.w4(32'h3bee37ae),
	.w5(32'h3cd2264d),
	.w6(32'hbc83f1c3),
	.w7(32'h3bb1e9d7),
	.w8(32'h3a8766b1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba078ad),
	.w1(32'hbb41cb86),
	.w2(32'hbc1c1e77),
	.w3(32'h3a19193e),
	.w4(32'h392c29db),
	.w5(32'hbad4dba6),
	.w6(32'h3bd468b6),
	.w7(32'h3ba23ae6),
	.w8(32'h3d06bb86),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2117e7),
	.w1(32'hbb006b2f),
	.w2(32'hbd3e414d),
	.w3(32'h3b8d6111),
	.w4(32'hbc874866),
	.w5(32'hbd35390e),
	.w6(32'h3b828a63),
	.w7(32'hbca15c91),
	.w8(32'hbd1a515e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd04ee3b),
	.w1(32'h3b08d976),
	.w2(32'h3d0ea146),
	.w3(32'hbbed8811),
	.w4(32'h3c9037d2),
	.w5(32'h3d049b41),
	.w6(32'hbc585ce6),
	.w7(32'h3c2dd935),
	.w8(32'hbc50ef55),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f0bdc),
	.w1(32'h3bbae8d1),
	.w2(32'h3d53b84b),
	.w3(32'h3d33e8b0),
	.w4(32'hbb4c2b4d),
	.w5(32'h3c915722),
	.w6(32'h3c3371e4),
	.w7(32'hbbdcb0ca),
	.w8(32'h3ca9a2d7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb11955),
	.w1(32'h3ad7c578),
	.w2(32'h3b9a7355),
	.w3(32'hbbe1b564),
	.w4(32'hbbe4e9fe),
	.w5(32'h3aca5f20),
	.w6(32'h3b4bbd00),
	.w7(32'hbb0cb53b),
	.w8(32'hba9113bc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb68829),
	.w1(32'hbac8cd8e),
	.w2(32'h3bb57af8),
	.w3(32'hbac7cdcc),
	.w4(32'h3a3a1b25),
	.w5(32'h3b13c4c7),
	.w6(32'hbbec43e3),
	.w7(32'h3a1336b6),
	.w8(32'h3b15f69b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc03f28),
	.w1(32'hbb1cde28),
	.w2(32'h3bab082c),
	.w3(32'h3b7f8823),
	.w4(32'hbab0785e),
	.w5(32'hbbf6bcde),
	.w6(32'h3c8e1d82),
	.w7(32'h3a3aa966),
	.w8(32'hbc52f73c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f88507),
	.w1(32'h3cc2fdde),
	.w2(32'h3c86f761),
	.w3(32'h3c3b963a),
	.w4(32'hbba7da6b),
	.w5(32'hbcc18855),
	.w6(32'h3d17853e),
	.w7(32'hbc0a101a),
	.w8(32'hbd1533e9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03818f),
	.w1(32'h3c681b8c),
	.w2(32'h3a31e29d),
	.w3(32'h3c1d0139),
	.w4(32'hbaab7342),
	.w5(32'hbc1a1c40),
	.w6(32'h3c45c5f0),
	.w7(32'hbb422ead),
	.w8(32'hbc61b74e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe18c35),
	.w1(32'hbb987852),
	.w2(32'hbbdfd7e2),
	.w3(32'h3b585a3b),
	.w4(32'h3abba7da),
	.w5(32'hbb89e557),
	.w6(32'hbba17135),
	.w7(32'hbb867848),
	.w8(32'hba6d8f2c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd3dfe),
	.w1(32'h3c233c9c),
	.w2(32'h3c64b49c),
	.w3(32'h3b2b7bc6),
	.w4(32'h3bb52b1b),
	.w5(32'hbc6dc514),
	.w6(32'h3d008550),
	.w7(32'h3bd3decb),
	.w8(32'hbcd709aa),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab01de8),
	.w1(32'h3abb8686),
	.w2(32'h3bcf8229),
	.w3(32'h3a9e4a06),
	.w4(32'h3a6d9c2d),
	.w5(32'h3be75765),
	.w6(32'h3bc9937b),
	.w7(32'h3c117e62),
	.w8(32'h3c0facab),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c653687),
	.w1(32'h3c55e5f3),
	.w2(32'h3a96941c),
	.w3(32'h3ca2f403),
	.w4(32'hbb54e884),
	.w5(32'hbc03d06f),
	.w6(32'h3c8ccec0),
	.w7(32'hbbe13953),
	.w8(32'hbc55c7b8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb0232),
	.w1(32'h3ce7ed99),
	.w2(32'h3d4773e1),
	.w3(32'h3866278a),
	.w4(32'h3d0562ae),
	.w5(32'h3d7776ea),
	.w6(32'hbbc54f86),
	.w7(32'h3d1d518b),
	.w8(32'h3d86ea44),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb138e1f),
	.w1(32'h3c4d287c),
	.w2(32'h3b4f1801),
	.w3(32'hb90d5666),
	.w4(32'hbc242dea),
	.w5(32'hbd016f0b),
	.w6(32'h3d1e09bc),
	.w7(32'hbd276d7d),
	.w8(32'hbd5798c3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0776d0),
	.w1(32'h3bd7a18f),
	.w2(32'h3b5bc7fa),
	.w3(32'hbb87e4ca),
	.w4(32'hba86843c),
	.w5(32'hbacac1c5),
	.w6(32'h3af5058a),
	.w7(32'hbb2290c4),
	.w8(32'h39a60ba2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb867b8),
	.w1(32'h3b6407bc),
	.w2(32'hbc902db5),
	.w3(32'h3c13ce3b),
	.w4(32'hbc5c94dd),
	.w5(32'hbd46a4ac),
	.w6(32'h3ae7f51e),
	.w7(32'hbc2604b5),
	.w8(32'hbd0ef665),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4da250),
	.w1(32'hba8c47fe),
	.w2(32'hbb01579c),
	.w3(32'hbad1c98e),
	.w4(32'h3b89c887),
	.w5(32'hbb0c4596),
	.w6(32'hbb5f5c40),
	.w7(32'hbac93320),
	.w8(32'h3bcf7d37),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c01b3),
	.w1(32'hbbb202e3),
	.w2(32'h3c996ad7),
	.w3(32'h3ce117e2),
	.w4(32'hbc82e91a),
	.w5(32'hbd349b2a),
	.w6(32'h3d5e0e58),
	.w7(32'h3cb41865),
	.w8(32'hbd40a71c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09f0a0),
	.w1(32'hbc28bfbf),
	.w2(32'hbc93ee12),
	.w3(32'hbbb77edd),
	.w4(32'hbc03103a),
	.w5(32'hbc6c1f28),
	.w6(32'hbafad31b),
	.w7(32'h3b125170),
	.w8(32'hbbc4948a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43dfb8),
	.w1(32'h3bb6b49a),
	.w2(32'hbb8da9a3),
	.w3(32'hbb845eab),
	.w4(32'hbc437262),
	.w5(32'hbc12f466),
	.w6(32'h3c9143be),
	.w7(32'hbc9fe96a),
	.w8(32'hbc78671b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb036f69),
	.w1(32'h3c066121),
	.w2(32'h3bbfb11e),
	.w3(32'h3bfbb651),
	.w4(32'h3c48742c),
	.w5(32'hbbb1d7f4),
	.w6(32'h3cc6ed95),
	.w7(32'h3c2af05d),
	.w8(32'hbc6ea3a0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bebe7),
	.w1(32'h3c31476c),
	.w2(32'h3c26b0d1),
	.w3(32'h3c5bd74c),
	.w4(32'h3c2e4f5d),
	.w5(32'h3bb78dd4),
	.w6(32'h3c9446ad),
	.w7(32'h3bf4ee31),
	.w8(32'h3c54464a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09019b),
	.w1(32'hbbb7b115),
	.w2(32'hba0c7315),
	.w3(32'h3ab6e295),
	.w4(32'hba6b844e),
	.w5(32'hb735e34a),
	.w6(32'hbb7f42c3),
	.w7(32'hbb8762ba),
	.w8(32'hbac3214e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bcdcb),
	.w1(32'h3b1b374c),
	.w2(32'h3b1c53ab),
	.w3(32'h38e56796),
	.w4(32'h39e2fd2d),
	.w5(32'hb9596ead),
	.w6(32'hba08c480),
	.w7(32'h399b793c),
	.w8(32'h38fe2828),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a50b1),
	.w1(32'h3c6b3bac),
	.w2(32'h3c9cc69b),
	.w3(32'h3cedb882),
	.w4(32'hbc025f75),
	.w5(32'hbc182b58),
	.w6(32'h3cb56a4e),
	.w7(32'h3af6ec9a),
	.w8(32'hbaef2707),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61d725),
	.w1(32'hbb42498a),
	.w2(32'hbba221b3),
	.w3(32'hbc4ce29a),
	.w4(32'hbc4406ea),
	.w5(32'hbb8aeef1),
	.w6(32'hbb614926),
	.w7(32'hbbdd38f2),
	.w8(32'hbb1ffac5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fbcce),
	.w1(32'h3b8b9aed),
	.w2(32'h3bc82794),
	.w3(32'h3aa7198c),
	.w4(32'h3b7f47df),
	.w5(32'h3be7fffc),
	.w6(32'h3bdfc85e),
	.w7(32'h3befbaf4),
	.w8(32'h3bd2688d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a81e1),
	.w1(32'hbb94939b),
	.w2(32'h3be99ca1),
	.w3(32'hbb5529b9),
	.w4(32'hbc044fd8),
	.w5(32'hba86ba16),
	.w6(32'h3b3d08ec),
	.w7(32'hbbac3943),
	.w8(32'h3a2b1908),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc098677),
	.w1(32'h3b543f92),
	.w2(32'h3c83f041),
	.w3(32'hbc0abaa9),
	.w4(32'h3ba9a5ae),
	.w5(32'h3c7d3ec2),
	.w6(32'hb8379236),
	.w7(32'h3bc02454),
	.w8(32'h3c3b0599),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a43b2),
	.w1(32'h3c0db994),
	.w2(32'h3c26394b),
	.w3(32'h3c2aec93),
	.w4(32'hbb0621c9),
	.w5(32'hbb7d7d2c),
	.w6(32'hbb0ecb59),
	.w7(32'hbb998eb3),
	.w8(32'hb88100b5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa19faa),
	.w1(32'h3a926625),
	.w2(32'h3b0aadd4),
	.w3(32'h3afc34e8),
	.w4(32'h3b03a895),
	.w5(32'h3b3ee623),
	.w6(32'h3b13ed7d),
	.w7(32'h3b281d92),
	.w8(32'hba60545a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee5b55),
	.w1(32'hbc2bfd17),
	.w2(32'h3c58cada),
	.w3(32'h3cbbe23a),
	.w4(32'h3ca1188b),
	.w5(32'hbd38c4fa),
	.w6(32'h3d95ddb4),
	.w7(32'h3c1492db),
	.w8(32'hbd9a26c5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cebd5),
	.w1(32'h3a1d72f1),
	.w2(32'h3a139a22),
	.w3(32'hba3e7a7f),
	.w4(32'hba2132e5),
	.w5(32'hb8844c74),
	.w6(32'h3a1b1b3d),
	.w7(32'hb935afdf),
	.w8(32'h3a554732),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4553f7),
	.w1(32'hbc254b81),
	.w2(32'h3b4189e6),
	.w3(32'hbb90df6d),
	.w4(32'hbbcaf009),
	.w5(32'h391a56ba),
	.w6(32'h3c7de931),
	.w7(32'h3c47a6c3),
	.w8(32'h3c32527d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d3de1),
	.w1(32'h3b2ef833),
	.w2(32'h3b622e28),
	.w3(32'h3b1894d0),
	.w4(32'h3ad5c532),
	.w5(32'h3b35b2ed),
	.w6(32'h3b32c9ac),
	.w7(32'h3aaef976),
	.w8(32'hba9625c0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25096d),
	.w1(32'hbc8df9d4),
	.w2(32'hbb5ec65a),
	.w3(32'h3c5fdf20),
	.w4(32'hbc51e553),
	.w5(32'hbc257647),
	.w6(32'h3c078112),
	.w7(32'h3bd7d3f5),
	.w8(32'h3bbca920),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1cf9f),
	.w1(32'h3a9115d4),
	.w2(32'h3a9fd36d),
	.w3(32'h39b7b1eb),
	.w4(32'h3a4b70b3),
	.w5(32'h3ab3c5be),
	.w6(32'h3a159827),
	.w7(32'h3a0bd3e9),
	.w8(32'h39a1e3d3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc61cf),
	.w1(32'hbc04dc23),
	.w2(32'hbc58e758),
	.w3(32'hbb138963),
	.w4(32'hbba5f5af),
	.w5(32'hbc895605),
	.w6(32'hbb08470a),
	.w7(32'hbbbc115a),
	.w8(32'hbc2edba3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6be1e1),
	.w1(32'h39e75b4f),
	.w2(32'h3a7dfdc4),
	.w3(32'hb9a6d0fb),
	.w4(32'h38f8bd74),
	.w5(32'h3a0e20e9),
	.w6(32'h3a15f0e4),
	.w7(32'h3a17df04),
	.w8(32'hbb339731),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82fc32),
	.w1(32'hbb6b787f),
	.w2(32'h3bb4a7fb),
	.w3(32'h3c212b39),
	.w4(32'h3a42cac0),
	.w5(32'hbca0db3e),
	.w6(32'h3cbe32fd),
	.w7(32'hbbf9a0d6),
	.w8(32'hbcdfa29b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c6484),
	.w1(32'h3b0fea31),
	.w2(32'hbb0cf32f),
	.w3(32'h3b3a4f1b),
	.w4(32'hbbdeeeee),
	.w5(32'hbc4fc807),
	.w6(32'h3af22eae),
	.w7(32'hbbab26e6),
	.w8(32'hbc2c7725),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68fb3f),
	.w1(32'hbb5dd3b5),
	.w2(32'hbb127876),
	.w3(32'hbb8abc76),
	.w4(32'hbaf6529f),
	.w5(32'hbb03907c),
	.w6(32'hbb42947a),
	.w7(32'hbb037ef3),
	.w8(32'h3ae59406),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cb4c4),
	.w1(32'h3a3ada3c),
	.w2(32'h3a07c06f),
	.w3(32'h3b6bf91d),
	.w4(32'h3949037d),
	.w5(32'hbb58d9c4),
	.w6(32'h3bbb8fbd),
	.w7(32'h3b68958a),
	.w8(32'h3a53ab20),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8025f0),
	.w1(32'hbc02c28b),
	.w2(32'h3a96e6b5),
	.w3(32'hbcb8a6c3),
	.w4(32'hbc37e041),
	.w5(32'h3bb7e48b),
	.w6(32'h3c4a184a),
	.w7(32'h3c3fb1fd),
	.w8(32'h3b9a5cdf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad87b22),
	.w1(32'h3c1cd928),
	.w2(32'h3ca47e05),
	.w3(32'h3c46d7a7),
	.w4(32'hbb013aee),
	.w5(32'hbb52301f),
	.w6(32'h3cdac272),
	.w7(32'h3b548900),
	.w8(32'hbc3e569a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d87c6f6),
	.w1(32'h3d85dda3),
	.w2(32'h3d254fd7),
	.w3(32'h3d765582),
	.w4(32'h3cc3ebb1),
	.w5(32'h3d32c5fd),
	.w6(32'h3a1470be),
	.w7(32'hbc8fa9de),
	.w8(32'h3d445265),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f4d6a),
	.w1(32'h3c955170),
	.w2(32'h3cd26bf9),
	.w3(32'h3d006012),
	.w4(32'hba9e7f6e),
	.w5(32'hbccfaa14),
	.w6(32'h3d654ad8),
	.w7(32'h3948fa6b),
	.w8(32'hbd0e175a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5be47b),
	.w1(32'h3b21857f),
	.w2(32'hbbc6ada6),
	.w3(32'hbacaaed9),
	.w4(32'hbc2bd9e5),
	.w5(32'hbb57bcda),
	.w6(32'h3c9b2626),
	.w7(32'h3b4d7a67),
	.w8(32'hbc60266b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905cc70),
	.w1(32'hb9c76f0a),
	.w2(32'h3abadf98),
	.w3(32'hba44a47d),
	.w4(32'hbac0d24c),
	.w5(32'h3a2a6641),
	.w6(32'h3a3717c7),
	.w7(32'h3afcd339),
	.w8(32'hbae8c266),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38750abd),
	.w1(32'hb9bd0b0e),
	.w2(32'h39845985),
	.w3(32'hba4bff10),
	.w4(32'h3a3e312c),
	.w5(32'h3a101ae9),
	.w6(32'hb9b09c96),
	.w7(32'hba2bd5a2),
	.w8(32'hba12e2fe),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b395db5),
	.w1(32'h3b2417f7),
	.w2(32'h3ade18b5),
	.w3(32'h3b1ab078),
	.w4(32'h3aedc5e4),
	.w5(32'h3b265e67),
	.w6(32'h3a48d50c),
	.w7(32'h3a26a67d),
	.w8(32'h3af8e9e5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea79bf),
	.w1(32'h3a76c896),
	.w2(32'h39148acd),
	.w3(32'h3c1b855a),
	.w4(32'h3b2c6c49),
	.w5(32'hbaefc38e),
	.w6(32'h3c7eb65d),
	.w7(32'h3c020920),
	.w8(32'h3a988e26),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45fa5c),
	.w1(32'h3ba79e6c),
	.w2(32'h3b3b4eab),
	.w3(32'h3afdb221),
	.w4(32'hb985f9c1),
	.w5(32'h3c0d71b7),
	.w6(32'h3a588fa8),
	.w7(32'h3c2671ef),
	.w8(32'h3bb97b7b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae95964),
	.w1(32'hb998ae5b),
	.w2(32'h399fbacb),
	.w3(32'hbad57210),
	.w4(32'hbae6d79c),
	.w5(32'hbb06694a),
	.w6(32'hba17b6df),
	.w7(32'hba487825),
	.w8(32'hbbfda097),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8d87e),
	.w1(32'hbc951489),
	.w2(32'hbbc44ff1),
	.w3(32'hbca7c8e5),
	.w4(32'hbbb01099),
	.w5(32'hbbbc58d7),
	.w6(32'h3b16f689),
	.w7(32'hbb50a147),
	.w8(32'h3c118259),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85b35a),
	.w1(32'h3b05d508),
	.w2(32'h3b85b54f),
	.w3(32'h38b0cc19),
	.w4(32'hbb67a6a1),
	.w5(32'hbb96e01f),
	.w6(32'h3bfa2080),
	.w7(32'h3960c3d4),
	.w8(32'hbb9abfb5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed4282),
	.w1(32'h3b987bfc),
	.w2(32'h3b850b15),
	.w3(32'h3ad9afcf),
	.w4(32'hbbe7c3ec),
	.w5(32'h3aa88752),
	.w6(32'h3b163333),
	.w7(32'h3bdd4b6d),
	.w8(32'h3c888ff4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab16b9),
	.w1(32'hbb86b2d3),
	.w2(32'h3b1b3ece),
	.w3(32'hbc827539),
	.w4(32'hbc78e5eb),
	.w5(32'hbc96bf0a),
	.w6(32'hbb98ecb3),
	.w7(32'hbc38e4cb),
	.w8(32'hbc96d38b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf175ff),
	.w1(32'h3c666563),
	.w2(32'h3c223339),
	.w3(32'hbb182c42),
	.w4(32'h3b1eddfb),
	.w5(32'h3b97af03),
	.w6(32'h3c68ef60),
	.w7(32'h3bc114d4),
	.w8(32'h3c8e0b14),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d03e6),
	.w1(32'hbb85d6e9),
	.w2(32'hbbec2d52),
	.w3(32'h3af0aaed),
	.w4(32'hb8ed64a6),
	.w5(32'hba9f8f12),
	.w6(32'hbaaeee6d),
	.w7(32'hbb388b71),
	.w8(32'hbb3795db),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a5fe1),
	.w1(32'h393f2990),
	.w2(32'hba52cf4c),
	.w3(32'hb9f76914),
	.w4(32'h3a8ba383),
	.w5(32'hb9237f8f),
	.w6(32'hbaab48e3),
	.w7(32'hbafe9d65),
	.w8(32'hba17991c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e1e50),
	.w1(32'hba278b2d),
	.w2(32'h3a192881),
	.w3(32'hba7b336f),
	.w4(32'h3a0d3093),
	.w5(32'h3a4d592a),
	.w6(32'hba374240),
	.w7(32'hb91fbb04),
	.w8(32'h3b052930),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b48a2),
	.w1(32'h3a3008cd),
	.w2(32'hb9d35af5),
	.w3(32'hba19dd65),
	.w4(32'hbaee38c7),
	.w5(32'hba37198f),
	.w6(32'hba8dd6fe),
	.w7(32'hbb2be68f),
	.w8(32'hba4efed2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ec3ba),
	.w1(32'hbbf01c2c),
	.w2(32'hbc00dd7a),
	.w3(32'hbc00c782),
	.w4(32'hbc224f11),
	.w5(32'hbb9507c7),
	.w6(32'h3b8620a9),
	.w7(32'h3ab90ba5),
	.w8(32'h39aebac5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb881a89),
	.w1(32'hb8c5780b),
	.w2(32'hbac61dbb),
	.w3(32'hbacf1ffd),
	.w4(32'h3b25a45a),
	.w5(32'hbaa8eb74),
	.w6(32'hba53be54),
	.w7(32'hbb1a61bd),
	.w8(32'hba924136),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23ebd0),
	.w1(32'hbc5542a7),
	.w2(32'hbb3537ea),
	.w3(32'hbccb0e76),
	.w4(32'hbc3316a7),
	.w5(32'h3bb3c66d),
	.w6(32'hbb8a97f8),
	.w7(32'h3aed228f),
	.w8(32'h3c62bdfc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f21c1),
	.w1(32'hbb805d22),
	.w2(32'hbb7fe4f8),
	.w3(32'hbb5b1bf2),
	.w4(32'hbb916f4c),
	.w5(32'h399c2a39),
	.w6(32'hb998596a),
	.w7(32'h3b1ebfdc),
	.w8(32'h3b97a1a7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8fef4),
	.w1(32'h3c1fd261),
	.w2(32'h3c996907),
	.w3(32'h3c5adfd2),
	.w4(32'h3c16592d),
	.w5(32'hbc368d9d),
	.w6(32'h3d25edd5),
	.w7(32'h3c544a3f),
	.w8(32'hbcc7a480),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385d53c0),
	.w1(32'h3b280e24),
	.w2(32'h3b25a470),
	.w3(32'h3b502899),
	.w4(32'h3b5b7a6c),
	.w5(32'h3b869fe5),
	.w6(32'h3c4af259),
	.w7(32'h3c20cb05),
	.w8(32'h3bdaa587),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc033d44),
	.w1(32'hbbc0136d),
	.w2(32'hbb382285),
	.w3(32'hbc1ab474),
	.w4(32'hbb7b088c),
	.w5(32'h3a6c18e6),
	.w6(32'h3b61b5ab),
	.w7(32'h3b81adc8),
	.w8(32'h3bf7f95b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b954d97),
	.w1(32'hbb15e156),
	.w2(32'hbc036100),
	.w3(32'h3b4e8542),
	.w4(32'h3ae1de20),
	.w5(32'hbb76bda6),
	.w6(32'h3b32a358),
	.w7(32'h3b89fd18),
	.w8(32'hbb03b12d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc817103),
	.w1(32'hbc1dbb54),
	.w2(32'hbc17788c),
	.w3(32'hbbac08c2),
	.w4(32'hbbfca17e),
	.w5(32'hbbc23f67),
	.w6(32'h3bc8dc22),
	.w7(32'h3b689819),
	.w8(32'h3b0ce63c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195f68),
	.w1(32'hbb70b684),
	.w2(32'h3b9ecc71),
	.w3(32'h3b650ad9),
	.w4(32'hbad23091),
	.w5(32'hba99cab8),
	.w6(32'h39fa6b4a),
	.w7(32'h3b3340e2),
	.w8(32'h3c5188bf),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b11a6),
	.w1(32'h3c23b58b),
	.w2(32'h3c7bd73d),
	.w3(32'h3b4ddb85),
	.w4(32'h3a8e504a),
	.w5(32'h3c4cb221),
	.w6(32'h3bbf2fb3),
	.w7(32'h3b45067c),
	.w8(32'h3c1c0460),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4a1b),
	.w1(32'hbc2ece33),
	.w2(32'hbc6ecf11),
	.w3(32'hbbd359ed),
	.w4(32'hbc7dff03),
	.w5(32'hbc075b1c),
	.w6(32'hbbc19084),
	.w7(32'hbc3ef11e),
	.w8(32'hbb0b5e34),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19094f),
	.w1(32'h39b533e7),
	.w2(32'hba1734b3),
	.w3(32'h3a3fe683),
	.w4(32'hb94cb942),
	.w5(32'hba8bbdbe),
	.w6(32'hb9fe29b0),
	.w7(32'hb9f03539),
	.w8(32'hbab59bc9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb062b),
	.w1(32'h3bb6409b),
	.w2(32'hb831d602),
	.w3(32'h3bab3556),
	.w4(32'h3b8dfd72),
	.w5(32'h3a9f0b8d),
	.w6(32'h3b87c78e),
	.w7(32'hb990c34d),
	.w8(32'h3ab59df0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc92aa),
	.w1(32'h3b12f1ee),
	.w2(32'hbaa3e7a3),
	.w3(32'h3b0a2395),
	.w4(32'h3b24773b),
	.w5(32'hbb5b9010),
	.w6(32'h3aed579a),
	.w7(32'hba17c473),
	.w8(32'h39766661),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fe5ab),
	.w1(32'hbbc8bff3),
	.w2(32'hbafd6fe6),
	.w3(32'hba234710),
	.w4(32'hbb9e21a9),
	.w5(32'hbb919086),
	.w6(32'h3b68ff06),
	.w7(32'h3bb6a81c),
	.w8(32'hbb77ab11),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af79963),
	.w1(32'h3c0bd93b),
	.w2(32'h3c7d71fc),
	.w3(32'h3c7b048c),
	.w4(32'h3bf374e2),
	.w5(32'hba8bc2c7),
	.w6(32'h3c989482),
	.w7(32'h3b91a44d),
	.w8(32'hbb9f5390),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3543e),
	.w1(32'hb74bd169),
	.w2(32'hba2adc75),
	.w3(32'hb95226cf),
	.w4(32'h3a52e3e0),
	.w5(32'hba85b61c),
	.w6(32'h3a24206c),
	.w7(32'hb9dc7424),
	.w8(32'hbb5f9652),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb853b3b),
	.w1(32'hbaddc28e),
	.w2(32'hbab75881),
	.w3(32'hbb4afc78),
	.w4(32'hbb2dbf4e),
	.w5(32'hbb1f8e5d),
	.w6(32'hbb270fd5),
	.w7(32'hbb2315dd),
	.w8(32'hbb9b6dd1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4302b3),
	.w1(32'hbc1a6cb9),
	.w2(32'hbc6e2d6e),
	.w3(32'h393ca996),
	.w4(32'hbb802fa7),
	.w5(32'hbc990b6b),
	.w6(32'h3c0d3cfa),
	.w7(32'h3c0c435e),
	.w8(32'hbb8ad8af),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02ee5e),
	.w1(32'hbb999225),
	.w2(32'hb93ccfaf),
	.w3(32'h3b5db6a1),
	.w4(32'hbb7e49bb),
	.w5(32'hba23d58f),
	.w6(32'hbb06f5aa),
	.w7(32'hbc27d23d),
	.w8(32'h3a960f8e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb284348),
	.w1(32'hbb4351e6),
	.w2(32'hbaae2f26),
	.w3(32'hbac7e51e),
	.w4(32'hbadfde68),
	.w5(32'hbad0016e),
	.w6(32'hbb1e37f3),
	.w7(32'hbaee36d3),
	.w8(32'hbbab7e05),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae603ce),
	.w1(32'hbb950cae),
	.w2(32'hbbe9dc49),
	.w3(32'hba799d16),
	.w4(32'hbbbef44f),
	.w5(32'hbbc322e2),
	.w6(32'hbbcf6294),
	.w7(32'hbbc6710c),
	.w8(32'hbb5e9796),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cf00b),
	.w1(32'hba4f3a8f),
	.w2(32'hbaf9c04d),
	.w3(32'hbb6ad583),
	.w4(32'hb8197bcb),
	.w5(32'h383140e5),
	.w6(32'h3b674209),
	.w7(32'h3bb380b0),
	.w8(32'h3b775674),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0d822),
	.w1(32'h3a0647cd),
	.w2(32'h3be1dfa0),
	.w3(32'h3b065142),
	.w4(32'h3bb5bb29),
	.w5(32'hbb1981a1),
	.w6(32'h3c362508),
	.w7(32'h3b955880),
	.w8(32'hbb9a02bf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a206c9b),
	.w1(32'hbb40fae0),
	.w2(32'hb9c3ce4f),
	.w3(32'h3b07bb22),
	.w4(32'hbc00b29d),
	.w5(32'h38be534f),
	.w6(32'h3aca0ab1),
	.w7(32'h37fd5fef),
	.w8(32'h3bc866ce),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf41fee),
	.w1(32'h3bd064b0),
	.w2(32'h3c1eb744),
	.w3(32'h3baa2f2b),
	.w4(32'h3c68e437),
	.w5(32'h3a078942),
	.w6(32'h3c45877b),
	.w7(32'h3bef9d5b),
	.w8(32'hbc106e08),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule