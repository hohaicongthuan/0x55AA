module layer_10_featuremap_60(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc163fe5),
	.w1(32'hbbc1fea9),
	.w2(32'hbc96d28f),
	.w3(32'h3bc1f3d3),
	.w4(32'h3c3144e2),
	.w5(32'hba26d298),
	.w6(32'h3c9a1726),
	.w7(32'h3c744102),
	.w8(32'h3c18d085),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9043f),
	.w1(32'hbd003540),
	.w2(32'hbb91f62f),
	.w3(32'hbac9c233),
	.w4(32'hba9c81de),
	.w5(32'hbb766c35),
	.w6(32'hbb963731),
	.w7(32'h3bd97ed9),
	.w8(32'h3c286238),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87e64f),
	.w1(32'h3bac3ae6),
	.w2(32'h3b9431f6),
	.w3(32'h3bc946e2),
	.w4(32'h3bb541f3),
	.w5(32'hbbe79b6d),
	.w6(32'h3c16d337),
	.w7(32'h3ba84d88),
	.w8(32'hbbdc7760),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d47e0),
	.w1(32'h3bed20db),
	.w2(32'hbc9a9dc3),
	.w3(32'hbb28c46d),
	.w4(32'hbb687941),
	.w5(32'hbbd7cd35),
	.w6(32'h3a955c69),
	.w7(32'h37733383),
	.w8(32'hbc8fec71),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad5f0e),
	.w1(32'h3bcd7afd),
	.w2(32'h3b527109),
	.w3(32'h3880e142),
	.w4(32'hbbd6f447),
	.w5(32'hbc1b9c26),
	.w6(32'hbc025d76),
	.w7(32'hbc00abe5),
	.w8(32'h3b875dd0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc222669),
	.w1(32'hbba0493b),
	.w2(32'h3b600e3c),
	.w3(32'hbd08845f),
	.w4(32'hbc02fb7a),
	.w5(32'hbb966d39),
	.w6(32'hbc778673),
	.w7(32'h3aea6aa4),
	.w8(32'hba06dfd7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07df30),
	.w1(32'h3bc32344),
	.w2(32'h3d0a48d5),
	.w3(32'hbbd84fc0),
	.w4(32'hbbaec9db),
	.w5(32'h3ccc180c),
	.w6(32'hbc4ca083),
	.w7(32'h3c98acb7),
	.w8(32'h3ca818e9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e9f6f),
	.w1(32'h3c1720ba),
	.w2(32'hba804b29),
	.w3(32'hbc558926),
	.w4(32'hbbd52895),
	.w5(32'hbbef032e),
	.w6(32'h3ac1ff54),
	.w7(32'hbccb56e2),
	.w8(32'h3be15301),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc929282),
	.w1(32'hbc225f4a),
	.w2(32'h3b9135d4),
	.w3(32'hbbb4edf1),
	.w4(32'hbad18e7f),
	.w5(32'h39b2bf32),
	.w6(32'h3bfffdaf),
	.w7(32'h3be81992),
	.w8(32'h3b91d54d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39b0e9),
	.w1(32'h3be5b8a1),
	.w2(32'h3c747604),
	.w3(32'hbc04356b),
	.w4(32'hbb873e0f),
	.w5(32'h3c0c6e1d),
	.w6(32'hbc6b227c),
	.w7(32'hbc2d725f),
	.w8(32'h3b33ea0c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9086b6),
	.w1(32'h3baf0741),
	.w2(32'hbb84f5e0),
	.w3(32'h3be9541a),
	.w4(32'h3ba69815),
	.w5(32'hbab70274),
	.w6(32'h3b7dac9c),
	.w7(32'h3b5411c6),
	.w8(32'h3a6e172c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bdc8f),
	.w1(32'h3c099280),
	.w2(32'h3d01c98b),
	.w3(32'h3b5595f6),
	.w4(32'hbbe70e33),
	.w5(32'h3cb6035a),
	.w6(32'h3a26bab0),
	.w7(32'h3b46ca69),
	.w8(32'h3c81e45f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a4870),
	.w1(32'h3ca10dd6),
	.w2(32'h3cba2cf2),
	.w3(32'h3829fbd2),
	.w4(32'h3c01d586),
	.w5(32'h3c47167e),
	.w6(32'hbb216095),
	.w7(32'h3b5c27ec),
	.w8(32'hbb8df352),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c653f0d),
	.w1(32'h3c3e9c7c),
	.w2(32'h3b935442),
	.w3(32'h3bf21b73),
	.w4(32'h3c13a1a4),
	.w5(32'h3c9fc848),
	.w6(32'hb92aa9a4),
	.w7(32'h3ab9634b),
	.w8(32'h3c546c3e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b800d27),
	.w1(32'hbaf4108c),
	.w2(32'hbc338012),
	.w3(32'h3caec2ce),
	.w4(32'h3c83563b),
	.w5(32'hbb8f0bf4),
	.w6(32'h3b820a15),
	.w7(32'h3ae6e4cc),
	.w8(32'hbc05cdc7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c733a1f),
	.w1(32'h3b0f83a3),
	.w2(32'h3b2dfbc6),
	.w3(32'hbb4068c8),
	.w4(32'hba8aea5d),
	.w5(32'h3a7f3a13),
	.w6(32'hbcc9605c),
	.w7(32'hbc2c62f5),
	.w8(32'hbbb6c026),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b712d02),
	.w1(32'h3b6272d5),
	.w2(32'hbc6c9dac),
	.w3(32'h3b8c4c24),
	.w4(32'h3b48b460),
	.w5(32'hbc2bdfe4),
	.w6(32'h3b239f78),
	.w7(32'h3a9f7c83),
	.w8(32'h3be85adc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec8ea1),
	.w1(32'hbc0e3602),
	.w2(32'h3c4419a7),
	.w3(32'hbcca8720),
	.w4(32'hbbfc1416),
	.w5(32'h3ab72794),
	.w6(32'hbc45fdfe),
	.w7(32'h3b74b279),
	.w8(32'hbc7a005b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcca5c),
	.w1(32'h3c69d1ef),
	.w2(32'h3c17fc30),
	.w3(32'hbafeaa62),
	.w4(32'h3b8fc1aa),
	.w5(32'h3bd6192e),
	.w6(32'h3a94a97b),
	.w7(32'h3a25adf1),
	.w8(32'hbc1aed73),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3952e),
	.w1(32'h3bdc38b0),
	.w2(32'h3b67e9d2),
	.w3(32'h3c7135e8),
	.w4(32'h3c63fc40),
	.w5(32'hbb93cfa3),
	.w6(32'h3aaaa471),
	.w7(32'h3bc7a116),
	.w8(32'hbb988b56),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c2b05),
	.w1(32'hbbc6ce06),
	.w2(32'hbb4188de),
	.w3(32'hbb6adc1a),
	.w4(32'hbb73aefc),
	.w5(32'h3b976f48),
	.w6(32'hbb2cd3d0),
	.w7(32'h39e4a727),
	.w8(32'h3bd68eb1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0f930),
	.w1(32'h3c0edbb6),
	.w2(32'hbc3c1e4b),
	.w3(32'h3c50f065),
	.w4(32'h3cb08556),
	.w5(32'h398e1b7d),
	.w6(32'h3cf0aee2),
	.w7(32'h3cfa0a41),
	.w8(32'hbb85e3dc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1288e),
	.w1(32'hbb777057),
	.w2(32'h3c1732a1),
	.w3(32'h3b700a87),
	.w4(32'hbcdba30a),
	.w5(32'h3c4fc7a3),
	.w6(32'hbce27941),
	.w7(32'hbbcefffa),
	.w8(32'h3c4eaaa3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb121ec1),
	.w1(32'h3b1b01ba),
	.w2(32'hbb21cf27),
	.w3(32'hb9d1222f),
	.w4(32'h39fd34e1),
	.w5(32'hbba909b7),
	.w6(32'hbbd70c40),
	.w7(32'hbbd21c73),
	.w8(32'hbc55e1d5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c9550),
	.w1(32'hbd032239),
	.w2(32'hbd6f9ec2),
	.w3(32'h3b08e5b6),
	.w4(32'hbbbb78eb),
	.w5(32'hbcc4f500),
	.w6(32'h3b99e881),
	.w7(32'h3c2ed665),
	.w8(32'h3a8ed317),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2198ff),
	.w1(32'hbbf8c50f),
	.w2(32'hbb5b9a53),
	.w3(32'h3c115239),
	.w4(32'h3c389fdb),
	.w5(32'hbb4dad5d),
	.w6(32'h3b954d7f),
	.w7(32'hbb411312),
	.w8(32'hbbf81d0b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb394d8e),
	.w1(32'h3bade7f9),
	.w2(32'hbba5f6cd),
	.w3(32'h3b750437),
	.w4(32'h3beece0b),
	.w5(32'hbc78d6e8),
	.w6(32'hbc358891),
	.w7(32'hbbff4800),
	.w8(32'hbc843f41),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca54d6a),
	.w1(32'h3cc4348d),
	.w2(32'h3c7b89ff),
	.w3(32'hbb68f696),
	.w4(32'h3d68933f),
	.w5(32'h3cc5e5a1),
	.w6(32'hbd03b074),
	.w7(32'h3cc55390),
	.w8(32'h3c9b6711),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36a0e0),
	.w1(32'h3bff1b51),
	.w2(32'hbac16d9f),
	.w3(32'h3bdd4bbe),
	.w4(32'h3bdb649a),
	.w5(32'hbbc29744),
	.w6(32'h3bfba724),
	.w7(32'h3b49e929),
	.w8(32'hbb9d5175),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a870c),
	.w1(32'hbc574934),
	.w2(32'hbcfb1ef2),
	.w3(32'h3c27f4ed),
	.w4(32'h3ce0b9ed),
	.w5(32'h3c66a39b),
	.w6(32'hbad342fe),
	.w7(32'h3cd04dc8),
	.w8(32'hba884bdb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca43faf),
	.w1(32'hbc5e7498),
	.w2(32'h394aab38),
	.w3(32'hbaa6daf4),
	.w4(32'hbcdbc75c),
	.w5(32'hb9be1982),
	.w6(32'h3c30432c),
	.w7(32'hbc087ed4),
	.w8(32'hb8f8ca53),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a6d03),
	.w1(32'hbc0911ae),
	.w2(32'hb93e2104),
	.w3(32'h3bcbd2b0),
	.w4(32'h3b6e7c34),
	.w5(32'h3b8d1a45),
	.w6(32'h3b8715b0),
	.w7(32'h3ae04a7f),
	.w8(32'h3b3a95f4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ecd00),
	.w1(32'hba899e31),
	.w2(32'h3caa2e72),
	.w3(32'h3be3563b),
	.w4(32'h3c016ec2),
	.w5(32'h3dc22464),
	.w6(32'h39bf43cd),
	.w7(32'hba473a9a),
	.w8(32'h3d998966),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1ab1b9),
	.w1(32'hbda9dd51),
	.w2(32'hbc04aee0),
	.w3(32'h3ce5666c),
	.w4(32'hbda52c96),
	.w5(32'hbc002e98),
	.w6(32'h3d9b3f05),
	.w7(32'hbcb2af98),
	.w8(32'h3b213e05),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb566c20),
	.w1(32'hbbc88e68),
	.w2(32'h3c394593),
	.w3(32'hba610baa),
	.w4(32'h3b382897),
	.w5(32'h3b5b959b),
	.w6(32'hbbb19555),
	.w7(32'h3c1030c2),
	.w8(32'h3c43ffa1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0535b5),
	.w1(32'hbbae92e4),
	.w2(32'h3c232117),
	.w3(32'hbbb35b6c),
	.w4(32'hbc056050),
	.w5(32'h3ca7718f),
	.w6(32'hbbf59afa),
	.w7(32'h3a5fa880),
	.w8(32'h3c15f1f4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c3059),
	.w1(32'hbd3f5df3),
	.w2(32'h3c103515),
	.w3(32'hbb423a0b),
	.w4(32'hbd41927f),
	.w5(32'h3d8e6c13),
	.w6(32'hb9f628c8),
	.w7(32'hbcf63276),
	.w8(32'h3dcd084c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd52c655),
	.w1(32'hbdd60d2d),
	.w2(32'hbd366ab4),
	.w3(32'h3cec2615),
	.w4(32'hbd988b1c),
	.w5(32'hbc83d8a8),
	.w6(32'h3db65a50),
	.w7(32'hbaaa77ac),
	.w8(32'h3aaa1a34),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd873b2),
	.w1(32'h3c2fedb0),
	.w2(32'hbc9096d2),
	.w3(32'h3c82f3f5),
	.w4(32'h3cce4668),
	.w5(32'hbc50d2d3),
	.w6(32'h3bd0b804),
	.w7(32'h3d03da3b),
	.w8(32'hbb19b890),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8941b5a),
	.w1(32'hbc07f7ec),
	.w2(32'hbc11d289),
	.w3(32'h3af440d9),
	.w4(32'hbbad74e0),
	.w5(32'hbb84b5aa),
	.w6(32'hbc016745),
	.w7(32'hbb9a3a21),
	.w8(32'hbc2fc51c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7ef1a),
	.w1(32'h3bb5f033),
	.w2(32'hb9cbd807),
	.w3(32'hbb86bbdb),
	.w4(32'h39324441),
	.w5(32'hba8d6ff3),
	.w6(32'h3a9f2895),
	.w7(32'h3b65213d),
	.w8(32'hb7ea2bc7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdba77),
	.w1(32'h3aee31cd),
	.w2(32'h3bc0733f),
	.w3(32'h3aa29bcc),
	.w4(32'h3b2f4ae5),
	.w5(32'h3b138314),
	.w6(32'h3b1d698a),
	.w7(32'hba6aa3e3),
	.w8(32'h3b87cdbc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefcf5b),
	.w1(32'hba3faa52),
	.w2(32'hbce8f968),
	.w3(32'h3adfb2f3),
	.w4(32'hb9ef5fa7),
	.w5(32'hbddbf7ce),
	.w6(32'h3b887b16),
	.w7(32'h3aa088ee),
	.w8(32'hbdc2424e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3da8f7c2),
	.w1(32'h3de7456f),
	.w2(32'h3ca8d252),
	.w3(32'hbc4a218e),
	.w4(32'h3ddfa39d),
	.w5(32'h3c52fc86),
	.w6(32'hbda54845),
	.w7(32'h3d119c4b),
	.w8(32'hbc84537f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2180b),
	.w1(32'hbc84505d),
	.w2(32'hbc4fed0c),
	.w3(32'h3c255540),
	.w4(32'hbb994c6b),
	.w5(32'hbb52ab61),
	.w6(32'h3bc865ef),
	.w7(32'h3aa23aba),
	.w8(32'hbc0650c3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb68406),
	.w1(32'hbc27cf16),
	.w2(32'hbc523a13),
	.w3(32'hbb6bc377),
	.w4(32'hbbefd2d2),
	.w5(32'hbbfc8f8b),
	.w6(32'hbb06806c),
	.w7(32'hba585bde),
	.w8(32'hbc128bca),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b517662),
	.w1(32'hbbb5f21b),
	.w2(32'hbc19065c),
	.w3(32'h3b286400),
	.w4(32'h3a9c9173),
	.w5(32'h3ad9802b),
	.w6(32'hbc20d296),
	.w7(32'hbae7cdcf),
	.w8(32'hbaaafeae),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab419f),
	.w1(32'h3d099d08),
	.w2(32'h3d2aad0d),
	.w3(32'hbca5c2fa),
	.w4(32'h3b549b64),
	.w5(32'hbbb5aede),
	.w6(32'hbcccc4fe),
	.w7(32'hbc7dca5a),
	.w8(32'hbb0e94b9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc7c970),
	.w1(32'h3c84480e),
	.w2(32'h3b569ddc),
	.w3(32'h39775e33),
	.w4(32'h3cebe17c),
	.w5(32'h3aac780e),
	.w6(32'hbc5e0f9f),
	.w7(32'h3c36782e),
	.w8(32'h3afbf173),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2645fb),
	.w1(32'hba899115),
	.w2(32'h3b4582af),
	.w3(32'hbb03a989),
	.w4(32'hbb5f97fb),
	.w5(32'h3bd0d0b2),
	.w6(32'hb9997808),
	.w7(32'hbbec1227),
	.w8(32'h3a7ee8f2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89735d),
	.w1(32'h3b122d6c),
	.w2(32'h3a8b1f06),
	.w3(32'h3bac7010),
	.w4(32'h3b41b8b9),
	.w5(32'h3bc977e0),
	.w6(32'h3af6b295),
	.w7(32'hbb311a1b),
	.w8(32'h3afddddb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabfb5b),
	.w1(32'h3a44af9c),
	.w2(32'h3b237f55),
	.w3(32'h3c2f5808),
	.w4(32'hbb0c6938),
	.w5(32'h3bcb4d14),
	.w6(32'hb9eee6a8),
	.w7(32'hbb648a6e),
	.w8(32'hbb1dd0e4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba877794),
	.w1(32'h3b857fb2),
	.w2(32'hbb6a791f),
	.w3(32'h3b8e8c4e),
	.w4(32'hbb9d25f5),
	.w5(32'hbab7f767),
	.w6(32'hbb62b62a),
	.w7(32'hbb78c2bd),
	.w8(32'h3b93f800),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca78026),
	.w1(32'h3cc078bf),
	.w2(32'h3cfdb568),
	.w3(32'hbbf49a5a),
	.w4(32'h3af59223),
	.w5(32'h3c9e82f6),
	.w6(32'hbc0c2daf),
	.w7(32'hbc23a906),
	.w8(32'hbbd7413e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb235d),
	.w1(32'h3c162f2d),
	.w2(32'h3b333d1d),
	.w3(32'hbb941333),
	.w4(32'h3b63fb68),
	.w5(32'hbb02afae),
	.w6(32'hba845b8f),
	.w7(32'hbb4e26ca),
	.w8(32'hbab9204e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bcfa4),
	.w1(32'h3a8ff8fb),
	.w2(32'hbb499b2c),
	.w3(32'hbb4f20d1),
	.w4(32'hb9a17312),
	.w5(32'hbbda1d0d),
	.w6(32'h3b224c52),
	.w7(32'h3a9f41a6),
	.w8(32'hbbe5fcfb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba887d47),
	.w1(32'hbaebe1c8),
	.w2(32'h3909ed92),
	.w3(32'h3afb1b8f),
	.w4(32'hbb837f83),
	.w5(32'hbaf3ce63),
	.w6(32'hbb83d19c),
	.w7(32'hba8dccbe),
	.w8(32'hbbcca09c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ae481),
	.w1(32'hbbc1bae3),
	.w2(32'hbb9274ec),
	.w3(32'hbc00a8fb),
	.w4(32'hbb4a093f),
	.w5(32'hba1b7781),
	.w6(32'hbc5c33a9),
	.w7(32'hbaddec24),
	.w8(32'hbbd2d540),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbace210),
	.w1(32'hbc2663b9),
	.w2(32'h3a8f5456),
	.w3(32'hbb8c003e),
	.w4(32'hbc609190),
	.w5(32'h3abf32d5),
	.w6(32'hbc07f8da),
	.w7(32'hbc735107),
	.w8(32'hba7b6ff1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe0c2a),
	.w1(32'h3bd3ec22),
	.w2(32'h3b0a52d4),
	.w3(32'h3b5a5b56),
	.w4(32'h3c16a8bf),
	.w5(32'h3ba7d848),
	.w6(32'hbaa37e06),
	.w7(32'h3b77fa48),
	.w8(32'hbb6c504a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc35fb4),
	.w1(32'hbaa316e8),
	.w2(32'h3ac97cbb),
	.w3(32'h3a86d243),
	.w4(32'h3a9fe512),
	.w5(32'hbc2a1f3b),
	.w6(32'hbb16fdff),
	.w7(32'h3b205388),
	.w8(32'hbbdec8e5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00ed19),
	.w1(32'hbba2e4e7),
	.w2(32'hbc131128),
	.w3(32'hb987ba72),
	.w4(32'h3c46f700),
	.w5(32'hba057751),
	.w6(32'hbbb4941f),
	.w7(32'h3c2fe568),
	.w8(32'hbc355082),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f734a),
	.w1(32'h3b639ceb),
	.w2(32'hbb4e2e68),
	.w3(32'hbb89ace3),
	.w4(32'h3b25246f),
	.w5(32'h3c191904),
	.w6(32'hbb2d56f1),
	.w7(32'hbb35139f),
	.w8(32'hbaa56d6a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ae283),
	.w1(32'h3b040029),
	.w2(32'hba8f2bee),
	.w3(32'h3c14967e),
	.w4(32'h3be2b3e4),
	.w5(32'h3b008415),
	.w6(32'h3b9ad22d),
	.w7(32'h3ba9fc6f),
	.w8(32'h3a96fb09),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6cb75),
	.w1(32'h3ae77ea5),
	.w2(32'h3bcc1387),
	.w3(32'h3b32753d),
	.w4(32'h3ae74cdc),
	.w5(32'h3c32f494),
	.w6(32'h3add918b),
	.w7(32'h39863445),
	.w8(32'h3bd96e0f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fb37a),
	.w1(32'h3a864684),
	.w2(32'hbc98e76f),
	.w3(32'h3c2c9f94),
	.w4(32'h3bd8b701),
	.w5(32'hbd83dd03),
	.w6(32'h3c2096a7),
	.w7(32'h3c16af7d),
	.w8(32'hbd97addb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6e88e1),
	.w1(32'h3de70691),
	.w2(32'h3c72f92f),
	.w3(32'h3ae53299),
	.w4(32'h3ddd5a42),
	.w5(32'h3c7b75a7),
	.w6(32'hbd65c353),
	.w7(32'h3ce41820),
	.w8(32'hbb981543),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3aa5e),
	.w1(32'hbbea61c1),
	.w2(32'h3ba8982b),
	.w3(32'hbc254ee0),
	.w4(32'h391b20e0),
	.w5(32'h3c168731),
	.w6(32'h3b8af155),
	.w7(32'h3b59f871),
	.w8(32'hbc9da072),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc7c3ce),
	.w1(32'h3b1eccb6),
	.w2(32'hbba46255),
	.w3(32'h3b66346e),
	.w4(32'hba280055),
	.w5(32'hbba8125a),
	.w6(32'hbb89a733),
	.w7(32'h3b876a60),
	.w8(32'hbc6b9103),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc005d94),
	.w1(32'hbcd3b132),
	.w2(32'hbd25ce0f),
	.w3(32'h3c334c23),
	.w4(32'h3c725715),
	.w5(32'hbbf8dec1),
	.w6(32'h3ce6bc2c),
	.w7(32'h3d0a9ac4),
	.w8(32'h3addea1f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b872c),
	.w1(32'h3bdec30e),
	.w2(32'h3a9e8afb),
	.w3(32'h3bd0fc63),
	.w4(32'h3bfc0713),
	.w5(32'h3b6e7554),
	.w6(32'hbaeac8ec),
	.w7(32'hba5b3006),
	.w8(32'h3bbfcc91),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972526c),
	.w1(32'hbbba594f),
	.w2(32'h3c1595b8),
	.w3(32'h3b40445a),
	.w4(32'hbaa63a42),
	.w5(32'h3bf6971f),
	.w6(32'h3c01ea97),
	.w7(32'h39cd915e),
	.w8(32'h3bc18b44),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf191a3),
	.w1(32'hbbca4f00),
	.w2(32'h3bcfe471),
	.w3(32'h3aa206be),
	.w4(32'hbb37ba42),
	.w5(32'hbb0998f6),
	.w6(32'h3ab5a628),
	.w7(32'h3b1cd419),
	.w8(32'hbba31eb5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a826a),
	.w1(32'h3c173125),
	.w2(32'h3b8e706b),
	.w3(32'hbc0694df),
	.w4(32'h3bc16237),
	.w5(32'hbd2094e7),
	.w6(32'hbbc28bea),
	.w7(32'hbb2ae497),
	.w8(32'hbd184d36),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50ec86),
	.w1(32'h3d2bcc56),
	.w2(32'h3bb1b819),
	.w3(32'hbc9c11a3),
	.w4(32'h3d227ae2),
	.w5(32'h3bab36f0),
	.w6(32'hbd17d0ea),
	.w7(32'h3ca550f6),
	.w8(32'h3bb7f306),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadf0f2),
	.w1(32'h3c858c4d),
	.w2(32'h3c999985),
	.w3(32'hbb53f9ad),
	.w4(32'hba003619),
	.w5(32'h3c4cb0a7),
	.w6(32'hbbcb78d5),
	.w7(32'hb9d34642),
	.w8(32'h3c1e795d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d2fb1),
	.w1(32'h3c1f94e5),
	.w2(32'h3cae2b78),
	.w3(32'hbc0f8451),
	.w4(32'h3a60fdbe),
	.w5(32'h3c19878a),
	.w6(32'hbb8c76e6),
	.w7(32'hbc07011f),
	.w8(32'h3c06d90a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89160d),
	.w1(32'hbc4ea573),
	.w2(32'hbc91edf7),
	.w3(32'h3c1bc099),
	.w4(32'h3ab199fe),
	.w5(32'hbc0287e7),
	.w6(32'h3c037554),
	.w7(32'hbb2573d2),
	.w8(32'hbaac1753),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d7f1),
	.w1(32'hba2f573a),
	.w2(32'hbc0363c7),
	.w3(32'hbc9f4ae2),
	.w4(32'hbbcf0119),
	.w5(32'hbcd2ffed),
	.w6(32'hbc15d55b),
	.w7(32'h39ad81ef),
	.w8(32'hbcfedc5d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7d0c1),
	.w1(32'h3d0d240b),
	.w2(32'h3c3e9e22),
	.w3(32'hbc4262ac),
	.w4(32'h3d04afde),
	.w5(32'h3ca4604f),
	.w6(32'hbcb38246),
	.w7(32'h3b814b6a),
	.w8(32'h3c5d3e24),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f4f90),
	.w1(32'h3ba08e94),
	.w2(32'hbc9d6697),
	.w3(32'hba6d0e34),
	.w4(32'h3c1dce78),
	.w5(32'hbd519a82),
	.w6(32'hbb3093d5),
	.w7(32'h3b91218d),
	.w8(32'hbd8ec1a0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8497cc),
	.w1(32'h3daf696a),
	.w2(32'h3c5e5f4d),
	.w3(32'hbc6a3fc3),
	.w4(32'h3d792015),
	.w5(32'h3c4cdc4e),
	.w6(32'hbd27933f),
	.w7(32'h3cefc860),
	.w8(32'h3bb72c50),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b52d5),
	.w1(32'h3c08096e),
	.w2(32'hba5a431e),
	.w3(32'h3bacaab0),
	.w4(32'h3b575db3),
	.w5(32'h394a55ba),
	.w6(32'h3b9bad58),
	.w7(32'h3bba62d6),
	.w8(32'h3b985467),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68f147),
	.w1(32'hbb330403),
	.w2(32'h3b4c9a6e),
	.w3(32'hbbaaa623),
	.w4(32'h3a04620b),
	.w5(32'h3b8bd38a),
	.w6(32'hbbc2c77b),
	.w7(32'hbb894b2f),
	.w8(32'h3ba909c7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38c972),
	.w1(32'hba110b7a),
	.w2(32'h3c1869df),
	.w3(32'h3c2e1f2a),
	.w4(32'h3b049e54),
	.w5(32'h3c22e5dd),
	.w6(32'h3ba7a392),
	.w7(32'h3b1afe09),
	.w8(32'h375f6bda),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba028d8),
	.w1(32'hba4ca8f9),
	.w2(32'hbbd5a930),
	.w3(32'h3c25b57c),
	.w4(32'hba669728),
	.w5(32'h3978c7c7),
	.w6(32'h3b5d43a5),
	.w7(32'h3ba7c07e),
	.w8(32'hb927d09e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4748b),
	.w1(32'hbc98e2ea),
	.w2(32'hbc3e086a),
	.w3(32'h3c282428),
	.w4(32'h385c3339),
	.w5(32'hbcea9c20),
	.w6(32'h3c87f8f9),
	.w7(32'h3be0295e),
	.w8(32'hbccb80f7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c578a54),
	.w1(32'h3cf213e3),
	.w2(32'hba787025),
	.w3(32'hbb31fd83),
	.w4(32'h3cf87feb),
	.w5(32'h3ae6ce7c),
	.w6(32'hbc9391aa),
	.w7(32'h3c4b0777),
	.w8(32'hbad82bd3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ee25c),
	.w1(32'hbc9cd7df),
	.w2(32'hbc8ed0a9),
	.w3(32'hbae1bcc3),
	.w4(32'hbc2bdac9),
	.w5(32'hbb8302ec),
	.w6(32'h3b426701),
	.w7(32'hbb27e4b0),
	.w8(32'hbb6ad793),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c60ec),
	.w1(32'h3b8c2ff4),
	.w2(32'h3ce3f88b),
	.w3(32'hbc5329a2),
	.w4(32'hbbe96b0e),
	.w5(32'h3ca3831a),
	.w6(32'hbc97d183),
	.w7(32'hbb478eee),
	.w8(32'hbc40c95c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d9b90),
	.w1(32'h3b91603b),
	.w2(32'h3c35b3ac),
	.w3(32'h3cc1dcd2),
	.w4(32'h3c9ece36),
	.w5(32'h3ce91454),
	.w6(32'hb9a2915a),
	.w7(32'h3c694803),
	.w8(32'h3ca900ad),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ce0df),
	.w1(32'h3ae7edcb),
	.w2(32'h3c98be48),
	.w3(32'h3c45f5ea),
	.w4(32'hbbdd9edb),
	.w5(32'h3b774c1c),
	.w6(32'hbbcefc9d),
	.w7(32'h3c9b721c),
	.w8(32'hbace89f6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6f372),
	.w1(32'h3c1bc7c4),
	.w2(32'hbcef35c3),
	.w3(32'h3c25aceb),
	.w4(32'h3bfa8de3),
	.w5(32'hbdaf0e39),
	.w6(32'h3c2bfff9),
	.w7(32'h3c34f410),
	.w8(32'hbdbf71da),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d37f1ad),
	.w1(32'h3dc88d10),
	.w2(32'h3b6fd651),
	.w3(32'hbcd58a57),
	.w4(32'h3dbc5467),
	.w5(32'h3a012c55),
	.w6(32'hbd8ce85e),
	.w7(32'h3d189f5e),
	.w8(32'hbbba6ceb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69eb64),
	.w1(32'hbbc6379e),
	.w2(32'hbb27aca2),
	.w3(32'h3a81a841),
	.w4(32'h3bffc27c),
	.w5(32'hbb68f780),
	.w6(32'hbc0ad6e7),
	.w7(32'h3a13b4fe),
	.w8(32'hbbc35b89),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af5fd),
	.w1(32'hbbcec5f1),
	.w2(32'hbcee4fe0),
	.w3(32'h3c689513),
	.w4(32'h3c8063ce),
	.w5(32'hbc21a19c),
	.w6(32'h3bb2be3c),
	.w7(32'h3c856d2d),
	.w8(32'hbc2c86f2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1978d8),
	.w1(32'hbbc93ca3),
	.w2(32'h3b91969f),
	.w3(32'hbbe69854),
	.w4(32'hbb9b9428),
	.w5(32'hbaecc85c),
	.w6(32'hbbaa3163),
	.w7(32'hbb0e3beb),
	.w8(32'hbb5f29f3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf68895),
	.w1(32'h3c3d6bb7),
	.w2(32'h3bb5c03f),
	.w3(32'hbb8981ca),
	.w4(32'h39bd1952),
	.w5(32'h3c709f0b),
	.w6(32'hbc5b4770),
	.w7(32'hbb9588d4),
	.w8(32'hbac005bd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30b2d7),
	.w1(32'h3c33fd18),
	.w2(32'h3ca99da6),
	.w3(32'h3b66d4e2),
	.w4(32'h3abc0e11),
	.w5(32'h3bb08219),
	.w6(32'hbb4882a6),
	.w7(32'hbb62dd3f),
	.w8(32'h3c83c69c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b4219),
	.w1(32'hbcbb98ee),
	.w2(32'hbcb4c93a),
	.w3(32'hbc17e751),
	.w4(32'hbd43cf8a),
	.w5(32'hbc00d75d),
	.w6(32'h390d20f3),
	.w7(32'hbca1f24e),
	.w8(32'h3c8e57ea),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14ff15),
	.w1(32'hbc3ae5f6),
	.w2(32'hbcce11d1),
	.w3(32'h3cbdff4e),
	.w4(32'h3bffbcd9),
	.w5(32'hbc97d029),
	.w6(32'h3cd016e2),
	.w7(32'h3ca75b14),
	.w8(32'hbc340a11),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba694303),
	.w1(32'hbcaa11a9),
	.w2(32'hbcaf063d),
	.w3(32'h3a1ddec4),
	.w4(32'hbbc7c0e3),
	.w5(32'hbbf58136),
	.w6(32'h3c59c78b),
	.w7(32'h3bdca401),
	.w8(32'hbc39ed49),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917ed6),
	.w1(32'h3c74be11),
	.w2(32'h3c91d959),
	.w3(32'hbba95181),
	.w4(32'hbc54dac1),
	.w5(32'h3becd0c6),
	.w6(32'hbc9fdf7f),
	.w7(32'hbc6a831a),
	.w8(32'hbb8241c9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad595b),
	.w1(32'h39e04587),
	.w2(32'h3b2a4e73),
	.w3(32'h3ac332d7),
	.w4(32'hbb0c918f),
	.w5(32'h3bc7e413),
	.w6(32'hbc73c4e3),
	.w7(32'hbb1c3ed4),
	.w8(32'h3b70a911),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7e6c9),
	.w1(32'hbc52bbbb),
	.w2(32'hbb892ea5),
	.w3(32'hbbd8e6ba),
	.w4(32'hbd05a793),
	.w5(32'hbc58d227),
	.w6(32'h3b2d05b7),
	.w7(32'hbcadf6a8),
	.w8(32'h3ca58507),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28d31d),
	.w1(32'h3bfeeccb),
	.w2(32'h3ca55063),
	.w3(32'h3c2dc3b8),
	.w4(32'hbb9e493b),
	.w5(32'h3c435b74),
	.w6(32'hbb3830a1),
	.w7(32'h3ae1756e),
	.w8(32'h3ca43e86),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac589c5),
	.w1(32'h3948e309),
	.w2(32'hbb761a0d),
	.w3(32'hbacf10f8),
	.w4(32'h3b4bb482),
	.w5(32'h3b4afd03),
	.w6(32'hbad03fef),
	.w7(32'h3964cabd),
	.w8(32'h3c1616ad),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba187e45),
	.w1(32'hbb4e675f),
	.w2(32'hbb392d0d),
	.w3(32'hba878a21),
	.w4(32'h3b15377a),
	.w5(32'hba278d25),
	.w6(32'h3be55531),
	.w7(32'h3bf6dc55),
	.w8(32'h3aa66cf4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4172a),
	.w1(32'h3c5063ac),
	.w2(32'h3c453da1),
	.w3(32'h39eae050),
	.w4(32'h3c5de5bd),
	.w5(32'h3c2db93d),
	.w6(32'hbc1c2383),
	.w7(32'h3b1737f2),
	.w8(32'h3ab949f7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaebe26),
	.w1(32'hbc3c4bcf),
	.w2(32'hbc3e9dac),
	.w3(32'h3bbe0edb),
	.w4(32'hba206fa2),
	.w5(32'hbb809b68),
	.w6(32'h3b8beb6f),
	.w7(32'h3bc26284),
	.w8(32'hbb86adf1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e1049),
	.w1(32'h3c2c5112),
	.w2(32'hbb8a430e),
	.w3(32'h3c41a17c),
	.w4(32'h3cbec75d),
	.w5(32'h3a7c7f0c),
	.w6(32'h3b6e0b69),
	.w7(32'h3c4ca972),
	.w8(32'h3ae32403),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51324d),
	.w1(32'hbc3ee370),
	.w2(32'hbc488027),
	.w3(32'hbc139054),
	.w4(32'hbc003f2f),
	.w5(32'hbac1c945),
	.w6(32'hbb478932),
	.w7(32'hbb084c13),
	.w8(32'hbb64fc8f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa169b),
	.w1(32'hbca80c80),
	.w2(32'hbc900528),
	.w3(32'hbb9736c0),
	.w4(32'hbc9cc05e),
	.w5(32'hbc15ae83),
	.w6(32'h3c1631b6),
	.w7(32'h3b1d7390),
	.w8(32'hbbbd7f76),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89588f),
	.w1(32'h3bb4c439),
	.w2(32'h3aede4a0),
	.w3(32'h3b83b6a4),
	.w4(32'h3b85b156),
	.w5(32'h3a7024ca),
	.w6(32'hbbf1792d),
	.w7(32'hbad4e256),
	.w8(32'hbaf14bd3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02bb5f),
	.w1(32'hba6a1742),
	.w2(32'hbb93132b),
	.w3(32'h3b127c61),
	.w4(32'h3ab45029),
	.w5(32'h3ab00907),
	.w6(32'hbbb4244c),
	.w7(32'h3ae74779),
	.w8(32'h3ae2d0dd),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa44bb4),
	.w1(32'h3b97daf9),
	.w2(32'h3adb72e2),
	.w3(32'h3a200fc3),
	.w4(32'hbbc0e2b5),
	.w5(32'hbb1df708),
	.w6(32'h3c244b0b),
	.w7(32'hb92830c5),
	.w8(32'hba184e85),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba264f1),
	.w1(32'hbb6d2f28),
	.w2(32'hbb8535ea),
	.w3(32'hbb1e4526),
	.w4(32'hb969d400),
	.w5(32'hba0e61b8),
	.w6(32'h3a7cfe08),
	.w7(32'h39cf0e7f),
	.w8(32'h3b176b2f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34a56a),
	.w1(32'h3a874d2e),
	.w2(32'h39636abc),
	.w3(32'hbb86479c),
	.w4(32'hbb77e774),
	.w5(32'hbaaac29e),
	.w6(32'h3a7fcf75),
	.w7(32'h3b04c0d9),
	.w8(32'h3b088da8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c1048),
	.w1(32'hbbf5282b),
	.w2(32'h3a83e895),
	.w3(32'h3b5f08d6),
	.w4(32'h3b1281b8),
	.w5(32'h3c1bfbfd),
	.w6(32'h3a91304d),
	.w7(32'hbb8ecdb2),
	.w8(32'h3bddfac5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68fb7d),
	.w1(32'hbc0c013a),
	.w2(32'hbba8debb),
	.w3(32'hbb11ba98),
	.w4(32'h3b09d131),
	.w5(32'hbbc0d7e6),
	.w6(32'h39847568),
	.w7(32'hbb2182fc),
	.w8(32'hba2836d9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abba3ae),
	.w1(32'h3844c1a6),
	.w2(32'hb97c4eec),
	.w3(32'hb990dbc0),
	.w4(32'hbb12faa0),
	.w5(32'h3cbc3375),
	.w6(32'h3a94aa6a),
	.w7(32'hbb550d6a),
	.w8(32'h3cc6cc1d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75b873),
	.w1(32'hbcade782),
	.w2(32'h3c5a1bdd),
	.w3(32'hbbd961d9),
	.w4(32'hbd013f97),
	.w5(32'h3ca509d1),
	.w6(32'h3c39867e),
	.w7(32'hbc8274f1),
	.w8(32'h3c0f9bb7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5180e),
	.w1(32'hbd31f0db),
	.w2(32'hbd2138a6),
	.w3(32'hba8109bf),
	.w4(32'hbca16d50),
	.w5(32'hbc84dd1e),
	.w6(32'h3caeb198),
	.w7(32'h3c1ec985),
	.w8(32'h39f7721b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35424a),
	.w1(32'hbb9d96c9),
	.w2(32'h38854025),
	.w3(32'hbbb25ad8),
	.w4(32'h3a82007e),
	.w5(32'h3afb8c4a),
	.w6(32'h3a7fdcd9),
	.w7(32'h3a9ce8d9),
	.w8(32'h3a380eb8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e5e5c),
	.w1(32'hbaefdd66),
	.w2(32'h3a5147a6),
	.w3(32'h3b441406),
	.w4(32'hbb150382),
	.w5(32'hba5b9fcf),
	.w6(32'hb9f31b04),
	.w7(32'h3a1f1a80),
	.w8(32'h3b8bde11),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70bdfd),
	.w1(32'hbad27c2e),
	.w2(32'h3ba2a4f7),
	.w3(32'h3bb4a42d),
	.w4(32'h3b5eab59),
	.w5(32'hba91d328),
	.w6(32'h3bb15b53),
	.w7(32'hbb166238),
	.w8(32'h3b245b49),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b4200),
	.w1(32'h397a8c1c),
	.w2(32'h38ad0bc3),
	.w3(32'h3c0d4932),
	.w4(32'h3b2f47c7),
	.w5(32'h3b34cb67),
	.w6(32'h3b875078),
	.w7(32'h3b519c03),
	.w8(32'h3b752b30),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd51e57),
	.w1(32'hbc86ced7),
	.w2(32'hbc02394f),
	.w3(32'hbb9ff69a),
	.w4(32'hbc0c793b),
	.w5(32'h3c79867c),
	.w6(32'h3c1886f7),
	.w7(32'h3ca4d041),
	.w8(32'h3ab07b3d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7945f3),
	.w1(32'h3c50785c),
	.w2(32'h3c7d609b),
	.w3(32'hbb9d3143),
	.w4(32'h3c1e872f),
	.w5(32'h3c2d6921),
	.w6(32'hbc18bf72),
	.w7(32'hbbc4e670),
	.w8(32'h3b50f613),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9aa20),
	.w1(32'h3be2f0af),
	.w2(32'h3b79fd2e),
	.w3(32'hbb933fb9),
	.w4(32'h3b11c4d8),
	.w5(32'h3babe1c6),
	.w6(32'hbbb759cd),
	.w7(32'h39f4d96f),
	.w8(32'h3b3c256d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3f568),
	.w1(32'hb9c55798),
	.w2(32'h3a8b8021),
	.w3(32'h3b5efd3d),
	.w4(32'h392abea5),
	.w5(32'h3aeb2af5),
	.w6(32'h3b8d2f5c),
	.w7(32'h3b4835a5),
	.w8(32'h3ac1269b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d403b),
	.w1(32'hba76b77b),
	.w2(32'hba82c08f),
	.w3(32'h3b36f8f4),
	.w4(32'hb93f20e6),
	.w5(32'h3b9a7e6c),
	.w6(32'hb820c4f6),
	.w7(32'h3a39c116),
	.w8(32'hbaade435),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b832553),
	.w1(32'hbb0d1f71),
	.w2(32'hbbc2308e),
	.w3(32'hbb04b85b),
	.w4(32'h3b5075c8),
	.w5(32'hbbe6ad33),
	.w6(32'hbc0dfe65),
	.w7(32'hbb70a098),
	.w8(32'hbc386a18),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd39543),
	.w1(32'hbc0f613d),
	.w2(32'hbd0f0c4e),
	.w3(32'h39c09d17),
	.w4(32'h3b808f80),
	.w5(32'hbdf4d464),
	.w6(32'hbc02e62d),
	.w7(32'hbb67848c),
	.w8(32'hbde364df),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1df61d),
	.w1(32'h3e013091),
	.w2(32'h3cc6e91c),
	.w3(32'hbd5c9786),
	.w4(32'h3dcf9ed0),
	.w5(32'h3c8c4e95),
	.w6(32'hbdd8ab89),
	.w7(32'h3d17ea86),
	.w8(32'h3ba4b179),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fee85),
	.w1(32'hbc24ee54),
	.w2(32'hbc83cfa7),
	.w3(32'hba112a43),
	.w4(32'hbbdd05a9),
	.w5(32'h3b1d2de6),
	.w6(32'h3bd8a871),
	.w7(32'h3b48301a),
	.w8(32'h3b187c25),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba09197),
	.w1(32'h3c07eb18),
	.w2(32'h39aeb0e3),
	.w3(32'hbbf2abfd),
	.w4(32'h3bdbb2d9),
	.w5(32'hbb2353f7),
	.w6(32'h39f16410),
	.w7(32'h3a9c7791),
	.w8(32'hbb8b85bc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc042d9),
	.w1(32'h3cae5276),
	.w2(32'h3c5839dd),
	.w3(32'hbc1aeacf),
	.w4(32'hbc68cf7f),
	.w5(32'h3bfcb240),
	.w6(32'hbcaaa3c3),
	.w7(32'hbc80f784),
	.w8(32'hbc6bb5bc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc841f72),
	.w1(32'hbc33c35e),
	.w2(32'hbc6e1a47),
	.w3(32'hbb2ebdfd),
	.w4(32'hbc2774ea),
	.w5(32'hbc16d429),
	.w6(32'h39f4b3b9),
	.w7(32'h390c93a7),
	.w8(32'hba857f91),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6e4dc),
	.w1(32'h3c0391c8),
	.w2(32'h3be90cb8),
	.w3(32'hbb5412d8),
	.w4(32'h3bdea4a1),
	.w5(32'hbb79da9c),
	.w6(32'h3a987b59),
	.w7(32'hbbcc7528),
	.w8(32'h3a47c554),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7586a6),
	.w1(32'h3b00eb4f),
	.w2(32'hbbef0817),
	.w3(32'hbbd5e054),
	.w4(32'hbade63c2),
	.w5(32'hbbc12e39),
	.w6(32'hbbe201b2),
	.w7(32'hbb4c536f),
	.w8(32'hbc1fb23a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51c4f3),
	.w1(32'hbb9f76e2),
	.w2(32'hbd03c2d2),
	.w3(32'hbae4cc8d),
	.w4(32'h3c542e54),
	.w5(32'hbc13ee33),
	.w6(32'hbbd1a531),
	.w7(32'h3c42679f),
	.w8(32'hbc8532b0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bdb73),
	.w1(32'hbbe69cd8),
	.w2(32'hbbd17538),
	.w3(32'h3b438954),
	.w4(32'h3b3c5e98),
	.w5(32'hbb41109b),
	.w6(32'h3ba4ffae),
	.w7(32'h3ac4b237),
	.w8(32'h3b512927),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf204c7),
	.w1(32'h39a68b68),
	.w2(32'hbc2a62e1),
	.w3(32'hbaefde61),
	.w4(32'h3b00de50),
	.w5(32'hbcf956b0),
	.w6(32'h3b9ebae7),
	.w7(32'hbb5f9587),
	.w8(32'hbd3338e3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b4604),
	.w1(32'h3d249ab8),
	.w2(32'hbb7d149b),
	.w3(32'hbb10ac9f),
	.w4(32'h3d0a431a),
	.w5(32'hb9e304a3),
	.w6(32'hbc941783),
	.w7(32'h3c8158a5),
	.w8(32'hbacf7e34),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9359fc),
	.w1(32'hbaa236d6),
	.w2(32'hbba28b86),
	.w3(32'h3baa3e1d),
	.w4(32'hba912e23),
	.w5(32'hbaf553e9),
	.w6(32'hbb9e455c),
	.w7(32'hbabfe7a5),
	.w8(32'hbb95f64c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10aea8),
	.w1(32'hbc8915f1),
	.w2(32'hbc21a0ed),
	.w3(32'h3b88fca9),
	.w4(32'h3be32fc8),
	.w5(32'hbb01ddcc),
	.w6(32'h3c2bde20),
	.w7(32'h3c624453),
	.w8(32'h3c2440b4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f9ba4),
	.w1(32'h3b6cc7da),
	.w2(32'h3b802b74),
	.w3(32'hbb366f24),
	.w4(32'h3afce1ee),
	.w5(32'h3bd51b2c),
	.w6(32'hbc132d17),
	.w7(32'hbb5ac4d8),
	.w8(32'hbb172342),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e52a2),
	.w1(32'hba6b6182),
	.w2(32'hbb08b462),
	.w3(32'h3ba054d2),
	.w4(32'h3b832928),
	.w5(32'h3af4d959),
	.w6(32'h3b527766),
	.w7(32'hbafb56b7),
	.w8(32'h3a96bcd2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c132c1d),
	.w1(32'h3c633cc3),
	.w2(32'h3c3879c0),
	.w3(32'h3c27fd6c),
	.w4(32'h3c19a054),
	.w5(32'h3b5ce3e4),
	.w6(32'hbbc08ea5),
	.w7(32'hbb11736e),
	.w8(32'hb94f8f6a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99a40d),
	.w1(32'hb9954483),
	.w2(32'h38502383),
	.w3(32'hbb825c58),
	.w4(32'hba8c4a3b),
	.w5(32'h3ce52a67),
	.w6(32'h3b567e6c),
	.w7(32'hbba9fed1),
	.w8(32'h3c8c7bc2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca581b5),
	.w1(32'hbc98e337),
	.w2(32'h3c3e5942),
	.w3(32'hbc89f13c),
	.w4(32'hbd60c933),
	.w5(32'hbab0ba23),
	.w6(32'h3a1e6040),
	.w7(32'hbcc93869),
	.w8(32'hbb9b8437),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9ccfe),
	.w1(32'h3bc8b2e1),
	.w2(32'hbc1dec81),
	.w3(32'hbbcb84b1),
	.w4(32'h3cdf0ee4),
	.w5(32'h3c3d4b5d),
	.w6(32'h3c063c01),
	.w7(32'h3d0b4714),
	.w8(32'h3c8deed9),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eb9ff),
	.w1(32'hbc2b32fb),
	.w2(32'hbba01c1c),
	.w3(32'hb9d60c76),
	.w4(32'hbb06966e),
	.w5(32'hbaba81d7),
	.w6(32'h3bcfe2f6),
	.w7(32'h3b4f451b),
	.w8(32'h3bf01239),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff443),
	.w1(32'hbaa058b3),
	.w2(32'h3bd61910),
	.w3(32'h3b485c34),
	.w4(32'hba9f0657),
	.w5(32'h3bee389f),
	.w6(32'h3be28114),
	.w7(32'h39c8244e),
	.w8(32'h3abf46fb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6949a),
	.w1(32'hbba1b8a0),
	.w2(32'hbccc1557),
	.w3(32'hbbe51d43),
	.w4(32'hbb2c8605),
	.w5(32'hbca7015c),
	.w6(32'hb9ae398e),
	.w7(32'hbb833671),
	.w8(32'hbc123ddc),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc679fa2),
	.w1(32'h3be2c254),
	.w2(32'h3b340bea),
	.w3(32'hbbcdf676),
	.w4(32'h3c871411),
	.w5(32'hbba19ae4),
	.w6(32'h3b0af62b),
	.w7(32'h3ca70cb4),
	.w8(32'hbbae64a2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0f3a2),
	.w1(32'hbbcb01d3),
	.w2(32'hbc9bf6f1),
	.w3(32'hbc1120c7),
	.w4(32'hbbef586a),
	.w5(32'hbca8e2ed),
	.w6(32'hbaf48104),
	.w7(32'hbb3e27de),
	.w8(32'hbc1ac345),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f4211),
	.w1(32'hba9fab41),
	.w2(32'h3c1ae3a7),
	.w3(32'hbd067dc2),
	.w4(32'hbcc58c7c),
	.w5(32'h3bf03350),
	.w6(32'hbcd937d2),
	.w7(32'hbc987b4a),
	.w8(32'hb8e8164a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9da873),
	.w1(32'h3b70aa3b),
	.w2(32'h3be0d306),
	.w3(32'h3c192c87),
	.w4(32'hbae77238),
	.w5(32'h3b36c939),
	.w6(32'h3bda04f1),
	.w7(32'h3b63cf06),
	.w8(32'h3c096c8c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c676337),
	.w1(32'h3c20bad2),
	.w2(32'h3be232f5),
	.w3(32'h3aa532c9),
	.w4(32'h3bc84193),
	.w5(32'h3b1d8b1b),
	.w6(32'h3a6c2d41),
	.w7(32'hbb84bcba),
	.w8(32'h3c89560a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33286b),
	.w1(32'h3c8fa9ba),
	.w2(32'h3bc4b6ce),
	.w3(32'h3b79accc),
	.w4(32'h3c900cd8),
	.w5(32'h3aa92ec8),
	.w6(32'h3c835b33),
	.w7(32'h3ccb4df5),
	.w8(32'h3b1f72f1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39b234),
	.w1(32'hba874e96),
	.w2(32'hbcba5c9c),
	.w3(32'h3c3a89cd),
	.w4(32'h3c2e62c9),
	.w5(32'hbc66a641),
	.w6(32'h3c3ae874),
	.w7(32'h3be846bf),
	.w8(32'hbc303a3c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95334a),
	.w1(32'hbbf3d905),
	.w2(32'hbb2f94b5),
	.w3(32'h3bac2248),
	.w4(32'h3b6d9724),
	.w5(32'hbb62ab28),
	.w6(32'h3badf50c),
	.w7(32'h3b0e26bd),
	.w8(32'hbb9b6e86),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87f048),
	.w1(32'hbb97c397),
	.w2(32'hbd5069dc),
	.w3(32'hbc28c7a0),
	.w4(32'h3b3f103e),
	.w5(32'hbd018142),
	.w6(32'hba4e64c4),
	.w7(32'h3bb50d6f),
	.w8(32'hbc6d5f45),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdaa983),
	.w1(32'hbcbbfcfa),
	.w2(32'hbb181a17),
	.w3(32'hbc2f3492),
	.w4(32'hbbdb767a),
	.w5(32'hbbacac51),
	.w6(32'h3bc6b87f),
	.w7(32'h3b6b0aac),
	.w8(32'h39dc9342),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e2663),
	.w1(32'hbba8a05d),
	.w2(32'hbb73b14a),
	.w3(32'hbbc22709),
	.w4(32'hbbfa7ce7),
	.w5(32'h3ba4119a),
	.w6(32'h3a3d745e),
	.w7(32'hbbaf7546),
	.w8(32'hb8a94406),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75e7bb),
	.w1(32'h3b767a37),
	.w2(32'hbbd3b66f),
	.w3(32'h3cba883c),
	.w4(32'h3cce9f99),
	.w5(32'hbb9bbd95),
	.w6(32'h3ca4d7c2),
	.w7(32'h3ca66206),
	.w8(32'hbb1e2c92),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba9629),
	.w1(32'hbbf2078c),
	.w2(32'h3c1adf60),
	.w3(32'hbcc3ace7),
	.w4(32'hbcd066ec),
	.w5(32'h3bd3b597),
	.w6(32'hbcab3470),
	.w7(32'hbcc4b6e8),
	.w8(32'hbbe821ba),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6f18b),
	.w1(32'hbb8f1349),
	.w2(32'h3b569e1c),
	.w3(32'h3b620b0e),
	.w4(32'h3b38fa0d),
	.w5(32'h3bd07ded),
	.w6(32'hbbc45670),
	.w7(32'hbc13a3bc),
	.w8(32'hba82b9a2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a77bf),
	.w1(32'hba8bf5b5),
	.w2(32'hbc9b560b),
	.w3(32'h3c3086b9),
	.w4(32'h3c2a72c6),
	.w5(32'hbc5a4ca8),
	.w6(32'h3bebdfdc),
	.w7(32'h3ba1b8db),
	.w8(32'hbc8793c4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eb85d),
	.w1(32'hbb9ab486),
	.w2(32'h3c366ab8),
	.w3(32'hbc87b306),
	.w4(32'hbc23f7d1),
	.w5(32'h3c9f145f),
	.w6(32'hbced29c5),
	.w7(32'hbcd456ca),
	.w8(32'h3bbe583a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cebddcb),
	.w1(32'h3c262d86),
	.w2(32'h3c081feb),
	.w3(32'h3abe59d2),
	.w4(32'h3b704866),
	.w5(32'hbb5028c4),
	.w6(32'hbc727670),
	.w7(32'h3b8c99cb),
	.w8(32'hbbfe91df),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb4114),
	.w1(32'h3ab3783e),
	.w2(32'h3b559061),
	.w3(32'hbc68da78),
	.w4(32'h3b46843f),
	.w5(32'h3bc38b31),
	.w6(32'h358a01e0),
	.w7(32'hbbd889d5),
	.w8(32'h3b0bb24d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44ceb0),
	.w1(32'h3c745df0),
	.w2(32'h3c0cc25d),
	.w3(32'hbb198cf9),
	.w4(32'h3bc8ba66),
	.w5(32'h3a4a0538),
	.w6(32'hbbd01f9c),
	.w7(32'h3ac0e1e6),
	.w8(32'hbb7f76c9),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91c746),
	.w1(32'hba599616),
	.w2(32'hbcf6772d),
	.w3(32'hbba229dc),
	.w4(32'hbbbdaa71),
	.w5(32'hbc742cb1),
	.w6(32'hbbab9de7),
	.w7(32'hbbe2bb04),
	.w8(32'hbc8e6ba0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc056eb7),
	.w1(32'hbc7bea08),
	.w2(32'h3b8dbd5f),
	.w3(32'h3bcb030e),
	.w4(32'h3b2e9d5b),
	.w5(32'h3b8c185e),
	.w6(32'hbafe4a87),
	.w7(32'hbbc4de17),
	.w8(32'h3c3e42e9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4924e9),
	.w1(32'h3c370a38),
	.w2(32'h3b9dbcf5),
	.w3(32'h3c9ba64c),
	.w4(32'h3c682d81),
	.w5(32'hbb1d7cbc),
	.w6(32'h3c874a10),
	.w7(32'h3c905203),
	.w8(32'hbbd626be),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3e6f9),
	.w1(32'h3b69b376),
	.w2(32'h3b245dcc),
	.w3(32'hbb3803b5),
	.w4(32'h3b5cefd2),
	.w5(32'hbb681819),
	.w6(32'hbbc25344),
	.w7(32'hbb93ad67),
	.w8(32'hbc20cc37),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dab07),
	.w1(32'hbb904812),
	.w2(32'h38ce2b60),
	.w3(32'hbbc44ba9),
	.w4(32'hbb347534),
	.w5(32'h3b7b9f00),
	.w6(32'hbaaa9c09),
	.w7(32'h3bd58c86),
	.w8(32'hbae75fe3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0646a),
	.w1(32'h3c63a07c),
	.w2(32'hb957d590),
	.w3(32'h3b6ea99f),
	.w4(32'h3beb7261),
	.w5(32'hbbfad1a6),
	.w6(32'hb9800142),
	.w7(32'h3b417f99),
	.w8(32'hbc05a812),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb587c43),
	.w1(32'hb9ec27fb),
	.w2(32'hba3acd7c),
	.w3(32'hba5f098a),
	.w4(32'hbb887def),
	.w5(32'h3c0dcbeb),
	.w6(32'h3b171c89),
	.w7(32'hbaf4180b),
	.w8(32'h3b6737c8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8b866),
	.w1(32'h3ad83989),
	.w2(32'h3aafb86d),
	.w3(32'h3c671939),
	.w4(32'h3c4c1b59),
	.w5(32'h3b0370b4),
	.w6(32'h3c7e411c),
	.w7(32'h3c1323ac),
	.w8(32'h3b84f7a0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbde1b7),
	.w1(32'hbbec1995),
	.w2(32'hbbbde298),
	.w3(32'hb98c8deb),
	.w4(32'h3bb31343),
	.w5(32'h3be73659),
	.w6(32'h3bc4703e),
	.w7(32'h3b08f4b2),
	.w8(32'h3bed3063),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ef543),
	.w1(32'h3c814d4e),
	.w2(32'hbc0a4b11),
	.w3(32'h3c5fe206),
	.w4(32'h3bf8aa48),
	.w5(32'h3bdf5605),
	.w6(32'h3c7c468c),
	.w7(32'h3c60f5b0),
	.w8(32'h3c267531),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc814f74),
	.w1(32'hbcfc6290),
	.w2(32'h3c40618f),
	.w3(32'hbb31acea),
	.w4(32'hbcfcd246),
	.w5(32'h3bfb9d73),
	.w6(32'hbb885f80),
	.w7(32'hbd123ec3),
	.w8(32'h3d21b1af),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a2534),
	.w1(32'h3cba2846),
	.w2(32'hbbea9abc),
	.w3(32'h3a3fc475),
	.w4(32'h3c9f364e),
	.w5(32'hbc3f3a66),
	.w6(32'h3cdc5821),
	.w7(32'h3d1e7672),
	.w8(32'hbcbbd6a0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11e89d),
	.w1(32'h3c447386),
	.w2(32'hbba8dd53),
	.w3(32'hbbe4bbfb),
	.w4(32'hbc0ba0ac),
	.w5(32'h3c16216b),
	.w6(32'hbd132eba),
	.w7(32'hbcadd74b),
	.w8(32'hbc1204c1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca86d56),
	.w1(32'h3b604864),
	.w2(32'hbca6291d),
	.w3(32'h3ccf3ebc),
	.w4(32'h3d4f1125),
	.w5(32'h3b24d400),
	.w6(32'h3bb44247),
	.w7(32'h3c8c35b6),
	.w8(32'hbc007c58),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc367a54),
	.w1(32'h3b208bba),
	.w2(32'h3b9e7827),
	.w3(32'hbc3a05b9),
	.w4(32'hbb665537),
	.w5(32'hbaec2c0e),
	.w6(32'hbc37112c),
	.w7(32'hbb48a42e),
	.w8(32'hba12ece7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade4fcf),
	.w1(32'hbb892c68),
	.w2(32'hbac4681c),
	.w3(32'hbba7255c),
	.w4(32'hbb4afb60),
	.w5(32'h3c16549d),
	.w6(32'hbc20ace7),
	.w7(32'hbbf62c7f),
	.w8(32'hbc148191),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa096d),
	.w1(32'hbb625bca),
	.w2(32'hbb52f6eb),
	.w3(32'h3bbabd7d),
	.w4(32'h3bc5624c),
	.w5(32'h3bd00fe9),
	.w6(32'hbc1ccaea),
	.w7(32'hbc46d179),
	.w8(32'hba56519c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7b5af),
	.w1(32'h3b7c48e0),
	.w2(32'hbb916c10),
	.w3(32'h3c0ca851),
	.w4(32'h3c558617),
	.w5(32'hbc0fca64),
	.w6(32'h3ab336e4),
	.w7(32'h3b24dc19),
	.w8(32'hbbf578af),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf660a0),
	.w1(32'h3b425396),
	.w2(32'h3cc105c5),
	.w3(32'hbbbdc33d),
	.w4(32'hbb580ec6),
	.w5(32'h3c3ee051),
	.w6(32'hbbeb3541),
	.w7(32'h3ba0c162),
	.w8(32'h3c01928c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49899c),
	.w1(32'hb8c1f994),
	.w2(32'h3bc65275),
	.w3(32'hbd025115),
	.w4(32'hbccf82f1),
	.w5(32'h3b3d00b5),
	.w6(32'hbcf9b64c),
	.w7(32'hbcb9ae1d),
	.w8(32'hba994150),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa4f9),
	.w1(32'hbc479c08),
	.w2(32'hbca46fd9),
	.w3(32'h3bd8520b),
	.w4(32'hbb0077a4),
	.w5(32'hbc0aeab2),
	.w6(32'h3c284283),
	.w7(32'h3c079ee5),
	.w8(32'hb9e8abc7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76dfbd),
	.w1(32'hbbb8e5d4),
	.w2(32'hbc1690d6),
	.w3(32'hbb3e3452),
	.w4(32'hbba7c9c4),
	.w5(32'hbc3f1724),
	.w6(32'hba92e572),
	.w7(32'hbb8e4b95),
	.w8(32'hbc3d43f7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2c27c),
	.w1(32'hbaf24f81),
	.w2(32'hbc9564d0),
	.w3(32'hbc9186f7),
	.w4(32'hbc70c4a7),
	.w5(32'hbcac90a2),
	.w6(32'hbcab774e),
	.w7(32'hbc6b96ed),
	.w8(32'hbcf7cd98),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7afb3),
	.w1(32'hbc07c0be),
	.w2(32'h3b0d5790),
	.w3(32'hbc3b894f),
	.w4(32'hba3ec5fe),
	.w5(32'h3c28a2a9),
	.w6(32'hbc8f6d9c),
	.w7(32'hbb327e3b),
	.w8(32'h3c2c4e8d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5f450),
	.w1(32'hbbf312e1),
	.w2(32'hbbb8c3f3),
	.w3(32'hbb8e9fbe),
	.w4(32'hbbb415aa),
	.w5(32'h3afb9327),
	.w6(32'hbaa1a0a1),
	.w7(32'h3881f763),
	.w8(32'h3b27966b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c858b97),
	.w1(32'h3bbce9f7),
	.w2(32'hbad39610),
	.w3(32'h3c26b5cc),
	.w4(32'h3b85463b),
	.w5(32'h3ba1b6b8),
	.w6(32'h3bd6598b),
	.w7(32'h3b6ad7be),
	.w8(32'h3bd9f9bb),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b194a05),
	.w1(32'hbb4c573e),
	.w2(32'hbc273f95),
	.w3(32'h3c376496),
	.w4(32'h3bd44d04),
	.w5(32'hbbf25398),
	.w6(32'h3c35102f),
	.w7(32'h38f70fe0),
	.w8(32'hbc14185c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba032ad1),
	.w1(32'hba274164),
	.w2(32'h3c2f6e66),
	.w3(32'hbb21ae33),
	.w4(32'hbae92dd4),
	.w5(32'h3c00686a),
	.w6(32'hbbf8154b),
	.w7(32'hbbb42501),
	.w8(32'h3bad86b7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92e20e),
	.w1(32'hbb24d981),
	.w2(32'hbcd8b401),
	.w3(32'h3c06f384),
	.w4(32'h3c602841),
	.w5(32'hbc20e905),
	.w6(32'h3c88f5b5),
	.w7(32'h3ca662a5),
	.w8(32'h3be0d21c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d499d),
	.w1(32'hbbd9662a),
	.w2(32'hbc621919),
	.w3(32'h3b1ecf54),
	.w4(32'hbb8ad5a1),
	.w5(32'hbc0653d2),
	.w6(32'h3b27f794),
	.w7(32'hbac6a232),
	.w8(32'hbb9d2a66),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1ee68),
	.w1(32'hb9bf84a3),
	.w2(32'h3b299ab3),
	.w3(32'h3a1999c9),
	.w4(32'h3bd018fd),
	.w5(32'h3c6c31ad),
	.w6(32'h3b6f3958),
	.w7(32'hbb06645b),
	.w8(32'h3c74d0b2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4575d),
	.w1(32'h3bbce9cc),
	.w2(32'hbba4e7cf),
	.w3(32'h3cb5a725),
	.w4(32'h3c438c96),
	.w5(32'hbb4917c5),
	.w6(32'h3c6cf371),
	.w7(32'h3c8896ce),
	.w8(32'hbb29fcac),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf14ac),
	.w1(32'h3c00c677),
	.w2(32'hba0d5e1f),
	.w3(32'hbcd4297e),
	.w4(32'hbbdfcc8f),
	.w5(32'hbbba4489),
	.w6(32'hbcb6e944),
	.w7(32'hbc003a69),
	.w8(32'hbb462afd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4cdd),
	.w1(32'hba4f19ca),
	.w2(32'h3c9a4cfc),
	.w3(32'h3a4a2e31),
	.w4(32'hbb28b324),
	.w5(32'h3b8be875),
	.w6(32'hbbd6d4ff),
	.w7(32'hbc186333),
	.w8(32'hbbe49544),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a4297),
	.w1(32'hbadd9221),
	.w2(32'h3c0532bd),
	.w3(32'hbd25c7d9),
	.w4(32'hbd11cd1b),
	.w5(32'h3ac9871c),
	.w6(32'hbd2a3577),
	.w7(32'hbd0a3f2f),
	.w8(32'h3b3944f8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5b023),
	.w1(32'hbaf59ed9),
	.w2(32'h3ad41f2f),
	.w3(32'hbbdf5344),
	.w4(32'hbc1593ed),
	.w5(32'hb9bd67d5),
	.w6(32'hbb7b2af0),
	.w7(32'hbbfbdfc4),
	.w8(32'hbb3e2895),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72be74),
	.w1(32'hba9da664),
	.w2(32'h3a27438a),
	.w3(32'hbbf30114),
	.w4(32'h3bcee75b),
	.w5(32'h3c43b5b3),
	.w6(32'hb9d97ea1),
	.w7(32'hbb5d7058),
	.w8(32'hbbfbb934),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e853e),
	.w1(32'h3b9f8b2a),
	.w2(32'h3c122813),
	.w3(32'h3bf47e6f),
	.w4(32'h3baa793e),
	.w5(32'h3c0ac31d),
	.w6(32'hb82de8b7),
	.w7(32'h3b8b2a1f),
	.w8(32'hbc42e7c6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15dbec),
	.w1(32'hbc59791c),
	.w2(32'hbc567c37),
	.w3(32'hbb6c2286),
	.w4(32'hbc2f1436),
	.w5(32'hbbc48b02),
	.w6(32'hbbb4bfbd),
	.w7(32'hbc4b57ce),
	.w8(32'hbb68231d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8fa4d),
	.w1(32'hbaa1e30d),
	.w2(32'h3bcd0df7),
	.w3(32'hb7efea00),
	.w4(32'hbaf0e47d),
	.w5(32'h3bcab54e),
	.w6(32'hbc156eb7),
	.w7(32'hbabe1f9a),
	.w8(32'hbb27160a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6059d2),
	.w1(32'hbc9b0d05),
	.w2(32'hba9f055f),
	.w3(32'hbcd6bc95),
	.w4(32'hbcd7d583),
	.w5(32'h3b9156cf),
	.w6(32'hbcb7bcf8),
	.w7(32'hbcba5996),
	.w8(32'hbbac13f5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dc15e),
	.w1(32'h3b435f89),
	.w2(32'hbaf41f03),
	.w3(32'h3c0cb8c5),
	.w4(32'h3b1e72c5),
	.w5(32'h3be5f778),
	.w6(32'h3b9ff1b0),
	.w7(32'h3b1f24a9),
	.w8(32'hb8f73bd7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3958db7e),
	.w1(32'h3b890dd7),
	.w2(32'h3c90b6e8),
	.w3(32'h3ccb7e88),
	.w4(32'hbb01d333),
	.w5(32'h3cbe2f7b),
	.w6(32'h3cbc9b24),
	.w7(32'h3c307673),
	.w8(32'hbb9ef607),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c946af2),
	.w1(32'h3cb97235),
	.w2(32'h3cc1e0f5),
	.w3(32'hba85c4b5),
	.w4(32'h3c09c60d),
	.w5(32'h3d3af6d2),
	.w6(32'hbcde1ca8),
	.w7(32'hbc497fca),
	.w8(32'h3d09769a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cee6fea),
	.w1(32'h3d2b92d7),
	.w2(32'hbc00c3db),
	.w3(32'h3d6e6c4e),
	.w4(32'h3d45657a),
	.w5(32'hbc830cb8),
	.w6(32'h3d5b2de8),
	.w7(32'h3d3de9c1),
	.w8(32'hbcb5ed53),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cc8cc),
	.w1(32'hbd05f21a),
	.w2(32'hbcd6646b),
	.w3(32'hbc883af3),
	.w4(32'hbcd414d4),
	.w5(32'hbccb6991),
	.w6(32'hbc15b712),
	.w7(32'hbca1734d),
	.w8(32'hbcc840f6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bccb7),
	.w1(32'hbcd545df),
	.w2(32'hbca9c062),
	.w3(32'hbd00b1da),
	.w4(32'hbcd8cf30),
	.w5(32'hbc49a948),
	.w6(32'hbd07d153),
	.w7(32'hbce2c75c),
	.w8(32'h39f029d1),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf51815),
	.w1(32'hbb189097),
	.w2(32'hba31d4b2),
	.w3(32'hbb7b5de1),
	.w4(32'hbb4cb026),
	.w5(32'hbb9d0e15),
	.w6(32'hbbf6418f),
	.w7(32'h3aca60cd),
	.w8(32'h3be87ba7),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b181df5),
	.w1(32'h3ad92522),
	.w2(32'h3c181cae),
	.w3(32'hbc0d9609),
	.w4(32'hbbb90dbf),
	.w5(32'h3c480a29),
	.w6(32'h3c676be3),
	.w7(32'h3c01f0fd),
	.w8(32'h3c7bb1ae),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f5f98),
	.w1(32'h3ca41634),
	.w2(32'hbaa09391),
	.w3(32'h3c92167e),
	.w4(32'h3cd58629),
	.w5(32'h3b831137),
	.w6(32'h3cc102e9),
	.w7(32'h3cfb2a0e),
	.w8(32'hbbf89e49),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc36ea7),
	.w1(32'h3b6398be),
	.w2(32'h39be6308),
	.w3(32'hb9909c5f),
	.w4(32'h3b42fe8f),
	.w5(32'hbb122c01),
	.w6(32'h3a187fd5),
	.w7(32'h3b79d150),
	.w8(32'hbb6d16bb),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8612b),
	.w1(32'h3c45d7ca),
	.w2(32'hbc13dff0),
	.w3(32'h3c1138c2),
	.w4(32'h3bf92712),
	.w5(32'hbadcef35),
	.w6(32'hbaa3eae1),
	.w7(32'h3a2a84ee),
	.w8(32'h3bccd185),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35942f),
	.w1(32'hbcf8efa3),
	.w2(32'hbc13cf3d),
	.w3(32'hbb883203),
	.w4(32'hbd0cfac5),
	.w5(32'h3a1dc7c2),
	.w6(32'h3acf2a6a),
	.w7(32'hbc4ffc6e),
	.w8(32'hbc29aa94),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b7d30),
	.w1(32'hbbd57025),
	.w2(32'hbbcd461b),
	.w3(32'hbbcd4e71),
	.w4(32'hbbf171f5),
	.w5(32'hbc213074),
	.w6(32'hbbb763eb),
	.w7(32'hbbd5d965),
	.w8(32'hbbb38ca4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ad58b),
	.w1(32'hbaeebc71),
	.w2(32'h3af13d62),
	.w3(32'h39d11931),
	.w4(32'hbc160e61),
	.w5(32'h3b3ae2bb),
	.w6(32'hb92f66ed),
	.w7(32'hbc090854),
	.w8(32'h3b9ba50e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07be23),
	.w1(32'h3c9482fa),
	.w2(32'h3c8fe034),
	.w3(32'hbc0e5fc3),
	.w4(32'hbc8990f9),
	.w5(32'h3adcc28b),
	.w6(32'hbb95c467),
	.w7(32'hbc886f14),
	.w8(32'hbb9c4661),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2cc23),
	.w1(32'h3b899c94),
	.w2(32'h3bf52b1a),
	.w3(32'h3a320cb8),
	.w4(32'hbbc44c3d),
	.w5(32'h3bc5338b),
	.w6(32'hbc8d3f77),
	.w7(32'hbc53e5d7),
	.w8(32'h3b866d6c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd35388),
	.w1(32'h3b634ae5),
	.w2(32'h3aa1cb6d),
	.w3(32'h3b54e37c),
	.w4(32'hbb8b9f05),
	.w5(32'h3b900f8a),
	.w6(32'hbbe96b2d),
	.w7(32'hbbba457a),
	.w8(32'h3bcb2b8d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25fb34),
	.w1(32'h3c4566d6),
	.w2(32'h3b8e14a0),
	.w3(32'hbc351a00),
	.w4(32'hbba32733),
	.w5(32'hbb10d57f),
	.w6(32'hbc45570a),
	.w7(32'hbbb9eca5),
	.w8(32'hbc1c35dc),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47e48c),
	.w1(32'hbb47c4f9),
	.w2(32'hbb907a92),
	.w3(32'hbc8fa7aa),
	.w4(32'hbc060107),
	.w5(32'hbc150bf0),
	.w6(32'hbca01c8d),
	.w7(32'hbbcdbb16),
	.w8(32'hbba6b399),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d6956),
	.w1(32'hbc59dc52),
	.w2(32'h394bccd4),
	.w3(32'hbc974fdc),
	.w4(32'hbca24bd0),
	.w5(32'h3b9c5454),
	.w6(32'hbc5aa41f),
	.w7(32'hbc16d7a7),
	.w8(32'h3ba5ed70),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8373fa),
	.w1(32'h3bf5063d),
	.w2(32'h3b55e141),
	.w3(32'hbba69166),
	.w4(32'hb9225083),
	.w5(32'hbb9b8029),
	.w6(32'h3af662c1),
	.w7(32'h3b439993),
	.w8(32'h3b4178d8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b12d3),
	.w1(32'h39c4660d),
	.w2(32'hbaabee71),
	.w3(32'hbbdba6c3),
	.w4(32'hbb4db0e3),
	.w5(32'h3bc59af8),
	.w6(32'hbb08be58),
	.w7(32'hba8e4540),
	.w8(32'hbac54783),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a963f43),
	.w1(32'hb851efc8),
	.w2(32'hbc7e935c),
	.w3(32'h3b56d0aa),
	.w4(32'hb8638eea),
	.w5(32'hbc02094c),
	.w6(32'h3af43643),
	.w7(32'h3b812f6e),
	.w8(32'hbbb6d46f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc23736),
	.w1(32'h3c8261d2),
	.w2(32'h3c9af3fc),
	.w3(32'h3c060c83),
	.w4(32'h3bd34741),
	.w5(32'h3c9e481c),
	.w6(32'hbc0aaa1e),
	.w7(32'h3a60b6d3),
	.w8(32'h3ba0557f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c102f95),
	.w1(32'h3c2df8e5),
	.w2(32'h3c3199dc),
	.w3(32'hbc143f76),
	.w4(32'h3bd8e6d1),
	.w5(32'h3c46d284),
	.w6(32'hbc2875a6),
	.w7(32'hbaae4b47),
	.w8(32'hbc27fe2c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc3449),
	.w1(32'h3cbe33f2),
	.w2(32'h3cd83272),
	.w3(32'h3c40f52d),
	.w4(32'h3c512018),
	.w5(32'h3cd3a68c),
	.w6(32'hbc2edd67),
	.w7(32'hbbd70ad8),
	.w8(32'h3b87b279),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c176e34),
	.w1(32'h3c23f06b),
	.w2(32'hbc6981e7),
	.w3(32'h3c9f1de5),
	.w4(32'h3c86ea52),
	.w5(32'hbc5f3afd),
	.w6(32'h3c3874f5),
	.w7(32'hbaa55acf),
	.w8(32'hbac62a4b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc824e1d),
	.w1(32'hbc5b201a),
	.w2(32'hbd1ceb7c),
	.w3(32'hbc486f0c),
	.w4(32'hbc04ce60),
	.w5(32'hbce10dfd),
	.w6(32'h3b3b3e2a),
	.w7(32'h3bb2c6a4),
	.w8(32'hbc6ce1d1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd07efa6),
	.w1(32'hbce11f9c),
	.w2(32'hbb18409b),
	.w3(32'hbcb4aa14),
	.w4(32'hbc8bd1c1),
	.w5(32'h38860c4e),
	.w6(32'hbbf5ab30),
	.w7(32'hbbfa27e3),
	.w8(32'hba9d3d23),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cea69),
	.w1(32'hbb16e971),
	.w2(32'hbb70ad53),
	.w3(32'h37c3d355),
	.w4(32'hba8aaaa4),
	.w5(32'h3993dba4),
	.w6(32'hbafb20f3),
	.w7(32'hbb77a833),
	.w8(32'hbb43b188),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e6465),
	.w1(32'h3b98008d),
	.w2(32'hbb3ef657),
	.w3(32'hbc0d6770),
	.w4(32'hbb29622b),
	.w5(32'hbc14f2c8),
	.w6(32'hbc12a412),
	.w7(32'h3a1c6147),
	.w8(32'hbbdc8a74),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75c095),
	.w1(32'hba89058e),
	.w2(32'hbaa93892),
	.w3(32'hbba13369),
	.w4(32'hbbdceb00),
	.w5(32'h3a6c3a0e),
	.w6(32'h3aaf2abd),
	.w7(32'h368b881b),
	.w8(32'hb9fd8e25),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21a0e4),
	.w1(32'hba73eb88),
	.w2(32'hbc7905a8),
	.w3(32'hbb478f80),
	.w4(32'h3b1a9178),
	.w5(32'hbc88085c),
	.w6(32'hbaa03d16),
	.w7(32'h3a600058),
	.w8(32'hbc35ad24),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29a816),
	.w1(32'hbc227f44),
	.w2(32'hbc76f5d8),
	.w3(32'hbbdd7b3a),
	.w4(32'hbc0f991c),
	.w5(32'hbcb9b42e),
	.w6(32'hbba3dd07),
	.w7(32'hbbcf33ac),
	.w8(32'hbc93e8e2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa3f3b),
	.w1(32'hbc76d3db),
	.w2(32'h3bb692e0),
	.w3(32'hbce378cf),
	.w4(32'hbcbac1bc),
	.w5(32'h3c1f0b41),
	.w6(32'hbcc0e21a),
	.w7(32'hbc97d1cd),
	.w8(32'h3b932c8c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bd6b0),
	.w1(32'h3b2c41ad),
	.w2(32'hbb18f946),
	.w3(32'h3c606067),
	.w4(32'hbc2fee63),
	.w5(32'hbb612ac8),
	.w6(32'h3b824014),
	.w7(32'hbc1119d2),
	.w8(32'hb9e50df3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb294ec5),
	.w1(32'hbb49b950),
	.w2(32'h3ad43196),
	.w3(32'hbb7c8340),
	.w4(32'h3aab6beb),
	.w5(32'hbbea3cba),
	.w6(32'hb92cc9df),
	.w7(32'h3b31afc1),
	.w8(32'hbb9bcd09),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d424ae7),
	.w1(32'h3c9ec9f2),
	.w2(32'hbb77f416),
	.w3(32'h3b14d20c),
	.w4(32'h3cb39ca3),
	.w5(32'hbba776ba),
	.w6(32'hbc9c952a),
	.w7(32'h3c33a839),
	.w8(32'hbcb352b7),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e42fcd),
	.w1(32'h3c0047a0),
	.w2(32'h3b1259d3),
	.w3(32'hba1125bf),
	.w4(32'h3be8bd7b),
	.w5(32'h3b57d3e3),
	.w6(32'hbc56f96b),
	.w7(32'h3b5e74af),
	.w8(32'hbb9b98ef),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc436959),
	.w1(32'hbc717e44),
	.w2(32'hbc9481d3),
	.w3(32'hba915464),
	.w4(32'hbc822fd2),
	.w5(32'hbc2f38db),
	.w6(32'h3c0122c7),
	.w7(32'hba0765dc),
	.w8(32'hbc222195),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule