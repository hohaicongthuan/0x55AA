module layer_8_featuremap_91(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd99601),
	.w1(32'hbb002890),
	.w2(32'h3c3aed79),
	.w3(32'hbc08841e),
	.w4(32'hbabb8982),
	.w5(32'h3bebd2da),
	.w6(32'hbb197295),
	.w7(32'h3c5eb1c3),
	.w8(32'h3c842814),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeb167),
	.w1(32'h3c033302),
	.w2(32'hbd244403),
	.w3(32'hbba82023),
	.w4(32'h3ba64e79),
	.w5(32'h3cd8b860),
	.w6(32'h3c39d425),
	.w7(32'hbc85a5fc),
	.w8(32'hbbb38c4a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da480),
	.w1(32'hbc6e6e88),
	.w2(32'hbc19d319),
	.w3(32'h3b9272eb),
	.w4(32'h3c106c69),
	.w5(32'hbc37b2f1),
	.w6(32'hbc76bce1),
	.w7(32'h3be1326c),
	.w8(32'hb79e4705),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd901ab),
	.w1(32'hbc4f011f),
	.w2(32'hbbbb0438),
	.w3(32'hbc07c8ec),
	.w4(32'hbc40f427),
	.w5(32'hbc33fb35),
	.w6(32'h3c0e870e),
	.w7(32'h3af1d3a2),
	.w8(32'h3c556d0f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1f1e5),
	.w1(32'hbc35856b),
	.w2(32'hbc207f30),
	.w3(32'h3c13f025),
	.w4(32'hbc3d8490),
	.w5(32'h3b51a116),
	.w6(32'hbc022748),
	.w7(32'h3c589011),
	.w8(32'hbc19f841),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f76cd),
	.w1(32'h3b2aec5b),
	.w2(32'hbcda305c),
	.w3(32'h3c1f5f41),
	.w4(32'h3bcec82d),
	.w5(32'hbd1e2a6c),
	.w6(32'h3c1fa0cb),
	.w7(32'hbc29ee23),
	.w8(32'hbc8d33e0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94a128),
	.w1(32'hbb82f539),
	.w2(32'h3c0d604c),
	.w3(32'hbcae93b4),
	.w4(32'h3af8f93c),
	.w5(32'h3a030ff8),
	.w6(32'h3d01b163),
	.w7(32'h3c4afb09),
	.w8(32'hbb130bfc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b5174),
	.w1(32'hbc834ff9),
	.w2(32'h3be72da8),
	.w3(32'h3d02be15),
	.w4(32'h3c0262b7),
	.w5(32'hba8f6568),
	.w6(32'h3c18c271),
	.w7(32'hbb8b00fe),
	.w8(32'h3c1cd35a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf119fd),
	.w1(32'hbc630ff8),
	.w2(32'h3b768930),
	.w3(32'hbcaf19e7),
	.w4(32'h3be17dc0),
	.w5(32'hbaeae366),
	.w6(32'h3cd01e05),
	.w7(32'h3bf821e1),
	.w8(32'h3b531adf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4a7f8),
	.w1(32'hbb95a609),
	.w2(32'h3ca38d4a),
	.w3(32'hbcc97db9),
	.w4(32'h3c843ac7),
	.w5(32'h3cd4817d),
	.w6(32'hbcf7c74a),
	.w7(32'h3cdf0203),
	.w8(32'h3ba613dd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e7db9),
	.w1(32'h3c7a8c59),
	.w2(32'h3c242dbc),
	.w3(32'hbc292dc9),
	.w4(32'hbc06028b),
	.w5(32'hbb984119),
	.w6(32'h3caa6c78),
	.w7(32'h3c17d892),
	.w8(32'h3be6b7b4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909aec),
	.w1(32'hbc8f14e2),
	.w2(32'h3bfacbce),
	.w3(32'h3cf4b1f7),
	.w4(32'h3c0406d5),
	.w5(32'h3c63e931),
	.w6(32'hbbd59487),
	.w7(32'hbbb5548e),
	.w8(32'hbb3f42a9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd090fe),
	.w1(32'hbb91fdd5),
	.w2(32'hbba2d881),
	.w3(32'hbc3f05bb),
	.w4(32'h3b051716),
	.w5(32'hbc677c53),
	.w6(32'hba8382e5),
	.w7(32'h3b6dfefe),
	.w8(32'hbca8115b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d66c0),
	.w1(32'hba1d8496),
	.w2(32'hbcd4f509),
	.w3(32'h3ba59ced),
	.w4(32'h3c83fc63),
	.w5(32'hbd359f54),
	.w6(32'h3cd7dfcc),
	.w7(32'hbb435691),
	.w8(32'h3d2ba02b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a6baf),
	.w1(32'hbc881865),
	.w2(32'hbda03099),
	.w3(32'hb7afc99b),
	.w4(32'h3c18042e),
	.w5(32'hbbe6dd96),
	.w6(32'h3bee4fe1),
	.w7(32'hbc49410c),
	.w8(32'hbd1c8810),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe19fd0),
	.w1(32'hbc10b273),
	.w2(32'h3d6f8a2c),
	.w3(32'hbc5f7095),
	.w4(32'hbd3db117),
	.w5(32'hbcda8991),
	.w6(32'hbcc3268a),
	.w7(32'hbc15ce31),
	.w8(32'hbc591c95),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b477931),
	.w1(32'h3cf1957d),
	.w2(32'hbce80e1e),
	.w3(32'hbbd2db09),
	.w4(32'hbc2236d0),
	.w5(32'hbba96183),
	.w6(32'hbd5cb73d),
	.w7(32'hbc1c9465),
	.w8(32'hbb794f58),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88316f),
	.w1(32'h3cac8b42),
	.w2(32'hbc59cd23),
	.w3(32'hbccfd707),
	.w4(32'h3d01e32f),
	.w5(32'h3c9cfac2),
	.w6(32'h3ca70c4f),
	.w7(32'h3aa03cb3),
	.w8(32'h399e74f5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd897b2a),
	.w1(32'hbd904f37),
	.w2(32'hbd2b8f04),
	.w3(32'h3d2006e9),
	.w4(32'h3c27d4d1),
	.w5(32'h3d90d9a7),
	.w6(32'hbb2901d8),
	.w7(32'h3d8e411a),
	.w8(32'h3de03d50),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabcf48),
	.w1(32'hbc6ab57d),
	.w2(32'h3b8bd727),
	.w3(32'h3c81bfdb),
	.w4(32'h3c25e4a5),
	.w5(32'h3c6f55fc),
	.w6(32'hbbf0b876),
	.w7(32'h3d37d0cb),
	.w8(32'h3be1df27),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c2245),
	.w1(32'hbbb7a239),
	.w2(32'hbc3a52f6),
	.w3(32'hbc030ab0),
	.w4(32'hbcb78231),
	.w5(32'hbc1afbf0),
	.w6(32'h3c174c17),
	.w7(32'hbb26176e),
	.w8(32'hbb2e3771),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8300a),
	.w1(32'h3ba6686d),
	.w2(32'h3ca210db),
	.w3(32'h3cacecc5),
	.w4(32'hbb0065d4),
	.w5(32'hbc6c472c),
	.w6(32'hbc5f3930),
	.w7(32'hbd23b9c5),
	.w8(32'hbb168dcf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce4ef58),
	.w1(32'hbcbbfae2),
	.w2(32'h3c205e21),
	.w3(32'hbd365617),
	.w4(32'h3c28d865),
	.w5(32'h3d97933c),
	.w6(32'hbd03ab66),
	.w7(32'h3cfb9b7c),
	.w8(32'h3d4f8571),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8ef7e),
	.w1(32'hbd4b47bd),
	.w2(32'h3c3eb3e7),
	.w3(32'hbbaa7259),
	.w4(32'h3c56b0f7),
	.w5(32'h3b676adf),
	.w6(32'hbc677c03),
	.w7(32'h3d0e4191),
	.w8(32'hbd458edd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c012c11),
	.w1(32'hbad08756),
	.w2(32'h3c42e71e),
	.w3(32'hbc28ff71),
	.w4(32'hbcba93f4),
	.w5(32'hbac05901),
	.w6(32'h3c260c08),
	.w7(32'h3c849ade),
	.w8(32'h3ba2877f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3445fa),
	.w1(32'hbccff380),
	.w2(32'h3a7acc6e),
	.w3(32'hba406b2d),
	.w4(32'hbbad6912),
	.w5(32'h3d1e9ee9),
	.w6(32'hbc524aa4),
	.w7(32'h3c0355e4),
	.w8(32'h3b0bb534),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c952bfe),
	.w1(32'hbc0fd470),
	.w2(32'h3bda7d30),
	.w3(32'h3c055248),
	.w4(32'h3d4e46cb),
	.w5(32'hbc0ec5a2),
	.w6(32'h3c141b6e),
	.w7(32'h3b1d7327),
	.w8(32'hbd057e94),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19087c),
	.w1(32'h3d01757c),
	.w2(32'hbd97a507),
	.w3(32'h3d1e89dc),
	.w4(32'hbb548834),
	.w5(32'hbd315210),
	.w6(32'hbd9280ce),
	.w7(32'h3c895ea3),
	.w8(32'h3e04cc11),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19fcc9),
	.w1(32'h3bcc31c0),
	.w2(32'h3c1dbbb8),
	.w3(32'hbbfe9c00),
	.w4(32'hba5dc3a6),
	.w5(32'h3c94e6d6),
	.w6(32'hbd24e01b),
	.w7(32'hbc0d99e5),
	.w8(32'h3caf1033),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d7a86),
	.w1(32'hbc3ea305),
	.w2(32'hbc9b70b7),
	.w3(32'h3abd5cf6),
	.w4(32'h3c1625cf),
	.w5(32'hbb43f6be),
	.w6(32'h3c45d750),
	.w7(32'h3c9812ee),
	.w8(32'hbc811689),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f32c11),
	.w1(32'hbb2b67f8),
	.w2(32'h3d6ee728),
	.w3(32'h3d178450),
	.w4(32'h3aeb9437),
	.w5(32'hbc39b7a6),
	.w6(32'h3c311aab),
	.w7(32'hbc37a032),
	.w8(32'h3b6e35ba),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf516d),
	.w1(32'hbc1e3369),
	.w2(32'h3b17dc04),
	.w3(32'hbb1021f7),
	.w4(32'hbc116683),
	.w5(32'hbd2cd96b),
	.w6(32'hbc9dba5c),
	.w7(32'hbc49181e),
	.w8(32'hbc1dd31e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ef25e),
	.w1(32'hbb88147c),
	.w2(32'h3b83dcbb),
	.w3(32'hbbf7cf9b),
	.w4(32'h3c10e38f),
	.w5(32'h3c06007c),
	.w6(32'hbb8d9929),
	.w7(32'h3b811b7a),
	.w8(32'h3ccd1f78),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1480a),
	.w1(32'hbc0a06e9),
	.w2(32'h3c3393fa),
	.w3(32'h39b7c6b2),
	.w4(32'h3c403ccd),
	.w5(32'h3cdc1aaa),
	.w6(32'h3b841ed8),
	.w7(32'hbcb4382c),
	.w8(32'hbc3a8231),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68d37b),
	.w1(32'h3cc10380),
	.w2(32'h3ba53307),
	.w3(32'hbb803dd8),
	.w4(32'h3c917fda),
	.w5(32'h3bb0a075),
	.w6(32'h3b11ee92),
	.w7(32'h3ab7c29e),
	.w8(32'hbc1d349a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e98dc),
	.w1(32'hbc91ed6c),
	.w2(32'hbcfda59c),
	.w3(32'hbbc6f298),
	.w4(32'h3b80d1e6),
	.w5(32'h3b2eb12b),
	.w6(32'hbc0960b1),
	.w7(32'hba5b69a0),
	.w8(32'h3b2ccc85),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21ee2a),
	.w1(32'hbc886771),
	.w2(32'hbb80ceda),
	.w3(32'h3cb292e4),
	.w4(32'hbb9999e6),
	.w5(32'h3c5736f9),
	.w6(32'h3cca6491),
	.w7(32'h3bde53ba),
	.w8(32'hbc732929),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43e693),
	.w1(32'hbaf9d2a7),
	.w2(32'h3c1b1875),
	.w3(32'hbc2d86e7),
	.w4(32'hbb5b6d0e),
	.w5(32'h3bb82e3d),
	.w6(32'hbabaab4b),
	.w7(32'h3c872682),
	.w8(32'hbca09ab3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6abe85),
	.w1(32'h3d225d16),
	.w2(32'h3c34057d),
	.w3(32'hbbd2fdca),
	.w4(32'hbb8aa782),
	.w5(32'h3c49564c),
	.w6(32'hbac3f346),
	.w7(32'h3c2731bc),
	.w8(32'h3a1a6a46),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1ba3f),
	.w1(32'hbbd299da),
	.w2(32'h3b7f8688),
	.w3(32'h3a0d9fa8),
	.w4(32'h3d085dfc),
	.w5(32'hbc090233),
	.w6(32'h3b68770f),
	.w7(32'h3b5e1c58),
	.w8(32'hbc11ff84),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2622f2),
	.w1(32'hba85575e),
	.w2(32'h3d087457),
	.w3(32'hbd03aff3),
	.w4(32'h3c457ed2),
	.w5(32'h3b0bce1c),
	.w6(32'hbbc5ff32),
	.w7(32'h3c93805a),
	.w8(32'hbb323d6e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced3dbe),
	.w1(32'h3c2e1a3a),
	.w2(32'hba97aa85),
	.w3(32'h3c161b4a),
	.w4(32'h3b8229c1),
	.w5(32'hbbe140ba),
	.w6(32'h3bf5aa66),
	.w7(32'h3ad82c96),
	.w8(32'hbbc65933),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba53320),
	.w1(32'hbb96c57a),
	.w2(32'hbb2ff633),
	.w3(32'h3cb84283),
	.w4(32'hbb10ff8d),
	.w5(32'hbc9d106a),
	.w6(32'h3a256b3e),
	.w7(32'h3cf1db21),
	.w8(32'hbc711c11),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0e9f5f),
	.w1(32'hbc9516ea),
	.w2(32'hbcfb97ab),
	.w3(32'hbb4fafcc),
	.w4(32'hbcecdca1),
	.w5(32'h3c47c3cb),
	.w6(32'hba1a5a3a),
	.w7(32'hbc97a155),
	.w8(32'hbc7e90ee),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a8ff7),
	.w1(32'hbd07c50a),
	.w2(32'hbc25a2a3),
	.w3(32'hbb9edca4),
	.w4(32'h389086c1),
	.w5(32'h3c85fddb),
	.w6(32'hbc4b06b7),
	.w7(32'h3c7989c7),
	.w8(32'h3c88df0b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0382b5),
	.w1(32'hbd022c3e),
	.w2(32'hbc30f357),
	.w3(32'h3b7d0178),
	.w4(32'hbb569556),
	.w5(32'h3be1e7a5),
	.w6(32'h3bc834b5),
	.w7(32'h3c621a32),
	.w8(32'hbcc6533e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d729056),
	.w1(32'hbcc7c3b4),
	.w2(32'hbb2a1d65),
	.w3(32'h3b922980),
	.w4(32'hbcba8971),
	.w5(32'hbca98a5c),
	.w6(32'hbd14656f),
	.w7(32'hbca1ac38),
	.w8(32'hbb211132),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57d640),
	.w1(32'hbce9f94d),
	.w2(32'hbcb29dae),
	.w3(32'hbc567275),
	.w4(32'hbbbf6cca),
	.w5(32'h3cc9736c),
	.w6(32'hbcc4c0e9),
	.w7(32'h3cb963b8),
	.w8(32'h3cc81239),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53918c),
	.w1(32'hbc5d150d),
	.w2(32'hbc008781),
	.w3(32'h3b9a3047),
	.w4(32'hb9e06a9f),
	.w5(32'h3b43067e),
	.w6(32'h3bcd970f),
	.w7(32'hbc243c1b),
	.w8(32'hbd080bc4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9040ea),
	.w1(32'hbc49c91e),
	.w2(32'hbc7898e3),
	.w3(32'h3c360b0d),
	.w4(32'hbc88c31e),
	.w5(32'h3c4a4b3d),
	.w6(32'h3cd38ad5),
	.w7(32'hbbb7249c),
	.w8(32'hbaaccf5b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdbaf7d),
	.w1(32'hbb14ca1f),
	.w2(32'hbbfcdcaf),
	.w3(32'hbba6a420),
	.w4(32'h3cf444be),
	.w5(32'hbc324c18),
	.w6(32'hbc52feb0),
	.w7(32'hbcadecc9),
	.w8(32'hbc4c201a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb03905),
	.w1(32'hbcbf1f93),
	.w2(32'hbbd8a91d),
	.w3(32'h3b8f1b12),
	.w4(32'hbd039083),
	.w5(32'hbd28fbb1),
	.w6(32'h3ca984e2),
	.w7(32'h3c442c32),
	.w8(32'hbc157d13),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd134e23),
	.w1(32'h3d501e62),
	.w2(32'hb91b836e),
	.w3(32'h3cdbdca9),
	.w4(32'h3bfc54bd),
	.w5(32'h3b2d24eb),
	.w6(32'h3c51d98e),
	.w7(32'h3c8c22dd),
	.w8(32'h3cf21d90),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20ec7f),
	.w1(32'hbaa59a23),
	.w2(32'h3cb343b9),
	.w3(32'hbd0ae633),
	.w4(32'hbadd935f),
	.w5(32'h3c2a06cb),
	.w6(32'hbc8e070d),
	.w7(32'h3cab604b),
	.w8(32'h3bc11187),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ef96e),
	.w1(32'h3c134d0a),
	.w2(32'hbaef1591),
	.w3(32'h3c3d54be),
	.w4(32'hbc14f498),
	.w5(32'h3c38b6fd),
	.w6(32'h3bc56d9e),
	.w7(32'hbc134cfc),
	.w8(32'h3d0ac217),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd84ad85),
	.w1(32'hbd511791),
	.w2(32'hbc4b3603),
	.w3(32'hbc8a1ce9),
	.w4(32'h3c2bddd6),
	.w5(32'h3c14477e),
	.w6(32'hbd87486b),
	.w7(32'hbd6f42da),
	.w8(32'h3b9e05c9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc7ac6),
	.w1(32'h3cbbb56e),
	.w2(32'h3d52791d),
	.w3(32'hbcca5905),
	.w4(32'h3b3877cd),
	.w5(32'hbd4f6d3e),
	.w6(32'hba0e5c52),
	.w7(32'hbbf2bab1),
	.w8(32'h3ba86db7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50c374),
	.w1(32'h3bc1ec27),
	.w2(32'hbc49eb7f),
	.w3(32'hbca00d03),
	.w4(32'h3b0c7b42),
	.w5(32'hbbecf0a2),
	.w6(32'h3bf2d631),
	.w7(32'hbc59d8d7),
	.w8(32'h3c18eac7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0ce41e),
	.w1(32'hbc1564a0),
	.w2(32'hbcc25424),
	.w3(32'hbd299891),
	.w4(32'hbc68d250),
	.w5(32'hbcfac0c6),
	.w6(32'hbbb30575),
	.w7(32'hbc6e4349),
	.w8(32'h3d0091f7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8da939),
	.w1(32'h39058516),
	.w2(32'hbb826697),
	.w3(32'hbca288a1),
	.w4(32'h3b912038),
	.w5(32'hbc19beec),
	.w6(32'hbd83d36f),
	.w7(32'h3cc4bc63),
	.w8(32'h3d03fb4e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf26f3),
	.w1(32'hbb0ab927),
	.w2(32'hbd202f36),
	.w3(32'h3c87d6e3),
	.w4(32'hbcab5c70),
	.w5(32'h3c800fe5),
	.w6(32'hbd0e9e76),
	.w7(32'hbd152563),
	.w8(32'hbc5d5385),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb3336),
	.w1(32'hbb1cb191),
	.w2(32'h3c113315),
	.w3(32'hbc179f49),
	.w4(32'h394fd9f9),
	.w5(32'h3c563d49),
	.w6(32'h3bcb187d),
	.w7(32'h3bcb32fc),
	.w8(32'hbaadeab7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba85acb),
	.w1(32'hbcbfc6c0),
	.w2(32'hbce34336),
	.w3(32'hbd1ce39b),
	.w4(32'h3c007c7b),
	.w5(32'hbc33b69c),
	.w6(32'hbce10a17),
	.w7(32'h3c921703),
	.w8(32'hbb520fbb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2eab56),
	.w1(32'hbd464422),
	.w2(32'h3cc94139),
	.w3(32'hbc33d4b1),
	.w4(32'h3adc7da4),
	.w5(32'h3c8a3dc4),
	.w6(32'hbd7ee701),
	.w7(32'h3b29079b),
	.w8(32'h3cae812a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdf24dd),
	.w1(32'hbd140f2f),
	.w2(32'hbd19009b),
	.w3(32'h3c893f5e),
	.w4(32'hbbe5caaf),
	.w5(32'hba716f3d),
	.w6(32'hbd42160f),
	.w7(32'h3be25d1a),
	.w8(32'hbc051316),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81cbe9),
	.w1(32'hbd71f51c),
	.w2(32'hbc2ecebe),
	.w3(32'hbc746631),
	.w4(32'hbcd9529a),
	.w5(32'h3b4439c2),
	.w6(32'hbd0b467d),
	.w7(32'h3c5acf02),
	.w8(32'h3c08f39b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab329d),
	.w1(32'h3bc5f748),
	.w2(32'hbd46102e),
	.w3(32'h3c6c32cd),
	.w4(32'hbc9dcdeb),
	.w5(32'hbc204fa0),
	.w6(32'h3d0a22ea),
	.w7(32'h3bea4502),
	.w8(32'hbc8f582f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05d48e),
	.w1(32'hbd0edcca),
	.w2(32'hbc457e7a),
	.w3(32'h3b15e284),
	.w4(32'h3b6defa7),
	.w5(32'h3cfa9e08),
	.w6(32'hbbdd503d),
	.w7(32'hbd1e6775),
	.w8(32'hbc45a3bd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb976e57),
	.w1(32'h3cab0c92),
	.w2(32'hbb15c059),
	.w3(32'h3bc18424),
	.w4(32'h3ab8d745),
	.w5(32'hbc0495d9),
	.w6(32'hbc13f009),
	.w7(32'h3be19c12),
	.w8(32'hbb5d3d3b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b994763),
	.w1(32'hbc951725),
	.w2(32'hbcc3eaee),
	.w3(32'hbcd1587a),
	.w4(32'hbd0fc8a5),
	.w5(32'hbc5874a0),
	.w6(32'hbd5dd985),
	.w7(32'h3d256c23),
	.w8(32'h3d74d342),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0162ca),
	.w1(32'hbbde2267),
	.w2(32'hbdc9d2d9),
	.w3(32'hbc0d75f0),
	.w4(32'h3ca98cc7),
	.w5(32'hbc3d067b),
	.w6(32'h3a769002),
	.w7(32'h3c5cac86),
	.w8(32'h3b6b7fee),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4e41e),
	.w1(32'hbc14898e),
	.w2(32'h3c204504),
	.w3(32'h3be6d66a),
	.w4(32'h3c8422cf),
	.w5(32'hbaa3cc1f),
	.w6(32'h3caee91b),
	.w7(32'hbc18ad9e),
	.w8(32'h3c62c61a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46e32c),
	.w1(32'h3c72397a),
	.w2(32'h3ce3697c),
	.w3(32'hbb8d3d4a),
	.w4(32'hbc0b302f),
	.w5(32'h3ae2c5e9),
	.w6(32'h3bf7e266),
	.w7(32'hbd32e1ce),
	.w8(32'hba00b307),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c986d60),
	.w1(32'hbc4ec94f),
	.w2(32'h3bb78a57),
	.w3(32'h3cbfdec5),
	.w4(32'hbc6fcbad),
	.w5(32'hbce9baa0),
	.w6(32'hbb829567),
	.w7(32'hbbc41084),
	.w8(32'hbb41e0de),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc210ad2),
	.w1(32'h3cda2352),
	.w2(32'h3c980fde),
	.w3(32'hbcbadd37),
	.w4(32'hbd17f9ef),
	.w5(32'h3c3fb091),
	.w6(32'hbc24fce8),
	.w7(32'hbb6bbbbf),
	.w8(32'hbaf13257),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca99adb),
	.w1(32'hbbc4d214),
	.w2(32'h3d81c4d4),
	.w3(32'h3ab46779),
	.w4(32'h3af91658),
	.w5(32'hbd1b233f),
	.w6(32'h3c944536),
	.w7(32'h3d0dad26),
	.w8(32'hbc8f22bb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bf43d),
	.w1(32'h3a21fd07),
	.w2(32'h3c6962a9),
	.w3(32'h3c372878),
	.w4(32'h3d32febd),
	.w5(32'hbb6c8639),
	.w6(32'h3bc7fa9a),
	.w7(32'h3b3a32cc),
	.w8(32'hbc72f2c6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4901c4),
	.w1(32'hb9cfe27b),
	.w2(32'hbd3ad458),
	.w3(32'h3a69403e),
	.w4(32'hbc3e4145),
	.w5(32'hbba14c1d),
	.w6(32'hbd1ead64),
	.w7(32'h3c047359),
	.w8(32'hbc890a05),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccb2909),
	.w1(32'hbcd7dd56),
	.w2(32'hbc4fc216),
	.w3(32'hbb2216e3),
	.w4(32'hbca588ae),
	.w5(32'h3d0c4cdc),
	.w6(32'h3c7a6df4),
	.w7(32'h3c805a34),
	.w8(32'hbc7fda41),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26fb4e),
	.w1(32'h3c552173),
	.w2(32'h3c2f279d),
	.w3(32'hb6969737),
	.w4(32'hbc846eef),
	.w5(32'hbc2bcb9d),
	.w6(32'h3bbb4ad6),
	.w7(32'hbc568612),
	.w8(32'hbc298bc5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb6d32a),
	.w1(32'h3c3d1603),
	.w2(32'hbc3455e3),
	.w3(32'hb99bd4be),
	.w4(32'hbd02d4b6),
	.w5(32'h3c557651),
	.w6(32'hbbdf3b7f),
	.w7(32'hbd7def5c),
	.w8(32'h3aad0ec1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb144db),
	.w1(32'h3b8fe9e8),
	.w2(32'hbbc3f3f9),
	.w3(32'hbd226fbc),
	.w4(32'hbc7250e8),
	.w5(32'hbc5105d9),
	.w6(32'hbc1a261d),
	.w7(32'h3cb631cb),
	.w8(32'h3bce3dcc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fee19),
	.w1(32'hbc0fdb59),
	.w2(32'hbd2aa8cf),
	.w3(32'h3c62dc75),
	.w4(32'h3bc7cca4),
	.w5(32'hbc96687d),
	.w6(32'hb9d4e0ea),
	.w7(32'h3cfe6a32),
	.w8(32'h3d1cbb26),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd750f29),
	.w1(32'hba877e74),
	.w2(32'hbca35646),
	.w3(32'hbcd331c8),
	.w4(32'h3c8ae55a),
	.w5(32'hbc61cb30),
	.w6(32'h3c88f0c1),
	.w7(32'h3d1f65d4),
	.w8(32'hbc2aa350),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd66942d),
	.w1(32'hbd16d50a),
	.w2(32'h3c28410e),
	.w3(32'hbd1442c2),
	.w4(32'h3c980555),
	.w5(32'h3d49541a),
	.w6(32'h3c27f86b),
	.w7(32'h3d17501c),
	.w8(32'h3cf481d2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc074a7a),
	.w1(32'hbb4f0c74),
	.w2(32'hbd720f19),
	.w3(32'h3bf52f03),
	.w4(32'h3b0c77a5),
	.w5(32'hbd1b15ad),
	.w6(32'hbd50e9fb),
	.w7(32'hbbb66949),
	.w8(32'h3c492515),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e61d03),
	.w1(32'h3c300405),
	.w2(32'h3c0528b1),
	.w3(32'h3c0b9e66),
	.w4(32'hbcbd0ff7),
	.w5(32'hbce342a8),
	.w6(32'hbc2f242a),
	.w7(32'h3bed10a7),
	.w8(32'h3c4ab9a7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb6f1e4),
	.w1(32'h3bc33857),
	.w2(32'h3c9f8e38),
	.w3(32'h3cadc54a),
	.w4(32'hbcbfdeec),
	.w5(32'hbc5732e4),
	.w6(32'h3914aa80),
	.w7(32'h3cfe2b9f),
	.w8(32'hbc3685f7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38526208),
	.w1(32'h3c247676),
	.w2(32'h3cba1975),
	.w3(32'h3c237394),
	.w4(32'hbd34ee29),
	.w5(32'h3bb08017),
	.w6(32'hbc359d7e),
	.w7(32'hbc3e9bc0),
	.w8(32'hbb877943),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cca6613),
	.w1(32'h3afb6dca),
	.w2(32'h3a2d37e4),
	.w3(32'h3c8a5a57),
	.w4(32'hbaf69b04),
	.w5(32'hbb25d728),
	.w6(32'hbcc5acc7),
	.w7(32'h3bfadbbe),
	.w8(32'hbca2cd02),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcebb1a3),
	.w1(32'h3c959d5e),
	.w2(32'h3c5eadb3),
	.w3(32'h3b0e62a0),
	.w4(32'hbd74b620),
	.w5(32'hbc27d7d1),
	.w6(32'hbbc4fe23),
	.w7(32'hbcfbab18),
	.w8(32'h3b8eaea5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a5bfb),
	.w1(32'hbcfbf8b7),
	.w2(32'hbcda9b99),
	.w3(32'h3c43d74a),
	.w4(32'h3b4739c3),
	.w5(32'hbcdee5a6),
	.w6(32'hbd1f3a10),
	.w7(32'hbbe09b59),
	.w8(32'h3c102a04),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e5e70),
	.w1(32'hbbdf4b17),
	.w2(32'hbc98b247),
	.w3(32'hbab898d8),
	.w4(32'h3c7103b2),
	.w5(32'hbd13747e),
	.w6(32'hbcd30af1),
	.w7(32'hbcc715d7),
	.w8(32'hbcdfdd36),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32a49b),
	.w1(32'hbc6bf98b),
	.w2(32'h3d2bf977),
	.w3(32'hbbca31e5),
	.w4(32'hbd28bca0),
	.w5(32'hbbacd90f),
	.w6(32'h3c684698),
	.w7(32'h3b4a6916),
	.w8(32'hbc0bd391),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dfca0),
	.w1(32'h3c01f7ed),
	.w2(32'hbc55ba80),
	.w3(32'h3866d698),
	.w4(32'h3cb99171),
	.w5(32'hbd776cd9),
	.w6(32'hbb32e978),
	.w7(32'h39c40ace),
	.w8(32'hbd316d60),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c904a),
	.w1(32'hbd0e0517),
	.w2(32'hbda2fd50),
	.w3(32'hbd27ceb7),
	.w4(32'h3a17688e),
	.w5(32'h3cd61414),
	.w6(32'hba392e5e),
	.w7(32'h3c174f58),
	.w8(32'h3c0bbf4c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1cde6e),
	.w1(32'hbc4d94ae),
	.w2(32'hbb460d47),
	.w3(32'h3cde7956),
	.w4(32'h3d03b30b),
	.w5(32'h3c1a6047),
	.w6(32'h3c6b6603),
	.w7(32'h3ca87998),
	.w8(32'h39a7ee85),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce6cd22),
	.w1(32'h3c86e8f0),
	.w2(32'h3ce96ee9),
	.w3(32'hbd257d68),
	.w4(32'h3c08329b),
	.w5(32'hbb708bf8),
	.w6(32'hbd25c05d),
	.w7(32'hbcd390a9),
	.w8(32'h3ba1f746),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc667c2),
	.w1(32'hbd137fac),
	.w2(32'hbc683c3a),
	.w3(32'hba6fb186),
	.w4(32'hbc599158),
	.w5(32'h3a4fabea),
	.w6(32'h3cd35990),
	.w7(32'h3cbf3224),
	.w8(32'hbc6f7c46),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9aa778),
	.w1(32'hbd02de5d),
	.w2(32'hbb0cb46b),
	.w3(32'h3cd86b69),
	.w4(32'h3d168b56),
	.w5(32'h3ba9cf5d),
	.w6(32'hbb2799eb),
	.w7(32'hbb196e05),
	.w8(32'hbc1b7528),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb93510),
	.w1(32'h3a35e873),
	.w2(32'h3bcc8b82),
	.w3(32'hbc76beba),
	.w4(32'h3cc071e5),
	.w5(32'hbc3ea979),
	.w6(32'h3d057b30),
	.w7(32'hba220f9b),
	.w8(32'h3bf447d3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc286180),
	.w1(32'hbac2290d),
	.w2(32'h3c69366f),
	.w3(32'hbbdf96ae),
	.w4(32'h3d362b00),
	.w5(32'hbbfc504a),
	.w6(32'h3bb6513f),
	.w7(32'hbb5acdf9),
	.w8(32'h3ca9e1db),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dca7c),
	.w1(32'h3cc3e3c5),
	.w2(32'hbb8404ce),
	.w3(32'hba7abde0),
	.w4(32'hbccf46a8),
	.w5(32'h3b831724),
	.w6(32'h3c623ae7),
	.w7(32'h3c3ed4a5),
	.w8(32'hbd1bb404),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9be902),
	.w1(32'h3c964429),
	.w2(32'h3b8ded9a),
	.w3(32'hbc26eb3f),
	.w4(32'hbc0b6b10),
	.w5(32'hbc4645fa),
	.w6(32'h3d47d978),
	.w7(32'hbc0211e5),
	.w8(32'h3c1da99d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10bd96),
	.w1(32'h3c6cc930),
	.w2(32'hbd87f1ac),
	.w3(32'hbb8dd586),
	.w4(32'h3b0ce7ac),
	.w5(32'hbbf5d4d9),
	.w6(32'h3d01be8f),
	.w7(32'h3c520f5b),
	.w8(32'hbba66fa4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbad53),
	.w1(32'hbc987ec2),
	.w2(32'hbc79c412),
	.w3(32'hbb39c6de),
	.w4(32'h3bd540bd),
	.w5(32'h3be540c2),
	.w6(32'h3cb0516a),
	.w7(32'h3cddfc03),
	.w8(32'h3d975348),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55d2e8),
	.w1(32'h3cf177e0),
	.w2(32'h3c1a7a21),
	.w3(32'h3cb39a64),
	.w4(32'h3bf1fe77),
	.w5(32'h3be32ca4),
	.w6(32'h3c6d534f),
	.w7(32'h3c60e046),
	.w8(32'hbc5856cf),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84094f),
	.w1(32'h3c4504e1),
	.w2(32'hbc12cf11),
	.w3(32'h3b94aa1e),
	.w4(32'hbbe6a29d),
	.w5(32'hbc3e4301),
	.w6(32'h3ad16a29),
	.w7(32'hb9be4627),
	.w8(32'h3d894597),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ae371),
	.w1(32'h3cac4c95),
	.w2(32'hbceb973d),
	.w3(32'h3c27c3a3),
	.w4(32'hbc7091dc),
	.w5(32'hbca2f4bc),
	.w6(32'hbb8f4137),
	.w7(32'hbc64e9d0),
	.w8(32'hbbd926b1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34ac1c),
	.w1(32'hbae9168e),
	.w2(32'h3b1bf724),
	.w3(32'hbc2021a1),
	.w4(32'hbce0ae16),
	.w5(32'h3cbeeb8e),
	.w6(32'hbcf6db7c),
	.w7(32'hbc3f2671),
	.w8(32'h3c888e75),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0d320),
	.w1(32'h3c885777),
	.w2(32'hbbe67919),
	.w3(32'h3c9fe86b),
	.w4(32'h3c52f8eb),
	.w5(32'hb9e44c5c),
	.w6(32'h3c9d37fd),
	.w7(32'h3c0f30d4),
	.w8(32'h3bd2c976),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0506a2),
	.w1(32'hbacd3a49),
	.w2(32'h3b723b62),
	.w3(32'h3d0b3a22),
	.w4(32'hbb4b454c),
	.w5(32'hbc65b382),
	.w6(32'h3b93e623),
	.w7(32'h3bb4736e),
	.w8(32'h3b0996f5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54a253),
	.w1(32'h3bab03bb),
	.w2(32'h3b5a9fc2),
	.w3(32'hbc9f6761),
	.w4(32'hbc222f3f),
	.w5(32'h3bc8a533),
	.w6(32'hbc0826c8),
	.w7(32'h3ae8bc54),
	.w8(32'hbbd5eaf0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bfe18),
	.w1(32'hbaa752e8),
	.w2(32'hbd374d47),
	.w3(32'h3c0bc1dc),
	.w4(32'hbc23249e),
	.w5(32'hbae938bb),
	.w6(32'h3cdbd859),
	.w7(32'hbbbc26eb),
	.w8(32'h3c914e55),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda40d7),
	.w1(32'hba6a403a),
	.w2(32'h3d334d36),
	.w3(32'hbd4d5969),
	.w4(32'hbc45cf5f),
	.w5(32'h3d491d1d),
	.w6(32'h3d1a24ce),
	.w7(32'h3c858799),
	.w8(32'h3beea0ec),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab3753),
	.w1(32'h3c13479d),
	.w2(32'h3ac58655),
	.w3(32'h3ba19de3),
	.w4(32'h3caccfcd),
	.w5(32'hbd09ed1e),
	.w6(32'hbc57b56f),
	.w7(32'hbbf89339),
	.w8(32'hbc3253c0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea36cd),
	.w1(32'h3c2bb5e9),
	.w2(32'hbc0c398f),
	.w3(32'hbd12fc3c),
	.w4(32'h3c918895),
	.w5(32'hbb05045a),
	.w6(32'h3af26714),
	.w7(32'h3bd7a2d1),
	.w8(32'hbc5440fb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9724e6),
	.w1(32'hbc972cae),
	.w2(32'hbcd22dd4),
	.w3(32'h3cb06fde),
	.w4(32'hbd1094e6),
	.w5(32'hbbbd7ece),
	.w6(32'hbba6cb6a),
	.w7(32'hbcebfc02),
	.w8(32'h3d23dd49),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03997d),
	.w1(32'hbd34d36c),
	.w2(32'hbb68fdc7),
	.w3(32'hbc269877),
	.w4(32'hbbefcb2d),
	.w5(32'h3d4cda7a),
	.w6(32'hbc56b00a),
	.w7(32'hbbbf052c),
	.w8(32'hbbbb3700),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba11b4d),
	.w1(32'hba9c2c14),
	.w2(32'hbc806907),
	.w3(32'hbc554d7d),
	.w4(32'h3c2444fa),
	.w5(32'hbd151b2e),
	.w6(32'hbc8e9dd6),
	.w7(32'h3c90e48b),
	.w8(32'hbb195ca6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3105c0),
	.w1(32'h3aedc7ab),
	.w2(32'h3c60734c),
	.w3(32'hbd2a1525),
	.w4(32'hbb13b426),
	.w5(32'h3c8f3e4a),
	.w6(32'hbd5fb041),
	.w7(32'hba9dbaa3),
	.w8(32'h3a476363),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd087843),
	.w1(32'h3c7752f3),
	.w2(32'h3c29ab07),
	.w3(32'h3c62fc12),
	.w4(32'hbbdf6533),
	.w5(32'h3b3d5c19),
	.w6(32'hbbf50fbb),
	.w7(32'hbcf580b3),
	.w8(32'h3c8235ea),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a552a),
	.w1(32'hbc49da05),
	.w2(32'h3b912d02),
	.w3(32'hbc9da7b8),
	.w4(32'hbb323bd3),
	.w5(32'h3b05f9bd),
	.w6(32'hbd0f3a7b),
	.w7(32'hbbfdaf63),
	.w8(32'h3d2e2015),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf29b6),
	.w1(32'hbc03485a),
	.w2(32'hbce0a6dd),
	.w3(32'h3cc5b24b),
	.w4(32'hbd79a223),
	.w5(32'hbbe5c8fa),
	.w6(32'hbd53f8e4),
	.w7(32'hbc1ca953),
	.w8(32'h3a48f702),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0b1743),
	.w1(32'h3a473c99),
	.w2(32'h3bde1964),
	.w3(32'hbd52caec),
	.w4(32'hbc950ee3),
	.w5(32'hbccf4cd0),
	.w6(32'h3c702312),
	.w7(32'h3b982d12),
	.w8(32'h3a8b0ba3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4ba40),
	.w1(32'hbce853b3),
	.w2(32'hbd12fe5e),
	.w3(32'h3cbf3a0c),
	.w4(32'h3b10916e),
	.w5(32'hbb7aa16b),
	.w6(32'hba9be413),
	.w7(32'hbcbcbce0),
	.w8(32'h3c02c2a1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c5274),
	.w1(32'hbccaeb09),
	.w2(32'h3c6868ed),
	.w3(32'hbcc0cbb1),
	.w4(32'h3bdfb169),
	.w5(32'hbbf97345),
	.w6(32'hbc016e46),
	.w7(32'h3c27bae1),
	.w8(32'hbbe0e116),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba628a9),
	.w1(32'hbc0bd4ee),
	.w2(32'hbc6aa1e9),
	.w3(32'hbc59c48a),
	.w4(32'hbc375bdf),
	.w5(32'h3a5322ec),
	.w6(32'h3b3825d7),
	.w7(32'hbccacecf),
	.w8(32'hbd504b37),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule