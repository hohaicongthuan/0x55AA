module layer_10_featuremap_300(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2d13d),
	.w1(32'hbb1d3ae5),
	.w2(32'h39ea4c41),
	.w3(32'h3b13ecef),
	.w4(32'h3a75b5a7),
	.w5(32'h3aaed3b3),
	.w6(32'hbb30ea6d),
	.w7(32'hbb344d06),
	.w8(32'h3a19c534),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69d701),
	.w1(32'hba47b3a8),
	.w2(32'hba3702a7),
	.w3(32'hba9b8ca8),
	.w4(32'hbb301a20),
	.w5(32'hba97e5da),
	.w6(32'h388b014d),
	.w7(32'h3987f728),
	.w8(32'hbb9012ff),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabce302),
	.w1(32'hba287b70),
	.w2(32'hba78f318),
	.w3(32'hbb1178a7),
	.w4(32'hbab51e56),
	.w5(32'hbad437c0),
	.w6(32'hba721237),
	.w7(32'h39abd4eb),
	.w8(32'h3a94b258),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02df08),
	.w1(32'h3b46eee7),
	.w2(32'h3b25a302),
	.w3(32'h392b0349),
	.w4(32'h3a743eb7),
	.w5(32'h3bcfb284),
	.w6(32'h3adc6034),
	.w7(32'h3b584f51),
	.w8(32'hbb32e2f9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b178d51),
	.w1(32'hbab0b514),
	.w2(32'hbab74925),
	.w3(32'h3ba9baa7),
	.w4(32'h3b8edc8c),
	.w5(32'h3b7a257e),
	.w6(32'hbb97ecfa),
	.w7(32'hbb27c623),
	.w8(32'h3a5d5561),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab215d0),
	.w1(32'h3a383cbf),
	.w2(32'h3a8e7476),
	.w3(32'h3ba1b2bf),
	.w4(32'h3b9f98aa),
	.w5(32'hbaa6e8a8),
	.w6(32'h390bcb1b),
	.w7(32'h39275be2),
	.w8(32'hba199066),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00e52d),
	.w1(32'h3a44fed9),
	.w2(32'hbab29fbc),
	.w3(32'h39d69ba3),
	.w4(32'hbad068d2),
	.w5(32'hbb34c556),
	.w6(32'h3aed2db1),
	.w7(32'hba006580),
	.w8(32'hbb8732fe),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dfc95),
	.w1(32'hbb8a3f25),
	.w2(32'hbb6ea17c),
	.w3(32'hbb94d38a),
	.w4(32'hbb5df5ec),
	.w5(32'h3b49b1cb),
	.w6(32'hbbd16a2e),
	.w7(32'hbb98a354),
	.w8(32'h3a81d4b6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fb12a),
	.w1(32'h3b1e7f07),
	.w2(32'h3b46a930),
	.w3(32'h3b89cde8),
	.w4(32'h3b6391c8),
	.w5(32'h3b5a2deb),
	.w6(32'h3ac95153),
	.w7(32'h3a890e9f),
	.w8(32'h3999bbb0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3244c1),
	.w1(32'h3775eeb9),
	.w2(32'hbb8330bc),
	.w3(32'h3b59a197),
	.w4(32'h3b982a5b),
	.w5(32'hbb962324),
	.w6(32'hb9bf5705),
	.w7(32'h3aff077f),
	.w8(32'hbb98c794),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08de4d),
	.w1(32'hb9cf337b),
	.w2(32'hba5036a8),
	.w3(32'h3b16e6db),
	.w4(32'h3b4168ec),
	.w5(32'hba4e4383),
	.w6(32'h3aa5718b),
	.w7(32'h3a6522a4),
	.w8(32'h39cf2d8d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05cc5d),
	.w1(32'h3a364116),
	.w2(32'hbb5166db),
	.w3(32'h38ddae84),
	.w4(32'hba8074d4),
	.w5(32'hbb527ea5),
	.w6(32'h3ae9b3a3),
	.w7(32'hb9d7bc18),
	.w8(32'hbb445b60),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb457495),
	.w1(32'hb9d15e3c),
	.w2(32'hbb80a106),
	.w3(32'hbaa7da0f),
	.w4(32'hbab24c12),
	.w5(32'hbb5bdfc6),
	.w6(32'h3a35a656),
	.w7(32'hb9f8f8fc),
	.w8(32'hbb39b86c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04af83),
	.w1(32'h3afc4511),
	.w2(32'h3b411360),
	.w3(32'hba97f53f),
	.w4(32'hba3e5d54),
	.w5(32'hbb0b14c9),
	.w6(32'h3a6d0b19),
	.w7(32'h3a898593),
	.w8(32'hba4dc909),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2e863),
	.w1(32'h3ac4fe79),
	.w2(32'hbb3822fa),
	.w3(32'hba96d627),
	.w4(32'h39989a3c),
	.w5(32'hba47b3b0),
	.w6(32'hba2e7caa),
	.w7(32'h3a8cfb25),
	.w8(32'hbb3ade88),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb772a1a),
	.w1(32'hbb640eb3),
	.w2(32'hbb7de76c),
	.w3(32'h3a3c149c),
	.w4(32'h3ab082a3),
	.w5(32'h39b1e364),
	.w6(32'hba92854f),
	.w7(32'hba003ec5),
	.w8(32'hb94b1f3b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addcb2f),
	.w1(32'hbaaa969f),
	.w2(32'h3a21aefd),
	.w3(32'h3aa89f31),
	.w4(32'h3b0f9ed3),
	.w5(32'hbb01b21e),
	.w6(32'h3a0d242e),
	.w7(32'hb9bed9b1),
	.w8(32'hbaeb26fe),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb97dc8),
	.w1(32'hbb8a3301),
	.w2(32'hbbadc96e),
	.w3(32'hbb9e7230),
	.w4(32'hbb9edc85),
	.w5(32'hbbf79546),
	.w6(32'hbb915182),
	.w7(32'hbba6c2c1),
	.w8(32'hbbf7c2ed),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05c9b6),
	.w1(32'hbadbce60),
	.w2(32'hbb07d5d6),
	.w3(32'hbb41cf48),
	.w4(32'hba86f09f),
	.w5(32'hbb65d954),
	.w6(32'hbb4dc6a6),
	.w7(32'hbb75ef1d),
	.w8(32'hbb6aeca7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9782c1),
	.w1(32'hbb2ce164),
	.w2(32'hbaf83c84),
	.w3(32'hbafdd0e2),
	.w4(32'hbad94323),
	.w5(32'hbb399276),
	.w6(32'hb9fdff73),
	.w7(32'hba4cd05a),
	.w8(32'hbb13932f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba444fd8),
	.w1(32'h3a3164fa),
	.w2(32'h3b3c8f7d),
	.w3(32'h3b10a692),
	.w4(32'h3af5f5c9),
	.w5(32'hba52ed66),
	.w6(32'h3af450a2),
	.w7(32'h3b4117e0),
	.w8(32'h3a03cc75),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a904bf7),
	.w1(32'h3b86c801),
	.w2(32'h3a6d4192),
	.w3(32'h39824b75),
	.w4(32'h39c5c74d),
	.w5(32'h3a71efce),
	.w6(32'h3b2d3eaf),
	.w7(32'h3b1b9b53),
	.w8(32'h39c83426),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89a085),
	.w1(32'h3a44b050),
	.w2(32'hbb8df9c6),
	.w3(32'h39d70662),
	.w4(32'h3aa4a620),
	.w5(32'hbbc8ffd4),
	.w6(32'hba94bea1),
	.w7(32'hba8a4c59),
	.w8(32'hbc16dd0b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac59fcc),
	.w1(32'h3aa8fefc),
	.w2(32'hbb53bba0),
	.w3(32'h3b59d47b),
	.w4(32'h3af6988d),
	.w5(32'hbb188763),
	.w6(32'hb8bc73e5),
	.w7(32'h3b447df7),
	.w8(32'hbbd1e0ec),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5295a3),
	.w1(32'h3a30873e),
	.w2(32'hbb40bd0f),
	.w3(32'hbae26619),
	.w4(32'h3b143e25),
	.w5(32'hbb91adf0),
	.w6(32'hbb9e23db),
	.w7(32'h397826d4),
	.w8(32'hbb257d86),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b214dbb),
	.w1(32'h3ac421d3),
	.w2(32'h3af003c7),
	.w3(32'hba86cce7),
	.w4(32'h3b0d1b3b),
	.w5(32'hba47cae4),
	.w6(32'h39bb1e28),
	.w7(32'h3a938e9e),
	.w8(32'hba9ff5f3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7262305),
	.w1(32'h3ad211c1),
	.w2(32'h368308e9),
	.w3(32'h3a483660),
	.w4(32'h3aca9c72),
	.w5(32'h3c1e2277),
	.w6(32'h3aac18f1),
	.w7(32'hb91d05d8),
	.w8(32'h3b401193),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc78a7c),
	.w1(32'h3aba161c),
	.w2(32'h3b93e242),
	.w3(32'h3bba6c16),
	.w4(32'h3bc4b16b),
	.w5(32'h3a9dff0a),
	.w6(32'hbb01609a),
	.w7(32'h3a93743b),
	.w8(32'h3a80a66e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae8288),
	.w1(32'h3a4d8e3b),
	.w2(32'h3b1c4e10),
	.w3(32'hbab02b48),
	.w4(32'h3ae3d5c9),
	.w5(32'hba8ee031),
	.w6(32'hb9802589),
	.w7(32'h3a8936b0),
	.w8(32'hbb18146d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70855c),
	.w1(32'hb80d0f93),
	.w2(32'hbb583498),
	.w3(32'hbb57e7aa),
	.w4(32'h378e62a5),
	.w5(32'hb9512af9),
	.w6(32'hbb4f9d7f),
	.w7(32'h3a64ff80),
	.w8(32'hbbb513f4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff8063),
	.w1(32'hbb19ed4b),
	.w2(32'h3a2182bd),
	.w3(32'hbabf017f),
	.w4(32'hba49a4c4),
	.w5(32'hb9eca0b6),
	.w6(32'hbb9556cb),
	.w7(32'hba035dc0),
	.w8(32'h3a8585e7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31da59),
	.w1(32'h3a06d8e5),
	.w2(32'h3a13829d),
	.w3(32'h397d2b06),
	.w4(32'hbaff4d89),
	.w5(32'hba10c179),
	.w6(32'h3af4c512),
	.w7(32'h3b05cedd),
	.w8(32'hba9c227d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3884a741),
	.w1(32'hbb5c87ff),
	.w2(32'h3a8f0db6),
	.w3(32'hbb668621),
	.w4(32'h3b954f8a),
	.w5(32'hbb8e4651),
	.w6(32'hbb50cd44),
	.w7(32'h3af0fef2),
	.w8(32'hbb90d946),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb627804),
	.w1(32'hbb0b9497),
	.w2(32'hbb121dd2),
	.w3(32'hbab498a2),
	.w4(32'hbb065dda),
	.w5(32'hb86fe095),
	.w6(32'hbb3ba33c),
	.w7(32'hbb648155),
	.w8(32'hbab2a73a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03a422),
	.w1(32'hba3401c2),
	.w2(32'hba974bc3),
	.w3(32'hb7f937a7),
	.w4(32'hb8f03b37),
	.w5(32'hbb13864c),
	.w6(32'h3af9cd16),
	.w7(32'hb8d84fc5),
	.w8(32'hbb3f82fa),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd471),
	.w1(32'hbb4a5b48),
	.w2(32'hbb30e66a),
	.w3(32'hb97b76fa),
	.w4(32'h3aa7fd49),
	.w5(32'hbb586ece),
	.w6(32'hbb0abb74),
	.w7(32'hbb12c8ab),
	.w8(32'hbb9bb31e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb377956),
	.w1(32'hbad07c57),
	.w2(32'hbb5aafa3),
	.w3(32'h38da78c4),
	.w4(32'hb6df45fb),
	.w5(32'hbabf871b),
	.w6(32'h3a49481a),
	.w7(32'h3a5e5d7d),
	.w8(32'hbb739005),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9808ce),
	.w1(32'h3b90cc4d),
	.w2(32'hba58ce28),
	.w3(32'h3b445665),
	.w4(32'h3c1c9d00),
	.w5(32'h3b092ed6),
	.w6(32'hbb2e1236),
	.w7(32'h39b3c0ae),
	.w8(32'hbb60d8c4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa2046),
	.w1(32'h3b6cf0fe),
	.w2(32'h3a0711af),
	.w3(32'hbb83334b),
	.w4(32'h3b00f509),
	.w5(32'h3a0a50d0),
	.w6(32'hbbb2fb21),
	.w7(32'hbad90975),
	.w8(32'hbaa57650),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0076e1),
	.w1(32'h3b3ed3d1),
	.w2(32'hbaa90d71),
	.w3(32'h3b2f950a),
	.w4(32'h3a9cf995),
	.w5(32'h3a7b31e9),
	.w6(32'h3b60b0d8),
	.w7(32'h3ad640d2),
	.w8(32'hb9809db0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b2d17),
	.w1(32'hb96ff91f),
	.w2(32'hba91df8b),
	.w3(32'hba83e9e2),
	.w4(32'hba32c28c),
	.w5(32'h3a4d7554),
	.w6(32'hba87bb2e),
	.w7(32'hbb05c06a),
	.w8(32'h3b01abe7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b828f1d),
	.w1(32'h3b65941b),
	.w2(32'h3b0d5e97),
	.w3(32'h3b2e4e3b),
	.w4(32'h3b516906),
	.w5(32'hbafe53cd),
	.w6(32'h3ba22a3f),
	.w7(32'h3b472705),
	.w8(32'hbad06265),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6327b7),
	.w1(32'hbb50cabe),
	.w2(32'hbb0ebb77),
	.w3(32'hbb672d75),
	.w4(32'hbb69c1bd),
	.w5(32'hbb25656d),
	.w6(32'hbb8106cf),
	.w7(32'hbb7e4a87),
	.w8(32'hbb649113),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2114fc),
	.w1(32'hbc12e6f0),
	.w2(32'hbc1abef4),
	.w3(32'hbbd5df10),
	.w4(32'hbb58cea7),
	.w5(32'hbbaa574b),
	.w6(32'hbc257769),
	.w7(32'hbc0ee441),
	.w8(32'hbbb2cf6c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399110fb),
	.w1(32'h3bbcb120),
	.w2(32'h3a27b4ce),
	.w3(32'h3aaa33ad),
	.w4(32'h3bb32c62),
	.w5(32'hbb9a8316),
	.w6(32'h3b860120),
	.w7(32'h3becee43),
	.w8(32'hbb58154e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d0924),
	.w1(32'hbb3a7302),
	.w2(32'hbc0273c4),
	.w3(32'hbb7506fa),
	.w4(32'hba8a8fd6),
	.w5(32'hbbb90308),
	.w6(32'hbbb191c5),
	.w7(32'hba2a6032),
	.w8(32'hbb956eca),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90c789),
	.w1(32'h3aa92894),
	.w2(32'hbb55b87a),
	.w3(32'hb95a4ee6),
	.w4(32'h3b703d85),
	.w5(32'h3a808965),
	.w6(32'hb97d9c49),
	.w7(32'h3ac46714),
	.w8(32'hb8bf699b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af793d0),
	.w1(32'h3b24949c),
	.w2(32'h39279d4e),
	.w3(32'h3ab464a3),
	.w4(32'hbac7eb6e),
	.w5(32'hbb8d604a),
	.w6(32'h3b325f21),
	.w7(32'hba35da46),
	.w8(32'hbb9c839b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfdf10),
	.w1(32'h3a226af2),
	.w2(32'h39fce48c),
	.w3(32'hb9920e5c),
	.w4(32'hb8649472),
	.w5(32'h39d5c36a),
	.w6(32'h3a114c0a),
	.w7(32'h39e048ad),
	.w8(32'h3a44d2fa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94661b),
	.w1(32'h3b4d4e0f),
	.w2(32'h3a29172a),
	.w3(32'h3a3df60f),
	.w4(32'hba179838),
	.w5(32'h3c17f2af),
	.w6(32'h3b40b6a0),
	.w7(32'h3a11eb3c),
	.w8(32'h3bbf459f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a4cf3),
	.w1(32'hb9920c69),
	.w2(32'h3af1d192),
	.w3(32'h3a697c21),
	.w4(32'h3b40d0f0),
	.w5(32'hb9ceefbe),
	.w6(32'hba1fc467),
	.w7(32'h3aa8ad09),
	.w8(32'hbaf2a5aa),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd3a8a),
	.w1(32'hbb5962cb),
	.w2(32'hbb767048),
	.w3(32'h39ee4e85),
	.w4(32'h3a1d2466),
	.w5(32'hba6ce33d),
	.w6(32'hbb1645b9),
	.w7(32'h39b1adb7),
	.w8(32'hba2fcf02),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba744019),
	.w1(32'hbae08d9c),
	.w2(32'hbb0af1c8),
	.w3(32'hba3dc822),
	.w4(32'h38b085bc),
	.w5(32'hbaff71e1),
	.w6(32'hba928dcc),
	.w7(32'h3a7d86d1),
	.w8(32'h39b01cc1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d1425),
	.w1(32'h3aa9a9ad),
	.w2(32'hbbecdbc0),
	.w3(32'h3b372d4c),
	.w4(32'hbae73541),
	.w5(32'hbc102ad4),
	.w6(32'h3b897337),
	.w7(32'hbaeaa0bd),
	.w8(32'hbbf0a866),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1349f2),
	.w1(32'hba794119),
	.w2(32'h390c807b),
	.w3(32'hbab41ccf),
	.w4(32'hb95347be),
	.w5(32'h3af205ce),
	.w6(32'hbacc2ade),
	.w7(32'h39eab25d),
	.w8(32'hba01b1ce),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9eced),
	.w1(32'hbad08fa7),
	.w2(32'h38eb6417),
	.w3(32'h3836cb27),
	.w4(32'hb89c6b5a),
	.w5(32'h396ba094),
	.w6(32'hba060785),
	.w7(32'hba0d1cdb),
	.w8(32'hb9a10376),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb811f456),
	.w1(32'hbaac0dbe),
	.w2(32'hbb060b6c),
	.w3(32'hbb066b76),
	.w4(32'hbaec392e),
	.w5(32'hba758cf9),
	.w6(32'hbaea7b70),
	.w7(32'hbb211313),
	.w8(32'h39a284a6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab1fa3),
	.w1(32'h39adce48),
	.w2(32'h39bfc072),
	.w3(32'h3aefcaff),
	.w4(32'h3b710c67),
	.w5(32'h3aa8627d),
	.w6(32'h3b463cc0),
	.w7(32'h3b35a553),
	.w8(32'h3ad27928),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11a993),
	.w1(32'h3b9a1970),
	.w2(32'h3b2cedd2),
	.w3(32'h3ac16d6d),
	.w4(32'h3b1ee514),
	.w5(32'h3b83e3c9),
	.w6(32'h3b649203),
	.w7(32'h3b246864),
	.w8(32'h3ae0aaef),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93f551),
	.w1(32'h3ad78b8a),
	.w2(32'hbba1dc3e),
	.w3(32'h3b014ceb),
	.w4(32'h3a887fb9),
	.w5(32'hb8bf6ad2),
	.w6(32'h3ab03f77),
	.w7(32'hbb5cbbdb),
	.w8(32'hb9d18cf7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88c0dc),
	.w1(32'hbb0b31b7),
	.w2(32'hbb3513bb),
	.w3(32'hbb1e61b0),
	.w4(32'hba8c030b),
	.w5(32'hbb72d24d),
	.w6(32'hba9f439e),
	.w7(32'hbadc1b13),
	.w8(32'hbadb387f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14c7ff),
	.w1(32'hba139577),
	.w2(32'hba416e9e),
	.w3(32'hbbbb6489),
	.w4(32'hbb81a10b),
	.w5(32'h3a5de257),
	.w6(32'hbb632c2b),
	.w7(32'hbb3ca531),
	.w8(32'hbb5a4522),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953807f),
	.w1(32'hba26c04a),
	.w2(32'hba509075),
	.w3(32'h3b0e1250),
	.w4(32'h3ad67fa3),
	.w5(32'h3ad14b37),
	.w6(32'hba97f5df),
	.w7(32'hbadd4023),
	.w8(32'h39dca255),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb854bc42),
	.w1(32'hb929e62e),
	.w2(32'hba2164a7),
	.w3(32'h3aa7ca2f),
	.w4(32'h3a1e2bd0),
	.w5(32'hbad50d38),
	.w6(32'h3a8910e5),
	.w7(32'hba603ff1),
	.w8(32'hb9ab888d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab950ea),
	.w1(32'h3a1bbad5),
	.w2(32'h3b3c8109),
	.w3(32'hbb3257c2),
	.w4(32'h3a8b2a58),
	.w5(32'hba24f5ca),
	.w6(32'h3acf0dee),
	.w7(32'h3b9670fd),
	.w8(32'hbace93c5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46592e),
	.w1(32'hbb318b36),
	.w2(32'hbb5e4ec7),
	.w3(32'h392f3365),
	.w4(32'hba0d12f5),
	.w5(32'hbae568f9),
	.w6(32'hbb616e05),
	.w7(32'hbb445280),
	.w8(32'hba72454e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac447b1),
	.w1(32'hbb06bb08),
	.w2(32'hbb4d746c),
	.w3(32'hbb26260e),
	.w4(32'hbb18d6de),
	.w5(32'h3adc2d87),
	.w6(32'hbb6b279c),
	.w7(32'hbb944530),
	.w8(32'h3a8702a5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b9dcc),
	.w1(32'h3b7edcbc),
	.w2(32'hb9a4882e),
	.w3(32'h3b700b6f),
	.w4(32'h3af91601),
	.w5(32'hbbdc3c74),
	.w6(32'h3b1e3d5d),
	.w7(32'h3b7fd2d1),
	.w8(32'hbb832cf7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabde6bc),
	.w1(32'hbb2efa3f),
	.w2(32'h3b4abccc),
	.w3(32'hbb9ab0bc),
	.w4(32'h3b967620),
	.w5(32'hbba29a5d),
	.w6(32'hbbb6d111),
	.w7(32'h3bbb2275),
	.w8(32'hbb855926),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ff91a),
	.w1(32'hbacd6e9a),
	.w2(32'hbc53ca91),
	.w3(32'h3a4dc95b),
	.w4(32'h3bc44025),
	.w5(32'hbb5e0dc6),
	.w6(32'hbb7ca997),
	.w7(32'h3aa4bb9c),
	.w8(32'hbb9be5e5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39634757),
	.w1(32'h3a882719),
	.w2(32'h3a7b727b),
	.w3(32'h3a7ee92f),
	.w4(32'h3a0c4699),
	.w5(32'hbb3959a1),
	.w6(32'h3987066d),
	.w7(32'hba2dc754),
	.w8(32'hbb01dc17),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e514f),
	.w1(32'hbac86a55),
	.w2(32'h3adde22c),
	.w3(32'h394d4f8f),
	.w4(32'h3b2ea0b7),
	.w5(32'h3abb397d),
	.w6(32'h3a123074),
	.w7(32'h3b914ea0),
	.w8(32'h3b376720),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0dbf7),
	.w1(32'h3aa44626),
	.w2(32'h3952b8fb),
	.w3(32'hb9dbb425),
	.w4(32'hbad4f96a),
	.w5(32'hbafce65b),
	.w6(32'h3ae8341e),
	.w7(32'hba1a6d12),
	.w8(32'hbb147a65),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e7e22),
	.w1(32'hbb32a70a),
	.w2(32'hbb0fe116),
	.w3(32'hbb2d8dd3),
	.w4(32'hbb76baeb),
	.w5(32'h394fa6bc),
	.w6(32'hbb1ae278),
	.w7(32'hbb8af299),
	.w8(32'h3ab7dd23),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb824c612),
	.w1(32'hbb424332),
	.w2(32'hbb6242c3),
	.w3(32'h3b601fc2),
	.w4(32'hb9e5342d),
	.w5(32'hbb5a7951),
	.w6(32'h3b086754),
	.w7(32'hbb775154),
	.w8(32'hbb0f01f5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae75ece),
	.w1(32'hbaa4ce79),
	.w2(32'hbb2de5ad),
	.w3(32'hbb7337b6),
	.w4(32'hbb8e7741),
	.w5(32'h3a631db7),
	.w6(32'hbb2ed5e2),
	.w7(32'hbb5ab54b),
	.w8(32'hbb161ae0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae9554),
	.w1(32'hbb380a18),
	.w2(32'hbbd27de9),
	.w3(32'hba2c3ddc),
	.w4(32'hba83e751),
	.w5(32'hbb3b1e1c),
	.w6(32'hbba915fc),
	.w7(32'hbb58c744),
	.w8(32'hbb7bdce5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb647716),
	.w1(32'hba530510),
	.w2(32'hbaa2daf0),
	.w3(32'hb929a251),
	.w4(32'h3aef5809),
	.w5(32'hbafae9ca),
	.w6(32'hbaee9599),
	.w7(32'h3a39788a),
	.w8(32'hbb30b55a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba697bad),
	.w1(32'h3a0a8f72),
	.w2(32'hbb3da857),
	.w3(32'hbab8843f),
	.w4(32'h3a50ab91),
	.w5(32'h3ad2138c),
	.w6(32'hbb1421d2),
	.w7(32'h387f1287),
	.w8(32'hbadcdd4e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43747d),
	.w1(32'hb9465007),
	.w2(32'hbab437b8),
	.w3(32'h3b24c9cc),
	.w4(32'h3a10559f),
	.w5(32'hbb8f65bb),
	.w6(32'hbac24330),
	.w7(32'hbb016c05),
	.w8(32'hbb429fa6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac385dd),
	.w1(32'h3a5b82fe),
	.w2(32'hbb9f5b1b),
	.w3(32'hbb2bb83e),
	.w4(32'hbb311623),
	.w5(32'hbae47c9b),
	.w6(32'hbaeba976),
	.w7(32'hbaaa101e),
	.w8(32'hbaa3b112),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6ca98),
	.w1(32'hbae98f7c),
	.w2(32'hbb8c90d1),
	.w3(32'hbaefb240),
	.w4(32'hbb39cf7d),
	.w5(32'hbadbdf91),
	.w6(32'hbacbb517),
	.w7(32'hbb25a7c3),
	.w8(32'hbaea1fa3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381f26a8),
	.w1(32'hbafc3ae6),
	.w2(32'h39d7bb00),
	.w3(32'hba38f2bb),
	.w4(32'hba2a3c51),
	.w5(32'hbab6f268),
	.w6(32'hbb0f2e53),
	.w7(32'h36f4aaad),
	.w8(32'h3a417bfe),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a620101),
	.w1(32'h3b38b67c),
	.w2(32'h39d47627),
	.w3(32'h3b78f81a),
	.w4(32'h3add7221),
	.w5(32'hb8f3059d),
	.w6(32'h3b9ee90c),
	.w7(32'h3b5347fc),
	.w8(32'hb78357f2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be912e),
	.w1(32'hb9f8a31e),
	.w2(32'h3a24349d),
	.w3(32'h39749fcd),
	.w4(32'hba0c1f21),
	.w5(32'h39017753),
	.w6(32'hba2b7aeb),
	.w7(32'hb9873aef),
	.w8(32'hb95b1850),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad752dd),
	.w1(32'hbba17ad6),
	.w2(32'hbb758125),
	.w3(32'hbb3be5f3),
	.w4(32'hbb27abb9),
	.w5(32'hbb522c07),
	.w6(32'hbbaa5afe),
	.w7(32'hbb2dfb6e),
	.w8(32'hbb02f7eb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa04ed6),
	.w1(32'hb9901ed6),
	.w2(32'hbbc21c2b),
	.w3(32'hbb2a08b6),
	.w4(32'h3a5f7b14),
	.w5(32'h3b55165a),
	.w6(32'hba347f9b),
	.w7(32'h395dfb9f),
	.w8(32'hbb3b494c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa3b5c),
	.w1(32'hba87cc0b),
	.w2(32'hbb101b83),
	.w3(32'h3b9148ae),
	.w4(32'h3b4bd53e),
	.w5(32'h3af69b20),
	.w6(32'hbb16a0d4),
	.w7(32'hbae1ceae),
	.w8(32'h39ae618f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812ad6a),
	.w1(32'h38b6c1d4),
	.w2(32'hbb2e937c),
	.w3(32'h3ae0e264),
	.w4(32'h3aa3b424),
	.w5(32'hbb451ac3),
	.w6(32'hba2d7566),
	.w7(32'hb9a1a17c),
	.w8(32'hbb7c4404),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0583d0),
	.w1(32'hbbc461eb),
	.w2(32'hbb4f71b5),
	.w3(32'hbc0e943e),
	.w4(32'hbb788b3e),
	.w5(32'h388e612c),
	.w6(32'hbc310db9),
	.w7(32'hbbb3a72c),
	.w8(32'hbad630c0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7a18c),
	.w1(32'h3b1a3bf2),
	.w2(32'h3b0a9497),
	.w3(32'h3aaeaa84),
	.w4(32'hbaa6c182),
	.w5(32'hba751632),
	.w6(32'h3a61ccc5),
	.w7(32'h3a71c250),
	.w8(32'hbae69cd8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558c82),
	.w1(32'hbb27986e),
	.w2(32'h3ab8018e),
	.w3(32'hbba60a40),
	.w4(32'h3aadf78a),
	.w5(32'hbb138ef3),
	.w6(32'hbb6bcef5),
	.w7(32'h3b2981df),
	.w8(32'hbbf86bd0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa909a9),
	.w1(32'h397c2e91),
	.w2(32'h3a820185),
	.w3(32'h3aceccd9),
	.w4(32'h3b0414fd),
	.w5(32'hbb03d125),
	.w6(32'h3910a726),
	.w7(32'h3ac93478),
	.w8(32'hbb0c3dbf),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7af79c),
	.w1(32'hbacec88a),
	.w2(32'h3ae814ca),
	.w3(32'hbb50b4f2),
	.w4(32'h3acc8582),
	.w5(32'hbb919d60),
	.w6(32'hbbbd2984),
	.w7(32'h3af22640),
	.w8(32'hbbf9773d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5417e8),
	.w1(32'hb9a73e97),
	.w2(32'hba3269f5),
	.w3(32'h3aca139b),
	.w4(32'h3b51c212),
	.w5(32'hbb5463f2),
	.w6(32'hba136a7e),
	.w7(32'h3b56b4e7),
	.w8(32'hbb74a60e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbbbbc),
	.w1(32'hbad4fd06),
	.w2(32'hbbe509c9),
	.w3(32'hba68f3ff),
	.w4(32'h38070708),
	.w5(32'hb9b4c236),
	.w6(32'hbadf000d),
	.w7(32'hbaab241b),
	.w8(32'hbaea65de),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb867a58d),
	.w1(32'h393acf82),
	.w2(32'hb9b838dc),
	.w3(32'h38a655fd),
	.w4(32'hb986aebf),
	.w5(32'h3afb70e7),
	.w6(32'hb9173e36),
	.w7(32'hb9b36122),
	.w8(32'hbb367dd6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ef590),
	.w1(32'hbb57e678),
	.w2(32'hbbd3abf0),
	.w3(32'hbb77517d),
	.w4(32'hbabdbdc6),
	.w5(32'hbbb50e85),
	.w6(32'hbb963b2f),
	.w7(32'hbb3f6acf),
	.w8(32'hbbdb245b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fb232),
	.w1(32'hbaff0c05),
	.w2(32'hbb5e6f93),
	.w3(32'hbae317a6),
	.w4(32'h398a9582),
	.w5(32'hbb1ba1cf),
	.w6(32'hbab108b0),
	.w7(32'hb90e490e),
	.w8(32'hbb863beb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e2a5c),
	.w1(32'hbacd7726),
	.w2(32'hbb983727),
	.w3(32'hba4b5ae1),
	.w4(32'hba9300b9),
	.w5(32'hbb9d02e9),
	.w6(32'h3a8d6e21),
	.w7(32'h3a447527),
	.w8(32'hbba266d1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9e404),
	.w1(32'hb99ce8e3),
	.w2(32'hbb17433a),
	.w3(32'hbb961b84),
	.w4(32'h3b501342),
	.w5(32'hba9f2a58),
	.w6(32'hbb975697),
	.w7(32'hb9c74c21),
	.w8(32'hbb8ff58a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab361b7),
	.w1(32'hb9a2eb4f),
	.w2(32'hbbb873ab),
	.w3(32'hb9b44432),
	.w4(32'hb81dac4d),
	.w5(32'hbb7867f4),
	.w6(32'hba43fc77),
	.w7(32'h3aa477aa),
	.w8(32'hbb7d3c04),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ae7bd),
	.w1(32'hbae45bd3),
	.w2(32'hbb7e12b2),
	.w3(32'hba9f208d),
	.w4(32'hbafec429),
	.w5(32'hbb8ad218),
	.w6(32'hb7172d69),
	.w7(32'hb8c40c78),
	.w8(32'hbb91296e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba287eda),
	.w1(32'h3a0c1449),
	.w2(32'hba65a62a),
	.w3(32'hb7320b6f),
	.w4(32'hb8f14701),
	.w5(32'hba04b0d0),
	.w6(32'h39eacd03),
	.w7(32'hb8b831a9),
	.w8(32'hbaccc827),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4562a),
	.w1(32'hbb95fdec),
	.w2(32'hbbef442c),
	.w3(32'hbaa779bf),
	.w4(32'hbb11df6a),
	.w5(32'hbbe7cfc2),
	.w6(32'hb90d0989),
	.w7(32'hb8c8e65f),
	.w8(32'hbb614c7c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72a0b2),
	.w1(32'hb9a43b13),
	.w2(32'hbb33bc72),
	.w3(32'hba00e3b1),
	.w4(32'h396e52b1),
	.w5(32'hbb530a22),
	.w6(32'h3a20197d),
	.w7(32'h3a8a6fb2),
	.w8(32'hbb1cb218),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a2834),
	.w1(32'hb9b2a6a1),
	.w2(32'hba76db4e),
	.w3(32'hba17fb8f),
	.w4(32'hba22a6b6),
	.w5(32'h38ace470),
	.w6(32'hbac1796a),
	.w7(32'hb9a40790),
	.w8(32'hba0b614d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cf46c),
	.w1(32'hba1d6fb5),
	.w2(32'hba023ad2),
	.w3(32'hb804b222),
	.w4(32'h39b1dd78),
	.w5(32'hbb01ae32),
	.w6(32'hba666ea8),
	.w7(32'hb8116684),
	.w8(32'hbb17ec36),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73ca56),
	.w1(32'hbb375706),
	.w2(32'hbb4bee47),
	.w3(32'hbb51d52f),
	.w4(32'hba8746e1),
	.w5(32'hbacf7a69),
	.w6(32'hbba5372f),
	.w7(32'hbb251706),
	.w8(32'hbb84b0a9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa46aea),
	.w1(32'hb9d8cc20),
	.w2(32'hbb4f95d9),
	.w3(32'h39be4115),
	.w4(32'h3afb77e0),
	.w5(32'hbafab096),
	.w6(32'hb9cb6fad),
	.w7(32'h3ae25af1),
	.w8(32'hbb0dcc83),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36159a),
	.w1(32'hb9847ae4),
	.w2(32'hbac7d79a),
	.w3(32'hbabfe784),
	.w4(32'hb7984971),
	.w5(32'hbaae289a),
	.w6(32'hbb0a992f),
	.w7(32'hbab8490b),
	.w8(32'hbb53502d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77c974),
	.w1(32'h38934b88),
	.w2(32'hbac68af9),
	.w3(32'hba41993c),
	.w4(32'h39d9098a),
	.w5(32'hba618acd),
	.w6(32'hba116e55),
	.w7(32'h3a24f2a7),
	.w8(32'hbab7b03b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d88946),
	.w1(32'h39c9c778),
	.w2(32'hb898dadf),
	.w3(32'hb9c1a879),
	.w4(32'h3a14393f),
	.w5(32'hba62ee5f),
	.w6(32'hba1a142d),
	.w7(32'hb99fae8b),
	.w8(32'hba38a7e2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba983c7a),
	.w1(32'hba3d1711),
	.w2(32'hbb344a6c),
	.w3(32'hba8b3a73),
	.w4(32'hba1b1687),
	.w5(32'hbaa2c1de),
	.w6(32'hba8a2bba),
	.w7(32'hb9566696),
	.w8(32'hba12a9f3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32159c),
	.w1(32'h3aec801a),
	.w2(32'hbae74e00),
	.w3(32'h39e60941),
	.w4(32'h3a76093e),
	.w5(32'hbac7a447),
	.w6(32'h39af5db3),
	.w7(32'h3a00b81a),
	.w8(32'hbb0550b0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7287916),
	.w1(32'hb80c2e75),
	.w2(32'h3a1b89b4),
	.w3(32'hb9c4155b),
	.w4(32'hb916001c),
	.w5(32'h39f5a507),
	.w6(32'hb9d469e5),
	.w7(32'h39967ba7),
	.w8(32'h39ac5dad),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3e57f),
	.w1(32'hb90a50ca),
	.w2(32'hb813776f),
	.w3(32'hb93896b0),
	.w4(32'hb998e6db),
	.w5(32'h38dc33e2),
	.w6(32'hb99632c4),
	.w7(32'h38a2f76f),
	.w8(32'hba0de500),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ec421b),
	.w1(32'hba2df01b),
	.w2(32'h3a0a4ff5),
	.w3(32'h3a0633f7),
	.w4(32'h395523de),
	.w5(32'hba143f64),
	.w6(32'hb9e61539),
	.w7(32'h39b2a2c2),
	.w8(32'hba4023c7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2c50b),
	.w1(32'hba4d80d8),
	.w2(32'hb936ab0d),
	.w3(32'hb9b7c24d),
	.w4(32'h39160911),
	.w5(32'hbb0506a8),
	.w6(32'hba7ab4ad),
	.w7(32'hb9976114),
	.w8(32'hbaf2e476),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39097f),
	.w1(32'hbad24a7c),
	.w2(32'hbb8ade10),
	.w3(32'hbb2013a9),
	.w4(32'h3a12b0ff),
	.w5(32'hbaf31582),
	.w6(32'hbba630e5),
	.w7(32'h39b42377),
	.w8(32'hba64d45f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77cb33),
	.w1(32'h3a1491b3),
	.w2(32'h389dcd52),
	.w3(32'h3a0def0f),
	.w4(32'h3500f3ae),
	.w5(32'hb9c36b3e),
	.w6(32'h39b4f32e),
	.w7(32'h39e29b31),
	.w8(32'hba967c81),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848b3e3),
	.w1(32'hba12d402),
	.w2(32'hbaab3ce4),
	.w3(32'h3a3491fa),
	.w4(32'hba537c68),
	.w5(32'hbb2817b3),
	.w6(32'h3a788deb),
	.w7(32'hb90fbbf0),
	.w8(32'hbb5014ee),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6329b2),
	.w1(32'hb932cebb),
	.w2(32'hba86137d),
	.w3(32'hbb3d4278),
	.w4(32'h39284c52),
	.w5(32'h3a36bf2d),
	.w6(32'hbb9de820),
	.w7(32'hbaaaf6a7),
	.w8(32'hbab6630b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e54685),
	.w1(32'h3a1573f5),
	.w2(32'h39cf18a9),
	.w3(32'h39f2bf98),
	.w4(32'hb765618a),
	.w5(32'h39605c7c),
	.w6(32'h3b083c9a),
	.w7(32'h38885789),
	.w8(32'hba1349d6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f5472b),
	.w1(32'hb9182f66),
	.w2(32'h38e9dfe8),
	.w3(32'h3a113733),
	.w4(32'h398f0954),
	.w5(32'h3a7228da),
	.w6(32'hb96f7f75),
	.w7(32'hb9d4c2b0),
	.w8(32'h3a4bcc74),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57c330),
	.w1(32'h3a86d479),
	.w2(32'h3a036aa7),
	.w3(32'h3a3f2318),
	.w4(32'h3a4fb6b0),
	.w5(32'h393a0d10),
	.w6(32'h3a8e521e),
	.w7(32'h3a01f304),
	.w8(32'hb95972f1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f398d5),
	.w1(32'hba6fac95),
	.w2(32'hba1eac8b),
	.w3(32'h3774c962),
	.w4(32'h39247d4d),
	.w5(32'hba350515),
	.w6(32'hb7c4733b),
	.w7(32'hb9f427e9),
	.w8(32'hba954670),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9e722),
	.w1(32'hbabb0d15),
	.w2(32'hbad44911),
	.w3(32'h38dd344d),
	.w4(32'hbafa8887),
	.w5(32'hbb1c61ba),
	.w6(32'hb91ae215),
	.w7(32'hba7672cf),
	.w8(32'hba93f0a1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa68dcd),
	.w1(32'hbaab7c21),
	.w2(32'hbb9360d3),
	.w3(32'h3a20ce8e),
	.w4(32'hba622e66),
	.w5(32'hbb8eebaf),
	.w6(32'h3a0259be),
	.w7(32'hb8b42d41),
	.w8(32'hbb954edc),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aef2ce),
	.w1(32'hb888d9b6),
	.w2(32'hb9e517c6),
	.w3(32'h394710ad),
	.w4(32'hb8a35460),
	.w5(32'h38d8f1e1),
	.w6(32'h3a73236f),
	.w7(32'hb95c87d1),
	.w8(32'hb9955182),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6fb68),
	.w1(32'hb9d8a87d),
	.w2(32'hba434fdd),
	.w3(32'hbb101589),
	.w4(32'hba8a5605),
	.w5(32'hba650a94),
	.w6(32'hbb1ccc93),
	.w7(32'hba784093),
	.w8(32'hbaf0cad8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7148b2),
	.w1(32'h390c89cd),
	.w2(32'hba337bd7),
	.w3(32'hba1e5a94),
	.w4(32'hb9c72149),
	.w5(32'hba990540),
	.w6(32'hbaceaf74),
	.w7(32'hb977a2ac),
	.w8(32'hbb2f98be),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb193082),
	.w1(32'hba4388df),
	.w2(32'hbaaad724),
	.w3(32'hbaaf4c3b),
	.w4(32'hba3e6b9e),
	.w5(32'hba4eefbc),
	.w6(32'hbb07e910),
	.w7(32'hbaac6610),
	.w8(32'hbae51efe),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b59fb),
	.w1(32'hba819f72),
	.w2(32'hbb32ce9e),
	.w3(32'hba43b866),
	.w4(32'h3a68abf7),
	.w5(32'hba890a96),
	.w6(32'hba22b933),
	.w7(32'h39dc60d6),
	.w8(32'hbac21699),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa86104),
	.w1(32'hba9aadd4),
	.w2(32'hbb882995),
	.w3(32'hba9f1574),
	.w4(32'hbb16aa25),
	.w5(32'hbb3b53ba),
	.w6(32'hb98b6709),
	.w7(32'hbaa73415),
	.w8(32'hbb93cbbb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae67b23),
	.w1(32'h3a02f15c),
	.w2(32'hba0ba5c5),
	.w3(32'hba72c46a),
	.w4(32'h3969ef60),
	.w5(32'hb9c8f9a3),
	.w6(32'hbaa7c289),
	.w7(32'h3a457d30),
	.w8(32'hbaef31f8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb1aa1),
	.w1(32'hbb022176),
	.w2(32'hbb5142f9),
	.w3(32'hb94d508b),
	.w4(32'hb8561fff),
	.w5(32'hbb04ed01),
	.w6(32'hb8855aad),
	.w7(32'hb79f2710),
	.w8(32'hbb168adf),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b269f),
	.w1(32'hbad44ed8),
	.w2(32'hbb51528c),
	.w3(32'hbad32d2d),
	.w4(32'hbac57fa4),
	.w5(32'hbb672e6e),
	.w6(32'hba8db533),
	.w7(32'hba64be84),
	.w8(32'hbb801ecd),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb064a0b),
	.w1(32'hba1e2236),
	.w2(32'hbaecc8d7),
	.w3(32'hba6ac420),
	.w4(32'hb9a72f10),
	.w5(32'hbad2ec5a),
	.w6(32'hba467b17),
	.w7(32'h39305b17),
	.w8(32'hbb048b62),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2c113),
	.w1(32'hba20e5a2),
	.w2(32'hbb32f8b1),
	.w3(32'hba3c9bd9),
	.w4(32'hba3a3b96),
	.w5(32'hba77cf4a),
	.w6(32'hbadbadb5),
	.w7(32'hba04520e),
	.w8(32'hbaf1d5e1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5df3dc9),
	.w1(32'h3a0099b1),
	.w2(32'hb96d647b),
	.w3(32'h39fb0105),
	.w4(32'h3a223e72),
	.w5(32'hb9910b91),
	.w6(32'hba15e51f),
	.w7(32'h39c238fa),
	.w8(32'hba7155ee),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8549b),
	.w1(32'h3b06d145),
	.w2(32'hba929b9d),
	.w3(32'hba9c21d6),
	.w4(32'h3ad6d798),
	.w5(32'hbad3504c),
	.w6(32'hba81b333),
	.w7(32'h3aa183ba),
	.w8(32'hbb74b913),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac35318),
	.w1(32'hba2d04a6),
	.w2(32'hba7ce470),
	.w3(32'hba8c5206),
	.w4(32'hb9fc473b),
	.w5(32'hbabc18e6),
	.w6(32'hbb102347),
	.w7(32'hba6ec1ef),
	.w8(32'hbb186e00),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e1bb6),
	.w1(32'hba717c01),
	.w2(32'hb9b68650),
	.w3(32'hb9dc0882),
	.w4(32'h3983df6d),
	.w5(32'h3a3cce4a),
	.w6(32'hba06d988),
	.w7(32'h37c29803),
	.w8(32'hb994d7db),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a380cb5),
	.w1(32'hb9f6678e),
	.w2(32'hb910bbf7),
	.w3(32'h3a356f6e),
	.w4(32'h3a6e8656),
	.w5(32'h3a24f45d),
	.w6(32'h39523972),
	.w7(32'h38efd522),
	.w8(32'h3a0fa28e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f78852),
	.w1(32'h39cc4488),
	.w2(32'hb9c14ef9),
	.w3(32'hb953d27c),
	.w4(32'h3a117694),
	.w5(32'hba3dd1ba),
	.w6(32'hb9ad4fc8),
	.w7(32'h39af1746),
	.w8(32'hba96fb39),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a9fd3),
	.w1(32'hba92b241),
	.w2(32'hbb603218),
	.w3(32'hba7a07ad),
	.w4(32'h391f165c),
	.w5(32'hbb128710),
	.w6(32'hbab1e642),
	.w7(32'h38cdbd4d),
	.w8(32'hbb27a7b9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d22e5),
	.w1(32'hbabec303),
	.w2(32'hbb3f8704),
	.w3(32'hbaf52650),
	.w4(32'hb89efb56),
	.w5(32'hbb7eb6a6),
	.w6(32'hba06e926),
	.w7(32'hb9905264),
	.w8(32'hbbb13988),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eae22e),
	.w1(32'hb9b51073),
	.w2(32'h38fa1bc5),
	.w3(32'hba647551),
	.w4(32'h39ca3c05),
	.w5(32'h3a2d681f),
	.w6(32'hb952cec6),
	.w7(32'h3a1a47ec),
	.w8(32'h39c5e93b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05417c),
	.w1(32'hba7509b1),
	.w2(32'hbb937e0e),
	.w3(32'hb8a7a721),
	.w4(32'h38d77ea9),
	.w5(32'hbb53ca8b),
	.w6(32'hba6361cf),
	.w7(32'hb8fca441),
	.w8(32'hbb6e788a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9205c),
	.w1(32'hb9b0fc4c),
	.w2(32'hbb0d064c),
	.w3(32'hba02695d),
	.w4(32'h392c6e06),
	.w5(32'hbb2baa1a),
	.w6(32'hba0005b8),
	.w7(32'h3a680abd),
	.w8(32'hbb4a6e22),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb466701),
	.w1(32'hbb29d5e0),
	.w2(32'hbb95ec1d),
	.w3(32'hba9789bc),
	.w4(32'hbb36ac2c),
	.w5(32'hbb1e8d3a),
	.w6(32'hba03f1f8),
	.w7(32'hbad8ea0b),
	.w8(32'hbb28f386),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13d942),
	.w1(32'h3b2eb7b1),
	.w2(32'hbb387708),
	.w3(32'h3b179b05),
	.w4(32'h3b719093),
	.w5(32'hbb12159b),
	.w6(32'h3a08f22b),
	.w7(32'h3b5ae691),
	.w8(32'hbb24e017),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71c874),
	.w1(32'hba3e4268),
	.w2(32'hba2d1f59),
	.w3(32'hba94bef6),
	.w4(32'hb72b14a2),
	.w5(32'hba428256),
	.w6(32'hbb205164),
	.w7(32'hba7e3f93),
	.w8(32'hbaffba95),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f4217),
	.w1(32'hba82a3f2),
	.w2(32'hb94bf77d),
	.w3(32'hba23371c),
	.w4(32'h3a5930bf),
	.w5(32'h3a8053bf),
	.w6(32'hba4f2ddb),
	.w7(32'hba0d6844),
	.w8(32'h39eb2504),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba789a71),
	.w1(32'h3a02f978),
	.w2(32'hba8485cc),
	.w3(32'h377ae6f3),
	.w4(32'h3b291fa5),
	.w5(32'h39922a2d),
	.w6(32'hbae41564),
	.w7(32'h3a963a3c),
	.w8(32'hba1b28ba),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a888b),
	.w1(32'h39ecec51),
	.w2(32'hba4e850f),
	.w3(32'hbabf8d94),
	.w4(32'h3a738159),
	.w5(32'hba7e25bb),
	.w6(32'hba673f85),
	.w7(32'h399ae477),
	.w8(32'hbb44b922),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b207b1),
	.w1(32'h3b07de6b),
	.w2(32'h3a1fea3e),
	.w3(32'h3a5824c1),
	.w4(32'h3ae423f5),
	.w5(32'h387b1713),
	.w6(32'hb8e24b03),
	.w7(32'h3aae294b),
	.w8(32'hb885ac25),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1d593),
	.w1(32'hba9d485c),
	.w2(32'hba07f681),
	.w3(32'hbb1b2b9d),
	.w4(32'hbb247f63),
	.w5(32'hb9c4fb1c),
	.w6(32'hba97e9de),
	.w7(32'hba5c79c7),
	.w8(32'h39e4873e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39998d4e),
	.w1(32'h3a661652),
	.w2(32'h399b5aba),
	.w3(32'h39fb608c),
	.w4(32'hb9d4dde7),
	.w5(32'hb981caa0),
	.w6(32'h3ab2de75),
	.w7(32'h3a2d3c1f),
	.w8(32'hb748b89c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eecc3),
	.w1(32'hba4806f3),
	.w2(32'hbaf1d01f),
	.w3(32'hb9e57f5b),
	.w4(32'hba0264a8),
	.w5(32'hbb0f68eb),
	.w6(32'hba985b59),
	.w7(32'h38ac5019),
	.w8(32'hbb2edef5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f5e4fb),
	.w1(32'h3a1ec786),
	.w2(32'h390e7d59),
	.w3(32'h3a23d57c),
	.w4(32'h3a1006d4),
	.w5(32'h39cb4a35),
	.w6(32'h38b54c14),
	.w7(32'h3a30f35f),
	.w8(32'h3a344709),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed6aea),
	.w1(32'h3a711d7b),
	.w2(32'h39518adc),
	.w3(32'h39cebbd6),
	.w4(32'h3ad115f9),
	.w5(32'hbabb947f),
	.w6(32'h38c9b12a),
	.w7(32'h3b059bea),
	.w8(32'hba90a674),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4148f),
	.w1(32'h39bd3587),
	.w2(32'h39e9d4b1),
	.w3(32'hb94946db),
	.w4(32'h393f8cb7),
	.w5(32'hba0644b7),
	.w6(32'h38db2b99),
	.w7(32'h39ad2444),
	.w8(32'hb9d45d01),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09d7cd),
	.w1(32'h3aa56498),
	.w2(32'h37c9669c),
	.w3(32'hba147f66),
	.w4(32'h3a159559),
	.w5(32'hb9e064c2),
	.w6(32'h397cdca3),
	.w7(32'h396d01b8),
	.w8(32'hba655c19),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a01b73),
	.w1(32'hba02f0f3),
	.w2(32'hb8cb49b9),
	.w3(32'h39259831),
	.w4(32'h39fc1a30),
	.w5(32'h39b3f2bc),
	.w6(32'h3a19c31f),
	.w7(32'h39b88707),
	.w8(32'h3996d172),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9861772),
	.w1(32'hba507aed),
	.w2(32'hb994c715),
	.w3(32'hba37a3f1),
	.w4(32'hb95c14cd),
	.w5(32'hba523670),
	.w6(32'h3aad237c),
	.w7(32'h3a5e774e),
	.w8(32'hba13146f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb257bcd),
	.w1(32'hba6eb1e1),
	.w2(32'hbb5776cd),
	.w3(32'hba696866),
	.w4(32'h398cdffe),
	.w5(32'hba1d84fd),
	.w6(32'hbace9ddf),
	.w7(32'hbaadda86),
	.w8(32'hbb0478df),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c2df0),
	.w1(32'hba2efa84),
	.w2(32'hbbab9075),
	.w3(32'hba9efea8),
	.w4(32'hbb2c3697),
	.w5(32'hbbf051e1),
	.w6(32'hba84f8db),
	.w7(32'h3a205ece),
	.w8(32'hbba2335d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a65445),
	.w1(32'h39b92af9),
	.w2(32'h39ccd5a6),
	.w3(32'hb97024c7),
	.w4(32'h3a41c815),
	.w5(32'hb8b522b2),
	.w6(32'hbaa8e78b),
	.w7(32'h39415beb),
	.w8(32'h393d61da),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa56bd),
	.w1(32'hb9bbcadb),
	.w2(32'hbb14e47b),
	.w3(32'hba8b06c9),
	.w4(32'h39b41874),
	.w5(32'hbb1138ec),
	.w6(32'hbad85efc),
	.w7(32'h39c2e5fb),
	.w8(32'hbb68478e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924dddb),
	.w1(32'hba6e595d),
	.w2(32'hb9ed483f),
	.w3(32'hb9ed7e04),
	.w4(32'h3a334fe5),
	.w5(32'hbac10e25),
	.w6(32'hb9b40b1b),
	.w7(32'hb8623339),
	.w8(32'hbac2efc0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb71d88),
	.w1(32'hbb311800),
	.w2(32'hbc15369d),
	.w3(32'hbb8a5ec7),
	.w4(32'hba42b12f),
	.w5(32'hbbb767b8),
	.w6(32'hbb8f7f32),
	.w7(32'hbaabf561),
	.w8(32'hbbe08444),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd40c4),
	.w1(32'hb8108194),
	.w2(32'hbb0a8bdb),
	.w3(32'hba990140),
	.w4(32'h3a96b4e4),
	.w5(32'hbb3b3875),
	.w6(32'hbaa9f285),
	.w7(32'h3a828923),
	.w8(32'hbb7a7928),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29f226),
	.w1(32'hbb2e9b8b),
	.w2(32'hbbd1838b),
	.w3(32'hbac52e1b),
	.w4(32'hbaad0b09),
	.w5(32'hbb626874),
	.w6(32'hbac6278b),
	.w7(32'hba371aa0),
	.w8(32'hbb3dc77b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eb975),
	.w1(32'h39ac2ef2),
	.w2(32'h397ac843),
	.w3(32'h3a219d19),
	.w4(32'h38bb780f),
	.w5(32'hb972c94c),
	.w6(32'h3a7535bd),
	.w7(32'h3980d230),
	.w8(32'hb9f7cdc0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03e031),
	.w1(32'hba63c4cd),
	.w2(32'hbb4c2859),
	.w3(32'hba59281e),
	.w4(32'hba776999),
	.w5(32'hbac09549),
	.w6(32'hba5ccb13),
	.w7(32'hb96c752a),
	.w8(32'hbaa35ee3),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb854deb8),
	.w1(32'hb9485121),
	.w2(32'hb9a6842b),
	.w3(32'h39129e10),
	.w4(32'h398ee1b7),
	.w5(32'hba4ca213),
	.w6(32'hb94c501d),
	.w7(32'h38069af2),
	.w8(32'hba32a43d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f298f9),
	.w1(32'hba4abd42),
	.w2(32'hbaa78583),
	.w3(32'h395cfb2f),
	.w4(32'h39088956),
	.w5(32'hb90eb7c8),
	.w6(32'hba0ee945),
	.w7(32'hb9ffa064),
	.w8(32'h38c28504),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398da747),
	.w1(32'h3a468915),
	.w2(32'h391d6a25),
	.w3(32'h38023c87),
	.w4(32'hb794f73b),
	.w5(32'hb838feef),
	.w6(32'hb9aa8a40),
	.w7(32'hb91ad537),
	.w8(32'hba331e0b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c0334),
	.w1(32'hba9294df),
	.w2(32'hbb328b7c),
	.w3(32'hbabecb73),
	.w4(32'hba8b6ffa),
	.w5(32'hbae5fb01),
	.w6(32'hbb105ffe),
	.w7(32'hbab1580d),
	.w8(32'hbb838d6d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f3c60),
	.w1(32'hb92f16ce),
	.w2(32'hba464fce),
	.w3(32'h399cb5d3),
	.w4(32'h385a5578),
	.w5(32'hb9e18d7d),
	.w6(32'hb97d24ae),
	.w7(32'hb9f900e9),
	.w8(32'hb99ba590),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e868f),
	.w1(32'hb99c7c15),
	.w2(32'hba2950ba),
	.w3(32'hb998b16a),
	.w4(32'h39347dbf),
	.w5(32'h38998017),
	.w6(32'h39021d5b),
	.w7(32'hb93e8b71),
	.w8(32'hb9a0128c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba399c8d),
	.w1(32'h3a26c92b),
	.w2(32'h398a2b48),
	.w3(32'h38b7fcc8),
	.w4(32'h3a87943a),
	.w5(32'h3a8622c0),
	.w6(32'hb9bec46a),
	.w7(32'h3a1c721d),
	.w8(32'h39fc58bc),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21cd3f),
	.w1(32'hb9a0f837),
	.w2(32'hbaaa67d5),
	.w3(32'hba1a0e9b),
	.w4(32'hb920d729),
	.w5(32'hbabe328a),
	.w6(32'hba374e3a),
	.w7(32'hb9ccb51d),
	.w8(32'hbb398d15),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac16aad),
	.w1(32'hba9ca6fb),
	.w2(32'hbaed8c3d),
	.w3(32'hba9b8db6),
	.w4(32'hba85a711),
	.w5(32'hb99f8705),
	.w6(32'hb95ce6c5),
	.w7(32'h3a1b6c9e),
	.w8(32'hba28d59d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5c00d),
	.w1(32'hba20b1da),
	.w2(32'hbaa736ff),
	.w3(32'hba4e38b6),
	.w4(32'hb9d0a67f),
	.w5(32'hb94cf0b9),
	.w6(32'hba5c4e0d),
	.w7(32'hb9877cf6),
	.w8(32'hba81c698),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc489f9),
	.w1(32'hbb5c5ea0),
	.w2(32'hbc288358),
	.w3(32'hbb6b6b37),
	.w4(32'hbae07b22),
	.w5(32'hbbee6d52),
	.w6(32'h3b0c7303),
	.w7(32'h39d43115),
	.w8(32'hbbcf914c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8063f9),
	.w1(32'hbabc4fee),
	.w2(32'hbb623f9f),
	.w3(32'hbb5c03e7),
	.w4(32'h3aad36ce),
	.w5(32'hb88d4538),
	.w6(32'hbb2ce170),
	.w7(32'h3a34fccd),
	.w8(32'hbb34e4ca),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928cb50),
	.w1(32'hba4f85f1),
	.w2(32'hb9d2ba67),
	.w3(32'h39bf58f2),
	.w4(32'hb984a74f),
	.w5(32'hba20c086),
	.w6(32'h39fce150),
	.w7(32'hb94a22fe),
	.w8(32'hb904ee44),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d955b6),
	.w1(32'hb7f3cc4d),
	.w2(32'h39cdf481),
	.w3(32'hb9058152),
	.w4(32'h3a085bc8),
	.w5(32'h38df1cb5),
	.w6(32'hb95d9234),
	.w7(32'h38e0a075),
	.w8(32'hb892e592),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac0875),
	.w1(32'h39bc7c1a),
	.w2(32'h39823141),
	.w3(32'h390b3f83),
	.w4(32'h3a48c779),
	.w5(32'hb895e283),
	.w6(32'hb868b94d),
	.w7(32'h3a569427),
	.w8(32'h3939ec36),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0fc9c),
	.w1(32'h3a0b3532),
	.w2(32'h3a06c773),
	.w3(32'h39b06b73),
	.w4(32'h39cb4b94),
	.w5(32'hba8df76b),
	.w6(32'h38e0a805),
	.w7(32'h3a69e287),
	.w8(32'hb9b00677),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952b4e2),
	.w1(32'hbaa7a628),
	.w2(32'hbab8bb54),
	.w3(32'hba39d789),
	.w4(32'hbaf0c747),
	.w5(32'hbaa01af8),
	.w6(32'hb9a380a6),
	.w7(32'hba9b499b),
	.w8(32'hbad6d6dd),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f3961),
	.w1(32'hba1c3ef6),
	.w2(32'hbb3af5eb),
	.w3(32'hbaddc303),
	.w4(32'hbb055786),
	.w5(32'hbb91002b),
	.w6(32'hba4f4d96),
	.w7(32'hba0ba4e4),
	.w8(32'hbb984058),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37456f),
	.w1(32'hbb29b0e4),
	.w2(32'hbb8affb1),
	.w3(32'hbb4ff198),
	.w4(32'hb9c94a73),
	.w5(32'hbb58d9a5),
	.w6(32'hbb58b91c),
	.w7(32'hba9457b9),
	.w8(32'hbb8e89eb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92d3ce),
	.w1(32'hba13233c),
	.w2(32'hb9bc748e),
	.w3(32'hbaaedebd),
	.w4(32'h39ea4170),
	.w5(32'hb99865ce),
	.w6(32'hba9ee672),
	.w7(32'h39d4daea),
	.w8(32'hb9b59514),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c4b63),
	.w1(32'hbad2ea18),
	.w2(32'hbb8539bf),
	.w3(32'hbac41ee5),
	.w4(32'hb9f8435a),
	.w5(32'hbb6736ae),
	.w6(32'hbab480a9),
	.w7(32'hba823d00),
	.w8(32'hbb9903ff),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba804b21),
	.w1(32'hbad1f1c8),
	.w2(32'hba90d6d0),
	.w3(32'hba7ba578),
	.w4(32'hba3949a2),
	.w5(32'hba554439),
	.w6(32'hbb096efa),
	.w7(32'hba922e94),
	.w8(32'hba728ec1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a285671),
	.w1(32'hb919ec78),
	.w2(32'h3a06ff16),
	.w3(32'hb9b634b1),
	.w4(32'hb9d87486),
	.w5(32'hb98ee714),
	.w6(32'hb94eaad2),
	.w7(32'h399fc1af),
	.w8(32'h3a96c26f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad413b),
	.w1(32'hb8a27e7a),
	.w2(32'h38c081e0),
	.w3(32'hbad08c98),
	.w4(32'hba35e1ae),
	.w5(32'h399f5087),
	.w6(32'h3a40f33f),
	.w7(32'h3a3de04f),
	.w8(32'h39a9e2fa),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b33d0),
	.w1(32'h3a30b0fd),
	.w2(32'h3a6b1766),
	.w3(32'h39faf333),
	.w4(32'h39d03018),
	.w5(32'h398bb79a),
	.w6(32'h3a91579a),
	.w7(32'h3a751fc0),
	.w8(32'h394bd41e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52dd7e),
	.w1(32'h3a601621),
	.w2(32'h396a228f),
	.w3(32'h39ead836),
	.w4(32'h3ac172cc),
	.w5(32'h393d5c79),
	.w6(32'h37f542d7),
	.w7(32'h39e6795d),
	.w8(32'hb9dcf900),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04b65f),
	.w1(32'h3aedcc2b),
	.w2(32'hba4eddbc),
	.w3(32'hbacc5271),
	.w4(32'h3b116262),
	.w5(32'hba002cd8),
	.w6(32'hbb126738),
	.w7(32'h3a9f1c11),
	.w8(32'hbaceac64),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01316b),
	.w1(32'hb86366cc),
	.w2(32'hbb214107),
	.w3(32'hba761e90),
	.w4(32'h39e81a73),
	.w5(32'hbb0a79fb),
	.w6(32'hbaae7f46),
	.w7(32'h3a89b7d8),
	.w8(32'hbb368eab),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab5151),
	.w1(32'hba203e6d),
	.w2(32'hb8feddee),
	.w3(32'hba85a454),
	.w4(32'h39439f4a),
	.w5(32'hb9c85260),
	.w6(32'hbb073b2d),
	.w7(32'hba582d1f),
	.w8(32'hba6a23fb),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb276f6b),
	.w1(32'h369fe2fa),
	.w2(32'hbb2469f4),
	.w3(32'hbad74e98),
	.w4(32'h39ca1789),
	.w5(32'hbab9e299),
	.w6(32'hbb2c2616),
	.w7(32'hb9ba9e07),
	.w8(32'hbb67bf7f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9a7cf),
	.w1(32'hba860a40),
	.w2(32'hbb1a6de6),
	.w3(32'hbac6cc75),
	.w4(32'hb9ec5ac0),
	.w5(32'hbae4408a),
	.w6(32'hba88ea79),
	.w7(32'hba1082a7),
	.w8(32'hbb37e4ad),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb976af4),
	.w1(32'hbaacdcb2),
	.w2(32'hbbb8d0c4),
	.w3(32'hbb25a70c),
	.w4(32'hba820ae4),
	.w5(32'hbb90b36e),
	.w6(32'hbaf3484a),
	.w7(32'hb95ed1cb),
	.w8(32'hbba0f1a1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25e771),
	.w1(32'h3a3f2213),
	.w2(32'h3a28ea95),
	.w3(32'hb7fe71e6),
	.w4(32'h394a85b8),
	.w5(32'h38e1f006),
	.w6(32'hb6a3e3f4),
	.w7(32'h38ee9fae),
	.w8(32'h39ae8b59),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387713a0),
	.w1(32'h399ea97a),
	.w2(32'h3a183f5e),
	.w3(32'h385abca3),
	.w4(32'h39296da5),
	.w5(32'hba26df39),
	.w6(32'hb8fc2421),
	.w7(32'h3a6b9293),
	.w8(32'hb9f98145),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12e7c4),
	.w1(32'h38478479),
	.w2(32'hbb3e9b91),
	.w3(32'hba2326ad),
	.w4(32'hb8e83a0d),
	.w5(32'hbb601c4c),
	.w6(32'h39ef8ca5),
	.w7(32'h38c97510),
	.w8(32'hbb3d8b77),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba902268),
	.w1(32'h3a932f7b),
	.w2(32'hbb85aa70),
	.w3(32'hb990f877),
	.w4(32'hb97013fd),
	.w5(32'hbbc061a2),
	.w6(32'hba7c3c2c),
	.w7(32'h3ac10e26),
	.w8(32'hbb516feb),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0082dc),
	.w1(32'hba41db96),
	.w2(32'hbb61cdf0),
	.w3(32'hb9b80ba8),
	.w4(32'h3a5442ba),
	.w5(32'hbb0fab00),
	.w6(32'hb9679972),
	.w7(32'h3b0640e8),
	.w8(32'hbb59eba9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d6fb9),
	.w1(32'hba6697a2),
	.w2(32'hba703eb6),
	.w3(32'hbaa7a794),
	.w4(32'hbac2c952),
	.w5(32'h39c86b04),
	.w6(32'hb9949900),
	.w7(32'hbabd108d),
	.w8(32'hba15d40e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38761d11),
	.w1(32'hb89627ba),
	.w2(32'hb818e89b),
	.w3(32'hb80e7dc8),
	.w4(32'h397a52dd),
	.w5(32'h3924ec0d),
	.w6(32'h39dac7e3),
	.w7(32'h3931789a),
	.w8(32'hb9bb39a9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9861ead),
	.w1(32'hba5aa32b),
	.w2(32'hba0266e0),
	.w3(32'hb988fb1a),
	.w4(32'hb9bd37c7),
	.w5(32'h3a0c5970),
	.w6(32'hb9ce8441),
	.w7(32'hba20b3c8),
	.w8(32'hb94f45a5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a350f1c),
	.w1(32'h39a4a2aa),
	.w2(32'hbb34d60d),
	.w3(32'h3a8c9f40),
	.w4(32'hbb5c266a),
	.w5(32'hbba35020),
	.w6(32'h3a9e4bb2),
	.w7(32'hbaf34cc7),
	.w8(32'hbb869481),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98a852),
	.w1(32'hbad22dec),
	.w2(32'hbb89fd52),
	.w3(32'hbb5539a0),
	.w4(32'hbb12327e),
	.w5(32'hbb9f4c5d),
	.w6(32'hbae10d80),
	.w7(32'hba6aa99e),
	.w8(32'hbb9407e6),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6784ec),
	.w1(32'hba9438a8),
	.w2(32'hbaac2cc7),
	.w3(32'h3966eca9),
	.w4(32'hba68f7c2),
	.w5(32'hbb2ec709),
	.w6(32'hb952eef8),
	.w7(32'hbad56335),
	.w8(32'hbb874a93),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba804543),
	.w1(32'h39ecbaab),
	.w2(32'hbabcf486),
	.w3(32'hba847e6b),
	.w4(32'h3a98b76a),
	.w5(32'hb9e490d9),
	.w6(32'hbb1056d4),
	.w7(32'hb7bfd2fc),
	.w8(32'hbacfca62),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa30d45),
	.w1(32'hba5beb73),
	.w2(32'hbb35db74),
	.w3(32'hbabfaba8),
	.w4(32'h3b06a729),
	.w5(32'hb9cd147f),
	.w6(32'hbb219ff0),
	.w7(32'h3a99c003),
	.w8(32'hba839422),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3899a),
	.w1(32'h3989d64b),
	.w2(32'h39e7bfd8),
	.w3(32'h39c36139),
	.w4(32'h3a04cc0b),
	.w5(32'h38f7f45d),
	.w6(32'h3a77a9eb),
	.w7(32'h3a8b9730),
	.w8(32'h38e90af1),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96081b8),
	.w1(32'hba78b010),
	.w2(32'hba08276d),
	.w3(32'h39f5f628),
	.w4(32'h3a40e14c),
	.w5(32'hba3a02b6),
	.w6(32'h394c6671),
	.w7(32'h38e36608),
	.w8(32'hb9983d58),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba192bc9),
	.w1(32'hb9630b93),
	.w2(32'hba4ec30e),
	.w3(32'hb9bb38f7),
	.w4(32'hba7759db),
	.w5(32'hb9596b3f),
	.w6(32'h3999b38a),
	.w7(32'hba809770),
	.w8(32'h3911ad29),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9672f59),
	.w1(32'hb919bd62),
	.w2(32'h39d08db7),
	.w3(32'hb93b1ef3),
	.w4(32'hba4499e9),
	.w5(32'h3aa7f20c),
	.w6(32'hb9dad44f),
	.w7(32'h3a15df9b),
	.w8(32'h3b1b59ca),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3e860),
	.w1(32'h3c18326e),
	.w2(32'h3bd04c07),
	.w3(32'h3bd4b784),
	.w4(32'h3bd6578c),
	.w5(32'h3aa4e1e2),
	.w6(32'h3c0ed076),
	.w7(32'h3bf18ffc),
	.w8(32'hbb3fed8e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47087f),
	.w1(32'hbc03423d),
	.w2(32'hbb7d9f86),
	.w3(32'hbb46493f),
	.w4(32'hbb0a0af9),
	.w5(32'hbc16f363),
	.w6(32'hbb8c921b),
	.w7(32'hbbf7708d),
	.w8(32'hbb3b8ff6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61865b),
	.w1(32'h3be01ebd),
	.w2(32'hbbe978c2),
	.w3(32'hbbac1066),
	.w4(32'hbada7db7),
	.w5(32'hbc05b64e),
	.w6(32'h3bee22c9),
	.w7(32'hb9c0f47a),
	.w8(32'hbc2c1b2f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe66614),
	.w1(32'h39056297),
	.w2(32'hba9c0162),
	.w3(32'hbb91c174),
	.w4(32'h3900cc62),
	.w5(32'h39547e66),
	.w6(32'hbada78b2),
	.w7(32'h3ad6e4d6),
	.w8(32'h3affb4fb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a6797),
	.w1(32'h39b7c0f2),
	.w2(32'hbbb9b3e7),
	.w3(32'hbba726e0),
	.w4(32'hbac3c55a),
	.w5(32'hbbd39716),
	.w6(32'hbaf21e51),
	.w7(32'h3a81da4a),
	.w8(32'hbbb8b1c1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62c87a),
	.w1(32'hbb3de896),
	.w2(32'hbc00ec92),
	.w3(32'hbbf18029),
	.w4(32'hbbb57c98),
	.w5(32'hbbeaf65d),
	.w6(32'hbb07094b),
	.w7(32'hbb69cc86),
	.w8(32'hbb69f345),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cced8),
	.w1(32'h3c103f72),
	.w2(32'h3b9ea9c8),
	.w3(32'h3bcfeb82),
	.w4(32'h3b43a43f),
	.w5(32'h3b85a97e),
	.w6(32'hbbd9a10e),
	.w7(32'hbbfc727e),
	.w8(32'h3ae5db4a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb044519),
	.w1(32'h3ae7bf11),
	.w2(32'hba1ba9ec),
	.w3(32'h3bb5c86a),
	.w4(32'h3aa6088f),
	.w5(32'hbc429506),
	.w6(32'h3ac196e1),
	.w7(32'h38b4d78b),
	.w8(32'hbbb3c4cb),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc089598),
	.w1(32'hbb54ee52),
	.w2(32'hb909f96e),
	.w3(32'hbbe26afb),
	.w4(32'hbad9b35a),
	.w5(32'hbbbe5b1a),
	.w6(32'hbc3d8a24),
	.w7(32'h3a7cf501),
	.w8(32'hb9a76a5e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf57c6),
	.w1(32'hbc32f225),
	.w2(32'hbb7cf4bb),
	.w3(32'hbb402c4c),
	.w4(32'h3b918f13),
	.w5(32'h3af5c528),
	.w6(32'h3ac25429),
	.w7(32'hbb5b1d1b),
	.w8(32'hba601efd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cdbed),
	.w1(32'h3ba44a76),
	.w2(32'h3a7db0fb),
	.w3(32'h3b87cfe5),
	.w4(32'h3bc6fc6d),
	.w5(32'h3b1bdd85),
	.w6(32'h3b79807f),
	.w7(32'h3b5a1e99),
	.w8(32'h3b8f4a16),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66ce0b),
	.w1(32'h3b5d40f0),
	.w2(32'hbb820f76),
	.w3(32'h3c19664b),
	.w4(32'h3c365086),
	.w5(32'h3b5bd825),
	.w6(32'h3c6f06e4),
	.w7(32'h3bb283cd),
	.w8(32'hb9b5de2f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23b314),
	.w1(32'h3bb30286),
	.w2(32'h3ab1d4f9),
	.w3(32'h3b10faec),
	.w4(32'h3a980897),
	.w5(32'hbad5a982),
	.w6(32'h3c0c85e2),
	.w7(32'hba236e21),
	.w8(32'h3941b6f0),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10de88),
	.w1(32'hb7569f15),
	.w2(32'hbb0a1d80),
	.w3(32'h39571431),
	.w4(32'h3a105cce),
	.w5(32'h3b903a35),
	.w6(32'h3af7f6a4),
	.w7(32'h3acbd697),
	.w8(32'h3b770960),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d03f9),
	.w1(32'h3c49e537),
	.w2(32'hbaa2ec5b),
	.w3(32'h3c29732b),
	.w4(32'h3abf34ef),
	.w5(32'hba43cee1),
	.w6(32'hbb05a1cc),
	.w7(32'hbaf6711e),
	.w8(32'hbb240cef),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0017de),
	.w1(32'hbc06e8b2),
	.w2(32'hbb610e96),
	.w3(32'h3ad87780),
	.w4(32'hba83d6f2),
	.w5(32'h3b08a3e4),
	.w6(32'hbaba2354),
	.w7(32'h3af48672),
	.w8(32'hbb28a304),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268d6f),
	.w1(32'hbbfad58b),
	.w2(32'hbb95952e),
	.w3(32'h3b549050),
	.w4(32'hbbded3e8),
	.w5(32'h3ae49377),
	.w6(32'hba8a8c40),
	.w7(32'hbc1716ca),
	.w8(32'hbad368f2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb968df0),
	.w1(32'hbb2f9c83),
	.w2(32'h3a4b333e),
	.w3(32'hbb09484e),
	.w4(32'h3b74e40b),
	.w5(32'hbc1c8edd),
	.w6(32'h3a43d90a),
	.w7(32'hba17f3b0),
	.w8(32'hbb7381cf),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ba3e4),
	.w1(32'h3ba997d3),
	.w2(32'h3c47e2d0),
	.w3(32'hb98468e5),
	.w4(32'h3b36e4f9),
	.w5(32'hbb8ac13d),
	.w6(32'h3c078150),
	.w7(32'h3c215748),
	.w8(32'h3ac1da3d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb266e61),
	.w1(32'hbbc4ca8f),
	.w2(32'hbc081ffb),
	.w3(32'hbbae7f30),
	.w4(32'hbc0e4f4a),
	.w5(32'h388d666a),
	.w6(32'hbbfd0f24),
	.w7(32'hbbcd2211),
	.w8(32'hbb00231a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae6c5f),
	.w1(32'h3a6ea12d),
	.w2(32'hbc15693d),
	.w3(32'hba7da955),
	.w4(32'hbb9bbf1c),
	.w5(32'h3a369625),
	.w6(32'hb9c13eb5),
	.w7(32'hb937cb7f),
	.w8(32'hbaf13f4f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f3c61),
	.w1(32'h3c85b9c2),
	.w2(32'h3c204744),
	.w3(32'h3b6a95b4),
	.w4(32'h3ba4f4c1),
	.w5(32'h3a3e59d3),
	.w6(32'h3bd8083a),
	.w7(32'h3c309cf6),
	.w8(32'h3b2b5be4),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a753569),
	.w1(32'h3b4bb332),
	.w2(32'hbb2295a9),
	.w3(32'hbb7abade),
	.w4(32'h3b46c390),
	.w5(32'h3b9459f0),
	.w6(32'hba8e634c),
	.w7(32'h3b5af135),
	.w8(32'hb882cb13),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae681f4),
	.w1(32'hbb3ce66a),
	.w2(32'hbb36d53c),
	.w3(32'h3a40f355),
	.w4(32'h3b7e1618),
	.w5(32'h3b0e4154),
	.w6(32'hbbc87b8e),
	.w7(32'hba16c04a),
	.w8(32'h3ab74837),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b67ef),
	.w1(32'h3ba064be),
	.w2(32'hbad90c1b),
	.w3(32'hbc3a9eaf),
	.w4(32'hbb77115a),
	.w5(32'h3c4a8b9c),
	.w6(32'hbbeb5589),
	.w7(32'hbb01cf72),
	.w8(32'h3c831175),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba947b62),
	.w1(32'hbc2cf92b),
	.w2(32'hbb86d2d6),
	.w3(32'h3bff9dab),
	.w4(32'h3bd90993),
	.w5(32'hb982de8f),
	.w6(32'h3b388661),
	.w7(32'hbb3d5d30),
	.w8(32'hbbb700f6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5596f0),
	.w1(32'h3a22ea23),
	.w2(32'h398c837c),
	.w3(32'hbba25c59),
	.w4(32'hbbd53ba0),
	.w5(32'h3aef055e),
	.w6(32'hbbc13a8d),
	.w7(32'hbc1a7e2d),
	.w8(32'hbc070545),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d8d3a),
	.w1(32'hbc559c91),
	.w2(32'hbbec7bad),
	.w3(32'h3b093b65),
	.w4(32'h3ac8cc61),
	.w5(32'h3bd1c80b),
	.w6(32'hbba862d2),
	.w7(32'hba304acd),
	.w8(32'h3b5b8fe3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9013f),
	.w1(32'hbb9a2843),
	.w2(32'hbc342840),
	.w3(32'h3b141ba6),
	.w4(32'h3acbfb70),
	.w5(32'hb925ad37),
	.w6(32'hbb46c407),
	.w7(32'hbb996c9c),
	.w8(32'hba266651),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d9fc),
	.w1(32'hbbe42e33),
	.w2(32'h3b393fc9),
	.w3(32'h3af88a93),
	.w4(32'hbae18068),
	.w5(32'h3c2a8889),
	.w6(32'hb9a37581),
	.w7(32'h3a931e56),
	.w8(32'h3b551338),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule