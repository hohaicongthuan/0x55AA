module layer_10_featuremap_413(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c1772),
	.w1(32'hba3fb62b),
	.w2(32'h3a8fafcd),
	.w3(32'hbb469c72),
	.w4(32'hbb8404fb),
	.w5(32'hbb8ac0c1),
	.w6(32'hbbf85b13),
	.w7(32'h3b0fa9c4),
	.w8(32'h39ae34b0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb39ecf),
	.w1(32'hbad8592a),
	.w2(32'hba4b30f8),
	.w3(32'hbc1fb296),
	.w4(32'hbb43184d),
	.w5(32'hbbf1e39f),
	.w6(32'h3a5eb9cb),
	.w7(32'hba189e5e),
	.w8(32'hbaa06c3f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0b4c9),
	.w1(32'hb94257aa),
	.w2(32'hbbbcb6ac),
	.w3(32'h3c4d35b3),
	.w4(32'h3bd751ef),
	.w5(32'hbb654f43),
	.w6(32'h3c2e7481),
	.w7(32'hbb3496dd),
	.w8(32'hbb3cbcec),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab1f07),
	.w1(32'hbbb044a9),
	.w2(32'hba89004d),
	.w3(32'hbbd9b547),
	.w4(32'hbb58632c),
	.w5(32'hbba62e24),
	.w6(32'hbb573d5c),
	.w7(32'hbbcad9ee),
	.w8(32'hbb9361dc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22ebb9),
	.w1(32'h3adf0b5d),
	.w2(32'hbb14838c),
	.w3(32'h3ab39d33),
	.w4(32'h3afb3c5d),
	.w5(32'hbbd441ff),
	.w6(32'h3b57300d),
	.w7(32'h3b542578),
	.w8(32'hba7d7ac3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26240e),
	.w1(32'hbaf3037c),
	.w2(32'hbb18089b),
	.w3(32'hbb6b88c8),
	.w4(32'hba24cba0),
	.w5(32'h3b5dc340),
	.w6(32'hbadee50b),
	.w7(32'hbb94892c),
	.w8(32'hbbe864e4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b866e54),
	.w1(32'h3b0c64c0),
	.w2(32'h3bf241de),
	.w3(32'h3bd61339),
	.w4(32'hbab2642b),
	.w5(32'h3c4ea989),
	.w6(32'hbba3e44a),
	.w7(32'h3a2049ef),
	.w8(32'h3ba8048f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc980c3e),
	.w1(32'hbbbb23d8),
	.w2(32'hbc648aaf),
	.w3(32'hbcc55b92),
	.w4(32'hbcf7f316),
	.w5(32'hbc985f29),
	.w6(32'hbc31d0a6),
	.w7(32'hbcb190be),
	.w8(32'hbbfd00bb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3ddc4),
	.w1(32'h3b06e540),
	.w2(32'h3a116780),
	.w3(32'hbb387c0e),
	.w4(32'hbb3148e7),
	.w5(32'hbb45b3b6),
	.w6(32'hbad5bdc7),
	.w7(32'h39dd6b6a),
	.w8(32'h39ef1233),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeedda),
	.w1(32'h3ba39060),
	.w2(32'h3bd799e4),
	.w3(32'hbb7da59c),
	.w4(32'hb97f95b0),
	.w5(32'hbbaba864),
	.w6(32'h3ba1c5bb),
	.w7(32'h3ac24515),
	.w8(32'hbab9d5dc),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97e845),
	.w1(32'hbb8f9d8d),
	.w2(32'hba68fecf),
	.w3(32'hbbe37985),
	.w4(32'hbb1df1c9),
	.w5(32'hbad2989b),
	.w6(32'h3b0f1a12),
	.w7(32'h3b45a6cd),
	.w8(32'h3b37bbd5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b9e27),
	.w1(32'hbb20c67b),
	.w2(32'h3bccaa69),
	.w3(32'h3b8607e1),
	.w4(32'hbadbeffd),
	.w5(32'h3c5f15aa),
	.w6(32'h3a164126),
	.w7(32'h39e64d02),
	.w8(32'h3bec5dc0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb115b15),
	.w1(32'hbc142e12),
	.w2(32'hbbda588b),
	.w3(32'h3a5d76ea),
	.w4(32'hbb121a3b),
	.w5(32'h3b625b5f),
	.w6(32'h38ba01ea),
	.w7(32'h3a419c9e),
	.w8(32'hba91832e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae576ea),
	.w1(32'hbb9c39d7),
	.w2(32'hbb92c277),
	.w3(32'h3b7d2211),
	.w4(32'hbb87d44f),
	.w5(32'hbb23b768),
	.w6(32'h3b3552ed),
	.w7(32'hbb60a352),
	.w8(32'hba2d9698),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb432d0c),
	.w1(32'h3a91c4b6),
	.w2(32'h3b35ac28),
	.w3(32'hbbbae241),
	.w4(32'hba74a7dc),
	.w5(32'h3bb08d9e),
	.w6(32'h3971d95e),
	.w7(32'hba75d347),
	.w8(32'hba0156c7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52ce1f),
	.w1(32'hbb9304f1),
	.w2(32'hbc14a167),
	.w3(32'hbc3c4ac2),
	.w4(32'h3b1d5a0e),
	.w5(32'h3b3185ac),
	.w6(32'hbc40cc0d),
	.w7(32'hb9cc64ec),
	.w8(32'hbbef006c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b99f5),
	.w1(32'h3a09a556),
	.w2(32'hba267f08),
	.w3(32'h3b2a6b1b),
	.w4(32'h3b7834a9),
	.w5(32'h3bbb022d),
	.w6(32'h3ad2ba76),
	.w7(32'h3be7698d),
	.w8(32'h3b0ce588),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc430d63),
	.w1(32'hbc42e5f8),
	.w2(32'hbb41030b),
	.w3(32'hbc034539),
	.w4(32'hbbf6d620),
	.w5(32'hbbc95029),
	.w6(32'hbbe5dc79),
	.w7(32'h3b6f8f9c),
	.w8(32'hbbca1619),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc64a8e),
	.w1(32'hbbd3e30d),
	.w2(32'hbb82c012),
	.w3(32'hbc0bcfeb),
	.w4(32'hbbbded96),
	.w5(32'hbb5d0e80),
	.w6(32'hbb9efdf5),
	.w7(32'hba3ffb18),
	.w8(32'hbbe2102c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68454b),
	.w1(32'h3ad31da6),
	.w2(32'h3b81c227),
	.w3(32'hbb41e368),
	.w4(32'h3ae3e253),
	.w5(32'h3b3a1839),
	.w6(32'hbbc5ab62),
	.w7(32'hba743178),
	.w8(32'h3af48350),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a024a),
	.w1(32'hb9838e2f),
	.w2(32'h3a66b180),
	.w3(32'h3bbca69f),
	.w4(32'hba4719d2),
	.w5(32'h3bb8a90c),
	.w6(32'h3b926397),
	.w7(32'hbbe457a6),
	.w8(32'hbb7314f1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b102dc8),
	.w1(32'h39b9a416),
	.w2(32'hba29a832),
	.w3(32'h3b8772bc),
	.w4(32'hbad016f4),
	.w5(32'h3bce7dbb),
	.w6(32'h3bb7165f),
	.w7(32'hbb3379b8),
	.w8(32'hbb0070c3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb921a56),
	.w1(32'hbcf45d53),
	.w2(32'hbb243130),
	.w3(32'hba23f900),
	.w4(32'hbc1b30f3),
	.w5(32'h3c99e159),
	.w6(32'hbc3be09f),
	.w7(32'h3c071423),
	.w8(32'h3c6ea3b0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b147893),
	.w1(32'h3c76bb6c),
	.w2(32'h3c6b7f20),
	.w3(32'h3bd525bd),
	.w4(32'h3c2cf6b9),
	.w5(32'h3cb5b743),
	.w6(32'h3c24db66),
	.w7(32'h3c77b556),
	.w8(32'h3b5c19e9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d0809),
	.w1(32'h3c40bb1c),
	.w2(32'h3c4344f8),
	.w3(32'hbb12a086),
	.w4(32'hba2b6db2),
	.w5(32'hbba42959),
	.w6(32'h3c87563c),
	.w7(32'h3ab1692c),
	.w8(32'h3bf1bde2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad733d),
	.w1(32'h3b9f210a),
	.w2(32'h3b934b84),
	.w3(32'hbc142f2f),
	.w4(32'h3b3a77ab),
	.w5(32'h3bedc6bd),
	.w6(32'hbbccb8e0),
	.w7(32'hba13f374),
	.w8(32'h3b9fb553),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac7418),
	.w1(32'hbb72a7f6),
	.w2(32'hbbddb99a),
	.w3(32'h3a085af3),
	.w4(32'hbc2704ca),
	.w5(32'hbbfdf3c3),
	.w6(32'h3bb1d96a),
	.w7(32'hba963072),
	.w8(32'h3c2e1b96),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d700466),
	.w1(32'hbc2e2882),
	.w2(32'hbc9335cb),
	.w3(32'h3d38c3d6),
	.w4(32'hbc674749),
	.w5(32'hbcb2b31d),
	.w6(32'h3d461cf1),
	.w7(32'hbc86fcc4),
	.w8(32'hbc9770d8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb899e0d),
	.w1(32'hbb2ad383),
	.w2(32'hbaa7ca62),
	.w3(32'hbbb0183d),
	.w4(32'h39925608),
	.w5(32'h39eda6b5),
	.w6(32'hbb382e2b),
	.w7(32'hba72d182),
	.w8(32'h39eb654f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d42d146),
	.w1(32'h3b6a8ff0),
	.w2(32'hbb2f8eb0),
	.w3(32'h3d16e013),
	.w4(32'hba1e4101),
	.w5(32'hbc966fd0),
	.w6(32'h3d2ccc19),
	.w7(32'h3bcb43d0),
	.w8(32'hbb61cdbc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc050a71),
	.w1(32'hbb262ef7),
	.w2(32'hbaea040f),
	.w3(32'hbc455077),
	.w4(32'hbb7035ae),
	.w5(32'hbbffd8d9),
	.w6(32'hbbdc7e33),
	.w7(32'hbb1caf35),
	.w8(32'h3b0d9222),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b057823),
	.w1(32'hba885709),
	.w2(32'h3b6a883e),
	.w3(32'h3a8e843d),
	.w4(32'hbb1476ac),
	.w5(32'hba0c14b0),
	.w6(32'h3b09e40f),
	.w7(32'h381cbc55),
	.w8(32'h3b6f3a21),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39340c),
	.w1(32'h39fa14f9),
	.w2(32'hb707136a),
	.w3(32'h3bf1f6b9),
	.w4(32'hbc0413ef),
	.w5(32'hbc076773),
	.w6(32'h3b124765),
	.w7(32'h3b398768),
	.w8(32'h3b89a05b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1c8c4),
	.w1(32'h3adca793),
	.w2(32'hbb2e84de),
	.w3(32'hbb16a4a9),
	.w4(32'h3af4404a),
	.w5(32'hbb24b949),
	.w6(32'h3bdb56b1),
	.w7(32'h3b6cc228),
	.w8(32'h3bbbda64),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395394d9),
	.w1(32'h3b61ef31),
	.w2(32'hbab8f06e),
	.w3(32'h3abf304e),
	.w4(32'hb9bf131e),
	.w5(32'hbb9b5a4b),
	.w6(32'h3be27f87),
	.w7(32'hbbd196eb),
	.w8(32'hbc3a910e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2102d0),
	.w1(32'hbb8bba35),
	.w2(32'h3a968eeb),
	.w3(32'hba1885a0),
	.w4(32'hbc5b1aeb),
	.w5(32'hbc168d65),
	.w6(32'hbbbda46c),
	.w7(32'hbbb0a2ea),
	.w8(32'hba20f374),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec4604),
	.w1(32'h3baf9d33),
	.w2(32'hbc4e9ac2),
	.w3(32'hbb3b1de7),
	.w4(32'hbac99b86),
	.w5(32'h3c387cf9),
	.w6(32'hbc6dc800),
	.w7(32'h3b9c0c5d),
	.w8(32'h3cb068ad),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad3ee7),
	.w1(32'hbbd49b76),
	.w2(32'hbbcd17e3),
	.w3(32'h3b9d5fb0),
	.w4(32'hbca4ca89),
	.w5(32'hbce136a4),
	.w6(32'h3cc7816f),
	.w7(32'hbc1f767f),
	.w8(32'hbc42dec4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d769295),
	.w1(32'hbc3c47a0),
	.w2(32'hb9afe564),
	.w3(32'h3d4e8ab1),
	.w4(32'hbc8de19b),
	.w5(32'hbca96076),
	.w6(32'h3d76fd4a),
	.w7(32'hbb8da45d),
	.w8(32'hbc4c36fb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8708d),
	.w1(32'hb8b4bedb),
	.w2(32'h3a1519d1),
	.w3(32'hbbda83fb),
	.w4(32'hbaddd234),
	.w5(32'hba4569a1),
	.w6(32'hbb2a3bfa),
	.w7(32'hbb4bf761),
	.w8(32'hba3291ff),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf9bbe),
	.w1(32'hbc2af906),
	.w2(32'hba2defd9),
	.w3(32'hbaca80f9),
	.w4(32'hbbe505bc),
	.w5(32'h3c1f5c13),
	.w6(32'h3a2bcc74),
	.w7(32'hbbaed672),
	.w8(32'hbb0e2e88),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c3c69),
	.w1(32'hbb44d33f),
	.w2(32'hbb2a121f),
	.w3(32'h3a98bf65),
	.w4(32'hbb317726),
	.w5(32'hbb20e9d3),
	.w6(32'hb9823570),
	.w7(32'hbb4c86c4),
	.w8(32'hbbbaba08),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc2547),
	.w1(32'h3a2aa6ea),
	.w2(32'h3b20b601),
	.w3(32'hbadf2b1b),
	.w4(32'h3b494461),
	.w5(32'h3b25c97a),
	.w6(32'hba84bc7e),
	.w7(32'h3a8fbe8e),
	.w8(32'hba9f84df),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fa85e),
	.w1(32'hbc712008),
	.w2(32'hbc5d547b),
	.w3(32'h39d87681),
	.w4(32'hbb07b016),
	.w5(32'hbb7e11a5),
	.w6(32'hba9c9f29),
	.w7(32'h3b222daf),
	.w8(32'h3ac34934),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd5c6d),
	.w1(32'h3c01965b),
	.w2(32'h3c0928fb),
	.w3(32'hbb1a543b),
	.w4(32'h3aa3108e),
	.w5(32'hbb89dc39),
	.w6(32'h3c0e450f),
	.w7(32'h3b7c378c),
	.w8(32'h3b66e8bb),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8004fa),
	.w1(32'h3bce5011),
	.w2(32'h3c387215),
	.w3(32'hbc2bf6bc),
	.w4(32'hbb97eda0),
	.w5(32'hbc01a210),
	.w6(32'h3b842feb),
	.w7(32'h3c8068e5),
	.w8(32'h3c48444f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb949bb9),
	.w1(32'hbb7a9a0b),
	.w2(32'hb9d4dde0),
	.w3(32'hbb92c7a3),
	.w4(32'hbb5ddf55),
	.w5(32'h3ab1ce2e),
	.w6(32'h3beb93b2),
	.w7(32'h3af477fb),
	.w8(32'h3b23910b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81476f),
	.w1(32'hbc3b01b1),
	.w2(32'hbbf021fa),
	.w3(32'hbba94541),
	.w4(32'hbc0e8d39),
	.w5(32'hbba91200),
	.w6(32'hbb553e19),
	.w7(32'h3b032f2d),
	.w8(32'h3adbe310),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad6c99),
	.w1(32'h3b588276),
	.w2(32'h3b103b6b),
	.w3(32'h3b9a9430),
	.w4(32'hbbf92413),
	.w5(32'hbb40196c),
	.w6(32'h3b7813e2),
	.w7(32'hbbb6a546),
	.w8(32'hbb1ec64c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30d89f),
	.w1(32'h3b8f36f3),
	.w2(32'h3bd10144),
	.w3(32'hbbdf983a),
	.w4(32'hbb75d2b6),
	.w5(32'hbbd510f1),
	.w6(32'hbb48f5d9),
	.w7(32'hbbb42120),
	.w8(32'hbb842075),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043a76),
	.w1(32'h3b58894b),
	.w2(32'hbc0288f5),
	.w3(32'hbbefe0bf),
	.w4(32'h3adc00e7),
	.w5(32'hbc4e613f),
	.w6(32'hbbca4b95),
	.w7(32'hbadca50f),
	.w8(32'hbc1d959c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11060d),
	.w1(32'hbb72f43a),
	.w2(32'h3c492881),
	.w3(32'h39e1a9c7),
	.w4(32'hbbc088f0),
	.w5(32'h3bb55bc5),
	.w6(32'hba6022bc),
	.w7(32'h3b1c4a31),
	.w8(32'h3bb386f6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b853c86),
	.w1(32'hbab99a82),
	.w2(32'hbb10dfbb),
	.w3(32'h3b89eb1e),
	.w4(32'hbba29796),
	.w5(32'hbba14bed),
	.w6(32'h3b86c752),
	.w7(32'hba0a62b9),
	.w8(32'h3aa82ebe),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1871a1),
	.w1(32'hbc611a67),
	.w2(32'hbc52bc13),
	.w3(32'hbc210b55),
	.w4(32'hbc17c21c),
	.w5(32'hbbdd8015),
	.w6(32'hbb9f7c10),
	.w7(32'hbbfa0e7e),
	.w8(32'hbbc6b212),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b509c67),
	.w1(32'hbb0ccad8),
	.w2(32'hba05c25b),
	.w3(32'hbbb9f038),
	.w4(32'hb96e3e63),
	.w5(32'hbc14eb61),
	.w6(32'h3b4a894b),
	.w7(32'h3be82f16),
	.w8(32'h3baca363),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb315575),
	.w1(32'h3bab2cbf),
	.w2(32'h3b59590c),
	.w3(32'hbc0cbcce),
	.w4(32'h3ba311c0),
	.w5(32'h3ad358af),
	.w6(32'hbba895d0),
	.w7(32'h3b522be5),
	.w8(32'h3b248b17),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c75da),
	.w1(32'hba1e02ca),
	.w2(32'hbba495d4),
	.w3(32'h3b83b4ba),
	.w4(32'hbb861fba),
	.w5(32'hbb8fbaf0),
	.w6(32'h3c557640),
	.w7(32'hbb8e12ab),
	.w8(32'hbbadcbfe),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacd533),
	.w1(32'hba18f113),
	.w2(32'h3a7850e0),
	.w3(32'hba585ae2),
	.w4(32'hb8e880e6),
	.w5(32'hba0345e4),
	.w6(32'h3ab58a07),
	.w7(32'hb98bfc70),
	.w8(32'hbae56b48),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ad2df),
	.w1(32'h3bb6eddc),
	.w2(32'h3b81cb9e),
	.w3(32'h3b6d2c17),
	.w4(32'h3afcc765),
	.w5(32'h3c2a179f),
	.w6(32'h3b4ac3f5),
	.w7(32'h3a8d2d59),
	.w8(32'hbaf392ff),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86544e),
	.w1(32'h396f557b),
	.w2(32'hbafaf226),
	.w3(32'hbbaf76d2),
	.w4(32'h3c0d6ff6),
	.w5(32'h3b153224),
	.w6(32'hbbc06c69),
	.w7(32'hbb842f31),
	.w8(32'hba216de8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc58fb7),
	.w1(32'hbbef61fc),
	.w2(32'h3a360290),
	.w3(32'hbb87d774),
	.w4(32'hbb26cfbc),
	.w5(32'hbabf25d1),
	.w6(32'hbc02dda3),
	.w7(32'h3a71091a),
	.w8(32'h3a9b6843),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b288da5),
	.w1(32'hbc16de61),
	.w2(32'hbae99402),
	.w3(32'hbba278e0),
	.w4(32'hbbffcc7f),
	.w5(32'hbc20fa4a),
	.w6(32'hbbc3ac4b),
	.w7(32'h3976d802),
	.w8(32'hbacbacb2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d762c),
	.w1(32'h3bf9c0be),
	.w2(32'h3bec0dcf),
	.w3(32'hbb97e804),
	.w4(32'h3c36e3fd),
	.w5(32'h3c33fadd),
	.w6(32'hba2b3f57),
	.w7(32'hbb09d466),
	.w8(32'hbb2c7e36),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15457d),
	.w1(32'hb8854802),
	.w2(32'hbb2068a9),
	.w3(32'hbb105357),
	.w4(32'hbb386bbe),
	.w5(32'hbb7e3129),
	.w6(32'hbaed3d55),
	.w7(32'h3bbea6cb),
	.w8(32'h3b8e48ec),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22b34b),
	.w1(32'h38be44bd),
	.w2(32'h3a97c4f0),
	.w3(32'h3ac0c524),
	.w4(32'hbaaef029),
	.w5(32'h3b5e03eb),
	.w6(32'h3ab9864b),
	.w7(32'hbbfc5e8b),
	.w8(32'hbbbf85a2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba557c2),
	.w1(32'hbb840a5d),
	.w2(32'hba6e002e),
	.w3(32'hbc09909f),
	.w4(32'hbbb7bc84),
	.w5(32'hbb4fde27),
	.w6(32'hbc192767),
	.w7(32'h39a98736),
	.w8(32'hbac4666d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65ba39),
	.w1(32'hbbdb6b18),
	.w2(32'hbcc64d7d),
	.w3(32'hbc29f598),
	.w4(32'h3c06ade3),
	.w5(32'h3b56ea67),
	.w6(32'hbc6426c1),
	.w7(32'hbadfcf1b),
	.w8(32'hbae6432d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40de7d),
	.w1(32'h3ca7fdcc),
	.w2(32'h3cc425a9),
	.w3(32'hbc745988),
	.w4(32'hbbaac235),
	.w5(32'hbcc1bec9),
	.w6(32'h3c312ec6),
	.w7(32'h3cea210b),
	.w8(32'h3cb4fea6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85c40f),
	.w1(32'h3c388638),
	.w2(32'h3bb862ab),
	.w3(32'hbc851cfb),
	.w4(32'h3bab869b),
	.w5(32'hbc41567c),
	.w6(32'hbbf375af),
	.w7(32'h3cbce45c),
	.w8(32'h3c22f35a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cec07e4),
	.w1(32'h3c49d959),
	.w2(32'h3c235235),
	.w3(32'h3a777b59),
	.w4(32'hbc2b0b04),
	.w5(32'hbc53d17c),
	.w6(32'h3cac740a),
	.w7(32'h3bfabdc7),
	.w8(32'h3b4d46fb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34f9eb),
	.w1(32'hbb3c5b7b),
	.w2(32'hbb2961b6),
	.w3(32'hbaa9ea18),
	.w4(32'hb9b1aeae),
	.w5(32'hbaecd0a5),
	.w6(32'h3af85bcb),
	.w7(32'hb9d53895),
	.w8(32'h3a8bb53c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbe0f0),
	.w1(32'h3b0bce21),
	.w2(32'hbb2635b8),
	.w3(32'hbad7d057),
	.w4(32'hbab16209),
	.w5(32'hbb06f3d0),
	.w6(32'hba9fe01a),
	.w7(32'hbb51a909),
	.w8(32'hba025202),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b3b82f),
	.w1(32'hbb2f2ca8),
	.w2(32'h3b6ecf11),
	.w3(32'hbb55ec9b),
	.w4(32'hbb8e7bab),
	.w5(32'h3af4a0af),
	.w6(32'hba5ccf65),
	.w7(32'hbbab6936),
	.w8(32'hbac6ec76),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb354509),
	.w1(32'hbb27c2d4),
	.w2(32'h39785bbf),
	.w3(32'h3b3d2dec),
	.w4(32'h3a321c4a),
	.w5(32'hbb0a2965),
	.w6(32'h3bb7c30b),
	.w7(32'h3ba45875),
	.w8(32'hbaf94dfb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77986a),
	.w1(32'hbbd566f7),
	.w2(32'hbc04b8c6),
	.w3(32'h3aa34b1a),
	.w4(32'hb7b84821),
	.w5(32'hbbdd6603),
	.w6(32'hbb2dbb9b),
	.w7(32'hbbb22e89),
	.w8(32'hbbda0722),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc755a03),
	.w1(32'hbba7283d),
	.w2(32'hbb83dc25),
	.w3(32'hbc5335a7),
	.w4(32'hbb989263),
	.w5(32'hbb9c6790),
	.w6(32'hbc2cb7ae),
	.w7(32'hbbfa2585),
	.w8(32'hbc015665),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d1a0c),
	.w1(32'h3af72f85),
	.w2(32'hbc0ccfe0),
	.w3(32'hbb4d1f6a),
	.w4(32'hbb9bfb6b),
	.w5(32'hbb95bfa2),
	.w6(32'hbb9b945c),
	.w7(32'hb990b94e),
	.w8(32'h3b26cf17),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a436b84),
	.w1(32'h3bf12993),
	.w2(32'h3c8484a6),
	.w3(32'h3b21dcbf),
	.w4(32'hbb4e2d06),
	.w5(32'h3b2334b1),
	.w6(32'h3c36ab87),
	.w7(32'h3c0865ce),
	.w8(32'h3c660312),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc31c38),
	.w1(32'h3b4483dc),
	.w2(32'hbb2b8f9f),
	.w3(32'h3b863084),
	.w4(32'h3a763587),
	.w5(32'h3b43865d),
	.w6(32'h3afdc335),
	.w7(32'h3bdf70b8),
	.w8(32'h3b07dc66),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01969e),
	.w1(32'hbb43d332),
	.w2(32'hbc0bdccc),
	.w3(32'hbb967484),
	.w4(32'hbb916376),
	.w5(32'hbb00f86a),
	.w6(32'hbac1a8d6),
	.w7(32'h3bb9ac46),
	.w8(32'hbb349f4f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94e644),
	.w1(32'h3b62cb8e),
	.w2(32'hba8a4f82),
	.w3(32'h3afd7479),
	.w4(32'h3bf44453),
	.w5(32'h3c2962bf),
	.w6(32'h3beecf10),
	.w7(32'h3c37c561),
	.w8(32'h3c230481),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24f61d),
	.w1(32'h3b74a968),
	.w2(32'h3bef8af8),
	.w3(32'hb8f8889a),
	.w4(32'h3ac57fcc),
	.w5(32'h3bdc5b98),
	.w6(32'h3b08b71e),
	.w7(32'h3bea29a1),
	.w8(32'h3c1ce48b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba45797),
	.w1(32'hb9a53ff9),
	.w2(32'h3b399d28),
	.w3(32'h3c4fff13),
	.w4(32'h3babe0a8),
	.w5(32'h3b907ec4),
	.w6(32'h3bd94ba5),
	.w7(32'h3b810dac),
	.w8(32'h3b00e4c2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf0c65),
	.w1(32'hbaf85623),
	.w2(32'hbb8c63fc),
	.w3(32'h3b91ff43),
	.w4(32'h3b17331f),
	.w5(32'hbb6755e8),
	.w6(32'hb995f048),
	.w7(32'hba99ab4b),
	.w8(32'hbb91da95),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd092fb),
	.w1(32'hba3180ea),
	.w2(32'h3ba09d87),
	.w3(32'hbb9c6d4a),
	.w4(32'hb9f8898d),
	.w5(32'h3b634fb8),
	.w6(32'hb6288210),
	.w7(32'h3aa1e3f3),
	.w8(32'h3ba3318e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90077c),
	.w1(32'hbbb4b2d3),
	.w2(32'hbc2b96a1),
	.w3(32'h3c214ed1),
	.w4(32'hbb0ea2d6),
	.w5(32'hbc8316a3),
	.w6(32'h3c2a1292),
	.w7(32'hbc4bd441),
	.w8(32'hbc0f22ab),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4acf8e),
	.w1(32'hbb94d497),
	.w2(32'hbba8a1ce),
	.w3(32'hbc8d3c00),
	.w4(32'hbb333c67),
	.w5(32'h39a29b6a),
	.w6(32'hbbe3022e),
	.w7(32'h3c25bf72),
	.w8(32'h3b46680f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b237678),
	.w1(32'h3902a373),
	.w2(32'hbb0016bb),
	.w3(32'hbba45f52),
	.w4(32'h3a54cbb7),
	.w5(32'hba2dd851),
	.w6(32'hbb1a88fe),
	.w7(32'h3b5c3237),
	.w8(32'h3b3144d6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb086f19),
	.w1(32'h3bc4d5cb),
	.w2(32'h3b596452),
	.w3(32'hbc5f6ab0),
	.w4(32'hbb4d9fe3),
	.w5(32'hbb7a9fe1),
	.w6(32'h3b7e512f),
	.w7(32'h3b8281f3),
	.w8(32'h3bce9e6e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc322566),
	.w1(32'h3b09c652),
	.w2(32'h3b4c0ee6),
	.w3(32'hbc9c21de),
	.w4(32'hbc29705b),
	.w5(32'h3af0310c),
	.w6(32'hbc136493),
	.w7(32'h3baadc6b),
	.w8(32'h39882e32),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca05270),
	.w1(32'hbaeec4cd),
	.w2(32'hbbd0fd23),
	.w3(32'h3c707529),
	.w4(32'hbbbc5cd1),
	.w5(32'hbc0ff4a9),
	.w6(32'h3c7be50b),
	.w7(32'h3b11bab9),
	.w8(32'hbb8607bc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cd344),
	.w1(32'hbca66b72),
	.w2(32'hbc774d0d),
	.w3(32'h3a4103b3),
	.w4(32'hbc04179c),
	.w5(32'h3c48ed25),
	.w6(32'hbc7472fb),
	.w7(32'hbbbbdb20),
	.w8(32'h3a570cb6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5a38c),
	.w1(32'hbbfd8a22),
	.w2(32'hbb65925e),
	.w3(32'hbc0c7c98),
	.w4(32'hbb6d5307),
	.w5(32'hbb576608),
	.w6(32'h3b41f67f),
	.w7(32'hbb0ac2b2),
	.w8(32'h3b07a9cf),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ec430),
	.w1(32'hbaf451f8),
	.w2(32'hbbed2904),
	.w3(32'hbc11603b),
	.w4(32'hbb3dd7d2),
	.w5(32'h3b8e250c),
	.w6(32'hbc1cbe32),
	.w7(32'hbabfb542),
	.w8(32'h3be65f70),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886aab),
	.w1(32'hbbbf5d39),
	.w2(32'h3b04e81a),
	.w3(32'hbb7f14e4),
	.w4(32'hbbd503c3),
	.w5(32'hbb8db16b),
	.w6(32'h3c1d9eaa),
	.w7(32'h3a92e563),
	.w8(32'h3bacc9d9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb57d16),
	.w1(32'h3afffd60),
	.w2(32'h3a8b399a),
	.w3(32'h3b8db7fb),
	.w4(32'hbba6ea5d),
	.w5(32'hbc3ecd85),
	.w6(32'h3c8e53ac),
	.w7(32'hba4ae1a6),
	.w8(32'hbbd103e5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c3b2a),
	.w1(32'h3b18c9c0),
	.w2(32'h3a23d3c8),
	.w3(32'hbbe21095),
	.w4(32'h3afa9d2e),
	.w5(32'hbbd2bbdb),
	.w6(32'hbbae2719),
	.w7(32'h386cb1e7),
	.w8(32'h3b2ae86b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae91257),
	.w1(32'hbc38b2a6),
	.w2(32'hbba784a9),
	.w3(32'h3b0fcb17),
	.w4(32'hbc30f6d2),
	.w5(32'hbbf724f0),
	.w6(32'h3bd9a4c9),
	.w7(32'hbaa185d5),
	.w8(32'hba8d9eb2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b368001),
	.w1(32'hbc4c35b1),
	.w2(32'hbc194aab),
	.w3(32'h3c1a6b5b),
	.w4(32'hbc0e7a88),
	.w5(32'h3b2ef88a),
	.w6(32'h3b814e4f),
	.w7(32'hbaa58089),
	.w8(32'hbbd8127b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e68f9),
	.w1(32'h3b79a4b0),
	.w2(32'hbb027667),
	.w3(32'hbc490983),
	.w4(32'hbcc5b849),
	.w5(32'h3c1dcced),
	.w6(32'hbcd169cd),
	.w7(32'hbaeaf524),
	.w8(32'h3cfca150),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ce614),
	.w1(32'hbbac995f),
	.w2(32'hbc11083c),
	.w3(32'hbbb57708),
	.w4(32'hbc000f53),
	.w5(32'hbc8c4d38),
	.w6(32'h3b04f41b),
	.w7(32'h3b1ad194),
	.w8(32'hba09d88e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b7ada),
	.w1(32'h3bf104ca),
	.w2(32'h3c75904a),
	.w3(32'hbac2e43d),
	.w4(32'hbb7ae4c0),
	.w5(32'hbb3d6d10),
	.w6(32'h3c441797),
	.w7(32'h3c00fbd7),
	.w8(32'h3c5f458d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4439),
	.w1(32'hbbe70893),
	.w2(32'hbc34ce15),
	.w3(32'h3c5e6550),
	.w4(32'hba955962),
	.w5(32'h3c523b2d),
	.w6(32'hba19936f),
	.w7(32'h39fc4ace),
	.w8(32'h3c46a66e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e43d0),
	.w1(32'hb9b1fbec),
	.w2(32'h3c11132d),
	.w3(32'hba588cde),
	.w4(32'hbbb68249),
	.w5(32'h3bed72f8),
	.w6(32'h3aae6254),
	.w7(32'h3b300152),
	.w8(32'h3b15b650),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab37ea),
	.w1(32'h3b428d05),
	.w2(32'hbc556583),
	.w3(32'hbb2137eb),
	.w4(32'h383877d1),
	.w5(32'h3c3d82ad),
	.w6(32'hbc2344c5),
	.w7(32'h3bb41dfa),
	.w8(32'h3ce0b4e1),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf096a3),
	.w1(32'h3bb4a92b),
	.w2(32'hbb12c915),
	.w3(32'hbb7cb233),
	.w4(32'h3c133e2d),
	.w5(32'h3a6333e6),
	.w6(32'hbbe1db70),
	.w7(32'h3b936036),
	.w8(32'h3c29c213),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ea4a0),
	.w1(32'hbb0d8160),
	.w2(32'h3ac68606),
	.w3(32'h3bfe8934),
	.w4(32'h390c6de4),
	.w5(32'h3bb6f23a),
	.w6(32'h3bca2500),
	.w7(32'hbaeadd18),
	.w8(32'h3b9b5127),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf67ce),
	.w1(32'hbb3664ec),
	.w2(32'h39c9e8d5),
	.w3(32'hba2a02f4),
	.w4(32'hbb44d645),
	.w5(32'h3bd2848e),
	.w6(32'hbb6e837a),
	.w7(32'hbb8da1ca),
	.w8(32'h3ab3ec2c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a732e),
	.w1(32'hbbf07998),
	.w2(32'hbad6ae7a),
	.w3(32'hba9f1c4d),
	.w4(32'hbb519982),
	.w5(32'hbb73a7c2),
	.w6(32'hbb1856e1),
	.w7(32'hb902ce1a),
	.w8(32'h3b46b240),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c245cdb),
	.w1(32'h3c0fba05),
	.w2(32'h3c556ef1),
	.w3(32'h3b09eabd),
	.w4(32'h3b9ded8d),
	.w5(32'h3b6c295b),
	.w6(32'h3c23d13f),
	.w7(32'h3bedfe84),
	.w8(32'h3c218b0b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d4e8b),
	.w1(32'hbc5cb614),
	.w2(32'hbb9fd317),
	.w3(32'h3c794012),
	.w4(32'hbc32fbbe),
	.w5(32'hbc5ea02b),
	.w6(32'h3d06e831),
	.w7(32'hbbebb23d),
	.w8(32'hbb8f70be),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbceeaf7),
	.w1(32'hbb7ebf57),
	.w2(32'h3c20ea8c),
	.w3(32'hbbee46ff),
	.w4(32'hbbff3d2d),
	.w5(32'hbbc39e85),
	.w6(32'hbb8ccee6),
	.w7(32'hbb931eb7),
	.w8(32'h3b4f6c07),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc748dc),
	.w1(32'h3b47825c),
	.w2(32'h3c9614b6),
	.w3(32'hbc074cd0),
	.w4(32'hbc6df3ea),
	.w5(32'hbb3fd820),
	.w6(32'hbbc5f257),
	.w7(32'hbb58c485),
	.w8(32'h3c9002b6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6032c4),
	.w1(32'hbbed8d42),
	.w2(32'hbc5965e0),
	.w3(32'hbaa1202f),
	.w4(32'h3b1eaab7),
	.w5(32'hb92d26a1),
	.w6(32'hbb379a0e),
	.w7(32'hbb2b66b6),
	.w8(32'hbc29da73),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8db5d9),
	.w1(32'hbb3590eb),
	.w2(32'hbb86ea81),
	.w3(32'hbb7922aa),
	.w4(32'h3917f306),
	.w5(32'hbac1d871),
	.w6(32'h3bd51380),
	.w7(32'h3a559aa1),
	.w8(32'hbb6d1cbe),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf37638),
	.w1(32'h3bd0fdd4),
	.w2(32'h3b5f54d1),
	.w3(32'h3bcc91a1),
	.w4(32'h3bae9d8a),
	.w5(32'h3b947045),
	.w6(32'h3b41fc5e),
	.w7(32'h3bb97337),
	.w8(32'h3b2d6efc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adda409),
	.w1(32'hbb4fe21a),
	.w2(32'h3a6a4c52),
	.w3(32'h3ac223b8),
	.w4(32'h3b636151),
	.w5(32'h3b17efc0),
	.w6(32'hbb72d65a),
	.w7(32'hb9482966),
	.w8(32'h37e8b456),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b07af),
	.w1(32'hbb27de91),
	.w2(32'hb950be13),
	.w3(32'h3c0942f3),
	.w4(32'hbbcbcd01),
	.w5(32'h3a5c7873),
	.w6(32'h3c1fa5ee),
	.w7(32'hb9a5489a),
	.w8(32'h3b1af52e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b654ab4),
	.w1(32'hba089e41),
	.w2(32'hb9d23ba7),
	.w3(32'h3bb7107b),
	.w4(32'h3b8e9a87),
	.w5(32'h399c9b35),
	.w6(32'h3bdcbe01),
	.w7(32'h3b0aff03),
	.w8(32'hba04fc88),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00e6b9),
	.w1(32'h3bee2bfa),
	.w2(32'h3c11aa7b),
	.w3(32'hbbaca3f4),
	.w4(32'h3acf9c2c),
	.w5(32'h3aca26ee),
	.w6(32'h3b1c703c),
	.w7(32'h3c013ffb),
	.w8(32'h3c4310a6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a90a7),
	.w1(32'h3b7467c4),
	.w2(32'hbc3c5de6),
	.w3(32'h3c31f495),
	.w4(32'h3b56dbdd),
	.w5(32'hbb204ce7),
	.w6(32'h3c1fed98),
	.w7(32'h3b0efe9a),
	.w8(32'hbbacd431),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3954ab),
	.w1(32'hbb48e814),
	.w2(32'hba0ebfac),
	.w3(32'hbbdff6d3),
	.w4(32'hbbc8864b),
	.w5(32'h3ab5a172),
	.w6(32'hbbde5c4c),
	.w7(32'hbc0786d1),
	.w8(32'hb89661a8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8dfc9),
	.w1(32'h3bdc22f5),
	.w2(32'h3be47df2),
	.w3(32'hbc40a147),
	.w4(32'hbb7fb231),
	.w5(32'hbc2150e0),
	.w6(32'h3be60ffd),
	.w7(32'hba09c5a4),
	.w8(32'h3b6d8bb4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971fa74),
	.w1(32'hbb91ee65),
	.w2(32'h3bb06639),
	.w3(32'hba0d1c32),
	.w4(32'hbb58da3a),
	.w5(32'hbbb6fa62),
	.w6(32'hba2a50bb),
	.w7(32'hba71f23f),
	.w8(32'h3ac19667),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6e870),
	.w1(32'hbbaf3190),
	.w2(32'h3b129c9d),
	.w3(32'h3bd2c8c4),
	.w4(32'hbbd2c185),
	.w5(32'hbbefcdd1),
	.w6(32'h3b7b0633),
	.w7(32'hbb744e48),
	.w8(32'hb94d3eaa),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42cb64),
	.w1(32'hbbaf8f29),
	.w2(32'h3ababf02),
	.w3(32'hbb674b49),
	.w4(32'hbae3d8d8),
	.w5(32'h3ab66238),
	.w6(32'hb8d51c30),
	.w7(32'hbbd7277c),
	.w8(32'hbb4915bd),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ce51b),
	.w1(32'hbb93fd53),
	.w2(32'hbb613d13),
	.w3(32'hbb6c3c42),
	.w4(32'hbc1d6fa2),
	.w5(32'hbc95697b),
	.w6(32'hbb332e5c),
	.w7(32'hbb9207be),
	.w8(32'hbc3977f8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c964b83),
	.w1(32'hbb1cf829),
	.w2(32'h3c3124d3),
	.w3(32'hbc6a7364),
	.w4(32'hbc837398),
	.w5(32'hbc48fd89),
	.w6(32'hbc515c5c),
	.w7(32'h3affca88),
	.w8(32'h39f5e535),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ca098),
	.w1(32'hbac50ee5),
	.w2(32'hbc42d26d),
	.w3(32'hbc6295ac),
	.w4(32'h3b3bc1a9),
	.w5(32'h3b0146ff),
	.w6(32'hbbfd31ae),
	.w7(32'h3a8cd639),
	.w8(32'hba603688),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc734883),
	.w1(32'hbb473be2),
	.w2(32'hbb95201d),
	.w3(32'hbc698cf9),
	.w4(32'hbb1aa0f3),
	.w5(32'hbaaac95b),
	.w6(32'hbc1e1d12),
	.w7(32'hba77dd83),
	.w8(32'hbbd60e9a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90e85f),
	.w1(32'h3b25f13d),
	.w2(32'h3b5daf57),
	.w3(32'hbc0c07cd),
	.w4(32'h38933218),
	.w5(32'h3bb95149),
	.w6(32'hbb192c02),
	.w7(32'h3b8b8e5a),
	.w8(32'h3ba3ab80),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85600f),
	.w1(32'hba7120cf),
	.w2(32'hbbd9f924),
	.w3(32'h3c146738),
	.w4(32'hbb321013),
	.w5(32'hba7710c5),
	.w6(32'h3c3ef2cd),
	.w7(32'hbb33e081),
	.w8(32'hbb7adf15),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07d3f8),
	.w1(32'hbbc22d7e),
	.w2(32'h3969f21c),
	.w3(32'hbc0f1d84),
	.w4(32'hbbf6fefe),
	.w5(32'hbb332840),
	.w6(32'hbbf9f39a),
	.w7(32'hbb200819),
	.w8(32'h3bfa6488),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40b948),
	.w1(32'hbb99b52c),
	.w2(32'hbbaf938d),
	.w3(32'hbbee6984),
	.w4(32'h3b82728e),
	.w5(32'hbbe38777),
	.w6(32'hbb68f98a),
	.w7(32'hbabbebf0),
	.w8(32'hbb433e96),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67fa00),
	.w1(32'hbc7cb1f7),
	.w2(32'hbc237877),
	.w3(32'h3b95d875),
	.w4(32'hbb4277c2),
	.w5(32'h3b06d8e1),
	.w6(32'hb9c1a9f2),
	.w7(32'hbbd51527),
	.w8(32'hbc194a5b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c7eb0),
	.w1(32'h3bbbf308),
	.w2(32'h3b577148),
	.w3(32'hbc2fb9bd),
	.w4(32'hbb512f1f),
	.w5(32'h3b3a79ce),
	.w6(32'hbaea24f6),
	.w7(32'h3b422145),
	.w8(32'h3bc6692c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe08ffe),
	.w1(32'hbb9abc7e),
	.w2(32'h3b7c1123),
	.w3(32'h39cf2865),
	.w4(32'hbb9bea0a),
	.w5(32'h3b9b0aa1),
	.w6(32'hbb2011c5),
	.w7(32'h3bf5b75e),
	.w8(32'h3be111cd),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86e021),
	.w1(32'hbcf0e5e2),
	.w2(32'hbc754bd0),
	.w3(32'h39c68f30),
	.w4(32'hbc588157),
	.w5(32'hbba24b7c),
	.w6(32'hbad6e7c4),
	.w7(32'hbc0fc164),
	.w8(32'hbb9c6a51),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59006b),
	.w1(32'h38188b20),
	.w2(32'hb79f4072),
	.w3(32'hbca6d9f8),
	.w4(32'hbbb62a64),
	.w5(32'hbc1def60),
	.w6(32'hbc5d4545),
	.w7(32'hb9e943c6),
	.w8(32'h3badf616),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedb17a),
	.w1(32'h3bc36f9e),
	.w2(32'h3b2f0a6e),
	.w3(32'hbb045e57),
	.w4(32'h3ba5c8e5),
	.w5(32'h3b97ee3a),
	.w6(32'h3a8ed42c),
	.w7(32'h3b0e0ee9),
	.w8(32'h3b2f60c1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22a52b),
	.w1(32'h3b92ec72),
	.w2(32'h3bf7acbf),
	.w3(32'h3c163d65),
	.w4(32'h3b8ea15a),
	.w5(32'h3bf6cd2d),
	.w6(32'h3bc4fa92),
	.w7(32'h3b596e8b),
	.w8(32'h3b3b86b2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d69767c),
	.w1(32'hbbdf8033),
	.w2(32'h3baa3333),
	.w3(32'h3d19cb72),
	.w4(32'hbcdfbbec),
	.w5(32'hbc9e0863),
	.w6(32'h3d3762a7),
	.w7(32'hbbf6d7d6),
	.w8(32'hbc1a604f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7ba7a),
	.w1(32'hbbeb659c),
	.w2(32'h3c11acbe),
	.w3(32'hbc08031d),
	.w4(32'hbbf48c12),
	.w5(32'hbbaec7de),
	.w6(32'h3aac3e95),
	.w7(32'hbbab119a),
	.w8(32'h3b17c9e0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befe2a0),
	.w1(32'h3b9a6d0f),
	.w2(32'h3b468f4e),
	.w3(32'h3c28b212),
	.w4(32'h3b83970c),
	.w5(32'h3b865f0d),
	.w6(32'h3b69960c),
	.w7(32'h3addab2c),
	.w8(32'h3b28e097),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae2707),
	.w1(32'h3b3ab4b9),
	.w2(32'h3ba697fc),
	.w3(32'h3b840602),
	.w4(32'h3bbc90af),
	.w5(32'h3b8e8bae),
	.w6(32'hbba81b8b),
	.w7(32'h3bbd6bc5),
	.w8(32'h3a296744),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b3051),
	.w1(32'h3b84c485),
	.w2(32'hbc56f398),
	.w3(32'hbb98a482),
	.w4(32'h3bb1a48e),
	.w5(32'h3a8f2b10),
	.w6(32'hbba7c487),
	.w7(32'h3badc931),
	.w8(32'h3bfcdf5a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18dd9d),
	.w1(32'h3ba68c97),
	.w2(32'h3beb1068),
	.w3(32'hbc926d31),
	.w4(32'h3afa7136),
	.w5(32'hbb9c93ec),
	.w6(32'hbc1aa010),
	.w7(32'h3b99eedc),
	.w8(32'h3bf8b006),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a7943),
	.w1(32'h3a30a233),
	.w2(32'hbb50f92c),
	.w3(32'h3bc5c26c),
	.w4(32'h3a8bcb5b),
	.w5(32'hb9fa99d0),
	.w6(32'h3be70143),
	.w7(32'h3bb96175),
	.w8(32'h3b4586c2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf30727),
	.w1(32'h3b4db5d6),
	.w2(32'h3b6cc2ef),
	.w3(32'h3c11caf0),
	.w4(32'h3b6a0f30),
	.w5(32'h3a7aacb3),
	.w6(32'hbb23692c),
	.w7(32'h3b2c0478),
	.w8(32'h39e19715),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be49a51),
	.w1(32'hbc311c28),
	.w2(32'hbc99ba2f),
	.w3(32'h3c3e99be),
	.w4(32'hbc326987),
	.w5(32'hbc6e56cd),
	.w6(32'h3c061609),
	.w7(32'hbc1a817c),
	.w8(32'hbc500ad6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b8f5b),
	.w1(32'hbaaed010),
	.w2(32'hbb06a57d),
	.w3(32'h3c07dcd3),
	.w4(32'hbbac4505),
	.w5(32'hbbc2f5ed),
	.w6(32'h3ba12420),
	.w7(32'hb9a86df0),
	.w8(32'h3a9c1bfe),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f83ae),
	.w1(32'hbc326afd),
	.w2(32'hbbc417ac),
	.w3(32'hbbfd67d8),
	.w4(32'hbbbc84f8),
	.w5(32'h3c0b6e30),
	.w6(32'hbbdbefd0),
	.w7(32'hbc1b7a1a),
	.w8(32'hbb88051b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0904e1),
	.w1(32'hbbd07c55),
	.w2(32'hbb3bd380),
	.w3(32'h3cd7e250),
	.w4(32'hbc66b3c8),
	.w5(32'hbbebda32),
	.w6(32'h3d1e08f0),
	.w7(32'h3b81c63a),
	.w8(32'hbb93f02f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8da1ee),
	.w1(32'hbaeaaf30),
	.w2(32'hb81267da),
	.w3(32'hbbea5f32),
	.w4(32'hbaf0b44b),
	.w5(32'hba380ab4),
	.w6(32'hbaebb24d),
	.w7(32'hbb1308f0),
	.w8(32'hbb956fba),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdbd81),
	.w1(32'hbb82619e),
	.w2(32'hbbf004b6),
	.w3(32'h3ba4b2f3),
	.w4(32'hbbfa1a4a),
	.w5(32'hbc0d135b),
	.w6(32'h384fec86),
	.w7(32'hbc2816b2),
	.w8(32'hbc0d71f9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac469ec),
	.w1(32'hbb91c720),
	.w2(32'h3af6df6b),
	.w3(32'hbc031cef),
	.w4(32'hbc0142a3),
	.w5(32'hba868b53),
	.w6(32'hbb432882),
	.w7(32'hbacc3bb0),
	.w8(32'h3b3a10c6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94843b),
	.w1(32'h3be35d37),
	.w2(32'hbb2d2782),
	.w3(32'hbb67427a),
	.w4(32'hba8cebae),
	.w5(32'hbbeb9249),
	.w6(32'h3b8fb6be),
	.w7(32'hbb3efc0b),
	.w8(32'h3a4adee9),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45900e),
	.w1(32'h3c07ae21),
	.w2(32'h3c04d244),
	.w3(32'hbb154b28),
	.w4(32'hbb63c989),
	.w5(32'hba075082),
	.w6(32'h3adc45ea),
	.w7(32'h3ac4a209),
	.w8(32'h3bb0de87),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1696aa),
	.w1(32'hbb63c66e),
	.w2(32'h3837b563),
	.w3(32'h3bbbe359),
	.w4(32'hbb1a7fe4),
	.w5(32'h3bf98e68),
	.w6(32'h3adda67a),
	.w7(32'hba343c90),
	.w8(32'h3b48f5ff),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb858712),
	.w1(32'h3b0ec38a),
	.w2(32'h3b8b18a5),
	.w3(32'hbb9a21fe),
	.w4(32'hb79c0341),
	.w5(32'h3bb4a331),
	.w6(32'hbc05ab1c),
	.w7(32'h3a4107f2),
	.w8(32'h3b6b3fd7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc8a50),
	.w1(32'hbbb7551a),
	.w2(32'hbbac4c66),
	.w3(32'h3b3424d0),
	.w4(32'hbba40059),
	.w5(32'hba24a358),
	.w6(32'hba376f6f),
	.w7(32'h3b3d4bf7),
	.w8(32'hb9ac96aa),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a918dab),
	.w1(32'hbb32b324),
	.w2(32'h39f00638),
	.w3(32'h3a2e4963),
	.w4(32'hbb1ad198),
	.w5(32'h3b799810),
	.w6(32'hbb315435),
	.w7(32'hba21edf7),
	.w8(32'h3a77e3a9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c6467),
	.w1(32'hbbad36a9),
	.w2(32'h3ba3c0ae),
	.w3(32'h3b6277d1),
	.w4(32'hbc4c83ff),
	.w5(32'hb8c7fbb9),
	.w6(32'h3baa7996),
	.w7(32'hbbc4285f),
	.w8(32'h3b5a4c26),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff9313),
	.w1(32'h39ff1581),
	.w2(32'hbbccce47),
	.w3(32'h3aa3a66c),
	.w4(32'h3a17ae5c),
	.w5(32'hba1d4b11),
	.w6(32'h3b6ce714),
	.w7(32'h3badf570),
	.w8(32'hbb84d9fa),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90058c),
	.w1(32'h3baa3a99),
	.w2(32'h3b98ff2c),
	.w3(32'h3a402080),
	.w4(32'hbb7b935c),
	.w5(32'hbc140a83),
	.w6(32'hbb03bf88),
	.w7(32'hb9d89b68),
	.w8(32'hbb492a1c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987a30e),
	.w1(32'hbb2cc29e),
	.w2(32'hbab816f9),
	.w3(32'h3ad2da9c),
	.w4(32'hbb981f45),
	.w5(32'h3ba00daa),
	.w6(32'h3b67679c),
	.w7(32'hbb372a1a),
	.w8(32'hbaca7f10),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c199e),
	.w1(32'h3a5c8c91),
	.w2(32'hbb9ad850),
	.w3(32'hbaa598d0),
	.w4(32'h3b9a8aaa),
	.w5(32'h3ab5ad72),
	.w6(32'hbba20d5f),
	.w7(32'h3bbf5a66),
	.w8(32'h3ae45d7d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91a311),
	.w1(32'hbbb6531c),
	.w2(32'hbba44f98),
	.w3(32'h3af6e83d),
	.w4(32'hbb922dfd),
	.w5(32'hb96871fe),
	.w6(32'h3c24385f),
	.w7(32'hba9aedc2),
	.w8(32'hbbffbd4d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c4eec),
	.w1(32'h3be0a7dc),
	.w2(32'h3bf13b41),
	.w3(32'hbbe611ee),
	.w4(32'hbc730e93),
	.w5(32'hbc0f0ca8),
	.w6(32'hbb05de30),
	.w7(32'h3bcce08e),
	.w8(32'h3c10b5e5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0cfe0),
	.w1(32'h3b28032e),
	.w2(32'h3b8523fc),
	.w3(32'h3a98d733),
	.w4(32'h3b5f8f88),
	.w5(32'hbbc3f7d7),
	.w6(32'hbaff11ca),
	.w7(32'hbb5ea55a),
	.w8(32'h3a50d62c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c368f24),
	.w1(32'h3c1f8d21),
	.w2(32'h3be6e5b7),
	.w3(32'h3baee30c),
	.w4(32'hbb3a412a),
	.w5(32'h3bd81be9),
	.w6(32'h3c5fe2bc),
	.w7(32'h3acd51a4),
	.w8(32'h3bbe971b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b609a8a),
	.w1(32'hbaeef974),
	.w2(32'hbc2d0829),
	.w3(32'h3b51bcf9),
	.w4(32'h3a07eea5),
	.w5(32'hbb542020),
	.w6(32'h3b7acdb5),
	.w7(32'hbb32b9b2),
	.w8(32'hbbfb71f1),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04f5be),
	.w1(32'hbc064e50),
	.w2(32'h3a4f8ead),
	.w3(32'hbc0d175f),
	.w4(32'hbacb1c6d),
	.w5(32'h3a9ee975),
	.w6(32'hbc0251bc),
	.w7(32'h3bb37e1c),
	.w8(32'h3bf30918),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b3ea5),
	.w1(32'h3bd1baf3),
	.w2(32'h3acedfef),
	.w3(32'h3b1b2b27),
	.w4(32'h3b50ed09),
	.w5(32'h3bf7b9a9),
	.w6(32'h3ae67db6),
	.w7(32'h3bb3de1c),
	.w8(32'h3c1f678b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca4b14),
	.w1(32'hbb5cc1b6),
	.w2(32'hbbc6c99d),
	.w3(32'h3ba88c4a),
	.w4(32'h3bd36fc0),
	.w5(32'hb836810e),
	.w6(32'hbb6830a9),
	.w7(32'hbaca98f3),
	.w8(32'hbbd29b09),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb76a8),
	.w1(32'hb8967659),
	.w2(32'hbb1f9fe4),
	.w3(32'hbb4dc8f8),
	.w4(32'h3a6486ba),
	.w5(32'hbb7f97fa),
	.w6(32'h36e6d556),
	.w7(32'hb9db77e4),
	.w8(32'hbbbcd8be),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ae6f8),
	.w1(32'hbbecb2c2),
	.w2(32'hbb847c1f),
	.w3(32'h3b820f6c),
	.w4(32'hbb35a36b),
	.w5(32'h396f0b4a),
	.w6(32'h3a9e4fd0),
	.w7(32'hbaec3b93),
	.w8(32'hbba66cf8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76419f),
	.w1(32'h3b6c6ade),
	.w2(32'hbba6c62a),
	.w3(32'hbba43dbd),
	.w4(32'hb996b461),
	.w5(32'hbb920bb4),
	.w6(32'hb9cd422a),
	.w7(32'h3b1caa54),
	.w8(32'hbb81b915),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922aa21),
	.w1(32'h3b912a68),
	.w2(32'h3b6153c7),
	.w3(32'hbaa74482),
	.w4(32'hba062883),
	.w5(32'h3b4bfec1),
	.w6(32'hba87f27f),
	.w7(32'h3ab7a05a),
	.w8(32'h3b61060e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bbab4),
	.w1(32'hbbc02a9f),
	.w2(32'hbba101be),
	.w3(32'h3bd4ac95),
	.w4(32'hbaa9b2a7),
	.w5(32'hbbba5c74),
	.w6(32'h3c09a547),
	.w7(32'hb8efd322),
	.w8(32'hbbbf04d6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1000a1),
	.w1(32'hbb15da20),
	.w2(32'hbb3fab78),
	.w3(32'hbbcb1e66),
	.w4(32'h3bda451c),
	.w5(32'h3c0d527b),
	.w6(32'hbbc3cb58),
	.w7(32'h3bae243b),
	.w8(32'hb9f05cff),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc71f15),
	.w1(32'h39bcb19b),
	.w2(32'hbb3d5c31),
	.w3(32'h3b86e67a),
	.w4(32'h3b44113a),
	.w5(32'h3bedc77d),
	.w6(32'h3acef1a6),
	.w7(32'h3af10c76),
	.w8(32'h3b38699e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ce04b),
	.w1(32'hbb24a9e8),
	.w2(32'hbb6267a3),
	.w3(32'hbbcc7af8),
	.w4(32'hbb484f13),
	.w5(32'hba2d5740),
	.w6(32'h3b80d7a1),
	.w7(32'hbaf717f2),
	.w8(32'hbb6e7d74),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0095fd),
	.w1(32'hbbcdc537),
	.w2(32'h3aa1e18c),
	.w3(32'hbaafbc3f),
	.w4(32'hbc37eb8f),
	.w5(32'h3998c9bc),
	.w6(32'hb9c71f78),
	.w7(32'h3b2d1bf4),
	.w8(32'h3aa3b75e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38669a),
	.w1(32'h3bb657fb),
	.w2(32'h3b90625d),
	.w3(32'hbbadf4bb),
	.w4(32'h3c06244c),
	.w5(32'h3c25f224),
	.w6(32'hbb1f5533),
	.w7(32'h3c80dffc),
	.w8(32'h3c95eb44),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe73b1b),
	.w1(32'hbc035f97),
	.w2(32'hbbb47ead),
	.w3(32'hbb909469),
	.w4(32'hbc659a7f),
	.w5(32'hbc74c288),
	.w6(32'hbc2b475a),
	.w7(32'hbc36cc87),
	.w8(32'hbad9588f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d8628),
	.w1(32'hb9a02e84),
	.w2(32'hbbb649de),
	.w3(32'h3bf44066),
	.w4(32'hbb8edb47),
	.w5(32'hbc1cd915),
	.w6(32'h3b058a48),
	.w7(32'hbc08db23),
	.w8(32'hbc2b66a9),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4893fd),
	.w1(32'hbc334732),
	.w2(32'hbba5b05f),
	.w3(32'hbcacc30d),
	.w4(32'hbc5a9969),
	.w5(32'hbbf55505),
	.w6(32'hbc874fff),
	.w7(32'h3c017c12),
	.w8(32'hba893da1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbf8b26),
	.w1(32'hbbd9e02d),
	.w2(32'hbbdb2b49),
	.w3(32'h3bdd3653),
	.w4(32'hbbc32ee9),
	.w5(32'hbbf0470a),
	.w6(32'h3c5f8311),
	.w7(32'hbbe34e88),
	.w8(32'hbb159a5f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60e652),
	.w1(32'hbb1df381),
	.w2(32'h3b878040),
	.w3(32'hbbbbe1c6),
	.w4(32'hbb3046ff),
	.w5(32'h38865c78),
	.w6(32'hbc016281),
	.w7(32'hbbe46915),
	.w8(32'h3b24fa87),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35d23c),
	.w1(32'h39cb9ec6),
	.w2(32'hbc01de3e),
	.w3(32'h3c01fb2d),
	.w4(32'hbb2e0061),
	.w5(32'h3a85cf7b),
	.w6(32'h3c050352),
	.w7(32'hbb2ff156),
	.w8(32'hbb30936f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeaffe),
	.w1(32'h3c011a2e),
	.w2(32'h3bed881a),
	.w3(32'hbb87417c),
	.w4(32'h3bcf94ad),
	.w5(32'h3bce2696),
	.w6(32'hbb0c862e),
	.w7(32'h3bcdbde4),
	.w8(32'h3c011863),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985a273),
	.w1(32'hb9335b6b),
	.w2(32'hbb7fb11a),
	.w3(32'h3af5a3a8),
	.w4(32'h3b9c0965),
	.w5(32'h3b8e03e5),
	.w6(32'hbba255f1),
	.w7(32'h3be4fb88),
	.w8(32'h3b7c4049),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbece56e),
	.w1(32'h3b4532ca),
	.w2(32'h3b9e8618),
	.w3(32'hbb8920d6),
	.w4(32'h3a75fd27),
	.w5(32'h3c0f33fc),
	.w6(32'hbb7d1ede),
	.w7(32'hbb1ee717),
	.w8(32'h3aec9769),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de418a),
	.w1(32'h3b858f78),
	.w2(32'hbafc7ccc),
	.w3(32'hba24ef7f),
	.w4(32'hba1238c8),
	.w5(32'hbb47ec07),
	.w6(32'h3bdded6b),
	.w7(32'h3c306af2),
	.w8(32'h3ba1c94b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94ecd4),
	.w1(32'h3c36511d),
	.w2(32'h3b4bbc78),
	.w3(32'hbb0c2051),
	.w4(32'h3af6ee9e),
	.w5(32'hbb94b223),
	.w6(32'h3b8c406d),
	.w7(32'h3b08d6a4),
	.w8(32'h3b77aa4b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b260ae8),
	.w1(32'hba1e1544),
	.w2(32'h387dbee8),
	.w3(32'hbab2ced1),
	.w4(32'hba6561e3),
	.w5(32'hbbea1819),
	.w6(32'hbacb3779),
	.w7(32'h3b308879),
	.w8(32'hbb792607),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c095c),
	.w1(32'hbc7fe1a2),
	.w2(32'h3ce00f53),
	.w3(32'h3ba8548e),
	.w4(32'hbb5d369b),
	.w5(32'h3bcbd1bb),
	.w6(32'h3b962a7e),
	.w7(32'h3bafbcdb),
	.w8(32'hbc89d1f7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b03e6),
	.w1(32'h3c41102a),
	.w2(32'h3c2d66ed),
	.w3(32'hbc1a9433),
	.w4(32'hbbe7b66e),
	.w5(32'h3bb769c4),
	.w6(32'hbc992f5b),
	.w7(32'hbbc7a9b3),
	.w8(32'hbc0cc135),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a0ff5),
	.w1(32'h3a969788),
	.w2(32'h3b7a629b),
	.w3(32'h3b8158af),
	.w4(32'hbb8efec5),
	.w5(32'h3c753330),
	.w6(32'hbc166f49),
	.w7(32'h3acfb910),
	.w8(32'hbbef21b0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99348e),
	.w1(32'h3c3343fe),
	.w2(32'hbbd2ad31),
	.w3(32'hbb65a9b4),
	.w4(32'hbb421ab9),
	.w5(32'hbc8092ba),
	.w6(32'h3a35d376),
	.w7(32'hbc62cae1),
	.w8(32'hbcb5c478),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1083b),
	.w1(32'hbacaa1ea),
	.w2(32'hbbc76ea2),
	.w3(32'hbb93350e),
	.w4(32'hbba988c1),
	.w5(32'hbafa81cc),
	.w6(32'hbbb8f88f),
	.w7(32'hbb6a5559),
	.w8(32'hbb3a2685),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46014d),
	.w1(32'hbc02579f),
	.w2(32'hbc6682d4),
	.w3(32'hbb5386ee),
	.w4(32'hbcfd3ac5),
	.w5(32'hbcd851ef),
	.w6(32'h3931c7ad),
	.w7(32'h3b35a2ef),
	.w8(32'hbb01a794),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad1f6d),
	.w1(32'h3bbd38d2),
	.w2(32'hbb0005ae),
	.w3(32'hbd23035f),
	.w4(32'h3b6260b9),
	.w5(32'h3c500591),
	.w6(32'h3bf00e6c),
	.w7(32'h3b20eb80),
	.w8(32'h3c05283f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d2aca),
	.w1(32'hbb5bc4ac),
	.w2(32'hbbed4713),
	.w3(32'h3bb30d35),
	.w4(32'hbbb8a70a),
	.w5(32'hbc6ee368),
	.w6(32'h3b2da7c4),
	.w7(32'hbbbfed82),
	.w8(32'h3b6244ed),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a57e8),
	.w1(32'h3c62799c),
	.w2(32'h3d11fbf4),
	.w3(32'hbbb7d239),
	.w4(32'h3c0913b8),
	.w5(32'h3bae79cb),
	.w6(32'h3aecaf95),
	.w7(32'hbc27cd8f),
	.w8(32'hbce299c3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e9c78),
	.w1(32'hbc171242),
	.w2(32'hbc896896),
	.w3(32'hbc940b27),
	.w4(32'h3a60a986),
	.w5(32'hbc08d6df),
	.w6(32'hbc42f808),
	.w7(32'h3c1b8400),
	.w8(32'h3c5ec5da),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc507074),
	.w1(32'h3c47981a),
	.w2(32'h3c856700),
	.w3(32'hbb22e2d2),
	.w4(32'h3abafdff),
	.w5(32'hbad2c15b),
	.w6(32'hbac4edbe),
	.w7(32'hbb7d1215),
	.w8(32'hbc1fddf0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d23cd),
	.w1(32'hbd02589c),
	.w2(32'hbd861784),
	.w3(32'hbc435a98),
	.w4(32'h3b6b8818),
	.w5(32'h3b8f5a5e),
	.w6(32'h3b1b9e5a),
	.w7(32'h3d3cc270),
	.w8(32'h3d8fed2b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1772ac),
	.w1(32'h392c0676),
	.w2(32'h3b867852),
	.w3(32'h3c809d07),
	.w4(32'h3b9b68ab),
	.w5(32'h3c0840b4),
	.w6(32'h3d3c9171),
	.w7(32'h3a1e0996),
	.w8(32'h3abeeb45),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41f7d7),
	.w1(32'hb8e5f1c7),
	.w2(32'hbc08a6d5),
	.w3(32'hba4624b5),
	.w4(32'h3b2ba56a),
	.w5(32'h3ab0247d),
	.w6(32'h3b3b962c),
	.w7(32'h38c7ce8d),
	.w8(32'hbb60a8b1),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abece15),
	.w1(32'h3bc3a295),
	.w2(32'h3c919e33),
	.w3(32'hbc272213),
	.w4(32'hbc4b29c0),
	.w5(32'h3a892bfc),
	.w6(32'h3ad34833),
	.w7(32'h3c1a25ae),
	.w8(32'h3cb9798e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2e370),
	.w1(32'h3c7108ba),
	.w2(32'h3c891ba2),
	.w3(32'hba57ee03),
	.w4(32'h3b23cafe),
	.w5(32'hbb146dab),
	.w6(32'h3beb2c73),
	.w7(32'h3c5f13b9),
	.w8(32'hb9d0d9e0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f3ac6),
	.w1(32'h3c7dce1b),
	.w2(32'h3cf0ee55),
	.w3(32'hbb88eba4),
	.w4(32'hbc478f41),
	.w5(32'hbc02b6f6),
	.w6(32'h38b47cc6),
	.w7(32'hbbd5b519),
	.w8(32'h3939dbae),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc011c60),
	.w1(32'h3c2776a5),
	.w2(32'h3c521951),
	.w3(32'hbad3dda7),
	.w4(32'h3a0f184b),
	.w5(32'h3be6d353),
	.w6(32'h3af34766),
	.w7(32'hbc4af813),
	.w8(32'hbc5d0b1f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e4cc7),
	.w1(32'h3c4899f9),
	.w2(32'hbbff395e),
	.w3(32'hb9dd692f),
	.w4(32'hbb230109),
	.w5(32'h3bfe3c2f),
	.w6(32'hbc2a3142),
	.w7(32'hbaf790e3),
	.w8(32'hbc0672a1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1de2d),
	.w1(32'h3bcb78d1),
	.w2(32'h3b005973),
	.w3(32'h3ab981a1),
	.w4(32'h3aa3decc),
	.w5(32'hbc030459),
	.w6(32'h3c14fc2a),
	.w7(32'hbb0aa985),
	.w8(32'hbb1851bc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f0f4f),
	.w1(32'h3c5421d7),
	.w2(32'h3c80988b),
	.w3(32'hb9608916),
	.w4(32'hbc8fbaf1),
	.w5(32'hbb09e9a9),
	.w6(32'hbc738f9f),
	.w7(32'hbcb8da74),
	.w8(32'h3b0a9c51),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cea3d),
	.w1(32'hbbd99371),
	.w2(32'h3cd18e56),
	.w3(32'hbca0ac68),
	.w4(32'hbc179d3b),
	.w5(32'hbadd5d91),
	.w6(32'hbccd5104),
	.w7(32'hbab0406d),
	.w8(32'hbcd4a067),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9f84e),
	.w1(32'hb88c5dd8),
	.w2(32'hbae1999b),
	.w3(32'hbc68a82b),
	.w4(32'h3b1fa663),
	.w5(32'hbb7ce5f8),
	.w6(32'hbcfee33f),
	.w7(32'hbbb15a83),
	.w8(32'hba01b090),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd5e37),
	.w1(32'hbc8abb71),
	.w2(32'hbcb5a993),
	.w3(32'hbad31257),
	.w4(32'h39f0ae39),
	.w5(32'h3ad1fd46),
	.w6(32'h3c04b9c6),
	.w7(32'h3c94f03b),
	.w8(32'h3cd661e2),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06eb14),
	.w1(32'hbb7a9a16),
	.w2(32'hbc883210),
	.w3(32'hba9e45e7),
	.w4(32'hb73bf060),
	.w5(32'hbc5b6c7c),
	.w6(32'h3cfb9af7),
	.w7(32'h3c48ed2e),
	.w8(32'h3ca0ae36),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd836df),
	.w1(32'h3b21e241),
	.w2(32'hbb2595dd),
	.w3(32'h3a187285),
	.w4(32'h3bcbeb8a),
	.w5(32'h3cc14355),
	.w6(32'h3c70380c),
	.w7(32'h38e79e44),
	.w8(32'hbcb4ecf2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09d90c),
	.w1(32'h3be214e8),
	.w2(32'h3cddac72),
	.w3(32'hbbdee1e0),
	.w4(32'hbc4c2c14),
	.w5(32'h3bb93dc9),
	.w6(32'hbc56188b),
	.w7(32'hbc702ecf),
	.w8(32'hbc4c83c5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2e571),
	.w1(32'h3c8da83e),
	.w2(32'h3cc5a868),
	.w3(32'h3aa02544),
	.w4(32'hbc21131e),
	.w5(32'hbb6b8731),
	.w6(32'hbc323b71),
	.w7(32'hbc26e4b3),
	.w8(32'hbc83cee2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f9268),
	.w1(32'h3bb19663),
	.w2(32'hba8dd6cc),
	.w3(32'hbbc1baa3),
	.w4(32'hba89e349),
	.w5(32'h3b6abe98),
	.w6(32'hbc71eb0a),
	.w7(32'hbc03f8bd),
	.w8(32'h3b9e8392),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecb077),
	.w1(32'h3b820e3e),
	.w2(32'h3c35caf3),
	.w3(32'hbbb9ba77),
	.w4(32'hbbbad6c3),
	.w5(32'hbcac7c67),
	.w6(32'hbbaf87ec),
	.w7(32'h3b07bf0a),
	.w8(32'hbc35a437),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44a4a8),
	.w1(32'h3beba6b7),
	.w2(32'h3c871764),
	.w3(32'hbca1b493),
	.w4(32'hbc0da302),
	.w5(32'hbc3276db),
	.w6(32'hbc6b9f19),
	.w7(32'h3b217427),
	.w8(32'h3bb0e500),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f644c),
	.w1(32'h3c01fa32),
	.w2(32'hb9ab2179),
	.w3(32'hbaf79f15),
	.w4(32'hb81d1930),
	.w5(32'h3b34969f),
	.w6(32'hbc763719),
	.w7(32'h3b9e7fb2),
	.w8(32'h3be2a7b6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d77c1),
	.w1(32'h3bff3e35),
	.w2(32'h3cf46e39),
	.w3(32'hbb315b72),
	.w4(32'h3b42f99b),
	.w5(32'h3bdbf704),
	.w6(32'h3bca9a11),
	.w7(32'hbc398c6c),
	.w8(32'hbc899f10),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4329d3),
	.w1(32'hbaea0975),
	.w2(32'hbbfa7a84),
	.w3(32'h3a6e97f8),
	.w4(32'hbbca8494),
	.w5(32'h3c92c2eb),
	.w6(32'hbcc389cd),
	.w7(32'hbb4f126f),
	.w8(32'hbbbbd295),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be785a1),
	.w1(32'hbb2e40ae),
	.w2(32'h3c90023d),
	.w3(32'h3c0f1029),
	.w4(32'hbc30f624),
	.w5(32'hbb8c13c4),
	.w6(32'hbc4f83e0),
	.w7(32'hbc3645ab),
	.w8(32'hbc9702fd),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c500aa7),
	.w1(32'hbb64a535),
	.w2(32'hbbf65f97),
	.w3(32'hbbc0460c),
	.w4(32'hbb18399b),
	.w5(32'h3c00ae7a),
	.w6(32'hbc5b5a62),
	.w7(32'h3c0e46da),
	.w8(32'h3be70b9d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86d4bc),
	.w1(32'hbb672d1b),
	.w2(32'h3a02bf0b),
	.w3(32'h3a6050c7),
	.w4(32'hbc2641e0),
	.w5(32'hbc957d1d),
	.w6(32'h3b93cbd5),
	.w7(32'hba39e3aa),
	.w8(32'hbb488856),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95bdee),
	.w1(32'h3bb8eb49),
	.w2(32'hbb41e064),
	.w3(32'hbc0e550b),
	.w4(32'hbb30782e),
	.w5(32'hbb56cf4e),
	.w6(32'hbab2d0f8),
	.w7(32'hbafd456a),
	.w8(32'h3badc885),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf0422),
	.w1(32'hbb24b2b0),
	.w2(32'h3c500c80),
	.w3(32'h3b1203d5),
	.w4(32'hbb7726b8),
	.w5(32'hbbca0962),
	.w6(32'h3bd97089),
	.w7(32'hbbb38492),
	.w8(32'hbc1aee00),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9fd24),
	.w1(32'hba48da91),
	.w2(32'hbc1a141b),
	.w3(32'hbbc7268b),
	.w4(32'hbbc2bf97),
	.w5(32'h3b7c6a7f),
	.w6(32'hbc47e1c6),
	.w7(32'hbbfcdf4a),
	.w8(32'hbc1439b8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dab2b),
	.w1(32'h3baa2a54),
	.w2(32'h3ca0ee5d),
	.w3(32'h3b292ed3),
	.w4(32'h3b9cd452),
	.w5(32'h3c22002f),
	.w6(32'hba1c6d2c),
	.w7(32'hbabf70d6),
	.w8(32'hbc630bd6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80115c),
	.w1(32'h3c11dbdb),
	.w2(32'h3c046983),
	.w3(32'hbc5ae60b),
	.w4(32'hba570eb4),
	.w5(32'hbbcd3692),
	.w6(32'hbbfa28e4),
	.w7(32'hbc0b864c),
	.w8(32'hb9343713),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc122c21),
	.w1(32'h3c5ec357),
	.w2(32'h3c8931eb),
	.w3(32'hbb8a29c6),
	.w4(32'hbb9ab617),
	.w5(32'hba232761),
	.w6(32'hbc6e3ec7),
	.w7(32'hbc879bdb),
	.w8(32'hbcecdd4e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa457e4),
	.w1(32'h3bc3ac4b),
	.w2(32'hbc12ec52),
	.w3(32'hbca263b6),
	.w4(32'hbbcd1e3b),
	.w5(32'hbc5ecff7),
	.w6(32'hbcc28e14),
	.w7(32'h3b37f2bb),
	.w8(32'hbb60d3df),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5ba6f),
	.w1(32'hbc196505),
	.w2(32'hbb28eac7),
	.w3(32'hba89f34b),
	.w4(32'hba051bfd),
	.w5(32'h3b764297),
	.w6(32'h3a241a1c),
	.w7(32'hbb89196e),
	.w8(32'hbaead995),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef891b),
	.w1(32'hba8660ef),
	.w2(32'h3b156b17),
	.w3(32'h3c22d6db),
	.w4(32'hbba40d97),
	.w5(32'h398e22a3),
	.w6(32'hbc571473),
	.w7(32'h3bf7b7f7),
	.w8(32'h3c28183d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fcaa9),
	.w1(32'h3c02e0ee),
	.w2(32'h3c39b0df),
	.w3(32'hbb21fd2b),
	.w4(32'hbaa8f684),
	.w5(32'hbb9528a6),
	.w6(32'h3c4f0337),
	.w7(32'hbbddbd1d),
	.w8(32'hbc6a5d83),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1340ba),
	.w1(32'hbbaf23bf),
	.w2(32'h3ba6fd5b),
	.w3(32'h3b96cce2),
	.w4(32'h3b5b3d05),
	.w5(32'h3bcbbd78),
	.w6(32'hbbb12508),
	.w7(32'hb7c64622),
	.w8(32'hba15116e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae74e27),
	.w1(32'h3b3a97f6),
	.w2(32'h39a3c1f6),
	.w3(32'hbbd22a7c),
	.w4(32'h3bd78007),
	.w5(32'h3b140a2d),
	.w6(32'hbb251d18),
	.w7(32'hbad60da7),
	.w8(32'hbb8ebb1f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31063d),
	.w1(32'hbbbcee87),
	.w2(32'hbb702348),
	.w3(32'hba60a11b),
	.w4(32'hbb6f117c),
	.w5(32'h3ccb143b),
	.w6(32'hbb464e0e),
	.w7(32'hbb21b862),
	.w8(32'hb9bf4d79),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d381b),
	.w1(32'h3bae114b),
	.w2(32'h3bcfaf7c),
	.w3(32'hbb8fee3e),
	.w4(32'hbb58aa0c),
	.w5(32'hbba0b53a),
	.w6(32'hbb385aeb),
	.w7(32'hbb9bc149),
	.w8(32'hbcb0ab21),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cd319),
	.w1(32'hbc5699dd),
	.w2(32'hbc83f48d),
	.w3(32'hbb1ed164),
	.w4(32'h3b8f3b83),
	.w5(32'hbbb1f303),
	.w6(32'hbc801f91),
	.w7(32'h3c4a5de6),
	.w8(32'h3c32dea5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0720c),
	.w1(32'hba97fede),
	.w2(32'hbbb1557f),
	.w3(32'hbb120080),
	.w4(32'h3ac01cad),
	.w5(32'h3b702135),
	.w6(32'h3bd129c0),
	.w7(32'hbc8b185e),
	.w8(32'hbcc9e37c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd38dbb),
	.w1(32'h3aa6f3a9),
	.w2(32'h3b3637dd),
	.w3(32'h3bf46379),
	.w4(32'h38c72f5e),
	.w5(32'h3aa6da31),
	.w6(32'hbcad8ddb),
	.w7(32'h3b15fb8c),
	.w8(32'hbbc2261e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a197c1c),
	.w1(32'hbc3b20d3),
	.w2(32'hbc5e5c05),
	.w3(32'hbb72a44a),
	.w4(32'hbacbca58),
	.w5(32'h3b022cae),
	.w6(32'h3a82835d),
	.w7(32'hb9a674ad),
	.w8(32'h3b1d20fd),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc405da2),
	.w1(32'h3bbd333a),
	.w2(32'h3c470d62),
	.w3(32'hba99e125),
	.w4(32'h3b7b3603),
	.w5(32'h3c759a56),
	.w6(32'h3bd18cc4),
	.w7(32'hbb950562),
	.w8(32'hbc38b49b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2af6e),
	.w1(32'hba09d752),
	.w2(32'hb924e70c),
	.w3(32'hbc5304c9),
	.w4(32'hbc308a9e),
	.w5(32'h3c275e57),
	.w6(32'hbc6e0d53),
	.w7(32'hbca5ed4b),
	.w8(32'hbc4ee888),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c537c5f),
	.w1(32'h3cbb5d5c),
	.w2(32'h3d4f5742),
	.w3(32'h3a60282c),
	.w4(32'hbc1b9f28),
	.w5(32'hbbffb505),
	.w6(32'hbb8fed04),
	.w7(32'hbce03f26),
	.w8(32'hbd17fdf0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c987654),
	.w1(32'h3ab917fe),
	.w2(32'h3cd3e8d8),
	.w3(32'hbd2d5478),
	.w4(32'hbcaa88c4),
	.w5(32'hbb840614),
	.w6(32'hbd4bc483),
	.w7(32'hbc1af6be),
	.w8(32'h3c546cbb),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule