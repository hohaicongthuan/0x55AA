module layer_10_featuremap_318(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e35d82),
	.w1(32'hb9631990),
	.w2(32'hb940d3ee),
	.w3(32'h3a2def49),
	.w4(32'h39ba22b5),
	.w5(32'hba9af01a),
	.w6(32'hba203439),
	.w7(32'hb9d0d76c),
	.w8(32'hbb0259c6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d9e0f),
	.w1(32'hbb0d6cc0),
	.w2(32'hbac113f1),
	.w3(32'hbabdc25d),
	.w4(32'hbb288a65),
	.w5(32'hbac2cc9d),
	.w6(32'hbac7a303),
	.w7(32'hbb2bdc9a),
	.w8(32'hbb14721b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf0a0c),
	.w1(32'hbb2cc9d6),
	.w2(32'hbac94223),
	.w3(32'hbb11a6cc),
	.w4(32'hba91d247),
	.w5(32'h3a9a1959),
	.w6(32'hbb147fd1),
	.w7(32'hbb088803),
	.w8(32'h3a9f8191),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a427ce3),
	.w1(32'h3a99ffe2),
	.w2(32'h3ab1d66e),
	.w3(32'h3a9e3ef3),
	.w4(32'h3a128e79),
	.w5(32'h3b190e1f),
	.w6(32'h3aefd1b2),
	.w7(32'h3a0cc63f),
	.w8(32'h3b034d32),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8843db),
	.w1(32'hba530d0c),
	.w2(32'h3a25381b),
	.w3(32'h3a7340c0),
	.w4(32'h3ae4ab29),
	.w5(32'h3a8f3777),
	.w6(32'hb94bcd2e),
	.w7(32'h3a9ac6f1),
	.w8(32'h3a5448d5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a5a041),
	.w1(32'hb912f9d8),
	.w2(32'hb9907ad2),
	.w3(32'h3a27d97e),
	.w4(32'h398146ff),
	.w5(32'h381e62b6),
	.w6(32'h3a602670),
	.w7(32'h385bb5f6),
	.w8(32'hba13303b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3045c7),
	.w1(32'hbaa3f3db),
	.w2(32'hba337003),
	.w3(32'hbb1e5c27),
	.w4(32'hbb07865d),
	.w5(32'hbaf33297),
	.w6(32'hb9a3c5ad),
	.w7(32'hba218e0d),
	.w8(32'hbaf1087a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf59f1),
	.w1(32'hb9de4a99),
	.w2(32'hbbb7d4e4),
	.w3(32'hbb815965),
	.w4(32'h3abaeb08),
	.w5(32'hbb82bd11),
	.w6(32'hbb7f824f),
	.w7(32'hbaeb5a50),
	.w8(32'h3b13a006),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2d6d3),
	.w1(32'hba89af5b),
	.w2(32'hba64fb6f),
	.w3(32'hb9fc058b),
	.w4(32'hba079cc8),
	.w5(32'h3ac218ba),
	.w6(32'hb996e452),
	.w7(32'hb90d6d33),
	.w8(32'h3a574405),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81c3d8e),
	.w1(32'hb9cb86da),
	.w2(32'hba262a44),
	.w3(32'h3a387a1f),
	.w4(32'hba9a030b),
	.w5(32'hba15a98d),
	.w6(32'h3aed28ca),
	.w7(32'h3aaaaecf),
	.w8(32'h3ab472a2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50d0c6),
	.w1(32'hb800eb94),
	.w2(32'hb99400a2),
	.w3(32'h3a6ff7c6),
	.w4(32'h388b93fd),
	.w5(32'hb8913f88),
	.w6(32'h3a8649bf),
	.w7(32'hb92178be),
	.w8(32'hb9cc80b3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd1962),
	.w1(32'h3a595700),
	.w2(32'h3a2dd354),
	.w3(32'hbb045697),
	.w4(32'hbaece953),
	.w5(32'hbb426e79),
	.w6(32'hba993f9b),
	.w7(32'hba8792de),
	.w8(32'hba15db22),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb765f50),
	.w1(32'hbb24e0a4),
	.w2(32'hbb57379c),
	.w3(32'hbbad1bbd),
	.w4(32'hbb58631b),
	.w5(32'hb9eb13c5),
	.w6(32'hbb9a9eaa),
	.w7(32'hbb18598a),
	.w8(32'hba40499b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba832e8f),
	.w1(32'hb996d458),
	.w2(32'hb9aa5109),
	.w3(32'h38e948da),
	.w4(32'h39a6c698),
	.w5(32'hba8e8163),
	.w6(32'hba9dd787),
	.w7(32'h3a867519),
	.w8(32'hb963817e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c1a55),
	.w1(32'hbaa134a5),
	.w2(32'hba3c1cec),
	.w3(32'hba1fb061),
	.w4(32'hbadea4f9),
	.w5(32'h3a514a9b),
	.w6(32'h3af14250),
	.w7(32'hb9c05180),
	.w8(32'h39d9879a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391455fb),
	.w1(32'h3a47dca3),
	.w2(32'h3ae5a902),
	.w3(32'hb9591920),
	.w4(32'hbb094949),
	.w5(32'h3a921fe3),
	.w6(32'h3b064de3),
	.w7(32'h39d9921b),
	.w8(32'hb8e59be2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9942723),
	.w1(32'hba3e5360),
	.w2(32'hb9cb69f7),
	.w3(32'h3a3a092e),
	.w4(32'h38bd53a1),
	.w5(32'hbb013419),
	.w6(32'h398093f4),
	.w7(32'hb9f11e48),
	.w8(32'hbabb1cf2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c09f),
	.w1(32'hb8b8a4f8),
	.w2(32'hb9f1c542),
	.w3(32'hbb50de93),
	.w4(32'hbaa2ee8a),
	.w5(32'hbae08fbd),
	.w6(32'hbaff774b),
	.w7(32'h3b3bc932),
	.w8(32'h3af728a5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3b2fc),
	.w1(32'h39bb7151),
	.w2(32'h3aa1c2ab),
	.w3(32'hbb2ca5b8),
	.w4(32'hb9f8f261),
	.w5(32'h39d08afb),
	.w6(32'hb806ecf2),
	.w7(32'h3aa08900),
	.w8(32'h3a9ec37e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec5f9b),
	.w1(32'h391196e0),
	.w2(32'h3ad4f245),
	.w3(32'h3a721b87),
	.w4(32'h3aa6183c),
	.w5(32'h39f06d1a),
	.w6(32'h3a27efc1),
	.w7(32'h3a84e86d),
	.w8(32'h39c4ec90),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce50fb),
	.w1(32'h39989035),
	.w2(32'h38781af2),
	.w3(32'h378fad7f),
	.w4(32'hba3b21cb),
	.w5(32'h3b0adae2),
	.w6(32'hb8a77715),
	.w7(32'hba294de6),
	.w8(32'h3af8c74b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d49f3),
	.w1(32'h3aee1a9d),
	.w2(32'h3b0bec23),
	.w3(32'h3b3ac119),
	.w4(32'h3b03a11a),
	.w5(32'h39ac388f),
	.w6(32'h3b3b8afe),
	.w7(32'h3ab9a801),
	.w8(32'h39225faf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab90978),
	.w1(32'hb8d95c8a),
	.w2(32'h3b792059),
	.w3(32'hbaedadd3),
	.w4(32'hbb0fc1b7),
	.w5(32'h3b744d28),
	.w6(32'h3b2b3f09),
	.w7(32'h3b57ff1e),
	.w8(32'h3b84ef27),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a584bea),
	.w1(32'hbafae069),
	.w2(32'hbb1ce422),
	.w3(32'h3a960af5),
	.w4(32'hbb304253),
	.w5(32'hba9d0133),
	.w6(32'h3ab6041c),
	.w7(32'hba8e1961),
	.w8(32'h3a9368ae),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92a494),
	.w1(32'h3a44c986),
	.w2(32'h3ad49745),
	.w3(32'h3b3685e0),
	.w4(32'h3a20c5c4),
	.w5(32'h3b2a2cfc),
	.w6(32'h3bc68ab5),
	.w7(32'h3aca61c6),
	.w8(32'h3adc2e10),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3745cf10),
	.w1(32'h39e1a883),
	.w2(32'h3a551a2d),
	.w3(32'h39c05585),
	.w4(32'h39cea391),
	.w5(32'h391c3ce7),
	.w6(32'h3ac7f86f),
	.w7(32'h3a5cc0c6),
	.w8(32'hb9e6ebab),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfe580),
	.w1(32'hbac8a71c),
	.w2(32'hb95dcab1),
	.w3(32'hb9c73dd9),
	.w4(32'h3a31ba20),
	.w5(32'hb862bcd1),
	.w6(32'hba8601ec),
	.w7(32'hb997bfbd),
	.w8(32'hba7a2556),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1031e9),
	.w1(32'h39e26358),
	.w2(32'h3ac34e88),
	.w3(32'h3b58f2d5),
	.w4(32'h39b7ce1a),
	.w5(32'h3876a416),
	.w6(32'h37829bf4),
	.w7(32'h38ecdd58),
	.w8(32'hba435b1f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a900bbb),
	.w1(32'h39f84108),
	.w2(32'h3b02720b),
	.w3(32'h3b139010),
	.w4(32'h3a7c4002),
	.w5(32'h3a1c8f07),
	.w6(32'h3a9efadf),
	.w7(32'h3a9b2733),
	.w8(32'h395a327c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba056b4),
	.w1(32'hb9c8d943),
	.w2(32'h3a0c4618),
	.w3(32'h3b8ae089),
	.w4(32'hb98fccc3),
	.w5(32'hbafe926b),
	.w6(32'h3b9e2b88),
	.w7(32'h396ce394),
	.w8(32'hbb05dccc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05a453),
	.w1(32'hb9c382af),
	.w2(32'h3a34a5d5),
	.w3(32'hb99422d3),
	.w4(32'h39b79701),
	.w5(32'hba411506),
	.w6(32'h3a8fd163),
	.w7(32'h3a9be68d),
	.w8(32'hb934b93e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a470e6d),
	.w1(32'h3a1b551a),
	.w2(32'h39d6f20f),
	.w3(32'hb9ae5ddc),
	.w4(32'hb8cdd412),
	.w5(32'hbb0050dd),
	.w6(32'hba27886b),
	.w7(32'hba4478d9),
	.w8(32'hbab1af90),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90a8f7),
	.w1(32'hb88a1638),
	.w2(32'h3a116832),
	.w3(32'hbacb518d),
	.w4(32'hba89a136),
	.w5(32'hbab1454e),
	.w6(32'h3a372524),
	.w7(32'h3a9bf382),
	.w8(32'hb97c1812),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37524204),
	.w1(32'hba4f0d12),
	.w2(32'hbaeb284e),
	.w3(32'hba4a45c4),
	.w4(32'hbb02c6e5),
	.w5(32'h3aea802a),
	.w6(32'h3a20e345),
	.w7(32'hbab0fe8d),
	.w8(32'h3b171261),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec5ca0),
	.w1(32'h3ad99584),
	.w2(32'h3a2d0f99),
	.w3(32'h3a342b17),
	.w4(32'h399db2f1),
	.w5(32'hba6826da),
	.w6(32'h3ad37fc6),
	.w7(32'h394b32e4),
	.w8(32'h37ff54d0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fec08),
	.w1(32'hbab03e62),
	.w2(32'hbad552d3),
	.w3(32'hbb635fbe),
	.w4(32'hba9c2b40),
	.w5(32'hba336aa2),
	.w6(32'hbadc5655),
	.w7(32'hbabe3ecf),
	.w8(32'hba713389),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fef3b),
	.w1(32'h3a0ca724),
	.w2(32'h3bca8c56),
	.w3(32'hbbae1456),
	.w4(32'hbb66f3b7),
	.w5(32'h3c1eeeac),
	.w6(32'hbae87403),
	.w7(32'hbab558b1),
	.w8(32'h3c1ec6f7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cf8d8),
	.w1(32'hbb256799),
	.w2(32'h3af40cc0),
	.w3(32'h3ba3df4e),
	.w4(32'hba137d26),
	.w5(32'h3a0e623a),
	.w6(32'h3bbddb8b),
	.w7(32'hbaea316e),
	.w8(32'hba35b32d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42ac8c),
	.w1(32'hbb80424a),
	.w2(32'hba695195),
	.w3(32'h396f5852),
	.w4(32'hbb8c2bb9),
	.w5(32'h3aaf7411),
	.w6(32'h3b0e6e73),
	.w7(32'hbb8d8ca3),
	.w8(32'h39037c0e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0dafa),
	.w1(32'h3aba1126),
	.w2(32'h3a3c6eca),
	.w3(32'h3b4c5f7c),
	.w4(32'h3a185d73),
	.w5(32'h3a64c2a2),
	.w6(32'h3b3fc077),
	.w7(32'h3a21a61d),
	.w8(32'h39c8a1b5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4cb711),
	.w1(32'h39e309ad),
	.w2(32'h39d17530),
	.w3(32'h3a827914),
	.w4(32'h3a0cd1f0),
	.w5(32'h3af30b38),
	.w6(32'hb9f17fb6),
	.w7(32'h38c3912f),
	.w8(32'h3a94e510),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82ba12),
	.w1(32'h3a5b9683),
	.w2(32'h3a61f24c),
	.w3(32'h3adee5d5),
	.w4(32'h3abb8fd7),
	.w5(32'hba9f25a3),
	.w6(32'h3b23734d),
	.w7(32'h3a97cdd0),
	.w8(32'hba9660a6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac59c94),
	.w1(32'hbb092401),
	.w2(32'h380e36f2),
	.w3(32'hba190d17),
	.w4(32'hb7cfe6cc),
	.w5(32'hbae53867),
	.w6(32'hba1ed24c),
	.w7(32'h3a20073a),
	.w8(32'hbb3ef6fb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb849b7f),
	.w1(32'hbb98f5c3),
	.w2(32'hbb2c289e),
	.w3(32'hbb9a34fc),
	.w4(32'hba4d220f),
	.w5(32'hbb981e58),
	.w6(32'hbb60926a),
	.w7(32'h3b1bbdc5),
	.w8(32'hbb5aeac3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaad532),
	.w1(32'hbab4eb71),
	.w2(32'hb9106e86),
	.w3(32'h3a9cfa23),
	.w4(32'hba431453),
	.w5(32'h3a9dff8c),
	.w6(32'h3b26226f),
	.w7(32'hb9b2dfa7),
	.w8(32'h3b00d599),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d12cdd),
	.w1(32'hba8a612c),
	.w2(32'hba81db84),
	.w3(32'hb9e528d4),
	.w4(32'hbaf627ce),
	.w5(32'h3aa1fe5b),
	.w6(32'h3b6a3207),
	.w7(32'h3a7b1048),
	.w8(32'h3b5d0c94),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba2e50),
	.w1(32'hb95f1346),
	.w2(32'h3a53e3ce),
	.w3(32'h3ab74f22),
	.w4(32'hba04f8bb),
	.w5(32'h3b205ff4),
	.w6(32'h3b4c858e),
	.w7(32'h3b0d99de),
	.w8(32'h3b65fb2d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14ad67),
	.w1(32'h3b189c58),
	.w2(32'h3bb37542),
	.w3(32'hba0e5b33),
	.w4(32'h3b215b4d),
	.w5(32'hbb1fcb03),
	.w6(32'hb9fcc95a),
	.w7(32'h3b887848),
	.w8(32'hba2a9f8d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f2d51),
	.w1(32'hbb6649ef),
	.w2(32'hbb837c45),
	.w3(32'hbb84a731),
	.w4(32'hbb6bd3dd),
	.w5(32'h3b0f530b),
	.w6(32'hbb750afb),
	.w7(32'hbb56b8ca),
	.w8(32'h3aee027d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e317a),
	.w1(32'h3aa96cbc),
	.w2(32'h3a9bdc17),
	.w3(32'h3afc3a60),
	.w4(32'h3add42a8),
	.w5(32'hba00e755),
	.w6(32'h3b0c3a76),
	.w7(32'h3a91d891),
	.w8(32'hba47ec21),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b1a1e1),
	.w1(32'hba730ad2),
	.w2(32'hba88881e),
	.w3(32'hba59fd1d),
	.w4(32'h3a114b45),
	.w5(32'hba385d8b),
	.w6(32'hba1c8a46),
	.w7(32'hb9bda360),
	.w8(32'hba4bdceb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cc007),
	.w1(32'hba9a03e9),
	.w2(32'h39220742),
	.w3(32'hba41c6c5),
	.w4(32'hb9a283dd),
	.w5(32'h3ad2926c),
	.w6(32'h3ad9b2b0),
	.w7(32'h3a8acdcb),
	.w8(32'h3a6a81e6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387ff897),
	.w1(32'hb9cc6320),
	.w2(32'hb9b87023),
	.w3(32'h3b00a550),
	.w4(32'h3ad2cfc0),
	.w5(32'h39c18164),
	.w6(32'h3a1c7cb6),
	.w7(32'h3997045b),
	.w8(32'h39965d79),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10bd7b),
	.w1(32'hba014d0a),
	.w2(32'h3a675f1b),
	.w3(32'hbb5aa7e7),
	.w4(32'hbaee8380),
	.w5(32'hba9b2a3e),
	.w6(32'hbb7e2225),
	.w7(32'h3a1c2e8b),
	.w8(32'h3b2eee9f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a408172),
	.w1(32'h3a9576be),
	.w2(32'h3aa89fd7),
	.w3(32'h3a7e1362),
	.w4(32'h3ac5b9dc),
	.w5(32'hb9447833),
	.w6(32'h3ac2e035),
	.w7(32'h3ab422e2),
	.w8(32'h3a867dcc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a3444),
	.w1(32'h39f47e20),
	.w2(32'hb9fa2dca),
	.w3(32'hb9b5f36e),
	.w4(32'hba3d533c),
	.w5(32'h39a2a449),
	.w6(32'h39d47b76),
	.w7(32'hba4978a2),
	.w8(32'h3a09d5bd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c298e4),
	.w1(32'h3a1ff82f),
	.w2(32'h3a48e4f9),
	.w3(32'hb953d916),
	.w4(32'h397e6abc),
	.w5(32'h39883e87),
	.w6(32'hb8cf2bd8),
	.w7(32'h399613ea),
	.w8(32'hb74e642f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bb947),
	.w1(32'h390a9618),
	.w2(32'hb8ecc6b1),
	.w3(32'h3a8cda0d),
	.w4(32'h3a331f4c),
	.w5(32'h3a7ee6a9),
	.w6(32'h3a09de51),
	.w7(32'hba048fd1),
	.w8(32'h3956e122),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00aa0a),
	.w1(32'h39e770ca),
	.w2(32'h3a83ddd5),
	.w3(32'h3b007107),
	.w4(32'h3acabcc6),
	.w5(32'h3b2c4e0b),
	.w6(32'h3b08af61),
	.w7(32'h3a85a6a9),
	.w8(32'h3b438c22),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9954c),
	.w1(32'h3a7d2cef),
	.w2(32'h3a781746),
	.w3(32'h3ab8fc01),
	.w4(32'h3ab4cd69),
	.w5(32'hba1094a7),
	.w6(32'h3aeab575),
	.w7(32'h3ad47161),
	.w8(32'hb9d5f79b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5442a),
	.w1(32'hba06cd1d),
	.w2(32'hba4f4499),
	.w3(32'hbaa0e3d8),
	.w4(32'hb9a0af65),
	.w5(32'hb9dff5eb),
	.w6(32'hba80bc71),
	.w7(32'h3a4d190a),
	.w8(32'h39aa0de3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ebf6d),
	.w1(32'h398f26a4),
	.w2(32'h3a1291e5),
	.w3(32'h38b195fd),
	.w4(32'hba6ff4c0),
	.w5(32'h39342f72),
	.w6(32'h3b31476c),
	.w7(32'h3ac3b46c),
	.w8(32'h39dc02c5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f57aa),
	.w1(32'hb98c0261),
	.w2(32'hb90fe986),
	.w3(32'hb9abf88e),
	.w4(32'h3a4e8a0b),
	.w5(32'h39fc8a23),
	.w6(32'h3a4f92c1),
	.w7(32'h3a0613ef),
	.w8(32'h3a4ba98f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dc72d),
	.w1(32'h395884a2),
	.w2(32'hb99d9ed1),
	.w3(32'hba51cd47),
	.w4(32'hba8ed66d),
	.w5(32'h3a729fbd),
	.w6(32'hba5c99a5),
	.w7(32'hbaacbcda),
	.w8(32'h3ac29ce3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9e70f),
	.w1(32'h37a45f9e),
	.w2(32'hb9fe0695),
	.w3(32'hb99f0bcd),
	.w4(32'hb9435e8c),
	.w5(32'h3a6ea6ae),
	.w6(32'hba0c8c6f),
	.w7(32'hba808157),
	.w8(32'h3aa36596),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a826de4),
	.w1(32'h3a68d3e4),
	.w2(32'h3aa7b661),
	.w3(32'h3a5a2608),
	.w4(32'h3ad78f4e),
	.w5(32'h3a2f3405),
	.w6(32'h3abad029),
	.w7(32'h3abfda23),
	.w8(32'h3a610caa),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab07a1d),
	.w1(32'h3b3257fc),
	.w2(32'h3b154d4d),
	.w3(32'hbac03c05),
	.w4(32'hb936ca05),
	.w5(32'hbb193183),
	.w6(32'h3a8cda8b),
	.w7(32'h3b876986),
	.w8(32'h3a922e16),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb100906),
	.w1(32'hbaf61150),
	.w2(32'hba2182df),
	.w3(32'hbb46ad4a),
	.w4(32'h3961615e),
	.w5(32'h3abd847c),
	.w6(32'hbaefbf0f),
	.w7(32'h3a85d0ce),
	.w8(32'h3b9261ec),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af73e32),
	.w1(32'hb908ef5f),
	.w2(32'hb885e6c9),
	.w3(32'h3b5a2bac),
	.w4(32'h3b250155),
	.w5(32'hbb43d7fd),
	.w6(32'h3b8a1c12),
	.w7(32'h3b8aca70),
	.w8(32'hb866d244),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38f403),
	.w1(32'hbb25835a),
	.w2(32'h385e92b0),
	.w3(32'h3a80ae7b),
	.w4(32'hbacf886e),
	.w5(32'h3b30f14f),
	.w6(32'h3ba99ca9),
	.w7(32'hb9c4bda1),
	.w8(32'h3aa5269d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39114273),
	.w1(32'h39581291),
	.w2(32'h3a3ff8b9),
	.w3(32'h391c8c3a),
	.w4(32'h39c3a4ef),
	.w5(32'hb94eb640),
	.w6(32'hb7e777dc),
	.w7(32'h39c3d305),
	.w8(32'hba5a3ea3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba469db2),
	.w1(32'h392f6b2c),
	.w2(32'hbae4997c),
	.w3(32'hba36c9d1),
	.w4(32'hba76bf8d),
	.w5(32'hbab1b381),
	.w6(32'hb939a9e9),
	.w7(32'hbaed21fe),
	.w8(32'hbb0d99b4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba757b5a),
	.w1(32'hbb13660b),
	.w2(32'hba68067f),
	.w3(32'hbaef3a00),
	.w4(32'hbabfccd8),
	.w5(32'hbb09fb28),
	.w6(32'hbb21bd0e),
	.w7(32'hbb280e86),
	.w8(32'hbb207b85),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33df59),
	.w1(32'hbb0965e4),
	.w2(32'hbad38255),
	.w3(32'hbb4d1b0e),
	.w4(32'hbb03a9b8),
	.w5(32'h3a88fffe),
	.w6(32'hbb3e540e),
	.w7(32'hbb1537f6),
	.w8(32'h3aa93201),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39740d38),
	.w1(32'hb9633328),
	.w2(32'hb889d2d7),
	.w3(32'h3a4daa08),
	.w4(32'h3a206069),
	.w5(32'hbb6149f8),
	.w6(32'h39077e24),
	.w7(32'hb978737d),
	.w8(32'hbb329ca8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947d2e),
	.w1(32'hbae6d5fa),
	.w2(32'hba13c681),
	.w3(32'hbb976421),
	.w4(32'hbb4d2ccc),
	.w5(32'h3a0ccdda),
	.w6(32'hbb7c0d25),
	.w7(32'hbb200653),
	.w8(32'h3b05c424),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb186870),
	.w1(32'hba0dac8e),
	.w2(32'h3aec63e3),
	.w3(32'hbab25a0c),
	.w4(32'h399c11f9),
	.w5(32'hb9c69044),
	.w6(32'hbabc98e5),
	.w7(32'h3a8af377),
	.w8(32'h3b410e10),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98db9f),
	.w1(32'h397b101a),
	.w2(32'h3b07c361),
	.w3(32'hb8ad857e),
	.w4(32'hb9d9a776),
	.w5(32'h3b5991d3),
	.w6(32'h3b05ba53),
	.w7(32'hb976a6b7),
	.w8(32'h3b4e0bf6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f13b5),
	.w1(32'h3a069357),
	.w2(32'hba616cf6),
	.w3(32'h3ae4e911),
	.w4(32'h399b85f2),
	.w5(32'hbac2d363),
	.w6(32'h3afe76cd),
	.w7(32'h3b006e48),
	.w8(32'hba2254a2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb338310),
	.w1(32'hba46d80f),
	.w2(32'hba10962d),
	.w3(32'hbb0e01e3),
	.w4(32'hbb163ee9),
	.w5(32'hba5b6d3f),
	.w6(32'hb98fec5b),
	.w7(32'h3a2042e4),
	.w8(32'h3a8bb432),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a007720),
	.w1(32'hba2fdaf9),
	.w2(32'hb91ac186),
	.w3(32'h3b1a3618),
	.w4(32'h3adb0c10),
	.w5(32'hbb114fc1),
	.w6(32'h3a368f87),
	.w7(32'h3a63a2b8),
	.w8(32'hbaa967a7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50eb22),
	.w1(32'hbabd1baf),
	.w2(32'hba1b9379),
	.w3(32'hbb6548ca),
	.w4(32'hbace312a),
	.w5(32'h39fe2969),
	.w6(32'hba87a42e),
	.w7(32'h39ffdd28),
	.w8(32'h3b028f13),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab66082),
	.w1(32'h3a9dcb6a),
	.w2(32'h3a82fb26),
	.w3(32'h3a65cfc7),
	.w4(32'h396ddf7e),
	.w5(32'h3b07653a),
	.w6(32'h3a5ad763),
	.w7(32'h399a151b),
	.w8(32'h3b070290),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ed25f),
	.w1(32'h3aaf6d7d),
	.w2(32'h3b105710),
	.w3(32'h3aff5c88),
	.w4(32'h3afa9e27),
	.w5(32'hba2b4fa1),
	.w6(32'h3a7ef382),
	.w7(32'h3a667138),
	.w8(32'hb7c8af23),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996c236),
	.w1(32'h3896632b),
	.w2(32'h39dc9b1e),
	.w3(32'hba2b283d),
	.w4(32'hba6ec4ca),
	.w5(32'h3a9748ac),
	.w6(32'hb8f564f2),
	.w7(32'hb9ed0bee),
	.w8(32'h3ab81fd2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab11083),
	.w1(32'h3a75ef92),
	.w2(32'h3a8539c3),
	.w3(32'h3a76909f),
	.w4(32'h3a8239c5),
	.w5(32'hbad60418),
	.w6(32'h3adf5e49),
	.w7(32'h3ab76f1e),
	.w8(32'hbb4b079d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba431d34),
	.w1(32'hbb7129ec),
	.w2(32'hbad7d280),
	.w3(32'hb9c69375),
	.w4(32'hb9fbbcdf),
	.w5(32'h3b26b197),
	.w6(32'h39a6a193),
	.w7(32'hbb0f94c9),
	.w8(32'h3ac3dfdb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88eb933),
	.w1(32'h3951cf93),
	.w2(32'h3ae31b66),
	.w3(32'h39fe367b),
	.w4(32'h3a1a6920),
	.w5(32'h39302e2a),
	.w6(32'h39fd6f2e),
	.w7(32'h3aa89c99),
	.w8(32'hb9ab1512),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcbe90),
	.w1(32'hbb2a0e98),
	.w2(32'hbab242f8),
	.w3(32'h3909c09c),
	.w4(32'hb9faf5b2),
	.w5(32'h3b247da3),
	.w6(32'h39ed2f9d),
	.w7(32'hb9ec91a9),
	.w8(32'h3b2ade5e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba394abf),
	.w1(32'h3b233695),
	.w2(32'h3ab0768e),
	.w3(32'h3ae2db06),
	.w4(32'h3b299310),
	.w5(32'hbab00aba),
	.w6(32'h3b2a1a8c),
	.w7(32'h3bb4320e),
	.w8(32'h3b02973d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33f8b9),
	.w1(32'hba177ede),
	.w2(32'h3a43d165),
	.w3(32'h3ac82545),
	.w4(32'hbac4bee6),
	.w5(32'h3aa11203),
	.w6(32'h3accece0),
	.w7(32'hba74616a),
	.w8(32'h3985c0e9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb970e97),
	.w1(32'h3b03e64a),
	.w2(32'h3be20ef8),
	.w3(32'hbbc49a76),
	.w4(32'hb9bd2455),
	.w5(32'h3b4429e0),
	.w6(32'hb9a5d807),
	.w7(32'h3b87b310),
	.w8(32'h3988babb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a16eb7),
	.w1(32'hbb9c0a82),
	.w2(32'hbb25e030),
	.w3(32'h3aaa020e),
	.w4(32'hba1c8585),
	.w5(32'hba9c6192),
	.w6(32'hbb3a9812),
	.w7(32'hbb41536c),
	.w8(32'hb9d5dee4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaca5e),
	.w1(32'hb6bb9dad),
	.w2(32'hbafdd1e5),
	.w3(32'hba7b5dfe),
	.w4(32'hbada43b5),
	.w5(32'hbacec338),
	.w6(32'h3b2917c3),
	.w7(32'h3b3a13a9),
	.w8(32'h39f1d064),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3faec3),
	.w1(32'h3b15184b),
	.w2(32'h3b00283a),
	.w3(32'h3ace1f73),
	.w4(32'h3b1a79df),
	.w5(32'h38aec4d0),
	.w6(32'h3b747e93),
	.w7(32'h3b4a488c),
	.w8(32'h3a5e994d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4cf47),
	.w1(32'hbafefcdd),
	.w2(32'h389f6cf3),
	.w3(32'h3adf04ca),
	.w4(32'hbadcd976),
	.w5(32'h3abd9e2c),
	.w6(32'h3b1a0ca3),
	.w7(32'hba62698b),
	.w8(32'h3adb0ba3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83bb47),
	.w1(32'h3b1b207c),
	.w2(32'h3ac1294c),
	.w3(32'h3b164a9f),
	.w4(32'h3a65d8bb),
	.w5(32'h3a2ddb30),
	.w6(32'h3b2c877e),
	.w7(32'h3aee1669),
	.w8(32'hba23aabc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba066ebb),
	.w1(32'hba439e5c),
	.w2(32'hba8b210b),
	.w3(32'hba8e24c5),
	.w4(32'hbac23ae5),
	.w5(32'hbb3adaec),
	.w6(32'hba943910),
	.w7(32'h3aefa0be),
	.w8(32'hbada63bc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d6f7),
	.w1(32'hbb0fbba8),
	.w2(32'h3a638a40),
	.w3(32'hbba8dc7c),
	.w4(32'hbb2ec79b),
	.w5(32'hbacb57c7),
	.w6(32'hbb4e2d28),
	.w7(32'hb880b711),
	.w8(32'h3a94258b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e2dc4),
	.w1(32'h3a002328),
	.w2(32'h3b016618),
	.w3(32'hbb92d01d),
	.w4(32'hba7b7247),
	.w5(32'h3c0351c3),
	.w6(32'hbbb91e43),
	.w7(32'hbbca5cd5),
	.w8(32'h3bc1f05c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f7a74),
	.w1(32'h3a26117d),
	.w2(32'hba889435),
	.w3(32'h3a641578),
	.w4(32'hbb90b716),
	.w5(32'h3a335fa2),
	.w6(32'h3b2b7cdc),
	.w7(32'hbb9310ef),
	.w8(32'h3b062e55),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2459d0),
	.w1(32'hba42aad1),
	.w2(32'hb75ff427),
	.w3(32'h3a9b5481),
	.w4(32'hba9e7e7e),
	.w5(32'h3add8e94),
	.w6(32'h3b19d6be),
	.w7(32'hb8a68d84),
	.w8(32'h3b003b73),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8231d5),
	.w1(32'h36df8cec),
	.w2(32'h3b17d55f),
	.w3(32'hbb503660),
	.w4(32'hba379f92),
	.w5(32'h3b283d3e),
	.w6(32'hba33652f),
	.w7(32'h39a67942),
	.w8(32'h3b9493e2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c70d3),
	.w1(32'h3b0285b0),
	.w2(32'h39f1fc53),
	.w3(32'h3b00f4e5),
	.w4(32'h3a10986e),
	.w5(32'hb9796be0),
	.w6(32'h3a8ac4f4),
	.w7(32'h3ab6b64c),
	.w8(32'h3a13874b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb8904),
	.w1(32'h3b6ea7fe),
	.w2(32'h3b5646ec),
	.w3(32'hbb819d19),
	.w4(32'h3baf2489),
	.w5(32'h3b4fbe83),
	.w6(32'hbaf760d4),
	.w7(32'h3a05c292),
	.w8(32'h3c011581),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8f49e),
	.w1(32'hba68a761),
	.w2(32'hbacb2191),
	.w3(32'hbaf884c4),
	.w4(32'hbad5ac72),
	.w5(32'hbabf4e98),
	.w6(32'hbb26f1d3),
	.w7(32'hbb129d4e),
	.w8(32'hbac30237),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e235e),
	.w1(32'hba1cd124),
	.w2(32'hba056a7e),
	.w3(32'hbaa373ff),
	.w4(32'hba92194f),
	.w5(32'h3a341ba3),
	.w6(32'hba6d5abc),
	.w7(32'hb8301323),
	.w8(32'hb9afb44b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910eff2),
	.w1(32'h39fcdf77),
	.w2(32'h3ab10d41),
	.w3(32'h3a35b632),
	.w4(32'h3a2ffba1),
	.w5(32'hbaac5f67),
	.w6(32'h3abd766c),
	.w7(32'h3a2c13c8),
	.w8(32'hbb3edb83),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4970d6),
	.w1(32'hbb5c9520),
	.w2(32'hbae28f28),
	.w3(32'hbb417ed3),
	.w4(32'hbb0aebdf),
	.w5(32'hba0c9926),
	.w6(32'hbb658b07),
	.w7(32'hba25e7ad),
	.w8(32'h3ad08697),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26493c),
	.w1(32'hba2537c2),
	.w2(32'h3a423d86),
	.w3(32'h3a66f63b),
	.w4(32'hb83f6049),
	.w5(32'hbb14cbfa),
	.w6(32'h3b067ee6),
	.w7(32'h3a90f522),
	.w8(32'h3924e606),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41af61),
	.w1(32'hbaf1df64),
	.w2(32'hbb24f88c),
	.w3(32'hbadb80e9),
	.w4(32'hbb05366d),
	.w5(32'hba78229c),
	.w6(32'h3a1e0bf6),
	.w7(32'hbb7b5ec6),
	.w8(32'hb8531bc0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a8989a),
	.w1(32'hbac8344a),
	.w2(32'h39b423da),
	.w3(32'h3914dd76),
	.w4(32'hbab7b527),
	.w5(32'h36dc9a82),
	.w6(32'h3ac484d0),
	.w7(32'hba6716e0),
	.w8(32'h3a87eb13),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf45aea),
	.w1(32'hbabe59d1),
	.w2(32'h3b19e7bb),
	.w3(32'hbb823f65),
	.w4(32'hba7b07dd),
	.w5(32'h3aaa9206),
	.w6(32'hbaba35c7),
	.w7(32'hba605892),
	.w8(32'h3b0df8b8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfa539),
	.w1(32'h3ac44cd4),
	.w2(32'h3b1ae176),
	.w3(32'h3a3bb7ba),
	.w4(32'h3a448e79),
	.w5(32'h3ab3dc43),
	.w6(32'h3b412a17),
	.w7(32'h3b6d3273),
	.w8(32'h3b20a14f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff1aa7),
	.w1(32'hba262bb5),
	.w2(32'h39da16e0),
	.w3(32'hbb0fd145),
	.w4(32'hba0e4a83),
	.w5(32'hba0c4f7f),
	.w6(32'h3a50eb6c),
	.w7(32'hba03c61b),
	.w8(32'h3a06f152),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2e42c),
	.w1(32'hbaa8d407),
	.w2(32'hb94d9056),
	.w3(32'hbaadfcfd),
	.w4(32'hb91852f0),
	.w5(32'hba5b3a19),
	.w6(32'hba5a86d6),
	.w7(32'hb9cb7295),
	.w8(32'hba383241),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a6b5e),
	.w1(32'h37ced518),
	.w2(32'h39b25728),
	.w3(32'hba9e9bc9),
	.w4(32'hba47b521),
	.w5(32'h3b42d290),
	.w6(32'h3938626c),
	.w7(32'hb9ce153d),
	.w8(32'h3b0952b9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67a500),
	.w1(32'h3a3ce0e3),
	.w2(32'h3a114052),
	.w3(32'h3aa6bb14),
	.w4(32'h3ac2e3d7),
	.w5(32'hb9d4255b),
	.w6(32'h3b1d4dc0),
	.w7(32'h3aad536c),
	.w8(32'h39eb4828),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398594a8),
	.w1(32'hba9dd9fe),
	.w2(32'hb964ab10),
	.w3(32'hba8cb254),
	.w4(32'h39c2965a),
	.w5(32'hbb418ef5),
	.w6(32'hba6e2fd4),
	.w7(32'hb9aa2a90),
	.w8(32'hbba2d79f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdbe74),
	.w1(32'hbb9d1c22),
	.w2(32'hbb966b7c),
	.w3(32'hbb8353ff),
	.w4(32'hbba19bcc),
	.w5(32'hbaa2ad53),
	.w6(32'hbba4b144),
	.w7(32'hbba5c46d),
	.w8(32'hb9fb6033),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba120d23),
	.w1(32'hb936a4fe),
	.w2(32'hb960d66e),
	.w3(32'h39d4c15e),
	.w4(32'h3a8ed7f7),
	.w5(32'hba9046b1),
	.w6(32'hba8a45f4),
	.w7(32'hb9ff011e),
	.w8(32'hbad984be),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33f8f8),
	.w1(32'hbaa4e43d),
	.w2(32'h3a84f6ff),
	.w3(32'hbab47a7d),
	.w4(32'hba5b545f),
	.w5(32'h39fc3b84),
	.w6(32'hbaa1ecb2),
	.w7(32'h3a0ae33b),
	.w8(32'h3ab33b5c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c99a2),
	.w1(32'hb9aa211b),
	.w2(32'h3ada71ea),
	.w3(32'h3b1f2af0),
	.w4(32'h39408390),
	.w5(32'h3b0dbc4a),
	.w6(32'h3a236bbc),
	.w7(32'hbb16de37),
	.w8(32'h3a0b6b3e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77f628),
	.w1(32'h3a504611),
	.w2(32'hb98fe5b3),
	.w3(32'h3a13e245),
	.w4(32'h39bc198a),
	.w5(32'h3a8af420),
	.w6(32'h39c32319),
	.w7(32'h39eaf990),
	.w8(32'h3ad30e2b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5507d5),
	.w1(32'h3a509072),
	.w2(32'h3ac7ee54),
	.w3(32'h39a30e6f),
	.w4(32'h3a146b0f),
	.w5(32'h3a8a98c2),
	.w6(32'hb9c0ebd2),
	.w7(32'h3a6fb58c),
	.w8(32'h398abc0c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2c70a),
	.w1(32'h3ab1dac8),
	.w2(32'h3ae139d5),
	.w3(32'h3ab8c558),
	.w4(32'h3af8d369),
	.w5(32'h3a798d8b),
	.w6(32'h39eba01f),
	.w7(32'h3b155519),
	.w8(32'hb9606cba),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5380fc),
	.w1(32'h38afdbaf),
	.w2(32'h3a1618f3),
	.w3(32'h3a3114ac),
	.w4(32'h3a5d863f),
	.w5(32'h3a0aefe0),
	.w6(32'h3ab617c5),
	.w7(32'h3a307492),
	.w8(32'hbab8a3be),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a5ab2),
	.w1(32'hbb958515),
	.w2(32'hbb4269c1),
	.w3(32'hbb9b2721),
	.w4(32'hbb339ee6),
	.w5(32'hb87d593a),
	.w6(32'hbb34fcd1),
	.w7(32'hbab11f40),
	.w8(32'h3b52bf06),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa6709),
	.w1(32'h3981f1a6),
	.w2(32'h39273246),
	.w3(32'hba1f82f3),
	.w4(32'h39970450),
	.w5(32'h39277d0d),
	.w6(32'hba5200dd),
	.w7(32'h3b314792),
	.w8(32'h3b1e6af4),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e8db8),
	.w1(32'h3a91f37e),
	.w2(32'h3ac7dd0d),
	.w3(32'h39be9b74),
	.w4(32'h3a47abcd),
	.w5(32'hba699e09),
	.w6(32'h3ac9536d),
	.w7(32'h3a8ad554),
	.w8(32'h393c8fe8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5df444),
	.w1(32'hba41580b),
	.w2(32'hba25b933),
	.w3(32'hba258c93),
	.w4(32'h39a1b8dd),
	.w5(32'h39858294),
	.w6(32'h39dbb7ea),
	.w7(32'hba4f39a7),
	.w8(32'h3afe8449),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98f5df),
	.w1(32'h38ea557d),
	.w2(32'hb9d2bd36),
	.w3(32'hba1de0fa),
	.w4(32'hba9d4969),
	.w5(32'h3a97645c),
	.w6(32'h3a1e109e),
	.w7(32'hbaa6f5f4),
	.w8(32'hb9c82f19),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0abd24),
	.w1(32'hbb3a8e2d),
	.w2(32'hbb1a6d94),
	.w3(32'hbb04a093),
	.w4(32'hbb04e9d3),
	.w5(32'hbad27e7b),
	.w6(32'hbb4d545d),
	.w7(32'hbae2e2b4),
	.w8(32'hb9f9d01e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cc0ba),
	.w1(32'h39a25aa4),
	.w2(32'h3a592988),
	.w3(32'hba135058),
	.w4(32'hba77ee07),
	.w5(32'h3a3472b1),
	.w6(32'h3b0378ae),
	.w7(32'hb7fd06bb),
	.w8(32'hb990049f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4295d4),
	.w1(32'h3994823a),
	.w2(32'h3adda9fa),
	.w3(32'hbb3aabb5),
	.w4(32'hba992218),
	.w5(32'hbadbe4bc),
	.w6(32'hbaa2a5db),
	.w7(32'h3a83832e),
	.w8(32'h3b309746),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e54e3),
	.w1(32'h399bd5c1),
	.w2(32'h3a1ddda0),
	.w3(32'hba0ed9a2),
	.w4(32'hbabfa32e),
	.w5(32'hb88c31d7),
	.w6(32'h3ae8aca8),
	.w7(32'h38def5e1),
	.w8(32'h3782ebe3),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb9cbe),
	.w1(32'h38c06ad7),
	.w2(32'h3af5fef5),
	.w3(32'hbb1ffee2),
	.w4(32'hb986bb77),
	.w5(32'h3a737660),
	.w6(32'h381cee57),
	.w7(32'h39b04120),
	.w8(32'h3ac76c46),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae52001),
	.w1(32'h39d11b19),
	.w2(32'h3a267328),
	.w3(32'hbb1e65c4),
	.w4(32'hb9405f25),
	.w5(32'hba9e4297),
	.w6(32'hba3ab173),
	.w7(32'h3a0a46cf),
	.w8(32'h3a8d8137),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39824ead),
	.w1(32'hb9b04047),
	.w2(32'h3a0a64b0),
	.w3(32'hba55dde4),
	.w4(32'hb9ce0b34),
	.w5(32'h3aa9dfdc),
	.w6(32'h39d739bc),
	.w7(32'hba2670c0),
	.w8(32'h3a4d7c2f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d41ec),
	.w1(32'hba49ad58),
	.w2(32'h3a2b47a6),
	.w3(32'hbad96586),
	.w4(32'hbb058ecb),
	.w5(32'hbb47d43d),
	.w6(32'hb9370ca1),
	.w7(32'hbaa1e73a),
	.w8(32'hbb4b5348),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e5b98),
	.w1(32'hbb258a38),
	.w2(32'hbb0c201e),
	.w3(32'h3a21be84),
	.w4(32'hba2da584),
	.w5(32'h3a986c15),
	.w6(32'hba0c2ae8),
	.w7(32'hba892e0d),
	.w8(32'hb9b84a9c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a95f5),
	.w1(32'hbb4107c8),
	.w2(32'h3a5f673c),
	.w3(32'h3b8d2f82),
	.w4(32'hba550408),
	.w5(32'hbaa54368),
	.w6(32'h3b97f892),
	.w7(32'hb98b0c75),
	.w8(32'hb8b79bda),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3617824d),
	.w1(32'hba8de6cf),
	.w2(32'hbb0508d1),
	.w3(32'hba5eb4c6),
	.w4(32'hba209970),
	.w5(32'h39373652),
	.w6(32'h3aa9964e),
	.w7(32'hb97fff26),
	.w8(32'h3a8200fb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6da9c14),
	.w1(32'hb9f59cfe),
	.w2(32'h38ed5e54),
	.w3(32'hb8d97a08),
	.w4(32'h39bc86a3),
	.w5(32'h3a80871b),
	.w6(32'h3828e4e6),
	.w7(32'hb92e3314),
	.w8(32'hb88c037e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39bfaa),
	.w1(32'h3a49b2d2),
	.w2(32'h3a48bf0a),
	.w3(32'h3a8a76bb),
	.w4(32'h3a6715b5),
	.w5(32'hb9a45871),
	.w6(32'h398ec18e),
	.w7(32'h388c9097),
	.w8(32'hb8f8e284),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c6074),
	.w1(32'hba4d1c52),
	.w2(32'hba575347),
	.w3(32'hbaa05688),
	.w4(32'hba0895bf),
	.w5(32'h3a89dbf3),
	.w6(32'hba3a4b14),
	.w7(32'hba4741be),
	.w8(32'h3b4315b6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab7302),
	.w1(32'hbaaf0c65),
	.w2(32'hba4d3db7),
	.w3(32'hb888ed18),
	.w4(32'hbb041f4e),
	.w5(32'h3b14f390),
	.w6(32'h3a5fe2a9),
	.w7(32'hbaec44c9),
	.w8(32'h3ae941d0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39248684),
	.w1(32'hb90d6757),
	.w2(32'h3a6941d2),
	.w3(32'h39ffd3e6),
	.w4(32'h3a8273cb),
	.w5(32'hba2acde8),
	.w6(32'h3a810c4f),
	.w7(32'h3b202aac),
	.w8(32'h3a3c3811),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c3175),
	.w1(32'hba1c2267),
	.w2(32'hba7093b8),
	.w3(32'h39672e08),
	.w4(32'hb5a0c3a8),
	.w5(32'hb9bedbb0),
	.w6(32'hb98a8b19),
	.w7(32'hb940634e),
	.w8(32'hb96283c7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3adbf),
	.w1(32'hba43b3b3),
	.w2(32'h39299d37),
	.w3(32'hba9162b9),
	.w4(32'hbac5352c),
	.w5(32'hbabba74a),
	.w6(32'hb9e39173),
	.w7(32'h3a924674),
	.w8(32'hb91baad3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43643e),
	.w1(32'hbb035fe6),
	.w2(32'hba53e4ef),
	.w3(32'h391da4f2),
	.w4(32'hba3a10a1),
	.w5(32'hba8971cf),
	.w6(32'h389a350f),
	.w7(32'h3a13b370),
	.w8(32'hba9822a8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b226a),
	.w1(32'hba220531),
	.w2(32'h3a92c5f1),
	.w3(32'hbb12186e),
	.w4(32'hba817f4f),
	.w5(32'h3b066877),
	.w6(32'h3a6cca7b),
	.w7(32'h3aa5f87e),
	.w8(32'h3b800f03),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82f6b1),
	.w1(32'hba1a64e7),
	.w2(32'h3b1fe8b5),
	.w3(32'h3b6b3386),
	.w4(32'h383d32ee),
	.w5(32'h387ebb68),
	.w6(32'h3b7ee0d7),
	.w7(32'h3a86ac8a),
	.w8(32'hba19388a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0023e2),
	.w1(32'hb9e38b45),
	.w2(32'hbaa817ed),
	.w3(32'h371e0e2e),
	.w4(32'hb9d9387c),
	.w5(32'hb91b7bfa),
	.w6(32'h3a98f6b1),
	.w7(32'hbaeabe31),
	.w8(32'hb9295ab1),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39efe668),
	.w1(32'h3a92e401),
	.w2(32'h3a9bcc14),
	.w3(32'hb520619d),
	.w4(32'h3a0a4e79),
	.w5(32'h38236940),
	.w6(32'h390e36ca),
	.w7(32'hb889b550),
	.w8(32'h39ee3154),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed693f),
	.w1(32'hba6fc76b),
	.w2(32'h3a31c5a5),
	.w3(32'h39c2464f),
	.w4(32'h39f83431),
	.w5(32'h3a9f40f8),
	.w6(32'h3a8f8a77),
	.w7(32'h3a9e1165),
	.w8(32'h3764d95a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a8f62),
	.w1(32'h3a9a57fc),
	.w2(32'h3a867aff),
	.w3(32'h3afd3c8c),
	.w4(32'h39ba5ada),
	.w5(32'hb8b634c7),
	.w6(32'h3b20e43b),
	.w7(32'hb867109c),
	.w8(32'hbaa9da48),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ef6a9),
	.w1(32'hbacfd509),
	.w2(32'hb9f72e50),
	.w3(32'h3ae29859),
	.w4(32'h394961b1),
	.w5(32'hbb15cbb0),
	.w6(32'h3a9a7e4d),
	.w7(32'hba4b29c6),
	.w8(32'h3a8f87ce),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba081d03),
	.w1(32'h3a9c8ce1),
	.w2(32'h3b0315bf),
	.w3(32'hbb6bfbfe),
	.w4(32'hbafe0258),
	.w5(32'h397eaafd),
	.w6(32'hbac04c84),
	.w7(32'hb9b24e8d),
	.w8(32'hb95c3139),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0aecda),
	.w1(32'h3a63de3d),
	.w2(32'h38828272),
	.w3(32'hba208083),
	.w4(32'hba8a8131),
	.w5(32'h3a93231b),
	.w6(32'h399214c8),
	.w7(32'hba17dd1a),
	.w8(32'h3a9cf99c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7d230),
	.w1(32'h39d32d8f),
	.w2(32'h39cc8999),
	.w3(32'hbb3b354b),
	.w4(32'hbb0ab5fd),
	.w5(32'hbaba28dc),
	.w6(32'h3b02743f),
	.w7(32'hba945d90),
	.w8(32'h3a1131c4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa32823),
	.w1(32'hb95f301e),
	.w2(32'hba518577),
	.w3(32'hb98d21bb),
	.w4(32'hba8a430c),
	.w5(32'h3b1fd55e),
	.w6(32'h39d76fc3),
	.w7(32'hb809e115),
	.w8(32'h3b4e1799),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b590fc5),
	.w1(32'h3b17a961),
	.w2(32'h3ae17bb6),
	.w3(32'h3b59b168),
	.w4(32'h3a9680ae),
	.w5(32'hbab5e913),
	.w6(32'h3b99cf5d),
	.w7(32'h3aee0cd8),
	.w8(32'hba81eb7c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2563a),
	.w1(32'hba8dfe6e),
	.w2(32'hbaf50263),
	.w3(32'hba22dcd8),
	.w4(32'hbadfcecf),
	.w5(32'h3aea09e7),
	.w6(32'hbaa619a0),
	.w7(32'hbb1bbf40),
	.w8(32'h3b168573),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9fc55),
	.w1(32'h3ac9eedf),
	.w2(32'h3b01ac73),
	.w3(32'h3aeef43d),
	.w4(32'h3a499be9),
	.w5(32'h39d77c69),
	.w6(32'h3a17347d),
	.w7(32'h3ace615e),
	.w8(32'h39f4328b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa93345),
	.w1(32'h3ad542e0),
	.w2(32'h3a601cc1),
	.w3(32'h3a06ff10),
	.w4(32'hba20f382),
	.w5(32'hb99e4b00),
	.w6(32'h3a883105),
	.w7(32'hb83dcd6a),
	.w8(32'h3a460235),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a078200),
	.w1(32'h3a74bc09),
	.w2(32'h39a22756),
	.w3(32'hba11eea2),
	.w4(32'h39f6a9be),
	.w5(32'hb978f46f),
	.w6(32'hba35c4cf),
	.w7(32'h39be9c4f),
	.w8(32'h3944746e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc9229),
	.w1(32'h37f2cd46),
	.w2(32'hba96d405),
	.w3(32'h3af6c825),
	.w4(32'hba6ea4d5),
	.w5(32'h3982f7b6),
	.w6(32'h3b4babfd),
	.w7(32'h39d41bc0),
	.w8(32'hb9ee3791),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e3ae6),
	.w1(32'hbb0cf9d5),
	.w2(32'h3aa32fab),
	.w3(32'hbab05755),
	.w4(32'hb9c8da1a),
	.w5(32'h3a807e2b),
	.w6(32'h392e2bb6),
	.w7(32'h3b094a0a),
	.w8(32'h3b26d90b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9188629),
	.w1(32'hb9fbf681),
	.w2(32'hb90932fc),
	.w3(32'h3a87838c),
	.w4(32'h38e8a56e),
	.w5(32'h3b7ded1f),
	.w6(32'h3a98ebf1),
	.w7(32'hbae06142),
	.w8(32'h3b908e17),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac86c7),
	.w1(32'h3a8e24e0),
	.w2(32'h3ad41485),
	.w3(32'h3aa50ad0),
	.w4(32'hba154802),
	.w5(32'hbad1ed3c),
	.w6(32'h3b812f2b),
	.w7(32'h3ace7bf8),
	.w8(32'hba0a7da7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c1549),
	.w1(32'hba4e9023),
	.w2(32'h395e849b),
	.w3(32'hbbaef3e5),
	.w4(32'hbb1df809),
	.w5(32'h3968ec82),
	.w6(32'hbb36e036),
	.w7(32'hbac8e9ea),
	.w8(32'hbacd6678),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99b00e),
	.w1(32'hba7ac42a),
	.w2(32'hbb1fc452),
	.w3(32'hb91e5412),
	.w4(32'hb9f6100d),
	.w5(32'hbb0288ca),
	.w6(32'hba65a2e2),
	.w7(32'h3a060a07),
	.w8(32'hbb244af3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90ed3f),
	.w1(32'h3a9eaaa0),
	.w2(32'hb9cefd2f),
	.w3(32'h3a5a8db7),
	.w4(32'h3a172f02),
	.w5(32'hbb0b9d3e),
	.w6(32'h3b38b5bd),
	.w7(32'h3af098a3),
	.w8(32'hba126075),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f4be5),
	.w1(32'hba564892),
	.w2(32'hbb42fb09),
	.w3(32'hbb4486dc),
	.w4(32'hbb313a1d),
	.w5(32'hba342807),
	.w6(32'hbb08bd96),
	.w7(32'hbabb2950),
	.w8(32'h3ac0d3ba),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ad0d0),
	.w1(32'h3a1e9429),
	.w2(32'h3af30b46),
	.w3(32'h39a84e54),
	.w4(32'h3a8432b1),
	.w5(32'hbb2db8e7),
	.w6(32'h3a52464a),
	.w7(32'h3a9d040d),
	.w8(32'hbae22fed),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b2a23),
	.w1(32'hb9beb784),
	.w2(32'hba883f1c),
	.w3(32'hb9fc6dc2),
	.w4(32'hb9720949),
	.w5(32'hb96ebdbd),
	.w6(32'h3a42d7a5),
	.w7(32'h3abbf8dc),
	.w8(32'h3a369609),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab67d7a),
	.w1(32'h3a98cf3e),
	.w2(32'h3a430987),
	.w3(32'h3a418bee),
	.w4(32'h38503f49),
	.w5(32'h3b20de24),
	.w6(32'h3a8a7178),
	.w7(32'hb92b5009),
	.w8(32'h3abac4be),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c198d),
	.w1(32'h3a901eec),
	.w2(32'h3af0f704),
	.w3(32'h3a940022),
	.w4(32'h3a99a60e),
	.w5(32'h3b1ece5d),
	.w6(32'h3a28b901),
	.w7(32'h3a91fb1f),
	.w8(32'h3b5c6913),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b239320),
	.w1(32'h3adefeda),
	.w2(32'h3a4af39d),
	.w3(32'hbaa1f32a),
	.w4(32'hba738f99),
	.w5(32'hbb01f029),
	.w6(32'h3ad5c6c5),
	.w7(32'hb8f552f6),
	.w8(32'hbaeba23c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac48d68),
	.w1(32'hba400028),
	.w2(32'h3ae62988),
	.w3(32'hb9e94c04),
	.w4(32'hb98cbd4c),
	.w5(32'hbb034f1c),
	.w6(32'hb91982e1),
	.w7(32'h3a1a9079),
	.w8(32'hba934b5c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba882bde),
	.w1(32'hb9db9341),
	.w2(32'hba8c409b),
	.w3(32'h3a82b7d4),
	.w4(32'hb9c24852),
	.w5(32'h3a037654),
	.w6(32'h3aa066fd),
	.w7(32'hbac57b21),
	.w8(32'hba276c4c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9846313),
	.w1(32'hba500f64),
	.w2(32'hba9e7b7c),
	.w3(32'hba30a88d),
	.w4(32'hb9975cdd),
	.w5(32'h3a295d03),
	.w6(32'hba56ff7a),
	.w7(32'hba185331),
	.w8(32'hba0a07eb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73a446c),
	.w1(32'h399485e2),
	.w2(32'h3a5c91c8),
	.w3(32'h3a973cee),
	.w4(32'h3a71825d),
	.w5(32'h3a8f5a0c),
	.w6(32'h3af42979),
	.w7(32'h3ab6492a),
	.w8(32'h39a1af27),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fd0be),
	.w1(32'h3923cb4f),
	.w2(32'h3b17f3e2),
	.w3(32'h3a9ae518),
	.w4(32'h3af7c6d1),
	.w5(32'h39af0bf1),
	.w6(32'h3b85a67d),
	.w7(32'h3b9b522f),
	.w8(32'h3a4a4133),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e1ed5),
	.w1(32'hba691642),
	.w2(32'h3ac0f238),
	.w3(32'hbb717316),
	.w4(32'h39579ffc),
	.w5(32'h3b2d1f20),
	.w6(32'hbb717e87),
	.w7(32'hb8abc733),
	.w8(32'h3b2d1092),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affb826),
	.w1(32'h3add69f9),
	.w2(32'h3a7e1a3c),
	.w3(32'h3aa185aa),
	.w4(32'h399011e6),
	.w5(32'h39eb40b4),
	.w6(32'h3b0c1f0f),
	.w7(32'h39018ef9),
	.w8(32'h3ac17b0f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986ffdf),
	.w1(32'h3a4a3722),
	.w2(32'hba876ee4),
	.w3(32'hbb423f73),
	.w4(32'h39d29696),
	.w5(32'hbb5696a0),
	.w6(32'hbb504d0f),
	.w7(32'h3b8a3b54),
	.w8(32'hba612feb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b992fe9),
	.w1(32'hb9de6fbf),
	.w2(32'h3afa34d1),
	.w3(32'h3ab9283d),
	.w4(32'hb830028d),
	.w5(32'h3a912ccc),
	.w6(32'h3b828920),
	.w7(32'h3b1c31b7),
	.w8(32'h3abaf6a0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd8053),
	.w1(32'hb923392a),
	.w2(32'h39eadcc5),
	.w3(32'hbb11d7c0),
	.w4(32'hb9661474),
	.w5(32'h3aaeca9e),
	.w6(32'hb9f3222b),
	.w7(32'hba6462ca),
	.w8(32'h3b20fc75),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd3417),
	.w1(32'h3afa9591),
	.w2(32'h3a97678c),
	.w3(32'hb96d7256),
	.w4(32'hb9990a9d),
	.w5(32'h3a93fcb5),
	.w6(32'hba56a4a5),
	.w7(32'hba5e11ca),
	.w8(32'hb8859012),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba064549),
	.w1(32'h39b6ad77),
	.w2(32'h3a6cc812),
	.w3(32'h3af1ca23),
	.w4(32'h39d514df),
	.w5(32'h3a8a4628),
	.w6(32'h3b276f39),
	.w7(32'h3a99fc32),
	.w8(32'h3a43ed69),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b169c57),
	.w1(32'h3a9d6cb0),
	.w2(32'hb9ef33ad),
	.w3(32'hb5439993),
	.w4(32'hba9903e1),
	.w5(32'hb95c4b29),
	.w6(32'h3a368a37),
	.w7(32'hbaae791b),
	.w8(32'hbaace296),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9876e18),
	.w1(32'hb9437f07),
	.w2(32'hb9613f18),
	.w3(32'hbb522c23),
	.w4(32'hbad038ed),
	.w5(32'hbaf5512e),
	.w6(32'hbb8fda7d),
	.w7(32'hbb47ccc1),
	.w8(32'h3a66960c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91296ce),
	.w1(32'h3a10942c),
	.w2(32'h3a9efdfe),
	.w3(32'hbaedd81d),
	.w4(32'hb9a6f363),
	.w5(32'h3b169098),
	.w6(32'h39fad752),
	.w7(32'h3a2aa7b0),
	.w8(32'h3b1fb69a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ccf55),
	.w1(32'h3a921ecd),
	.w2(32'h3b4c4e9f),
	.w3(32'h3b236496),
	.w4(32'h3b437f57),
	.w5(32'h3a2ed55d),
	.w6(32'h3b89929c),
	.w7(32'h3b8113aa),
	.w8(32'hb9e69d64),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39ab54),
	.w1(32'hba8fcee6),
	.w2(32'hb94d0040),
	.w3(32'hba71e86e),
	.w4(32'hb9c35247),
	.w5(32'hbb0f28f8),
	.w6(32'h3a81745d),
	.w7(32'hb91782ca),
	.w8(32'hb87e41d4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab912ff),
	.w1(32'hb9bc3173),
	.w2(32'hbaf208ff),
	.w3(32'hbba788c1),
	.w4(32'hbb581f7d),
	.w5(32'h3ab3484c),
	.w6(32'hbaf5ab9b),
	.w7(32'hbb2d3fe1),
	.w8(32'h3b8b45da),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af91c02),
	.w1(32'h3a178069),
	.w2(32'h3a2c0cfe),
	.w3(32'h39a91a02),
	.w4(32'h38976607),
	.w5(32'hba5340c0),
	.w6(32'hb858eb12),
	.w7(32'hb89ced9d),
	.w8(32'hbaca1cd6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabae678),
	.w1(32'h385b0f46),
	.w2(32'hb9ae59ca),
	.w3(32'hba9a5434),
	.w4(32'hba20a2cd),
	.w5(32'h3a7610b9),
	.w6(32'hba12f617),
	.w7(32'h394ab550),
	.w8(32'h3b0a54c8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad92bf2),
	.w1(32'h3b0a1b01),
	.w2(32'h3abe02b2),
	.w3(32'h3a54505e),
	.w4(32'h3ac42d15),
	.w5(32'h3ac0c02f),
	.w6(32'h3ab3cda3),
	.w7(32'h3b4625fe),
	.w8(32'h3b0f5bda),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fa12f),
	.w1(32'h39414c39),
	.w2(32'h3a8824b4),
	.w3(32'h3acd7294),
	.w4(32'h3a2f4dd1),
	.w5(32'hb92dd064),
	.w6(32'h3b2a9bcb),
	.w7(32'h3adbda0f),
	.w8(32'hb93eba53),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8684a55),
	.w1(32'h3a6b2b4d),
	.w2(32'h3ac9084d),
	.w3(32'h3a2a4c08),
	.w4(32'h397e4a71),
	.w5(32'hbad3bdd2),
	.w6(32'h3acf37df),
	.w7(32'h3ad46a5c),
	.w8(32'hba323ef9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91eba56),
	.w1(32'hba7c9f66),
	.w2(32'h3a32fa8a),
	.w3(32'h3b16ae93),
	.w4(32'h39fd3514),
	.w5(32'h3abb14ad),
	.w6(32'h3b582997),
	.w7(32'h3aa3094d),
	.w8(32'h3a3147f9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ccc5b),
	.w1(32'hbad4ec1b),
	.w2(32'hb6b37ba2),
	.w3(32'h3ac2111e),
	.w4(32'h39e37517),
	.w5(32'hb8b8158f),
	.w6(32'h3a996089),
	.w7(32'h39a5807b),
	.w8(32'hba278821),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa1a50),
	.w1(32'hbafe063e),
	.w2(32'hbaf58630),
	.w3(32'hbb21da5b),
	.w4(32'hbadee350),
	.w5(32'hbae3c7b2),
	.w6(32'hbb3e7556),
	.w7(32'hbb3d9b0c),
	.w8(32'hba543bdf),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf2853),
	.w1(32'hba8e9f4c),
	.w2(32'h3896421f),
	.w3(32'hba9c5300),
	.w4(32'hba816132),
	.w5(32'h39aa682f),
	.w6(32'h3adc5771),
	.w7(32'h3a4f8a56),
	.w8(32'h3a9dcaec),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7f656),
	.w1(32'h37a751f2),
	.w2(32'h3a4a1e47),
	.w3(32'hbb05a07c),
	.w4(32'hba1c73ae),
	.w5(32'hba8ddb1b),
	.w6(32'h3943925e),
	.w7(32'h3ac34180),
	.w8(32'hba3e78a1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0814a5),
	.w1(32'hbb45ed7f),
	.w2(32'hbb0a5317),
	.w3(32'hb70db336),
	.w4(32'h37c2db59),
	.w5(32'hba5eea17),
	.w6(32'h3a5b1de0),
	.w7(32'h3a9faefb),
	.w8(32'h3abb73ad),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939ea84),
	.w1(32'hba6bc305),
	.w2(32'hb9c18b2f),
	.w3(32'h381574bd),
	.w4(32'hb82bf7a1),
	.w5(32'hb9d06925),
	.w6(32'h39a21b09),
	.w7(32'hb7b446a6),
	.w8(32'hb8e7c35b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a57d1b),
	.w1(32'h3910b4f4),
	.w2(32'h3a932a46),
	.w3(32'h3a81aca7),
	.w4(32'h37f8103d),
	.w5(32'h3b048932),
	.w6(32'h3a4f044a),
	.w7(32'h39c4391a),
	.w8(32'h3aec66d2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf8396),
	.w1(32'h3b28d0e9),
	.w2(32'h3b856493),
	.w3(32'h3a6cf21b),
	.w4(32'h3b27f8e2),
	.w5(32'h3a9f25dd),
	.w6(32'h3b92e129),
	.w7(32'h3b7b05a1),
	.w8(32'h3b49df74),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369bbe3c),
	.w1(32'hbaafb630),
	.w2(32'h3a040c84),
	.w3(32'h39aa781c),
	.w4(32'hba301cb1),
	.w5(32'hba142f91),
	.w6(32'h3b08a9cd),
	.w7(32'h3b684756),
	.w8(32'h3b1f8b3c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44b3de),
	.w1(32'h3a89cc2e),
	.w2(32'h3a968c5a),
	.w3(32'h3ab1aa35),
	.w4(32'h3a2ea56a),
	.w5(32'hbacc56ba),
	.w6(32'h3b1e0a76),
	.w7(32'h3b1d1984),
	.w8(32'h3ad53b33),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb717602),
	.w1(32'h3a8b8d98),
	.w2(32'h3a76b274),
	.w3(32'hbba5f55b),
	.w4(32'hbb1acb9e),
	.w5(32'h3ae8d052),
	.w6(32'hba372d70),
	.w7(32'hbab5d1ab),
	.w8(32'h3b643573),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6a770),
	.w1(32'h3a247663),
	.w2(32'h3a66ec43),
	.w3(32'h39ca6fe7),
	.w4(32'h3a99a440),
	.w5(32'hba200b80),
	.w6(32'hba8d9fb6),
	.w7(32'h3a309079),
	.w8(32'hb9f5953d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f2a08),
	.w1(32'h39ff2fb0),
	.w2(32'h3995aa05),
	.w3(32'hbabca572),
	.w4(32'hba04062c),
	.w5(32'h3a076fad),
	.w6(32'h391c775d),
	.w7(32'hb879ad44),
	.w8(32'hba207f18),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb542c1),
	.w1(32'hbaec607a),
	.w2(32'h3b0e4483),
	.w3(32'hbabe0f8c),
	.w4(32'hba7d5917),
	.w5(32'h3b69e420),
	.w6(32'hbb2bd4bf),
	.w7(32'hbba2b6ed),
	.w8(32'h3b0342f1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb804bbb),
	.w1(32'h38c3ba1a),
	.w2(32'hba60dd2e),
	.w3(32'hba1d6c6a),
	.w4(32'hba657419),
	.w5(32'hbab1b91b),
	.w6(32'h36debd96),
	.w7(32'h3b006418),
	.w8(32'hbaa02a12),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba29aba),
	.w1(32'hbb6fbb06),
	.w2(32'h3a83c23f),
	.w3(32'hbb9fff57),
	.w4(32'h3a85ec93),
	.w5(32'h3b63f846),
	.w6(32'hbb9675be),
	.w7(32'hba86abb3),
	.w8(32'h3b22f0aa),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17e58c),
	.w1(32'hba88b8a3),
	.w2(32'h386b3b0c),
	.w3(32'h399782f4),
	.w4(32'hba19d8f2),
	.w5(32'h3aaaf7dd),
	.w6(32'h3a68882c),
	.w7(32'hbb22268c),
	.w8(32'h3af0af8e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b756a),
	.w1(32'hb9d56087),
	.w2(32'h3a40dcf8),
	.w3(32'h3aaae155),
	.w4(32'hba3fc61e),
	.w5(32'h3b118616),
	.w6(32'h3b6ac690),
	.w7(32'h398e0eb4),
	.w8(32'h3a9f9bc6),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43c895),
	.w1(32'h3a7cd1f3),
	.w2(32'h39a8a72b),
	.w3(32'h3a563ab9),
	.w4(32'h3a088f71),
	.w5(32'h3b84e921),
	.w6(32'h3ae22b6a),
	.w7(32'h39488d85),
	.w8(32'h3b2ed745),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44ef02),
	.w1(32'h3b8b8f54),
	.w2(32'h3b824e23),
	.w3(32'hba4043d9),
	.w4(32'hbaa5477d),
	.w5(32'h39b2f667),
	.w6(32'h3a748ec5),
	.w7(32'hb6e33563),
	.w8(32'h3ab085ef),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849de68),
	.w1(32'h3a8c3992),
	.w2(32'h3b171b9a),
	.w3(32'hb9815eb1),
	.w4(32'h39898671),
	.w5(32'h3a9ce048),
	.w6(32'h35b69daa),
	.w7(32'h3b4f8911),
	.w8(32'h38a38a44),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39919e55),
	.w1(32'h3a107ba0),
	.w2(32'h3919293e),
	.w3(32'h3973fa15),
	.w4(32'hbaad9cbd),
	.w5(32'hb68ce581),
	.w6(32'h3aae046b),
	.w7(32'hba9b5610),
	.w8(32'h336b3d7d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40970a),
	.w1(32'hb9c74cc9),
	.w2(32'hb9fecc06),
	.w3(32'hba75a37f),
	.w4(32'hb991af75),
	.w5(32'hba8ca75f),
	.w6(32'hba49767f),
	.w7(32'hb9d64d23),
	.w8(32'hb9aa3b17),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fbb40),
	.w1(32'hba747818),
	.w2(32'hb9344ddb),
	.w3(32'hb9863d7e),
	.w4(32'hba6d8f12),
	.w5(32'hb786a3a0),
	.w6(32'h3a614c27),
	.w7(32'h3a9a6c5b),
	.w8(32'h3b06a267),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967e164),
	.w1(32'hba7006c0),
	.w2(32'hba3d648e),
	.w3(32'h39c8fb50),
	.w4(32'hb965495d),
	.w5(32'h357065da),
	.w6(32'h3a5f6fcb),
	.w7(32'h39bf9023),
	.w8(32'h3a822023),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3622baf0),
	.w1(32'h3545c3b2),
	.w2(32'h3615bba4),
	.w3(32'hb7216944),
	.w4(32'hb640fbe7),
	.w5(32'h37631fd0),
	.w6(32'hb71937c8),
	.w7(32'hb7b4d2df),
	.w8(32'h36c9b0f1),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba48d8b),
	.w1(32'h3749e70f),
	.w2(32'h3b3c532d),
	.w3(32'hbba2d2af),
	.w4(32'hba2bb0ef),
	.w5(32'h3b53135e),
	.w6(32'hbb5d889b),
	.w7(32'h3a21f5ca),
	.w8(32'h3b8d341b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab95dda),
	.w1(32'hb9e37161),
	.w2(32'h39714e4b),
	.w3(32'hbaa6c994),
	.w4(32'hb9f59515),
	.w5(32'hb92e24e2),
	.w6(32'hb9fd04d2),
	.w7(32'h3a643b94),
	.w8(32'h3a2602ce),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb812e4e5),
	.w1(32'hb77d731c),
	.w2(32'h378631b1),
	.w3(32'hb8a19611),
	.w4(32'hb84be9b3),
	.w5(32'h373d4330),
	.w6(32'hb89568b0),
	.w7(32'hb7ac08f7),
	.w8(32'h38044800),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae81487),
	.w1(32'h393a3e7c),
	.w2(32'h3a25283b),
	.w3(32'hbae463b8),
	.w4(32'hb9c04d50),
	.w5(32'h38875cee),
	.w6(32'hbab92660),
	.w7(32'h3a10b88c),
	.w8(32'h3a80bbac),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3876d66c),
	.w1(32'h37cf8445),
	.w2(32'h37e59096),
	.w3(32'h3752ae08),
	.w4(32'hb7c82967),
	.w5(32'hb583d3c4),
	.w6(32'h37c515dd),
	.w7(32'h3733c85b),
	.w8(32'h3810140e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385e174b),
	.w1(32'h3908f0e4),
	.w2(32'h3873dcb4),
	.w3(32'hb8becf0b),
	.w4(32'hb8143fa8),
	.w5(32'h38b9867f),
	.w6(32'hb9886a0b),
	.w7(32'hb5a195dc),
	.w8(32'h390afbbf),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bf4220),
	.w1(32'h370372d9),
	.w2(32'h369d80a7),
	.w3(32'h373ccca5),
	.w4(32'h37bee58a),
	.w5(32'h3772caf8),
	.w6(32'h36e8da42),
	.w7(32'h3779b957),
	.w8(32'h36800ade),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b3c329),
	.w1(32'hb807f690),
	.w2(32'h3759cbc7),
	.w3(32'hb72f697e),
	.w4(32'hb73c9c2d),
	.w5(32'hb762e0e6),
	.w6(32'hb768c092),
	.w7(32'hb74453cc),
	.w8(32'hb7c326e5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d49496),
	.w1(32'hb9a47b56),
	.w2(32'h3a07bc58),
	.w3(32'h3a094640),
	.w4(32'hb9aa49a5),
	.w5(32'h39bd8833),
	.w6(32'h38e81a5c),
	.w7(32'hb9f1f324),
	.w8(32'h3992d61f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39580cad),
	.w1(32'h3a4b46ba),
	.w2(32'h3a23f6b7),
	.w3(32'h380b0608),
	.w4(32'hb91ef7df),
	.w5(32'hbaa1d2f0),
	.w6(32'h3b0af59f),
	.w7(32'h3b4d85d6),
	.w8(32'hb9a61311),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5f1cb),
	.w1(32'hba6e6c4b),
	.w2(32'hba9b6a7d),
	.w3(32'hbaa139e8),
	.w4(32'hba8c784f),
	.w5(32'hbaeb4508),
	.w6(32'hb9d5186d),
	.w7(32'h3a4f3169),
	.w8(32'hb7bd9e17),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac80a06),
	.w1(32'h38d78f77),
	.w2(32'h38ab446c),
	.w3(32'hbaab6e13),
	.w4(32'hba407479),
	.w5(32'hbb0130a6),
	.w6(32'hba280450),
	.w7(32'h3aac3f1f),
	.w8(32'hb9601283),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ba1cc9),
	.w1(32'h38a4a784),
	.w2(32'h38f9dd47),
	.w3(32'h37e7cfea),
	.w4(32'h38eb2472),
	.w5(32'h39135a30),
	.w6(32'hb6211204),
	.w7(32'h3887d9f7),
	.w8(32'h38b42dcc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90bc603),
	.w1(32'h38ae5495),
	.w2(32'h38dd42cc),
	.w3(32'h388d1f51),
	.w4(32'h391a546c),
	.w5(32'h38ba2ffb),
	.w6(32'h38909e8f),
	.w7(32'h392d0c82),
	.w8(32'h397a049e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a24418),
	.w1(32'hb6fc7422),
	.w2(32'hb729b569),
	.w3(32'h368a4325),
	.w4(32'hb782d536),
	.w5(32'hb73b7f44),
	.w6(32'hb68df6a1),
	.w7(32'hb79b279f),
	.w8(32'hb7c65bff),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb48671ea),
	.w1(32'h36abf561),
	.w2(32'hb5d8fe31),
	.w3(32'h34ddec9a),
	.w4(32'h370a692f),
	.w5(32'h37701ecc),
	.w6(32'h367b6bfe),
	.w7(32'h3723ed4c),
	.w8(32'h373afd57),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383a3288),
	.w1(32'h38cb0865),
	.w2(32'hba710657),
	.w3(32'h3a01324e),
	.w4(32'hb984d89e),
	.w5(32'hbaae23a6),
	.w6(32'h3aa02ffe),
	.w7(32'h3ae95122),
	.w8(32'h39226683),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a01de),
	.w1(32'hb8808a5f),
	.w2(32'hb78ed7dc),
	.w3(32'hb886adf6),
	.w4(32'hb8a59650),
	.w5(32'hb8480a19),
	.w6(32'hb87056be),
	.w7(32'hb8919b6f),
	.w8(32'hb81830c1),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38953f46),
	.w1(32'h39ae0d03),
	.w2(32'h3a26fa90),
	.w3(32'h3943ff2c),
	.w4(32'h39ef107d),
	.w5(32'h3a544d14),
	.w6(32'h39388f22),
	.w7(32'h395603d8),
	.w8(32'h3a10c6b4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f28b50),
	.w1(32'hb96a265c),
	.w2(32'h3976244b),
	.w3(32'hb9c4dff5),
	.w4(32'h35fedf7c),
	.w5(32'h38e0106e),
	.w6(32'hb923552e),
	.w7(32'hb99aca1b),
	.w8(32'h3912337d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b1abea),
	.w1(32'h3786088e),
	.w2(32'h3789f40d),
	.w3(32'hb7e10a88),
	.w4(32'h3723704c),
	.w5(32'hb6a6715e),
	.w6(32'hb65cd99a),
	.w7(32'h37c51e67),
	.w8(32'hb70ed5c5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a7047),
	.w1(32'h3906cd16),
	.w2(32'h38cf311d),
	.w3(32'hb9c81165),
	.w4(32'h38875f55),
	.w5(32'h37b51421),
	.w6(32'hb95ab8ee),
	.w7(32'h39d8d80b),
	.w8(32'h39ba2bc1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ef14c6),
	.w1(32'h38915077),
	.w2(32'hb741aa41),
	.w3(32'h391a134b),
	.w4(32'h389740a7),
	.w5(32'hb8942cb2),
	.w6(32'h39c64943),
	.w7(32'h3951f36e),
	.w8(32'hb925e14c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13f3f1),
	.w1(32'h3b3ab50c),
	.w2(32'h3b2715ad),
	.w3(32'hb97a3f0c),
	.w4(32'h39f89674),
	.w5(32'hba737c53),
	.w6(32'h3b228b8e),
	.w7(32'h3b49777f),
	.w8(32'hb9ff54f0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94620b1),
	.w1(32'hb8a31264),
	.w2(32'hb8475d68),
	.w3(32'hb931f687),
	.w4(32'hb7f78cd2),
	.w5(32'hb83ba3f7),
	.w6(32'hb863acf0),
	.w7(32'h382de3e7),
	.w8(32'h35a2d60a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9995cf3),
	.w1(32'hba44b567),
	.w2(32'hb98c1c0a),
	.w3(32'h39a73f41),
	.w4(32'h3a85fcd6),
	.w5(32'h3a92df1c),
	.w6(32'h3b30fcba),
	.w7(32'h3aeb0bfd),
	.w8(32'h3b2ca3f8),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule