module layer_10_featuremap_238(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91941bf),
	.w1(32'hbac5b9ca),
	.w2(32'hbb946b75),
	.w3(32'h3ab18747),
	.w4(32'h398d6ed5),
	.w5(32'h39fcbb5a),
	.w6(32'h3a605576),
	.w7(32'hbb91e9d4),
	.w8(32'h3bb88560),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb784f),
	.w1(32'h3af33834),
	.w2(32'h3a323ecc),
	.w3(32'hbb037553),
	.w4(32'hba2a6f0e),
	.w5(32'hbbb5f210),
	.w6(32'h3bb2283d),
	.w7(32'h3a1c12a9),
	.w8(32'hbb0d41d8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dae86),
	.w1(32'hbb22ccbb),
	.w2(32'h3b494590),
	.w3(32'h398c0c6d),
	.w4(32'hbb177781),
	.w5(32'h3b59fde9),
	.w6(32'hbb02e056),
	.w7(32'h3b062c53),
	.w8(32'h3bf88d35),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1f8ff),
	.w1(32'h3b0e2d06),
	.w2(32'hbacafe13),
	.w3(32'hba965182),
	.w4(32'hba9c5fc8),
	.w5(32'hbbf71920),
	.w6(32'hb9116120),
	.w7(32'hbb3886af),
	.w8(32'h3ab2bfbb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02a3e8),
	.w1(32'h39dbcf5e),
	.w2(32'h3c6ad844),
	.w3(32'hbc0190a3),
	.w4(32'h3c28fcbc),
	.w5(32'h3b96b50d),
	.w6(32'hba5a4fb9),
	.w7(32'h3cd60718),
	.w8(32'h3b7cfb49),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5450de),
	.w1(32'h3a3c773f),
	.w2(32'hbae6dd21),
	.w3(32'h3af470fa),
	.w4(32'hba1b3559),
	.w5(32'hbaf87952),
	.w6(32'h3b0360c7),
	.w7(32'hbb3ef62b),
	.w8(32'hb9caf8cf),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965073b),
	.w1(32'hba36659d),
	.w2(32'hbb1cf516),
	.w3(32'hbb97c550),
	.w4(32'hbb1b97f7),
	.w5(32'hbaf233ce),
	.w6(32'hbb02029c),
	.w7(32'hbb7459f9),
	.w8(32'hbb66ac73),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae52f19),
	.w1(32'hbb426cc7),
	.w2(32'hba1b6cc7),
	.w3(32'h39a9b084),
	.w4(32'h3abac11a),
	.w5(32'h3b45f83e),
	.w6(32'hbab939ff),
	.w7(32'hba9935c9),
	.w8(32'h3b54c20e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e4551),
	.w1(32'h3ae09599),
	.w2(32'h387839fc),
	.w3(32'h3a0d6b49),
	.w4(32'h3a929d4c),
	.w5(32'h3b78d2ef),
	.w6(32'h3b01e1c5),
	.w7(32'hba26550d),
	.w8(32'h3b7f1d04),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12ff0c),
	.w1(32'h3a440a0f),
	.w2(32'hbb17907c),
	.w3(32'hb684da4b),
	.w4(32'hbab951b6),
	.w5(32'h3a40479e),
	.w6(32'hb9d61054),
	.w7(32'hbb7095bc),
	.w8(32'h3b51c822),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b256232),
	.w1(32'hba4e6402),
	.w2(32'hbb0cf9b4),
	.w3(32'h3a213312),
	.w4(32'hbafc05eb),
	.w5(32'h3ae70dfc),
	.w6(32'h3b5fddf0),
	.w7(32'hbb11d5ec),
	.w8(32'h3b296064),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b192bf),
	.w1(32'hbb544374),
	.w2(32'hbae06c5f),
	.w3(32'h3ad0ad3f),
	.w4(32'h39567b0d),
	.w5(32'hbc0905ed),
	.w6(32'h3b109d78),
	.w7(32'hb82ddf95),
	.w8(32'hbb19e876),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cce31),
	.w1(32'h3b3615b4),
	.w2(32'h3c104605),
	.w3(32'h3a2108a2),
	.w4(32'h3bce15d2),
	.w5(32'h39d95760),
	.w6(32'h3b99bcb1),
	.w7(32'h3c1de15f),
	.w8(32'hbba4a902),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8e221),
	.w1(32'h3ba1b6f1),
	.w2(32'h3b2f4a32),
	.w3(32'h3c0b5c9d),
	.w4(32'h3b7bb82f),
	.w5(32'h3a1c59b5),
	.w6(32'h3c3b1fcd),
	.w7(32'h3c601d9b),
	.w8(32'h3b7057ee),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4e24b),
	.w1(32'hbb2d173d),
	.w2(32'hba7b96ba),
	.w3(32'h3aee41f8),
	.w4(32'hbb3a3a79),
	.w5(32'h3a2c90c1),
	.w6(32'h3b87baa0),
	.w7(32'hbba51781),
	.w8(32'h38a7ff67),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f2d964),
	.w1(32'hbb33f78c),
	.w2(32'h3afaaab8),
	.w3(32'hba780af4),
	.w4(32'hba21275b),
	.w5(32'h39f1ef4a),
	.w6(32'h3a66cd8d),
	.w7(32'h3aac88d7),
	.w8(32'h3abb8d65),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d0ff3),
	.w1(32'h3a7e93d7),
	.w2(32'h3b4b542a),
	.w3(32'h3a207d05),
	.w4(32'h3afdf129),
	.w5(32'hbc0e5732),
	.w6(32'h3b56829b),
	.w7(32'h3ab1beb4),
	.w8(32'hbc144bcc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf57752),
	.w1(32'h3b8d3195),
	.w2(32'h3c8c763d),
	.w3(32'hbb4c0965),
	.w4(32'h3c30f30a),
	.w5(32'hbac98690),
	.w6(32'hbb25e702),
	.w7(32'h3c7591e3),
	.w8(32'hbb528d9d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a817895),
	.w1(32'h3bc3a12e),
	.w2(32'h3bd637bf),
	.w3(32'h3a539bab),
	.w4(32'hba3d979b),
	.w5(32'hb9cfd378),
	.w6(32'h3b3eb617),
	.w7(32'h3c2013aa),
	.w8(32'hbb46b7d5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0accd1),
	.w1(32'hbba21b3a),
	.w2(32'hb88493b0),
	.w3(32'h3bdb86e0),
	.w4(32'h3bf32105),
	.w5(32'h3b919b69),
	.w6(32'hbb603bdf),
	.w7(32'h3c274d9f),
	.w8(32'h3b71d5ae),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bcbd1),
	.w1(32'h3b3d8e76),
	.w2(32'h3b23c69e),
	.w3(32'h3b28e98b),
	.w4(32'hba88dc3b),
	.w5(32'h3a127de8),
	.w6(32'h3ad0c30f),
	.w7(32'h3b9e02e6),
	.w8(32'hb8989ab1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3157f8),
	.w1(32'hb9c9822b),
	.w2(32'hbbd3216e),
	.w3(32'hbb27c488),
	.w4(32'hbb42e5b5),
	.w5(32'hbb72d8b3),
	.w6(32'hbbac914b),
	.w7(32'hbbf2ce43),
	.w8(32'hb9db4800),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921da2f),
	.w1(32'h3a47d97a),
	.w2(32'hb916df09),
	.w3(32'h3a861f40),
	.w4(32'h3ab1eea1),
	.w5(32'h398b8322),
	.w6(32'h3bc5c155),
	.w7(32'h3b45589b),
	.w8(32'h398db806),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b325e),
	.w1(32'hbbd8d592),
	.w2(32'h3b869772),
	.w3(32'hbc0f4132),
	.w4(32'hbaec00a5),
	.w5(32'h3ad5f7e6),
	.w6(32'hbc82c85b),
	.w7(32'h3b4637c9),
	.w8(32'hbab866f5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8932b4),
	.w1(32'h3b9e3766),
	.w2(32'h3b8eee77),
	.w3(32'hbae828b9),
	.w4(32'hbb5ddb27),
	.w5(32'hb8e24eb2),
	.w6(32'hbaac1c37),
	.w7(32'h3b399002),
	.w8(32'hb7bae707),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeba660),
	.w1(32'h3a982b5a),
	.w2(32'hba18436c),
	.w3(32'h3b6a3986),
	.w4(32'hbacc672f),
	.w5(32'h3b312eb2),
	.w6(32'h3be21ed2),
	.w7(32'hbb52f8e3),
	.w8(32'hbaa0a001),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f646a9),
	.w1(32'hbb73842c),
	.w2(32'hbb743feb),
	.w3(32'hba9fb335),
	.w4(32'hbb0c29c4),
	.w5(32'h3a90d172),
	.w6(32'h3a09d7d4),
	.w7(32'hbbc0faa3),
	.w8(32'hba3d21ca),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba2b0d),
	.w1(32'h3a9c1634),
	.w2(32'hba3f4ed2),
	.w3(32'hb95ee781),
	.w4(32'h39a56bb2),
	.w5(32'h3b357779),
	.w6(32'hba33bb64),
	.w7(32'hbb27f758),
	.w8(32'hbbce6232),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86da5f),
	.w1(32'hbb9f9b7a),
	.w2(32'hbbfafc7b),
	.w3(32'h3adc40b1),
	.w4(32'hbb9d301f),
	.w5(32'hbb41cf98),
	.w6(32'h39b08fa2),
	.w7(32'h3b318b30),
	.w8(32'hbb715502),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a3f9a),
	.w1(32'hbb7872cd),
	.w2(32'hb84d0096),
	.w3(32'h38a54328),
	.w4(32'hbb100167),
	.w5(32'hbb66c332),
	.w6(32'hbbbc1413),
	.w7(32'h3b9a421b),
	.w8(32'hbb26c9a7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a1999),
	.w1(32'hbbe1229c),
	.w2(32'hbbb74ecd),
	.w3(32'hbbb0f8da),
	.w4(32'h3bc2d63c),
	.w5(32'hbc073344),
	.w6(32'hbbb27801),
	.w7(32'h3b17f236),
	.w8(32'hbb6819d6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd84317),
	.w1(32'hbc0e2bfb),
	.w2(32'h3b2765ba),
	.w3(32'h3a8c70c0),
	.w4(32'hbb044b26),
	.w5(32'hbb391c10),
	.w6(32'h3a9d8b83),
	.w7(32'h37a00573),
	.w8(32'hb73f1464),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba50c38),
	.w1(32'h38ac9cb2),
	.w2(32'h3ba37185),
	.w3(32'hbb284b7e),
	.w4(32'h3c35e7ab),
	.w5(32'hbc2aee99),
	.w6(32'hb9fb37be),
	.w7(32'h3c466e94),
	.w8(32'hbc51009f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cef4d),
	.w1(32'h38a32343),
	.w2(32'h3c8593f5),
	.w3(32'hbc1657df),
	.w4(32'h3c38df41),
	.w5(32'h3ba6fda8),
	.w6(32'hbb45ca41),
	.w7(32'h3c99b19f),
	.w8(32'h3b1e62e7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e3c2d),
	.w1(32'hba6a6dd2),
	.w2(32'h398726f3),
	.w3(32'h3b14e9c7),
	.w4(32'h3b646c53),
	.w5(32'hbbeebc47),
	.w6(32'h3be27096),
	.w7(32'h3b78f1f1),
	.w8(32'hbbc0f30b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ebdb2),
	.w1(32'h3b40a939),
	.w2(32'h3c8c23b4),
	.w3(32'hbaf1267a),
	.w4(32'h3c18384e),
	.w5(32'hba597577),
	.w6(32'hbc00744f),
	.w7(32'h3cb0b935),
	.w8(32'h3ae7e25b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba556d4a),
	.w1(32'h3af20b74),
	.w2(32'hbb9c11c5),
	.w3(32'h383bbb7c),
	.w4(32'h3ab6de2a),
	.w5(32'h3b2793dd),
	.w6(32'h3c44cdf6),
	.w7(32'h3bce321b),
	.w8(32'hbb246c8e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51ae16),
	.w1(32'hbac282ad),
	.w2(32'hbbf28499),
	.w3(32'hbaad0578),
	.w4(32'hbbe77a7e),
	.w5(32'h3a08ace5),
	.w6(32'h3a43d43e),
	.w7(32'hbbf4f697),
	.w8(32'h3a1c1899),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87fc929),
	.w1(32'h3c12f785),
	.w2(32'h3c0edf06),
	.w3(32'hb91fe6ab),
	.w4(32'h3ae88f78),
	.w5(32'h3b9e99e7),
	.w6(32'h3b540dce),
	.w7(32'h3afe29a6),
	.w8(32'h3b866a99),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf720cc),
	.w1(32'hbaf51a45),
	.w2(32'hbc10bee2),
	.w3(32'hb976d5a3),
	.w4(32'hb96f9843),
	.w5(32'hba78ff2f),
	.w6(32'hbb61fe71),
	.w7(32'hbc1a69d5),
	.w8(32'hbb1c8889),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3c191),
	.w1(32'hbac159d5),
	.w2(32'h3b5b0ede),
	.w3(32'h3aa1cc7f),
	.w4(32'h3b3b4724),
	.w5(32'h3a06456c),
	.w6(32'hbaa13796),
	.w7(32'h3c096c31),
	.w8(32'h3a46b4c8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac345db),
	.w1(32'h3ab686aa),
	.w2(32'hbb398b06),
	.w3(32'h3a74c600),
	.w4(32'hbabcb159),
	.w5(32'h3bbed14d),
	.w6(32'h3b8cd43c),
	.w7(32'hbbcee710),
	.w8(32'h3bd33576),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be08797),
	.w1(32'h3aaaabfa),
	.w2(32'hba3af6c3),
	.w3(32'hbaf3411f),
	.w4(32'hbbbf2561),
	.w5(32'h3b7b0acb),
	.w6(32'h3b8ec7f5),
	.w7(32'hbbbd4fda),
	.w8(32'h3beac4ce),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8deaa6),
	.w1(32'h3b31ddf9),
	.w2(32'hba4df5e9),
	.w3(32'hbac05484),
	.w4(32'hbbaf8237),
	.w5(32'hbb6b0e79),
	.w6(32'h3c4bcef0),
	.w7(32'h3bec48aa),
	.w8(32'h3ba750fb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65d627),
	.w1(32'h3aa4b810),
	.w2(32'hbc190c20),
	.w3(32'hbb9323b5),
	.w4(32'hbb74007c),
	.w5(32'h3a40e059),
	.w6(32'hbb4d402a),
	.w7(32'hbbf076c9),
	.w8(32'hb7b00576),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c3a8b),
	.w1(32'hbaf7bca9),
	.w2(32'hbacdb3eb),
	.w3(32'h3a088d3e),
	.w4(32'h39fc9c2d),
	.w5(32'h38d7c008),
	.w6(32'h3ba6063c),
	.w7(32'hbb65ddf2),
	.w8(32'h3b42cd20),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cfbd9),
	.w1(32'h3a3cecb6),
	.w2(32'hbb0f74d3),
	.w3(32'h38aa3fa3),
	.w4(32'hbab449fd),
	.w5(32'hba6cdb15),
	.w6(32'h3b7b6161),
	.w7(32'hbb566620),
	.w8(32'hba8579d0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f35f2),
	.w1(32'hbb958378),
	.w2(32'hbc23c930),
	.w3(32'hbba6f036),
	.w4(32'hbc24f1c3),
	.w5(32'hbbfbd218),
	.w6(32'hbb9364e0),
	.w7(32'hbc5fefc6),
	.w8(32'hbb9f4075),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc94ae5),
	.w1(32'hbaf82023),
	.w2(32'hbb1871af),
	.w3(32'hbb877bb8),
	.w4(32'hbbc6e2cb),
	.w5(32'h3a596e05),
	.w6(32'h3988229b),
	.w7(32'hbbc4b917),
	.w8(32'h39bd813a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ca197),
	.w1(32'hba344018),
	.w2(32'hbb6ec65a),
	.w3(32'hba80db08),
	.w4(32'hbad86978),
	.w5(32'hbb33eea7),
	.w6(32'hbb70f9a1),
	.w7(32'hbbcf14b2),
	.w8(32'hbbb21e52),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05eba6),
	.w1(32'hbbcec3a0),
	.w2(32'h3bf11987),
	.w3(32'hbaeafb53),
	.w4(32'h3c50d102),
	.w5(32'h3a94d3a2),
	.w6(32'hbcb1acef),
	.w7(32'h3c7693e2),
	.w8(32'hbb7115d0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93734d),
	.w1(32'hbb193a2c),
	.w2(32'h3a7e363f),
	.w3(32'h3a703d60),
	.w4(32'h3beecdfd),
	.w5(32'hbb4a097a),
	.w6(32'hbac7028b),
	.w7(32'h3b6834b6),
	.w8(32'hbaa6fc46),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b581f7a),
	.w1(32'h3b086abc),
	.w2(32'hbaab9483),
	.w3(32'hbb4be521),
	.w4(32'h3b1a722b),
	.w5(32'hbb2596aa),
	.w6(32'hbb699a61),
	.w7(32'h3bf92d88),
	.w8(32'hbb6ee0ee),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860b47),
	.w1(32'hba698398),
	.w2(32'hbb440f5e),
	.w3(32'h3b211410),
	.w4(32'h371ef421),
	.w5(32'hbb84bd9a),
	.w6(32'hb83a0266),
	.w7(32'h3b5d2c6d),
	.w8(32'hbb4cbe40),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8929a2),
	.w1(32'hbb9a6da8),
	.w2(32'h3b16ec1c),
	.w3(32'h3b9e603c),
	.w4(32'h3c445b06),
	.w5(32'hb993d4fe),
	.w6(32'hbba902b9),
	.w7(32'h3c3f1b79),
	.w8(32'hbb48bfdd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca9cb1),
	.w1(32'hbb9a4a10),
	.w2(32'hba8373bb),
	.w3(32'hbbc74158),
	.w4(32'h3a506f7b),
	.w5(32'hb906ce90),
	.w6(32'hbb85660e),
	.w7(32'h3c059369),
	.w8(32'hbb112a51),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61dab2),
	.w1(32'hbabd32ed),
	.w2(32'hba47cbe6),
	.w3(32'hba556a4b),
	.w4(32'hba1c65d2),
	.w5(32'h3aaa39dd),
	.w6(32'hbb53b938),
	.w7(32'h3ad8f5bb),
	.w8(32'hbaf3fa62),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a4e83),
	.w1(32'hbb984495),
	.w2(32'hbc3abdf8),
	.w3(32'h3b8e6a27),
	.w4(32'hbbccfe3b),
	.w5(32'hbb0fbfd3),
	.w6(32'h3b6cccb4),
	.w7(32'hb9c921c0),
	.w8(32'hbac36b05),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de1d91),
	.w1(32'hba52a9dc),
	.w2(32'hbb0a0aaa),
	.w3(32'hbb1eaeeb),
	.w4(32'hbacad1f1),
	.w5(32'h3b27077e),
	.w6(32'hbb233ecb),
	.w7(32'hbbb1e6b9),
	.w8(32'hbb2c1e43),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa7a6b),
	.w1(32'h3b02d2de),
	.w2(32'hbc24ff1a),
	.w3(32'h3a544478),
	.w4(32'hbb02597b),
	.w5(32'hb785d99d),
	.w6(32'h3be9c2a8),
	.w7(32'hbc27e3be),
	.w8(32'h3b3337d2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb050ccb),
	.w1(32'h3b8bf7a2),
	.w2(32'h3b16f1c7),
	.w3(32'h398a6320),
	.w4(32'h3a9eefb0),
	.w5(32'hb99f2f72),
	.w6(32'h3b85447a),
	.w7(32'h39a88424),
	.w8(32'h3b8a3057),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17a0a7),
	.w1(32'h3b5a23e2),
	.w2(32'h3ba2bfa3),
	.w3(32'hbae4e3c8),
	.w4(32'hb80f571e),
	.w5(32'h3bb97d11),
	.w6(32'h3b92efc7),
	.w7(32'hbac35eed),
	.w8(32'h3bcfd161),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10f6f5),
	.w1(32'h3ae3e2bd),
	.w2(32'h3b1b15b0),
	.w3(32'h39d5626d),
	.w4(32'h3b9a2cdf),
	.w5(32'hbb149119),
	.w6(32'h3c06ac9c),
	.w7(32'h3bf7d7e1),
	.w8(32'hbba9bef6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc76d0),
	.w1(32'hbb30ff5c),
	.w2(32'h3b3251c7),
	.w3(32'h398b1a6f),
	.w4(32'h3b82f29f),
	.w5(32'h3b7eb0b5),
	.w6(32'hb8bc3d26),
	.w7(32'h3c1afca7),
	.w8(32'hba22803e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3d119),
	.w1(32'hbbec0c90),
	.w2(32'hbb5a3681),
	.w3(32'h3b8c64e7),
	.w4(32'hbb192466),
	.w5(32'hbb0686f9),
	.w6(32'hbaecb34a),
	.w7(32'h3b5f2cd2),
	.w8(32'hbb1f8f4b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa35a9),
	.w1(32'hbbe48a5e),
	.w2(32'hba8ee864),
	.w3(32'h3b1459e6),
	.w4(32'h3bf1f781),
	.w5(32'h3af40233),
	.w6(32'hbaac7301),
	.w7(32'h3bc79457),
	.w8(32'h3a1c53af),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0f147),
	.w1(32'hba91aa01),
	.w2(32'h39aec922),
	.w3(32'h3ba78117),
	.w4(32'hbb06ab2f),
	.w5(32'h3c142d47),
	.w6(32'h3bd6387e),
	.w7(32'hbb0387c4),
	.w8(32'h3c2b0545),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2eb598),
	.w1(32'hbb9e5d03),
	.w2(32'hbc1903d4),
	.w3(32'hbaa98820),
	.w4(32'hbc5bfe40),
	.w5(32'hbb934cdf),
	.w6(32'h3bce112b),
	.w7(32'hbc4afd1a),
	.w8(32'hbb648b7a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaf0a1),
	.w1(32'hbbc9fa4b),
	.w2(32'h3be90713),
	.w3(32'hb9942f86),
	.w4(32'h3bcd24e9),
	.w5(32'h3b974e3c),
	.w6(32'hbc63fe37),
	.w7(32'h3c747b69),
	.w8(32'h3a20f0fb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1647e4),
	.w1(32'hbab30f4a),
	.w2(32'h3bc8f229),
	.w3(32'hb90b9b01),
	.w4(32'h3ab7e213),
	.w5(32'h3b5e79cf),
	.w6(32'h3b71751d),
	.w7(32'h3acbbf8e),
	.w8(32'h3bff79b6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf102),
	.w1(32'h3a7c0384),
	.w2(32'hbb8a901d),
	.w3(32'h3b0f8049),
	.w4(32'hbbbf6362),
	.w5(32'h3b91aad9),
	.w6(32'h3c106dae),
	.w7(32'hbba6a761),
	.w8(32'h3b7c5fd0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb35bb3),
	.w1(32'hba344e73),
	.w2(32'hbb2f0479),
	.w3(32'h3be76a15),
	.w4(32'hbacd73ac),
	.w5(32'hb981e1c6),
	.w6(32'h3b5b7ac6),
	.w7(32'h3a7cfa2d),
	.w8(32'hbb0fb260),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8579c),
	.w1(32'h3b415447),
	.w2(32'h3b18e85e),
	.w3(32'hb93ff7c8),
	.w4(32'hba8da7e9),
	.w5(32'hbb2fe5e3),
	.w6(32'hbb005d91),
	.w7(32'hbb16ac6f),
	.w8(32'hba0431e3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e9d28),
	.w1(32'hbb9af55e),
	.w2(32'h39c99dc3),
	.w3(32'hbbcb62ef),
	.w4(32'h3ae18339),
	.w5(32'h3b0cf79f),
	.w6(32'h3aabd8f8),
	.w7(32'h3b2118c2),
	.w8(32'h3b371d5f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b519910),
	.w1(32'hb990142b),
	.w2(32'hbb72490b),
	.w3(32'h3b9aa53c),
	.w4(32'hbb472cb2),
	.w5(32'hbc08d532),
	.w6(32'h3c1da6c3),
	.w7(32'hbb8c13d1),
	.w8(32'hbbdb930c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf99a8a),
	.w1(32'h3b71d9ba),
	.w2(32'h3c53774c),
	.w3(32'h3abf0f08),
	.w4(32'h3c235e7e),
	.w5(32'h3ab5313a),
	.w6(32'h3b74657a),
	.w7(32'h3c83d5fb),
	.w8(32'h3ac397e2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaad7bc),
	.w1(32'hbb858060),
	.w2(32'hbacebb8e),
	.w3(32'hb9ea3745),
	.w4(32'hb9203952),
	.w5(32'hbb97bc11),
	.w6(32'hba1f5f8a),
	.w7(32'h38496d92),
	.w8(32'hbbc11095),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba562528),
	.w1(32'hba2ac047),
	.w2(32'h3c258c57),
	.w3(32'hbb8aaaf7),
	.w4(32'h3c487542),
	.w5(32'h38e2220e),
	.w6(32'hbbfc8e23),
	.w7(32'h3c89a152),
	.w8(32'h3ac3ba60),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d2c6),
	.w1(32'hbb89a6d6),
	.w2(32'hbbd5781c),
	.w3(32'hb88dede8),
	.w4(32'hb94ef2d0),
	.w5(32'h3bb23836),
	.w6(32'hbaeee869),
	.w7(32'hbbbc3704),
	.w8(32'h3bac0fd0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cc8fe),
	.w1(32'h3b281937),
	.w2(32'h3b84deb0),
	.w3(32'h3b35e359),
	.w4(32'hb83ce278),
	.w5(32'h39050b3e),
	.w6(32'h3be28d28),
	.w7(32'h3a1aff76),
	.w8(32'h3ac2c2dc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56c310),
	.w1(32'hbba05c2a),
	.w2(32'hbc739f62),
	.w3(32'h3976420a),
	.w4(32'hbc18b1ec),
	.w5(32'hbc1b17be),
	.w6(32'hbb334cf2),
	.w7(32'hbc4dd929),
	.w8(32'hbbee84e8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecc2ff),
	.w1(32'h3b1c2aaa),
	.w2(32'h3c283046),
	.w3(32'hbaf8deb7),
	.w4(32'h3b3ad8d8),
	.w5(32'hbb62ee6a),
	.w6(32'h3a8718ea),
	.w7(32'h3c341d40),
	.w8(32'hbaf4ac35),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05c270),
	.w1(32'hbb32f38d),
	.w2(32'hbafe28a2),
	.w3(32'hbb5a9fbd),
	.w4(32'hbbad8d0b),
	.w5(32'h3c3892d1),
	.w6(32'hbba44220),
	.w7(32'h3b9f6224),
	.w8(32'h3c59a99e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f8362),
	.w1(32'hbb69a67f),
	.w2(32'hbba0ba37),
	.w3(32'h3b3aec3b),
	.w4(32'hbc1e0bbc),
	.w5(32'hbb63bb9c),
	.w6(32'h3b7fac22),
	.w7(32'hbb3147d9),
	.w8(32'h3b51a464),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b525cc3),
	.w1(32'hba89f17b),
	.w2(32'h39985fcf),
	.w3(32'hbb25be85),
	.w4(32'hbb3bf07a),
	.w5(32'hbba72ee5),
	.w6(32'h3b0daba3),
	.w7(32'h3adcd6ae),
	.w8(32'hba0fa670),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb841e97),
	.w1(32'h3a5fc2f3),
	.w2(32'h3baee54f),
	.w3(32'h3ac8bf36),
	.w4(32'hbb2bc567),
	.w5(32'hb9df6f4a),
	.w6(32'h3ba467ee),
	.w7(32'h3ab2dc64),
	.w8(32'hba0b3a0e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a687ffd),
	.w1(32'hba441b8c),
	.w2(32'h3b04c098),
	.w3(32'h3ac5b71d),
	.w4(32'h3b12d50c),
	.w5(32'h3b6e6c73),
	.w6(32'h3b314b5c),
	.w7(32'h3b4c9d0f),
	.w8(32'h3b8d0755),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ba84c),
	.w1(32'hbb8e7f12),
	.w2(32'hbb9a6eb9),
	.w3(32'h3b81bd88),
	.w4(32'h3bc9481f),
	.w5(32'h398ac020),
	.w6(32'h3a83f623),
	.w7(32'h3b9e2f78),
	.w8(32'h38ea4aee),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ff3ce),
	.w1(32'h3a9619ea),
	.w2(32'h3b3f2ab1),
	.w3(32'hbb18ed44),
	.w4(32'h3a827a5b),
	.w5(32'hbb1ca31e),
	.w6(32'hb8e70079),
	.w7(32'hbb07a3f7),
	.w8(32'hbb1c7536),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4701a5),
	.w1(32'hbbfcf7cb),
	.w2(32'h3c0580e3),
	.w3(32'hbb9ba5a7),
	.w4(32'h39f356a0),
	.w5(32'h3a8a8f35),
	.w6(32'hbc2a255d),
	.w7(32'h3beb2d63),
	.w8(32'h3bc341b1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6ab61),
	.w1(32'hbb421105),
	.w2(32'h3aeb1ce6),
	.w3(32'hbbb249e4),
	.w4(32'hba28a8ba),
	.w5(32'hbb91750d),
	.w6(32'hbb330cc1),
	.w7(32'hbadbf691),
	.w8(32'hbbf04551),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f1a8b),
	.w1(32'hbbdadec3),
	.w2(32'h3b9047f0),
	.w3(32'hbbdaa8b2),
	.w4(32'hbb9612ef),
	.w5(32'hbc0a9b55),
	.w6(32'hbc5388a6),
	.w7(32'h3c049f35),
	.w8(32'hbb30899d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98afe97),
	.w1(32'hbb8c2d81),
	.w2(32'h3c3c5992),
	.w3(32'hbc10a2b8),
	.w4(32'h3c223890),
	.w5(32'h3a1f0261),
	.w6(32'hbbf6d229),
	.w7(32'h3c4d42c7),
	.w8(32'hbb628518),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a57f1),
	.w1(32'hbbb4139d),
	.w2(32'hbc3c78a9),
	.w3(32'h3aca7f47),
	.w4(32'hbc1648a6),
	.w5(32'h3b4f88b2),
	.w6(32'hb953a771),
	.w7(32'hbbe92b6d),
	.w8(32'h3b08301e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab4c68),
	.w1(32'hbacf69b0),
	.w2(32'hbb66083b),
	.w3(32'h3a703d83),
	.w4(32'hbbada2ef),
	.w5(32'h3b9d70aa),
	.w6(32'hbb194e96),
	.w7(32'hbbb3b083),
	.w8(32'h39d72b3b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb050d1f),
	.w1(32'hbbba0126),
	.w2(32'hbbc8ecb4),
	.w3(32'h3b1f1d45),
	.w4(32'hbc0d2591),
	.w5(32'h3b4bcf30),
	.w6(32'h3b5da5ee),
	.w7(32'hbbefa63d),
	.w8(32'h3bb6b28a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7253),
	.w1(32'hbacdf6c0),
	.w2(32'hbc05e897),
	.w3(32'hbabd0bd6),
	.w4(32'h3b0b7d3b),
	.w5(32'hbbc86acf),
	.w6(32'hbad59f2d),
	.w7(32'hbbc6be21),
	.w8(32'hbc146619),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f13f3),
	.w1(32'hbc2c5eee),
	.w2(32'h3b161917),
	.w3(32'hbc31cb48),
	.w4(32'h3bb9fd30),
	.w5(32'hbaacb236),
	.w6(32'hbc8b9b7b),
	.w7(32'h3c11c2cc),
	.w8(32'hba988079),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacae45d),
	.w1(32'hbb01eebb),
	.w2(32'hbab35b8b),
	.w3(32'hbacb68f4),
	.w4(32'hbac06ec4),
	.w5(32'hb9c39257),
	.w6(32'hbad37868),
	.w7(32'hba94488e),
	.w8(32'hbac56b2b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93377ed),
	.w1(32'hb9c2e562),
	.w2(32'h3a96b4d4),
	.w3(32'hbad4e44a),
	.w4(32'h38a857a6),
	.w5(32'hba6a977e),
	.w6(32'hbb033625),
	.w7(32'h383effa2),
	.w8(32'hb892092d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa03429),
	.w1(32'h3a515c7a),
	.w2(32'h3b5d8478),
	.w3(32'h3a1ae59a),
	.w4(32'h3b7454f9),
	.w5(32'hbb04a42a),
	.w6(32'h3aa31bff),
	.w7(32'h3b5a5184),
	.w8(32'hbadec8e1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1afd66),
	.w1(32'hba9d4db0),
	.w2(32'hba6498f6),
	.w3(32'hbb1107e1),
	.w4(32'hbb07719f),
	.w5(32'hbac0cb0a),
	.w6(32'hba75828b),
	.w7(32'hba759fb3),
	.w8(32'hbab05089),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab38b16),
	.w1(32'hb9fe2c2e),
	.w2(32'h3a7a9fb8),
	.w3(32'hbad7f582),
	.w4(32'hb9f1e125),
	.w5(32'hba83be9c),
	.w6(32'hba99b98a),
	.w7(32'h3a3618ed),
	.w8(32'hba49dba3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c28e5),
	.w1(32'hba5bdac7),
	.w2(32'h39c6f2e6),
	.w3(32'hb9e20e5b),
	.w4(32'hba0da273),
	.w5(32'hbb21576a),
	.w6(32'hbad7f80b),
	.w7(32'h38f16d7d),
	.w8(32'hbb2a22aa),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98e9ee),
	.w1(32'hbae252c3),
	.w2(32'hba9c7093),
	.w3(32'hbb0f7994),
	.w4(32'hbafb98d9),
	.w5(32'hba2d9d03),
	.w6(32'hbb81a0c5),
	.w7(32'hbb307274),
	.w8(32'hb9c5d688),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a855bf3),
	.w1(32'h3a899ac9),
	.w2(32'h3a00e8af),
	.w3(32'h39b49564),
	.w4(32'h39a4aee6),
	.w5(32'h3a191fe1),
	.w6(32'hb89e4dfa),
	.w7(32'h39b7f178),
	.w8(32'h3846bd1f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c907cb),
	.w1(32'hb9b23e7b),
	.w2(32'h39dc38d1),
	.w3(32'hb919cc4a),
	.w4(32'hba665f01),
	.w5(32'h3aab1362),
	.w6(32'hba8cbdcc),
	.w7(32'hba9e1996),
	.w8(32'h3a2f0d99),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba156df3),
	.w1(32'h3adb26f0),
	.w2(32'h3a5f070a),
	.w3(32'h3b289826),
	.w4(32'h3afd39c9),
	.w5(32'hbaa5efd9),
	.w6(32'h3b489b5b),
	.w7(32'h3b267aed),
	.w8(32'hb959dd31),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab56799),
	.w1(32'hbaac645b),
	.w2(32'hba8c5f60),
	.w3(32'hbaa588f0),
	.w4(32'hba854a66),
	.w5(32'hb9eb63fe),
	.w6(32'hba4c08d8),
	.w7(32'hba095002),
	.w8(32'hb917fac5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdf196),
	.w1(32'h3a5ef52f),
	.w2(32'h3b0b1339),
	.w3(32'h3a39e4a8),
	.w4(32'h3b24a995),
	.w5(32'h3af04fdc),
	.w6(32'h3b289094),
	.w7(32'h3b807095),
	.w8(32'h3ab0cf14),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8aad9e),
	.w1(32'h392dfe97),
	.w2(32'h3a9efac3),
	.w3(32'h3a357347),
	.w4(32'h3a6e5fa5),
	.w5(32'hbab58191),
	.w6(32'h3a456f3f),
	.w7(32'h3ad49b57),
	.w8(32'hbb2cce18),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248e18),
	.w1(32'hb994b726),
	.w2(32'h39cbe63f),
	.w3(32'hba3be6ff),
	.w4(32'hba177dc1),
	.w5(32'h3b0308ca),
	.w6(32'hba95647e),
	.w7(32'h38f94143),
	.w8(32'h3b023f22),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeff14d),
	.w1(32'h3a848d7d),
	.w2(32'h3a694e80),
	.w3(32'h3a717c44),
	.w4(32'h3aba31b8),
	.w5(32'hba92fec7),
	.w6(32'h3a67a510),
	.w7(32'h3a3db876),
	.w8(32'hba4372e1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99af4ea),
	.w1(32'hb9d506dd),
	.w2(32'h395ec910),
	.w3(32'hba27dc53),
	.w4(32'hba5e4987),
	.w5(32'hb8d7285b),
	.w6(32'hba7a3bda),
	.w7(32'hba631c05),
	.w8(32'hbb2bd83a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb523b2c),
	.w1(32'hbb2219a0),
	.w2(32'hbb527a76),
	.w3(32'hbad9aa86),
	.w4(32'hbb0e3389),
	.w5(32'hba80b8a4),
	.w6(32'h3a05b74f),
	.w7(32'hbb20d86c),
	.w8(32'hbb204115),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fd565),
	.w1(32'hbab900f6),
	.w2(32'hb961d0eb),
	.w3(32'hba2ed583),
	.w4(32'hba90e829),
	.w5(32'h3a14d448),
	.w6(32'hbb12a369),
	.w7(32'hba0c2d68),
	.w8(32'h3a879d57),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a890e),
	.w1(32'h3abe3311),
	.w2(32'h3abd8008),
	.w3(32'h3a4b1521),
	.w4(32'h3a17702b),
	.w5(32'hbb5f919f),
	.w6(32'h3a761d32),
	.w7(32'h3a364e38),
	.w8(32'hbb30e352),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78fd61),
	.w1(32'hba1e21f9),
	.w2(32'hba905c8c),
	.w3(32'hbb28f348),
	.w4(32'hbb2a1ad2),
	.w5(32'hba4ed3d2),
	.w6(32'hbb5500af),
	.w7(32'hbab8a0fd),
	.w8(32'hba26fac8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385548bd),
	.w1(32'hba16f98f),
	.w2(32'h3b22e6e6),
	.w3(32'hbadd39d8),
	.w4(32'h3aa53b8e),
	.w5(32'hbb5ea8dc),
	.w6(32'hbabaf84b),
	.w7(32'h3aaf572c),
	.w8(32'hbb2af1c6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8df2c4),
	.w1(32'hbb93a781),
	.w2(32'hbb1ea792),
	.w3(32'hbb895fba),
	.w4(32'hbb81a743),
	.w5(32'hba5048a8),
	.w6(32'hbb8919d4),
	.w7(32'hbb59328d),
	.w8(32'hba8f24e6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf99f6d),
	.w1(32'hba528076),
	.w2(32'hb9097eb5),
	.w3(32'h385c727d),
	.w4(32'hb81fbb66),
	.w5(32'h38026abb),
	.w6(32'hbac863e4),
	.w7(32'hb98a9e63),
	.w8(32'h383b50d6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c4c32),
	.w1(32'hba948cca),
	.w2(32'hba1c7215),
	.w3(32'hba3ae17d),
	.w4(32'h3a6439c8),
	.w5(32'hba090066),
	.w6(32'hba9c2ea5),
	.w7(32'h3a5cb5aa),
	.w8(32'hb9ebebb1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a6539),
	.w1(32'hba423347),
	.w2(32'hb9fd0ae8),
	.w3(32'hb988a7b2),
	.w4(32'hbb314887),
	.w5(32'hba24408c),
	.w6(32'hba24a1e2),
	.w7(32'hba974ead),
	.w8(32'h3809e138),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f27d00),
	.w1(32'hba8a3510),
	.w2(32'hba8283cc),
	.w3(32'hbaca568c),
	.w4(32'h385b9577),
	.w5(32'hb9bb7ba2),
	.w6(32'hba736d51),
	.w7(32'hba802485),
	.w8(32'h3a3fdde6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa76ede),
	.w1(32'h3a0447e1),
	.w2(32'h3aa63894),
	.w3(32'hba8f2fa1),
	.w4(32'hbb13f2a9),
	.w5(32'hbaeb27d5),
	.w6(32'h3a29688f),
	.w7(32'hb96157ed),
	.w8(32'hb92a0e77),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f783a),
	.w1(32'h391298f3),
	.w2(32'h38e1080e),
	.w3(32'hba11e857),
	.w4(32'hb972475f),
	.w5(32'hba5b7cc7),
	.w6(32'h3a53d738),
	.w7(32'h3a0df615),
	.w8(32'hba1e8848),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0195a),
	.w1(32'hbaa1d894),
	.w2(32'hb9efa4aa),
	.w3(32'h397bef31),
	.w4(32'h39e9c590),
	.w5(32'h39491c92),
	.w6(32'h39de93c0),
	.w7(32'h39f9874a),
	.w8(32'hb8f31a62),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab70557),
	.w1(32'hb9f49919),
	.w2(32'hb9bc74a7),
	.w3(32'hba5bdf7a),
	.w4(32'hba4885bf),
	.w5(32'h3b114ba2),
	.w6(32'hb91aca21),
	.w7(32'h3878bc0f),
	.w8(32'h3adb0a70),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987e37f),
	.w1(32'h3b4cfa76),
	.w2(32'h3b861820),
	.w3(32'h3b8fb407),
	.w4(32'h3bb85fbd),
	.w5(32'hb906f636),
	.w6(32'h3ba2f0a6),
	.w7(32'h3bd1dd3a),
	.w8(32'hbaa64dd5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11284a),
	.w1(32'hbad86c3b),
	.w2(32'hba2463b6),
	.w3(32'hba89aa8e),
	.w4(32'hbae3df38),
	.w5(32'hb99e99e2),
	.w6(32'hba8c7b15),
	.w7(32'hbae53793),
	.w8(32'hb94a8392),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba968886),
	.w1(32'hba7431d6),
	.w2(32'h3afbd092),
	.w3(32'hb9055e76),
	.w4(32'h3920bf22),
	.w5(32'hbac5027c),
	.w6(32'hbacefe71),
	.w7(32'h3a28bc65),
	.w8(32'hbaddf20f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2a36b),
	.w1(32'hbb06fb98),
	.w2(32'hbaf33756),
	.w3(32'hbad90275),
	.w4(32'hbb108d4c),
	.w5(32'hba8e60fb),
	.w6(32'hbaa424df),
	.w7(32'hbb21edb8),
	.w8(32'hbaeaee83),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba513a42),
	.w1(32'hbb209e8a),
	.w2(32'hbac43d14),
	.w3(32'hbab5d3a3),
	.w4(32'h39c6ddca),
	.w5(32'hbb146315),
	.w6(32'hbb34fcd0),
	.w7(32'hbaaacdad),
	.w8(32'hbabe84c7),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb286359),
	.w1(32'hba875a68),
	.w2(32'hba3f7f38),
	.w3(32'hba75b72b),
	.w4(32'hba6eee6e),
	.w5(32'hba4f51d3),
	.w6(32'h3a40d6b3),
	.w7(32'h39793423),
	.w8(32'hba470a38),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ea8f6),
	.w1(32'h3981ec95),
	.w2(32'h3a4ae72c),
	.w3(32'hb7b0e02a),
	.w4(32'h39f4d998),
	.w5(32'hba7bbba7),
	.w6(32'h3a08fac4),
	.w7(32'h383ebb37),
	.w8(32'hbadf59b2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae78eed),
	.w1(32'hba65dcee),
	.w2(32'hbb18a987),
	.w3(32'hb977e302),
	.w4(32'hb8cde565),
	.w5(32'h3a75ace7),
	.w6(32'h39a900b2),
	.w7(32'hba61e74e),
	.w8(32'h3a98a1c5),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a124063),
	.w1(32'h3aca4674),
	.w2(32'h3aa78722),
	.w3(32'h3aa10f86),
	.w4(32'h3a99f884),
	.w5(32'hbb0a8705),
	.w6(32'h3ae75cee),
	.w7(32'h3ab98820),
	.w8(32'hbabf640a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25e291),
	.w1(32'hba464e18),
	.w2(32'hb9f186a6),
	.w3(32'hba3ed02e),
	.w4(32'hba2670cb),
	.w5(32'hbb30238c),
	.w6(32'h3a2a9d30),
	.w7(32'h39c8a262),
	.w8(32'hbae6e951),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1da08d),
	.w1(32'hba9a2228),
	.w2(32'hba446faf),
	.w3(32'hbaf22144),
	.w4(32'hba9c47d0),
	.w5(32'h3ac24bab),
	.w6(32'hb861c652),
	.w7(32'hb9cfce8b),
	.w8(32'h39bf6821),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392dea8a),
	.w1(32'hbab9524b),
	.w2(32'hbaa95c03),
	.w3(32'h3a0a8cce),
	.w4(32'hba124a50),
	.w5(32'hba8549f0),
	.w6(32'hb9eb9203),
	.w7(32'hba8ab8d4),
	.w8(32'hbafb0b59),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a4ea8),
	.w1(32'hba861b19),
	.w2(32'hba08b81e),
	.w3(32'hb9fe7408),
	.w4(32'hb995d734),
	.w5(32'h3a00dd10),
	.w6(32'hbaf3e7df),
	.w7(32'hba89d608),
	.w8(32'h393cb436),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eb809),
	.w1(32'hb7e87d57),
	.w2(32'h3a4eb169),
	.w3(32'hbaa5b1e3),
	.w4(32'hba95c359),
	.w5(32'h3a502b97),
	.w6(32'hb9cf3ecd),
	.w7(32'hb78fca6c),
	.w8(32'h39ed6df7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914a446),
	.w1(32'hb93cf1db),
	.w2(32'h38bf68a3),
	.w3(32'h39dbe02d),
	.w4(32'hb982dcf6),
	.w5(32'h381243bd),
	.w6(32'h39ec4f2d),
	.w7(32'hb8e60565),
	.w8(32'h37c4fff6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fcbd0),
	.w1(32'hb9c1b858),
	.w2(32'hb9787650),
	.w3(32'h39d463e1),
	.w4(32'h39c3ce22),
	.w5(32'h3a3bb179),
	.w6(32'h38814f7a),
	.w7(32'h3a8d15a8),
	.w8(32'h390bd8ec),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f7a06),
	.w1(32'h39f05911),
	.w2(32'h3887d890),
	.w3(32'h3b01ba67),
	.w4(32'h3a1cbbb0),
	.w5(32'hba5e51e2),
	.w6(32'h3b1a7a0c),
	.w7(32'h3a1156a7),
	.w8(32'hba1ac3ed),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9baadf3),
	.w1(32'hb92f59ae),
	.w2(32'h389614a2),
	.w3(32'hba43abc2),
	.w4(32'hb8f70020),
	.w5(32'hb93e9b99),
	.w6(32'hba1b177f),
	.w7(32'hb993497e),
	.w8(32'h3aa9071f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafc5bd),
	.w1(32'h3a9f0eb6),
	.w2(32'h3ad3693a),
	.w3(32'hb875ae5f),
	.w4(32'h3a99d17a),
	.w5(32'hbb0d411c),
	.w6(32'h3ab253ac),
	.w7(32'h3b143229),
	.w8(32'hba84d1f8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7251cc),
	.w1(32'hba521521),
	.w2(32'hbaa974a9),
	.w3(32'hba5aa9a5),
	.w4(32'h39dae53f),
	.w5(32'hb84414bd),
	.w6(32'hb83cf4c0),
	.w7(32'hba22a485),
	.w8(32'h3a81d218),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdf03d),
	.w1(32'h3a7bc9dd),
	.w2(32'h3a9e3a52),
	.w3(32'h3a1aa2b7),
	.w4(32'h3adbef3b),
	.w5(32'h3a8f8d7e),
	.w6(32'h3a30688f),
	.w7(32'h3b44b3fc),
	.w8(32'h3ae57d40),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab17317),
	.w1(32'h3b03b7b0),
	.w2(32'h3b00639c),
	.w3(32'h3aa78554),
	.w4(32'h3aa0a6fb),
	.w5(32'hbac6ff06),
	.w6(32'h3b0485ca),
	.w7(32'h3aac2240),
	.w8(32'hba96c7da),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf68ebf),
	.w1(32'hbb124500),
	.w2(32'hba5a7de4),
	.w3(32'hbb32467a),
	.w4(32'hbae96980),
	.w5(32'hb9c0dc67),
	.w6(32'hbb086ffc),
	.w7(32'hba8a4ebb),
	.w8(32'hba7d693e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae47bf),
	.w1(32'hba420fd8),
	.w2(32'hbb1036d0),
	.w3(32'h3a49487d),
	.w4(32'hbb1b7d4f),
	.w5(32'hbac5202a),
	.w6(32'h3a5460b9),
	.w7(32'hbae75bbb),
	.w8(32'hbadb6734),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7f24),
	.w1(32'hbab65f0f),
	.w2(32'hba0b8b55),
	.w3(32'hba801adb),
	.w4(32'hbab61c60),
	.w5(32'h3a995c5e),
	.w6(32'hbaa0ff0f),
	.w7(32'hbac7d6ed),
	.w8(32'h3aa11225),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0aa430),
	.w1(32'h3b4baf6d),
	.w2(32'h3b1b29d3),
	.w3(32'h3b66b095),
	.w4(32'h3b951bca),
	.w5(32'h39836226),
	.w6(32'h3b7f9280),
	.w7(32'h3b8a0c4a),
	.w8(32'h3a229430),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391788a6),
	.w1(32'h3ac0d506),
	.w2(32'h3aff73de),
	.w3(32'h3a9ef343),
	.w4(32'h3ae50e28),
	.w5(32'h3a3c2b8c),
	.w6(32'h3ab675e7),
	.w7(32'h3ae58562),
	.w8(32'h3a6e663a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944929a),
	.w1(32'h3abe6b1e),
	.w2(32'h3b1a89db),
	.w3(32'h3aafe10e),
	.w4(32'h3b37b8fd),
	.w5(32'hbb06f38e),
	.w6(32'h3b0720c6),
	.w7(32'h3b6e6d95),
	.w8(32'hba7eda94),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85bafb2),
	.w1(32'hba57b238),
	.w2(32'hbabef424),
	.w3(32'hbb36d0c0),
	.w4(32'hbb3b6bc5),
	.w5(32'hbac597fb),
	.w6(32'hbac88e25),
	.w7(32'hbb080421),
	.w8(32'hba1587e5),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba7492),
	.w1(32'hb9b2a458),
	.w2(32'hb88f4114),
	.w3(32'hba63cfc5),
	.w4(32'h39a9bb8b),
	.w5(32'hb93ab9bd),
	.w6(32'hba18f194),
	.w7(32'h38f02324),
	.w8(32'h3850b072),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c00ba),
	.w1(32'h39dc7bbb),
	.w2(32'hba86b861),
	.w3(32'hbb1a9e53),
	.w4(32'h39c87aed),
	.w5(32'h3a4bd05c),
	.w6(32'hb9d7ecea),
	.w7(32'hb86e3719),
	.w8(32'hba66c8cb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77923a),
	.w1(32'hbadd092d),
	.w2(32'hb74b9a56),
	.w3(32'h3b1566a2),
	.w4(32'h3a1d9ca3),
	.w5(32'hb95720f4),
	.w6(32'h38a0d155),
	.w7(32'hb983d7bc),
	.w8(32'h3990a2a5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa21d2c),
	.w1(32'h3af41f82),
	.w2(32'h3b0c9ba2),
	.w3(32'h39b352e8),
	.w4(32'h3b58dc9f),
	.w5(32'hba5cacd7),
	.w6(32'h3a447890),
	.w7(32'h3b805798),
	.w8(32'hba807f84),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f538a),
	.w1(32'hb97c378d),
	.w2(32'h399ccb02),
	.w3(32'hba489f6c),
	.w4(32'hba73b7d5),
	.w5(32'hba272bf2),
	.w6(32'hba350fd3),
	.w7(32'hba3a8355),
	.w8(32'hb950fe3b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984256a),
	.w1(32'hba0e02df),
	.w2(32'hb9b29c9c),
	.w3(32'hba2556e7),
	.w4(32'h39367cf4),
	.w5(32'hba917d1d),
	.w6(32'h399b8170),
	.w7(32'hba80b069),
	.w8(32'hbaa23c3b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e1a67),
	.w1(32'hbaba73a1),
	.w2(32'hba4461ec),
	.w3(32'hbb024882),
	.w4(32'hba9b5558),
	.w5(32'hbad2dc79),
	.w6(32'hbb05338f),
	.w7(32'hba4a5e56),
	.w8(32'h3a02efd0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6125c),
	.w1(32'h3aea6d18),
	.w2(32'h3987ca2d),
	.w3(32'hb9fc06b3),
	.w4(32'h39d0b598),
	.w5(32'hbb0afc6f),
	.w6(32'hb935e01b),
	.w7(32'hba857c47),
	.w8(32'hba5ae9c5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe73d0),
	.w1(32'h3a0480b4),
	.w2(32'h3a7c69f9),
	.w3(32'h36ed54e9),
	.w4(32'h392fa876),
	.w5(32'hba22cf06),
	.w6(32'h3a6e5a81),
	.w7(32'h3b0154d2),
	.w8(32'hba3595d5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaada301),
	.w1(32'hbb0664c9),
	.w2(32'hbad04938),
	.w3(32'hbac9e4a6),
	.w4(32'hbad06533),
	.w5(32'hba59d64f),
	.w6(32'hba110dc8),
	.w7(32'hbb221fb1),
	.w8(32'hb9f09f1b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bc21b4),
	.w1(32'h39e39e5a),
	.w2(32'h3ab7c35d),
	.w3(32'h3a874df9),
	.w4(32'h3aea711a),
	.w5(32'hb8dbb553),
	.w6(32'h39cc8917),
	.w7(32'h3a5d3448),
	.w8(32'hba52f4b0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb23ce),
	.w1(32'hbac7a1cf),
	.w2(32'hba8ad82d),
	.w3(32'hbb2150b9),
	.w4(32'hbae09b9f),
	.w5(32'h3a3cd40d),
	.w6(32'hbb098e68),
	.w7(32'hba9d0b71),
	.w8(32'h3a990993),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc0468),
	.w1(32'h3b216789),
	.w2(32'h3b108cd4),
	.w3(32'h3b3b74f6),
	.w4(32'h3b70a14a),
	.w5(32'hbb42d7a4),
	.w6(32'h3b58391f),
	.w7(32'h3b51c525),
	.w8(32'hbae07933),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9a97f),
	.w1(32'hbab69188),
	.w2(32'hbaea9346),
	.w3(32'hbb4c6504),
	.w4(32'hbb305372),
	.w5(32'hbb830b49),
	.w6(32'hbafbe90c),
	.w7(32'hba8fddd6),
	.w8(32'hbbba02dc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb697cb9),
	.w1(32'hbb8ebcd6),
	.w2(32'hbaf95b38),
	.w3(32'hbbc222dd),
	.w4(32'hbb57c738),
	.w5(32'hba2952ac),
	.w6(32'hbb9127c4),
	.w7(32'hbb0d07c9),
	.w8(32'hb93bdd34),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820d91),
	.w1(32'h3a2d3eeb),
	.w2(32'h3abf1da5),
	.w3(32'hba236ae3),
	.w4(32'h3aa6e55a),
	.w5(32'h3b13f46b),
	.w6(32'hb9faf87c),
	.w7(32'h3a3ea2b7),
	.w8(32'h3b297bd8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15726c),
	.w1(32'h3ab7a604),
	.w2(32'h3b063795),
	.w3(32'h3afd930d),
	.w4(32'h3b15849b),
	.w5(32'h39ffcc80),
	.w6(32'h3b1c3fdd),
	.w7(32'h3b603a25),
	.w8(32'h379d90b6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff5155),
	.w1(32'h38b5c5e3),
	.w2(32'h3ad437ee),
	.w3(32'h3a300f5d),
	.w4(32'hba15f650),
	.w5(32'h3b6df7d9),
	.w6(32'h39a3049e),
	.w7(32'h3a65283e),
	.w8(32'h3b69a5a8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3483c4),
	.w1(32'h3b44b749),
	.w2(32'h3b0debc4),
	.w3(32'h3b590c35),
	.w4(32'h3b09b3fc),
	.w5(32'hba16a096),
	.w6(32'h3b69f36a),
	.w7(32'h3affe176),
	.w8(32'hb9c9f048),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e0f315),
	.w1(32'hb97974d6),
	.w2(32'hba63959a),
	.w3(32'hb998c8a5),
	.w4(32'h38e677db),
	.w5(32'h3b1ede0f),
	.w6(32'hb99ac958),
	.w7(32'hb9ccfa7f),
	.w8(32'h3b55cea0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c84e4),
	.w1(32'h3b53cec8),
	.w2(32'h3b5f3b2b),
	.w3(32'h3b3d5e58),
	.w4(32'h3b5a529a),
	.w5(32'h398fa74d),
	.w6(32'h3b5f3963),
	.w7(32'h3b24d882),
	.w8(32'hbac205a5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaece49a),
	.w1(32'h38a32aca),
	.w2(32'hba237e44),
	.w3(32'h3aa4a134),
	.w4(32'hba0d10de),
	.w5(32'hbab3e88a),
	.w6(32'h39fcd119),
	.w7(32'h39761159),
	.w8(32'hbb10818d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70f995),
	.w1(32'hb9f358b0),
	.w2(32'hbab0b96e),
	.w3(32'hbae00819),
	.w4(32'hba9563bb),
	.w5(32'h398a416a),
	.w6(32'hb9a5ecdf),
	.w7(32'hba345eb8),
	.w8(32'hb7a92c60),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba891891),
	.w1(32'hba92c40c),
	.w2(32'hbab55e97),
	.w3(32'hb9a2aefe),
	.w4(32'hb9e2edd7),
	.w5(32'hb70aa1f4),
	.w6(32'hb996f2e6),
	.w7(32'hba89e460),
	.w8(32'h39260aed),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af32f9),
	.w1(32'hba480a0c),
	.w2(32'hba05985a),
	.w3(32'hb8dd3698),
	.w4(32'h3a924c5f),
	.w5(32'hbb08cdb8),
	.w6(32'hbafe651d),
	.w7(32'hb95817c6),
	.w8(32'hbae72a90),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba606adf),
	.w1(32'hbab5880c),
	.w2(32'hbb25555f),
	.w3(32'hba737d86),
	.w4(32'hba1d3972),
	.w5(32'hbaf9930e),
	.w6(32'hba8d00b7),
	.w7(32'hbafbf205),
	.w8(32'hbaa421e8),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba571760),
	.w1(32'hbadef608),
	.w2(32'hbb0f8d20),
	.w3(32'hbae2dc6a),
	.w4(32'hbb2843d0),
	.w5(32'h39e20cb3),
	.w6(32'hb9f04941),
	.w7(32'hbafd5c26),
	.w8(32'h3a060840),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab854f3),
	.w1(32'hb909bf7c),
	.w2(32'hb9bec196),
	.w3(32'hba3aa4c4),
	.w4(32'hba41293a),
	.w5(32'h3930c320),
	.w6(32'hb9ebbd95),
	.w7(32'h367cdc6a),
	.w8(32'hb8e6c64b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac448c),
	.w1(32'hb9b565c1),
	.w2(32'hb76fffee),
	.w3(32'hba2c8a39),
	.w4(32'h3a638a4d),
	.w5(32'h3b0083ca),
	.w6(32'hba5b5c15),
	.w7(32'h3a0ef83a),
	.w8(32'h3b1d83dc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace40c5),
	.w1(32'h3b51cb27),
	.w2(32'h3b53e007),
	.w3(32'h3b3d40a4),
	.w4(32'h3b6d76a0),
	.w5(32'h3a1a2b72),
	.w6(32'h3b4d6aab),
	.w7(32'h3b2dc60b),
	.w8(32'h3af9d6ee),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21ce04),
	.w1(32'h3a88e8ee),
	.w2(32'h3aa2ebad),
	.w3(32'h39b8bfc4),
	.w4(32'h39c6ef12),
	.w5(32'h39ded9d8),
	.w6(32'h399107ba),
	.w7(32'h3a86a323),
	.w8(32'h37f3f7eb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972e588),
	.w1(32'hbaaabf25),
	.w2(32'h37645c6e),
	.w3(32'hb9945b79),
	.w4(32'h3a75fc72),
	.w5(32'h3a1ee057),
	.w6(32'hb9c29921),
	.w7(32'h3847df4c),
	.w8(32'h39432d1a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdfbba),
	.w1(32'hba597fd2),
	.w2(32'hbad23b07),
	.w3(32'h3aa4b4b9),
	.w4(32'h3ad2f674),
	.w5(32'hb9e0dea5),
	.w6(32'h3aa29ee2),
	.w7(32'h39aafd05),
	.w8(32'hb9cd4a71),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7bf5f),
	.w1(32'hbabd0dbb),
	.w2(32'hba209ee0),
	.w3(32'hb9963f65),
	.w4(32'h3a91fcfd),
	.w5(32'hba888be5),
	.w6(32'hba1e4092),
	.w7(32'hb9c1658a),
	.w8(32'hba4fe3fc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81616a),
	.w1(32'hba9c74c1),
	.w2(32'hba086cc0),
	.w3(32'hbadd41f1),
	.w4(32'hba86d5ca),
	.w5(32'hbb38d0a9),
	.w6(32'hba2bb9a5),
	.w7(32'hba0fe08d),
	.w8(32'hbae609d7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f9d68),
	.w1(32'hba191723),
	.w2(32'hba17b141),
	.w3(32'hba97e1ab),
	.w4(32'hb9e4dd3e),
	.w5(32'hbae6c43f),
	.w6(32'hba264a7f),
	.w7(32'hba6a10c8),
	.w8(32'hbb0181d9),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabefb83),
	.w1(32'hbb35d6af),
	.w2(32'hbb3cd66c),
	.w3(32'hba878f78),
	.w4(32'hb8b3fecf),
	.w5(32'h3a1a4a7c),
	.w6(32'hbb0663ad),
	.w7(32'hbb13e0f7),
	.w8(32'h3a08b55d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fceec),
	.w1(32'hba880cdb),
	.w2(32'hba1ef0a3),
	.w3(32'h398b40a1),
	.w4(32'h3ae832f6),
	.w5(32'hbab4fa0e),
	.w6(32'h3a1bc37b),
	.w7(32'h3a79e880),
	.w8(32'hba51a291),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf6886),
	.w1(32'hba5e2dc8),
	.w2(32'hbade0c3d),
	.w3(32'hbad79a32),
	.w4(32'hbb2eb2ec),
	.w5(32'hbaace45c),
	.w6(32'hba85b2a0),
	.w7(32'hbaf25381),
	.w8(32'hbae50de1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb089eef),
	.w1(32'h3a287ca4),
	.w2(32'hbae296d9),
	.w3(32'h36c79add),
	.w4(32'hbab3e785),
	.w5(32'hba53bc1f),
	.w6(32'h3995863b),
	.w7(32'hba70dd24),
	.w8(32'hbab668bc),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9495e73),
	.w1(32'hba3b55ea),
	.w2(32'hba311a1d),
	.w3(32'hbb0f57a4),
	.w4(32'hbaf69ae3),
	.w5(32'hbaecda33),
	.w6(32'hbac6ed9f),
	.w7(32'hba5e972c),
	.w8(32'hba960a6d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1ed21),
	.w1(32'hba6a7797),
	.w2(32'hba6cbdec),
	.w3(32'hbaa52caa),
	.w4(32'hba83f6ba),
	.w5(32'h3a4750e5),
	.w6(32'hba6de8e7),
	.w7(32'hba9728fe),
	.w8(32'hba48dcda),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a34402),
	.w1(32'h37f45a22),
	.w2(32'h3acf8d08),
	.w3(32'h3b12e68e),
	.w4(32'h3af1a996),
	.w5(32'h3a8b27f8),
	.w6(32'h3b0b6f9c),
	.w7(32'h3b4ed850),
	.w8(32'h37d5e40c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba536a97),
	.w1(32'hb99055e3),
	.w2(32'hbac198ba),
	.w3(32'h3a75a9be),
	.w4(32'h39cd111e),
	.w5(32'hbb1c6f91),
	.w6(32'h3984abc5),
	.w7(32'hbab0ebbf),
	.w8(32'hbac4717c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd412b),
	.w1(32'hb9f937ec),
	.w2(32'h378c1eda),
	.w3(32'hbab8c325),
	.w4(32'hba5d6940),
	.w5(32'h3aabe028),
	.w6(32'hbaddda6b),
	.w7(32'hb9db490c),
	.w8(32'h3b1fe9d5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94c263),
	.w1(32'hb8028bcf),
	.w2(32'h39cc783a),
	.w3(32'h3a29e703),
	.w4(32'h3a469b3e),
	.w5(32'hbb13eab0),
	.w6(32'h3a9685de),
	.w7(32'h3abd7f2b),
	.w8(32'hbae18b47),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5aca7),
	.w1(32'hba395d85),
	.w2(32'hba7a7e45),
	.w3(32'hbb01669e),
	.w4(32'hbb0934b6),
	.w5(32'hbaba34a5),
	.w6(32'hbad279ba),
	.w7(32'hbac62e49),
	.w8(32'hbaf2410f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1200a9),
	.w1(32'hbb1417b8),
	.w2(32'hb9ff3ef9),
	.w3(32'hbafd59a1),
	.w4(32'hba0a4137),
	.w5(32'hb9d751f1),
	.w6(32'hbb1396c6),
	.w7(32'hba69be24),
	.w8(32'hbaf5564e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ace0fc),
	.w1(32'h382ff8e6),
	.w2(32'hb8ce9905),
	.w3(32'hbaa55103),
	.w4(32'hba5a8c56),
	.w5(32'h3a54efad),
	.w6(32'hba87606d),
	.w7(32'hb982980b),
	.w8(32'hb9274589),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b9f58),
	.w1(32'hba9e954d),
	.w2(32'h389d8333),
	.w3(32'h38b6ced9),
	.w4(32'h39bb3f47),
	.w5(32'h3a34b892),
	.w6(32'hba8becc4),
	.w7(32'h3a4da69b),
	.w8(32'h39b0db8f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387df72b),
	.w1(32'hba6461f2),
	.w2(32'hba997043),
	.w3(32'h39c3d73b),
	.w4(32'h3a574ad6),
	.w5(32'h3a876186),
	.w6(32'h3a6fc69e),
	.w7(32'h3a0a07d4),
	.w8(32'h381b9563),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2029a6),
	.w1(32'h395437d8),
	.w2(32'h39ff1ad0),
	.w3(32'h3aba7761),
	.w4(32'hb9ce3c9e),
	.w5(32'hb9bb0a9d),
	.w6(32'h37982e7a),
	.w7(32'h39e72a17),
	.w8(32'h3a8c2627),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c9b3d),
	.w1(32'h39f68499),
	.w2(32'h39a3ea18),
	.w3(32'hb9601563),
	.w4(32'h399d629f),
	.w5(32'hba208e8a),
	.w6(32'h3a30a2f2),
	.w7(32'h3a4fe7d0),
	.w8(32'hba2e2c7a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba648797),
	.w1(32'hb9d621e5),
	.w2(32'h3a1afc46),
	.w3(32'hb9845285),
	.w4(32'hba782297),
	.w5(32'hba581b80),
	.w6(32'hb9f29264),
	.w7(32'h39d751ef),
	.w8(32'h3a445e30),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc5830),
	.w1(32'hb9042f91),
	.w2(32'hba7013cd),
	.w3(32'h3906f8e5),
	.w4(32'hbac64f74),
	.w5(32'hba933394),
	.w6(32'h3a94030a),
	.w7(32'hb91a8f8b),
	.w8(32'hb9beb6d4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ccb14),
	.w1(32'hba888387),
	.w2(32'h395bd68d),
	.w3(32'hbaabb3e2),
	.w4(32'hbab5733f),
	.w5(32'h39a6ad1a),
	.w6(32'hbab99de4),
	.w7(32'hb9dbad9a),
	.w8(32'h39cf2852),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85e673),
	.w1(32'hbaa64c84),
	.w2(32'hb9e213be),
	.w3(32'h3a1d480b),
	.w4(32'h3acb031c),
	.w5(32'h3aa650c9),
	.w6(32'h39af6f85),
	.w7(32'h3b11e682),
	.w8(32'h3ad878c0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bf6af),
	.w1(32'h3ac6da2d),
	.w2(32'h3b2c234a),
	.w3(32'h3b28ca50),
	.w4(32'h3b4a0b76),
	.w5(32'hba8338d8),
	.w6(32'h3a65a004),
	.w7(32'h3acafa4d),
	.w8(32'hb9c71f9c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8367d),
	.w1(32'hba5a9908),
	.w2(32'hba51df79),
	.w3(32'hb99f18c4),
	.w4(32'h3a517efe),
	.w5(32'hb8bb63dd),
	.w6(32'hb9880704),
	.w7(32'hb8cd1206),
	.w8(32'hb9c6bd42),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32158a),
	.w1(32'hb9553629),
	.w2(32'hb9803639),
	.w3(32'h39fe8db8),
	.w4(32'h39364c5d),
	.w5(32'hbadc7864),
	.w6(32'h3a242d37),
	.w7(32'hb8780a5d),
	.w8(32'hba8930eb),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15d4b8),
	.w1(32'h39b07ca1),
	.w2(32'hb9cca127),
	.w3(32'hba76c848),
	.w4(32'h3a32c1b7),
	.w5(32'h39bae6f6),
	.w6(32'h3a594980),
	.w7(32'h3a97383a),
	.w8(32'hba84e783),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1f1ba),
	.w1(32'hbaa6bc92),
	.w2(32'hba8de7ae),
	.w3(32'h3a78385a),
	.w4(32'hba893428),
	.w5(32'hbad17a5e),
	.w6(32'hb98ea01c),
	.w7(32'hba7ba56a),
	.w8(32'hbae2b8d7),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae87124),
	.w1(32'h39b70ade),
	.w2(32'h3b0c150f),
	.w3(32'hba4b1c40),
	.w4(32'h3b0980f2),
	.w5(32'hbaea74ba),
	.w6(32'h3a3759c4),
	.w7(32'h3b21d18c),
	.w8(32'hbb6f39d6),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5049d7),
	.w1(32'hbad9124c),
	.w2(32'h3ab41566),
	.w3(32'hbb088aac),
	.w4(32'hba05a216),
	.w5(32'hba90abd9),
	.w6(32'hba582d3f),
	.w7(32'hbab756e8),
	.w8(32'hba32bc59),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f0632),
	.w1(32'h39fda3ce),
	.w2(32'h3b8d289b),
	.w3(32'hba902188),
	.w4(32'h3b01b4b9),
	.w5(32'hb9575b7c),
	.w6(32'hb9c2eed6),
	.w7(32'h3b3f13eb),
	.w8(32'hba09243a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba054600),
	.w1(32'h3b1f8b1b),
	.w2(32'h3b47480e),
	.w3(32'h3b0443f3),
	.w4(32'h3b835a2f),
	.w5(32'hbb1d0b24),
	.w6(32'h3b2c9f72),
	.w7(32'h3ba54679),
	.w8(32'hbac33edf),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9b451),
	.w1(32'hbaa4a655),
	.w2(32'h39ff2704),
	.w3(32'h378b69fa),
	.w4(32'hb9d21351),
	.w5(32'hba227bf3),
	.w6(32'h3aebee00),
	.w7(32'h3a94b277),
	.w8(32'hbab51cc6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb115c67),
	.w1(32'hbb48108d),
	.w2(32'hbac683ba),
	.w3(32'hbaa4bf2c),
	.w4(32'hbafc1c41),
	.w5(32'h39903ae2),
	.w6(32'hbb35ea67),
	.w7(32'hbab44b6e),
	.w8(32'hbadfe124),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb003d58),
	.w1(32'h3994f050),
	.w2(32'h392016bd),
	.w3(32'h39c9359a),
	.w4(32'h3a9474b7),
	.w5(32'hbc3ebb5a),
	.w6(32'h3a058178),
	.w7(32'h3ac9bc7d),
	.w8(32'hbc077d5f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1b810),
	.w1(32'h3b280050),
	.w2(32'h3c2d3a4e),
	.w3(32'hbc2bc48d),
	.w4(32'h3af9857a),
	.w5(32'hbbd84b4f),
	.w6(32'hbc4e2a29),
	.w7(32'h3c406025),
	.w8(32'hbba483a0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc322f),
	.w1(32'hb931051c),
	.w2(32'hbbd02f8c),
	.w3(32'hb9cb2cd6),
	.w4(32'hbb3fa85b),
	.w5(32'hbb86240d),
	.w6(32'h3a2864c4),
	.w7(32'hbbe03d23),
	.w8(32'hbc29fc6d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e0151),
	.w1(32'h3c0a8b7a),
	.w2(32'h3c121839),
	.w3(32'hbc54fe95),
	.w4(32'hbb80565c),
	.w5(32'hba1debe8),
	.w6(32'hbb0c8855),
	.w7(32'h3c5acc3c),
	.w8(32'hbb0217b3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc064a2b),
	.w1(32'hbbc3e693),
	.w2(32'hbb3c80d0),
	.w3(32'h3b157e56),
	.w4(32'h3b56152a),
	.w5(32'hbbc1c6ce),
	.w6(32'hbb675f8d),
	.w7(32'h3a24a811),
	.w8(32'hbbc389b8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64214b),
	.w1(32'hbbf5779d),
	.w2(32'hbb8a58c5),
	.w3(32'hbb6fb258),
	.w4(32'hbb7e6216),
	.w5(32'hbd16fc46),
	.w6(32'h3c24152c),
	.w7(32'hbb9364af),
	.w8(32'hbd3e0cbb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcd723),
	.w1(32'h3d1ed771),
	.w2(32'h3d31d109),
	.w3(32'hbd2c53b0),
	.w4(32'h3be8292a),
	.w5(32'h3aadf5ba),
	.w6(32'hbbf3551a),
	.w7(32'h3d62b2a4),
	.w8(32'h3c9837af),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d7913),
	.w1(32'h3adc7409),
	.w2(32'hbc01742a),
	.w3(32'hbbb4bd0a),
	.w4(32'h3c1c17fc),
	.w5(32'h3b2385fb),
	.w6(32'h3bc692c5),
	.w7(32'h3c217436),
	.w8(32'h3b8608ef),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd17eec),
	.w1(32'hbbaa6161),
	.w2(32'hba46dc6c),
	.w3(32'hba6855f7),
	.w4(32'hbbeb7713),
	.w5(32'h3bf48971),
	.w6(32'hbb0b63d5),
	.w7(32'hbbd1ddc8),
	.w8(32'h3b646bcc),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe097db),
	.w1(32'hbc2479ee),
	.w2(32'h3c387972),
	.w3(32'h3c133fb8),
	.w4(32'hbad23847),
	.w5(32'hbb5fa861),
	.w6(32'hbb238233),
	.w7(32'hb8f875f3),
	.w8(32'hbbb6e8f5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0328e5),
	.w1(32'hbb151182),
	.w2(32'h3bb165a3),
	.w3(32'h3b45d392),
	.w4(32'hba32a6da),
	.w5(32'hb836f29d),
	.w6(32'hbb67df21),
	.w7(32'h3b2ea0a0),
	.w8(32'hbba627bd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acebdc8),
	.w1(32'h3bd1a547),
	.w2(32'h3caa1625),
	.w3(32'hbbfbc0a2),
	.w4(32'h3bd520a7),
	.w5(32'hbc1105c4),
	.w6(32'hbc3edcdb),
	.w7(32'h3c723dbe),
	.w8(32'hbbac6042),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e99f8),
	.w1(32'hbc130c50),
	.w2(32'hbc0c34a6),
	.w3(32'hbb9ac1b6),
	.w4(32'hbbbf4602),
	.w5(32'hbbbe7f9c),
	.w6(32'hbbd1219a),
	.w7(32'hbba9843d),
	.w8(32'h3c0bd6c6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5c8a8),
	.w1(32'hbbf25941),
	.w2(32'hbb805a0e),
	.w3(32'h3bdfc962),
	.w4(32'h3b9e376c),
	.w5(32'hbacfcd61),
	.w6(32'hbb317cec),
	.w7(32'hb95f8483),
	.w8(32'hbb807c38),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b821fab),
	.w1(32'h3ac08700),
	.w2(32'hbbf26357),
	.w3(32'hb9bc051b),
	.w4(32'hbb679ee5),
	.w5(32'h3c9401ca),
	.w6(32'h3cb186d7),
	.w7(32'hbb0062a2),
	.w8(32'h3ca628e3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0d4dc),
	.w1(32'hbccb4b51),
	.w2(32'hbca4f76d),
	.w3(32'h3bc69fdc),
	.w4(32'hbc2528c4),
	.w5(32'hbb1ea4d6),
	.w6(32'hbc495c3b),
	.w7(32'hbcb95a9a),
	.w8(32'hba8d9d34),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01575b),
	.w1(32'hbba84a4c),
	.w2(32'hbbf9b479),
	.w3(32'hb9ce8bff),
	.w4(32'hbaf789ff),
	.w5(32'hbb56d796),
	.w6(32'h3bf6faef),
	.w7(32'hbb8946b3),
	.w8(32'h3b54660c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66aaa0),
	.w1(32'h3b1a3f49),
	.w2(32'hbb016eda),
	.w3(32'hbc45f73a),
	.w4(32'hb8fc2d97),
	.w5(32'h3ada6396),
	.w6(32'hbb8f076c),
	.w7(32'h3c8a54eb),
	.w8(32'hbb87dd19),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34e0b7),
	.w1(32'hb9bdd0b1),
	.w2(32'hbc06dfd5),
	.w3(32'hbb8748e0),
	.w4(32'hbb701fd2),
	.w5(32'hbb8ee609),
	.w6(32'h3c81d8d3),
	.w7(32'h3b417993),
	.w8(32'hb95c9a22),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8288da),
	.w1(32'h3b1e7d6c),
	.w2(32'hbbdc762d),
	.w3(32'hbb2cbe30),
	.w4(32'hb9bed932),
	.w5(32'h3b1a61bc),
	.w6(32'h3b61abcc),
	.w7(32'hbb5c5713),
	.w8(32'hb9c9833e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd59143),
	.w1(32'hb9e60bf8),
	.w2(32'h3af097a3),
	.w3(32'hbb34ec45),
	.w4(32'hba7870ff),
	.w5(32'hbc9c0a0d),
	.w6(32'hbc7fe20c),
	.w7(32'h3b4def1a),
	.w8(32'hbc606f1f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce0dca),
	.w1(32'hb69bce3e),
	.w2(32'h3ad56fbe),
	.w3(32'hbc3bef31),
	.w4(32'hbbd3ffe0),
	.w5(32'hbcc1031c),
	.w6(32'hbbe68628),
	.w7(32'h3b314b45),
	.w8(32'hbd104e3e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb557daf),
	.w1(32'h3ceab6e5),
	.w2(32'h3ce2f830),
	.w3(32'hbcaaa7d3),
	.w4(32'h3bbf8be0),
	.w5(32'h3c03a65f),
	.w6(32'hbc5855f3),
	.w7(32'h3cec3d18),
	.w8(32'hbbf3380b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab45f9a),
	.w1(32'h3be5c6bb),
	.w2(32'hbb592c23),
	.w3(32'h3874a7bd),
	.w4(32'hba57b89a),
	.w5(32'hbb545e0e),
	.w6(32'h3c696e36),
	.w7(32'h3b04c86c),
	.w8(32'h3c07557e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84c482),
	.w1(32'hbc049d68),
	.w2(32'hbaa949f7),
	.w3(32'h3bc43f33),
	.w4(32'h3b40181a),
	.w5(32'h3bfbfe0a),
	.w6(32'h3beabda1),
	.w7(32'h3b94710e),
	.w8(32'h3bd5d87e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828b8c),
	.w1(32'hbb63834f),
	.w2(32'h3a20d2e8),
	.w3(32'h3c5d2767),
	.w4(32'hbb956b62),
	.w5(32'h3bd0449e),
	.w6(32'hbc385317),
	.w7(32'hbc94e2c0),
	.w8(32'h3c56e90e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad79e8e),
	.w1(32'hbc3b0725),
	.w2(32'hbc02b517),
	.w3(32'h3ba08de0),
	.w4(32'h3b0fad8e),
	.w5(32'h3c089603),
	.w6(32'hbba25e6f),
	.w7(32'hbb1cb94d),
	.w8(32'h3c5541c0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b867250),
	.w1(32'hbba14ba4),
	.w2(32'hbae216bd),
	.w3(32'h3bf5315f),
	.w4(32'hbbe88729),
	.w5(32'hbb75d2cc),
	.w6(32'h3baa8f5d),
	.w7(32'hbc2bfa8e),
	.w8(32'hbbf346ca),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab27e07),
	.w1(32'hbc17c684),
	.w2(32'hbc479d6d),
	.w3(32'hbbc260a7),
	.w4(32'h3a72e9af),
	.w5(32'hb8cd7b1c),
	.w6(32'hbbd13f16),
	.w7(32'h3ad27c74),
	.w8(32'h3b4f3096),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c8d91),
	.w1(32'hbb4bee91),
	.w2(32'h3b3c4005),
	.w3(32'h3b78eb26),
	.w4(32'h3b52d520),
	.w5(32'h3b8d01b1),
	.w6(32'h3b510c7c),
	.w7(32'h3be3ad72),
	.w8(32'h39bacee4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb97d),
	.w1(32'hbb8c63b6),
	.w2(32'h37ab86d0),
	.w3(32'hbc2a287f),
	.w4(32'hbaac2750),
	.w5(32'h3ad94eaa),
	.w6(32'hb9b7d1e5),
	.w7(32'h3b9cb289),
	.w8(32'hba7a4f6e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule