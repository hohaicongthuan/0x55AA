module layer_10_featuremap_437(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf1a43),
	.w1(32'h3ab8dfd0),
	.w2(32'h3b5d6d6d),
	.w3(32'h3992b96c),
	.w4(32'h3a3d38b2),
	.w5(32'hbb2e195f),
	.w6(32'hbbb917c4),
	.w7(32'hbae5b917),
	.w8(32'hbbb375b3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd7f28),
	.w1(32'h3b621b2b),
	.w2(32'h3b10ee97),
	.w3(32'hba59c235),
	.w4(32'hbab8f2b1),
	.w5(32'hbbb82fc8),
	.w6(32'hbbc1761d),
	.w7(32'h39c36574),
	.w8(32'hbb8149d6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c5179),
	.w1(32'h3bcd7023),
	.w2(32'h3b4d8539),
	.w3(32'h3b35e8e1),
	.w4(32'h3c292ae4),
	.w5(32'hbb9678b0),
	.w6(32'h3b84c0c3),
	.w7(32'hb9f51250),
	.w8(32'hbbd23643),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc10083),
	.w1(32'h3b9756a1),
	.w2(32'h3b74cfdd),
	.w3(32'h3a03f4da),
	.w4(32'hbacd2f6d),
	.w5(32'h3c781aba),
	.w6(32'hb9ef5d4b),
	.w7(32'h3b31a966),
	.w8(32'h3b245bf4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27aa36),
	.w1(32'h3ab8d846),
	.w2(32'hbb5e2a41),
	.w3(32'hbb65173b),
	.w4(32'hba3396c6),
	.w5(32'h3ac5b901),
	.w6(32'hbb4f3c04),
	.w7(32'hbb27d794),
	.w8(32'hba865d8a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2d11f),
	.w1(32'hbbcef2c6),
	.w2(32'h3b51a75f),
	.w3(32'h3ba0c0f5),
	.w4(32'h3c50cfe3),
	.w5(32'h3bc95996),
	.w6(32'h3b254878),
	.w7(32'hba36cc0f),
	.w8(32'hbb79e33f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20725c),
	.w1(32'h3bc2fabe),
	.w2(32'h3b98abdc),
	.w3(32'h3c321dc9),
	.w4(32'hbbbb01a0),
	.w5(32'h3a7bf771),
	.w6(32'h3c2efa27),
	.w7(32'hbb6c97c7),
	.w8(32'hba69a497),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb795a7),
	.w1(32'hbaa3cd65),
	.w2(32'hba945c5b),
	.w3(32'hbb792020),
	.w4(32'h3a8e7305),
	.w5(32'hbbacbb5a),
	.w6(32'hbb19c76f),
	.w7(32'hbb0d33be),
	.w8(32'h3bbc25ba),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3d99d),
	.w1(32'h3b2e018a),
	.w2(32'h3acb9bc1),
	.w3(32'h3ab14115),
	.w4(32'h3a7fd8a1),
	.w5(32'h395b8cb2),
	.w6(32'h3c0964bb),
	.w7(32'hbb91d606),
	.w8(32'hbb3e4db2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e92da),
	.w1(32'hbbdba99e),
	.w2(32'hba1195ae),
	.w3(32'hbb7509d7),
	.w4(32'h391ae55f),
	.w5(32'h3bbdca9d),
	.w6(32'hbbb4b89e),
	.w7(32'hbba2bd6d),
	.w8(32'hbbba773a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab26612),
	.w1(32'hbb819750),
	.w2(32'h39bcc3f5),
	.w3(32'h3b290146),
	.w4(32'hba99ef10),
	.w5(32'h3b44ca8b),
	.w6(32'hbae0d601),
	.w7(32'h3ab8563e),
	.w8(32'h3a18f614),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dd55a),
	.w1(32'hbb3c110d),
	.w2(32'hbb4ec2e0),
	.w3(32'h3b441d8a),
	.w4(32'hbb143b27),
	.w5(32'hbbb573dc),
	.w6(32'h39ff549a),
	.w7(32'hbbb3d5f9),
	.w8(32'hbb3c8ebf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcc5a9),
	.w1(32'hbaae6c98),
	.w2(32'hbb811167),
	.w3(32'hbbd9c52c),
	.w4(32'hbbd26a29),
	.w5(32'hbb64b283),
	.w6(32'hbb83bae5),
	.w7(32'hbbaa8c01),
	.w8(32'hbae01db8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb451996),
	.w1(32'h3b19907f),
	.w2(32'h3ae0bf93),
	.w3(32'hbab81180),
	.w4(32'hbaa80906),
	.w5(32'hba97526f),
	.w6(32'hbb9fc403),
	.w7(32'h3b808cbe),
	.w8(32'hbb2de49a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70cb4b),
	.w1(32'hbb8dfbe1),
	.w2(32'hbb05fef0),
	.w3(32'h3b586775),
	.w4(32'hbc0e6bef),
	.w5(32'hba865029),
	.w6(32'h3b1eccd1),
	.w7(32'hba426fc9),
	.w8(32'hbb129796),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6ae61),
	.w1(32'hbbf37a1c),
	.w2(32'hbbe30dfb),
	.w3(32'hbac02d9e),
	.w4(32'hbb7fd4ef),
	.w5(32'hbbe606e1),
	.w6(32'h3aa3e5b9),
	.w7(32'hbbe48781),
	.w8(32'hbb65f68e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31bd24),
	.w1(32'h3a6f7606),
	.w2(32'hbb0bd0d3),
	.w3(32'hbbe17f20),
	.w4(32'hbb456716),
	.w5(32'hbbb193b1),
	.w6(32'hbbb776e2),
	.w7(32'hbba3bb33),
	.w8(32'hbac5ed3f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd53f1d),
	.w1(32'hbb9bfc49),
	.w2(32'hbc05ae38),
	.w3(32'hbb6a1d56),
	.w4(32'h3b058db5),
	.w5(32'hbaebd8d0),
	.w6(32'hba821be8),
	.w7(32'hbb7b7b09),
	.w8(32'hbb19cd3b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bcfad),
	.w1(32'hbb0cfe22),
	.w2(32'hba9ef9b7),
	.w3(32'h3982f49d),
	.w4(32'hbb41d005),
	.w5(32'hbbd0aa2b),
	.w6(32'hbb902620),
	.w7(32'hbc0f69fc),
	.w8(32'hbbb5912e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69ada1),
	.w1(32'h3bbc66aa),
	.w2(32'hb9a8aafd),
	.w3(32'hba72f554),
	.w4(32'hbb5f9bf1),
	.w5(32'hbc43ee37),
	.w6(32'hbb509cf2),
	.w7(32'hbb9a1b04),
	.w8(32'hbc210bbe),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07c705),
	.w1(32'h3a680406),
	.w2(32'h3ac8d36f),
	.w3(32'h3bea4ed5),
	.w4(32'h3b56d16d),
	.w5(32'hbb5186a7),
	.w6(32'h3a68dd87),
	.w7(32'h3ae38345),
	.w8(32'h39067905),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa2daf),
	.w1(32'hbad1afc1),
	.w2(32'h3b15ef21),
	.w3(32'h3bc0e40d),
	.w4(32'hbb4626f5),
	.w5(32'hbc39b96c),
	.w6(32'h3bceece5),
	.w7(32'h3b60c9cf),
	.w8(32'hbba86417),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08acf3),
	.w1(32'hbb09c2ed),
	.w2(32'hbb487dcf),
	.w3(32'hbb99efee),
	.w4(32'h3b88a348),
	.w5(32'h3ccb9374),
	.w6(32'hbaa810a0),
	.w7(32'h3bdfc8c6),
	.w8(32'hbc280a6d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba558469),
	.w1(32'hba6da5d7),
	.w2(32'hbbf6dbcd),
	.w3(32'hbbfdf6c7),
	.w4(32'hbb93f79c),
	.w5(32'hbc2dbb9e),
	.w6(32'h3ba532e6),
	.w7(32'hbc0539ad),
	.w8(32'hbc314bdf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab23a88),
	.w1(32'h3ac8bd5c),
	.w2(32'h3c882903),
	.w3(32'hbc038fe0),
	.w4(32'h3c2f7b70),
	.w5(32'h3c9c50a5),
	.w6(32'hbbed2e1b),
	.w7(32'h3c3e279a),
	.w8(32'h3b739538),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29395c),
	.w1(32'hbae01d4b),
	.w2(32'h3b71586e),
	.w3(32'h3b27f2a9),
	.w4(32'h3bcfb881),
	.w5(32'h3c6f36e5),
	.w6(32'hb998fb49),
	.w7(32'h3b146200),
	.w8(32'hb9f25eff),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa4525),
	.w1(32'h3b482f9a),
	.w2(32'h3b113ae2),
	.w3(32'h3bb817c1),
	.w4(32'hba9f5d48),
	.w5(32'hbad43b19),
	.w6(32'h3ba1648c),
	.w7(32'h3a3d16e4),
	.w8(32'hbbb7df04),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada123a),
	.w1(32'h3b2d94e8),
	.w2(32'h3bb29188),
	.w3(32'hbb6fc2f4),
	.w4(32'hbb915de8),
	.w5(32'h3c715fc4),
	.w6(32'hbb678737),
	.w7(32'h3b4de697),
	.w8(32'h3c24c2f4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc387d),
	.w1(32'hb7a75bb0),
	.w2(32'h39a69303),
	.w3(32'hbafe7d25),
	.w4(32'h3b5024f6),
	.w5(32'h3bfd320e),
	.w6(32'hbb093e18),
	.w7(32'hbb472248),
	.w8(32'hbac1a82c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e3072),
	.w1(32'h3b670b1d),
	.w2(32'hbbb81656),
	.w3(32'hbc041724),
	.w4(32'h3b6a1421),
	.w5(32'h3a0bc4db),
	.w6(32'h3b2c0a00),
	.w7(32'hbba322fa),
	.w8(32'hbb24d84d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05672e),
	.w1(32'h3ba5ad98),
	.w2(32'hb92118e5),
	.w3(32'h3b8d59fc),
	.w4(32'hbb6b6f56),
	.w5(32'hbb520055),
	.w6(32'h3c0b2f6f),
	.w7(32'hbb31cce1),
	.w8(32'hbb956ace),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82c879),
	.w1(32'h3bdd599e),
	.w2(32'h3b41dd27),
	.w3(32'hbbbf8548),
	.w4(32'hbaf5997e),
	.w5(32'h3b0c7a7b),
	.w6(32'hbb813857),
	.w7(32'hbbf19e00),
	.w8(32'hbb5520d9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3231db),
	.w1(32'hbbcb2cf2),
	.w2(32'hbb0a2e86),
	.w3(32'h3ada2f76),
	.w4(32'hbb78b4bb),
	.w5(32'hbbe5e2a4),
	.w6(32'hb89c67a8),
	.w7(32'hbbcfa969),
	.w8(32'hbb9ba613),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bd421),
	.w1(32'h3ab93728),
	.w2(32'h3b90f0b2),
	.w3(32'hba9db3ed),
	.w4(32'h3a77c106),
	.w5(32'h3c6584d5),
	.w6(32'h3a265d88),
	.w7(32'h3a9a1e1d),
	.w8(32'hbb44ff13),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b110c38),
	.w1(32'h3a07fb28),
	.w2(32'hbb31aa7d),
	.w3(32'h3b918010),
	.w4(32'hbb513767),
	.w5(32'hbc1f9b6f),
	.w6(32'h3ae423b5),
	.w7(32'h3c1390b2),
	.w8(32'h3b267a30),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8855fa),
	.w1(32'h399079a8),
	.w2(32'h3a20066b),
	.w3(32'hba52ec8a),
	.w4(32'hbb3f74fc),
	.w5(32'hbbc79ce7),
	.w6(32'h3bedc7f7),
	.w7(32'hbb0459c6),
	.w8(32'hba1f468e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992bbac),
	.w1(32'hbb6a2e6b),
	.w2(32'hbb44fb96),
	.w3(32'hbb9eaaad),
	.w4(32'hb85ac790),
	.w5(32'hb9a35b9c),
	.w6(32'hbaa242ac),
	.w7(32'h3bd2a0b2),
	.w8(32'h3a973dd9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb12ed6),
	.w1(32'h3b20afbb),
	.w2(32'h3b6ec33f),
	.w3(32'hbba39bba),
	.w4(32'h3bbe1d36),
	.w5(32'hb9f5b5c1),
	.w6(32'hbba04304),
	.w7(32'h3b5feafc),
	.w8(32'h3beca910),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ef03c),
	.w1(32'h3c08b56d),
	.w2(32'h3c16e195),
	.w3(32'hba874b61),
	.w4(32'h3ba3314f),
	.w5(32'h3ae3b6c9),
	.w6(32'hb8caedfc),
	.w7(32'h3ad803f2),
	.w8(32'hbb19d3a2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8a130),
	.w1(32'h3b6bf622),
	.w2(32'h3bcd91d2),
	.w3(32'hbb38b3e3),
	.w4(32'h39c91ac6),
	.w5(32'h3c316886),
	.w6(32'hbc240d25),
	.w7(32'h3b88480b),
	.w8(32'h3b8a8c9e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ae072),
	.w1(32'hb9fa43cd),
	.w2(32'hba3d47f9),
	.w3(32'hba8ef856),
	.w4(32'hbb28bc1f),
	.w5(32'h3b8906bb),
	.w6(32'hbbadd09b),
	.w7(32'hbaecd58b),
	.w8(32'h3b08164f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1759c7),
	.w1(32'hbaee9718),
	.w2(32'h3b43432a),
	.w3(32'h3c1db567),
	.w4(32'h3b8ebdf6),
	.w5(32'h39a102bc),
	.w6(32'h3a9be7dd),
	.w7(32'h3b263a85),
	.w8(32'h3a2f1e2e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba868621),
	.w1(32'h3bbb9c7b),
	.w2(32'h3c032753),
	.w3(32'h3a138100),
	.w4(32'hb82c58d2),
	.w5(32'h3be0df63),
	.w6(32'h36e0cf99),
	.w7(32'h3b1202f6),
	.w8(32'h3b3204d6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16bf79),
	.w1(32'hbb51c5cc),
	.w2(32'hbb73d4d1),
	.w3(32'h38f6b960),
	.w4(32'hbb632120),
	.w5(32'h3ad8b8e1),
	.w6(32'hbb7bbbca),
	.w7(32'hbc009913),
	.w8(32'hbc49b648),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb990cf5),
	.w1(32'hbbf71f8a),
	.w2(32'hbab32456),
	.w3(32'hbb8f6a74),
	.w4(32'hbbf33f56),
	.w5(32'h3ab4dd2b),
	.w6(32'hbc0a9f0d),
	.w7(32'hbb648456),
	.w8(32'hbb1fe4f9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277a59),
	.w1(32'hbb65bff5),
	.w2(32'hbc401010),
	.w3(32'hbb69575f),
	.w4(32'hbb476b1d),
	.w5(32'hbc0f9a55),
	.w6(32'hbb77e818),
	.w7(32'hbb972fff),
	.w8(32'hbb811c6c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c467e),
	.w1(32'h3891d52a),
	.w2(32'hb9c96bb3),
	.w3(32'hbbc649fa),
	.w4(32'h3ba6f211),
	.w5(32'hbc577a79),
	.w6(32'hbb1a50ed),
	.w7(32'h3bf67821),
	.w8(32'h3be57715),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a442170),
	.w1(32'hbb59484c),
	.w2(32'hba941125),
	.w3(32'h3bdaad32),
	.w4(32'hbbc3a833),
	.w5(32'hbbbf7a34),
	.w6(32'h3bb9a78f),
	.w7(32'hbbd203fb),
	.w8(32'hbb8e87b0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac1347),
	.w1(32'hbb156724),
	.w2(32'h3a96211a),
	.w3(32'hbaa1d45a),
	.w4(32'h3b21c0a1),
	.w5(32'hbb95c24d),
	.w6(32'hbac3dbc0),
	.w7(32'h3c1af879),
	.w8(32'h3b9bfe75),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81f785),
	.w1(32'h3a695f78),
	.w2(32'h3b9f6ebf),
	.w3(32'h3afff688),
	.w4(32'h3b9ff63a),
	.w5(32'h3af51f66),
	.w6(32'h3b2e8da6),
	.w7(32'h3b8d1771),
	.w8(32'h3b99b38f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dbc79),
	.w1(32'hbad305de),
	.w2(32'hba9451c4),
	.w3(32'hbad8e847),
	.w4(32'h39e4501b),
	.w5(32'hbbb4a070),
	.w6(32'h3bc48507),
	.w7(32'h3aebd6d1),
	.w8(32'hbb3c5108),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb846c090),
	.w1(32'h3b9b5776),
	.w2(32'hbc0feffa),
	.w3(32'h392578c2),
	.w4(32'hbb984d49),
	.w5(32'hbc6db600),
	.w6(32'h3b32c1bf),
	.w7(32'hbb453ee1),
	.w8(32'hbafbe96a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48edee),
	.w1(32'hbb2e95dc),
	.w2(32'h3b43ae74),
	.w3(32'h3aa6f02e),
	.w4(32'h3bc80354),
	.w5(32'h3b116994),
	.w6(32'hbb1927f7),
	.w7(32'h3b2d9ca4),
	.w8(32'h3a2a2e06),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3367d),
	.w1(32'hbb479cd7),
	.w2(32'hbc112208),
	.w3(32'h3a12da62),
	.w4(32'h3b814195),
	.w5(32'hbbb5840e),
	.w6(32'h3bcc350d),
	.w7(32'h3bb4f0e0),
	.w8(32'h3b8ec850),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b102c92),
	.w1(32'hbb360d51),
	.w2(32'h3c0d131f),
	.w3(32'h3b778e10),
	.w4(32'hbb8273d6),
	.w5(32'h3a605d14),
	.w6(32'h3bd7f9f0),
	.w7(32'hbaa4ecce),
	.w8(32'h3bfef9fd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babe571),
	.w1(32'h3b08eac1),
	.w2(32'h3bb56b5c),
	.w3(32'hba793485),
	.w4(32'hbb5ab67f),
	.w5(32'hbb57704e),
	.w6(32'hbb5751ae),
	.w7(32'hbb5c8a8b),
	.w8(32'hba92ed94),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d50c),
	.w1(32'h3bae9b8b),
	.w2(32'h3bb3361e),
	.w3(32'h39178e84),
	.w4(32'h3ba09a29),
	.w5(32'h3b8d5faa),
	.w6(32'hbbd42759),
	.w7(32'hbafb239e),
	.w8(32'h39df21a1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd4332),
	.w1(32'hbacab399),
	.w2(32'hbbded1a4),
	.w3(32'h3b9e238e),
	.w4(32'hbb98b919),
	.w5(32'hbab832b1),
	.w6(32'h3b5623f6),
	.w7(32'hbb3d953a),
	.w8(32'hbbf9a818),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d06277),
	.w1(32'hbb59bba0),
	.w2(32'hbb36a6c6),
	.w3(32'hbb0557f0),
	.w4(32'hbbd71dc0),
	.w5(32'hb9e0090a),
	.w6(32'h3a8bcbba),
	.w7(32'hbbbf0a01),
	.w8(32'hbb26f588),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53a1e8),
	.w1(32'hbad14749),
	.w2(32'h3ac09f11),
	.w3(32'hbb4510fc),
	.w4(32'hb9e83fdf),
	.w5(32'hbc748d7a),
	.w6(32'hbbbb4f9a),
	.w7(32'hbb3a1726),
	.w8(32'h3b9f8446),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15ca01),
	.w1(32'hbbb3c869),
	.w2(32'hbb080462),
	.w3(32'h39fb189d),
	.w4(32'hb9e3152f),
	.w5(32'hbbc8c4ac),
	.w6(32'hbb303bfa),
	.w7(32'hbbabad8c),
	.w8(32'h3bcfac94),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf87c7),
	.w1(32'hbac2ff40),
	.w2(32'h39d3a004),
	.w3(32'h3b829dd1),
	.w4(32'hbbca4d47),
	.w5(32'hb8128dec),
	.w6(32'hbb470a48),
	.w7(32'hbab203ce),
	.w8(32'h3bc5287e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8128e4),
	.w1(32'h3b9361fc),
	.w2(32'h3aaf1a19),
	.w3(32'h3ae35216),
	.w4(32'hb9591471),
	.w5(32'h3b994ddd),
	.w6(32'h3b6796a6),
	.w7(32'h3b4c2094),
	.w8(32'hba9ef26c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc34f7),
	.w1(32'hb9a38897),
	.w2(32'hba341dbf),
	.w3(32'hba469866),
	.w4(32'hbbcbd960),
	.w5(32'hbb09472e),
	.w6(32'hbba3d1b8),
	.w7(32'hbb8db4dc),
	.w8(32'hbb21ed7c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86c570),
	.w1(32'h3a0dd641),
	.w2(32'hbb6b7d1c),
	.w3(32'h39460d8e),
	.w4(32'hba3ca85c),
	.w5(32'hbb874a02),
	.w6(32'hbb238e23),
	.w7(32'hba3f2b0e),
	.w8(32'h3a841e88),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4af12),
	.w1(32'h3ab57d94),
	.w2(32'h3bdcdf38),
	.w3(32'h3b4beefc),
	.w4(32'h3b749695),
	.w5(32'hba094ffc),
	.w6(32'h3a5319e8),
	.w7(32'h3b26b618),
	.w8(32'hbb24c4fa),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7beca2),
	.w1(32'h3b7ac699),
	.w2(32'h3bd18623),
	.w3(32'hbbe6f4a2),
	.w4(32'h3b22416b),
	.w5(32'hba8dae07),
	.w6(32'hbb7da89b),
	.w7(32'hb9c4f119),
	.w8(32'h3ad71878),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba948184),
	.w1(32'h3ab28ee6),
	.w2(32'hba8a606a),
	.w3(32'h3c455cd0),
	.w4(32'h3c1196b3),
	.w5(32'hba400e8c),
	.w6(32'h3bf39f23),
	.w7(32'h3ba0817c),
	.w8(32'h3bc5c271),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67b419),
	.w1(32'hbb961ade),
	.w2(32'hbb64e6a0),
	.w3(32'h3c13d192),
	.w4(32'hbadd791d),
	.w5(32'hbba474f0),
	.w6(32'h3c1d6a66),
	.w7(32'h3c04268d),
	.w8(32'hba8cb8ca),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e26e3),
	.w1(32'h39a1b872),
	.w2(32'hbb63795c),
	.w3(32'hbbaa6a5b),
	.w4(32'h3aec2fbc),
	.w5(32'hba7bbe86),
	.w6(32'hbaed1400),
	.w7(32'h3b97b494),
	.w8(32'h3a9aecb6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70f499),
	.w1(32'h3a1b86fd),
	.w2(32'h393c5b26),
	.w3(32'h3a34122e),
	.w4(32'h3a42cd4e),
	.w5(32'hb8900d6b),
	.w6(32'h3a07eac5),
	.w7(32'h39c75279),
	.w8(32'hb821ffc0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e09a95),
	.w1(32'h394dc508),
	.w2(32'hb9a007f3),
	.w3(32'hba006688),
	.w4(32'hb9a932d8),
	.w5(32'hba2a87ae),
	.w6(32'hb98ee7da),
	.w7(32'hba289bd2),
	.w8(32'hba8d8bc2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d725fb),
	.w1(32'hba80cdc4),
	.w2(32'hb9d42768),
	.w3(32'hba22f564),
	.w4(32'hba9a57bf),
	.w5(32'hba8f62c1),
	.w6(32'hba3ade83),
	.w7(32'hbacee671),
	.w8(32'hba4dba24),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fa48b7),
	.w1(32'h39593ab7),
	.w2(32'h3994a17e),
	.w3(32'h39052f09),
	.w4(32'h38b81d55),
	.w5(32'hb88f7abe),
	.w6(32'hba4bc357),
	.w7(32'hb9e2556e),
	.w8(32'hb8fb6d8b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918747a),
	.w1(32'hba702ab6),
	.w2(32'hba5a17fd),
	.w3(32'hb8b0bea3),
	.w4(32'hba196ca4),
	.w5(32'hb9b9fb97),
	.w6(32'hb95fd5b0),
	.w7(32'h3a06e1ee),
	.w8(32'hb9ac33c8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae48a0e),
	.w1(32'hb87bb1ab),
	.w2(32'hba0deae9),
	.w3(32'hbabbc176),
	.w4(32'h3a66034f),
	.w5(32'h39d7a180),
	.w6(32'h3997e7c9),
	.w7(32'h3a8656ac),
	.w8(32'h3a618fe1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a179d),
	.w1(32'hbb33587e),
	.w2(32'hbb55ff61),
	.w3(32'hbaedc6f2),
	.w4(32'hbb147c84),
	.w5(32'hbb34e517),
	.w6(32'h39935e5b),
	.w7(32'hb9678fa2),
	.w8(32'hbaf54c12),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a8939),
	.w1(32'hbb07d280),
	.w2(32'hbb45ad9a),
	.w3(32'hbb9965b8),
	.w4(32'hbb0db9fe),
	.w5(32'hbb236d9b),
	.w6(32'hbb64e6e1),
	.w7(32'hbabdf6ec),
	.w8(32'hbb0ccc3a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b8e7c),
	.w1(32'hba5059c2),
	.w2(32'hbabec0c0),
	.w3(32'h3920a7d9),
	.w4(32'h3a2bdb89),
	.w5(32'hba04d1b3),
	.w6(32'hba04dcc3),
	.w7(32'h393e37c0),
	.w8(32'hba899e52),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3867d016),
	.w1(32'hba8d7a47),
	.w2(32'hbaa48286),
	.w3(32'h39bb69ac),
	.w4(32'hb94ef63e),
	.w5(32'hba9fa7c0),
	.w6(32'h3a08b99c),
	.w7(32'hb9be89df),
	.w8(32'hbaa15367),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbb8e1),
	.w1(32'h3ae3550e),
	.w2(32'hb99d915d),
	.w3(32'hba5edd42),
	.w4(32'h3aca9d80),
	.w5(32'hb99469f0),
	.w6(32'hb9e6d782),
	.w7(32'h3b17cf71),
	.w8(32'h3a52a4b2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4acbb),
	.w1(32'hba592664),
	.w2(32'hbaa5db1e),
	.w3(32'h3ac3e5df),
	.w4(32'hb95fb5ad),
	.w5(32'hba87fb9e),
	.w6(32'h3af878c8),
	.w7(32'hb98d88f7),
	.w8(32'hba29929b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2875a),
	.w1(32'h38f18c6c),
	.w2(32'hb961c5b9),
	.w3(32'hb9874e74),
	.w4(32'hb882a567),
	.w5(32'hb951c654),
	.w6(32'h39d4e841),
	.w7(32'h3a1bc7a1),
	.w8(32'h3a237a38),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd3199),
	.w1(32'hba781d5d),
	.w2(32'hb9f03cd7),
	.w3(32'hb90e8b29),
	.w4(32'hba8f8e68),
	.w5(32'hba2e497c),
	.w6(32'h3a1f32a1),
	.w7(32'hba04ed76),
	.w8(32'hba1fcc45),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c87107),
	.w1(32'hba53b038),
	.w2(32'hba10a36d),
	.w3(32'h393f7f11),
	.w4(32'hba0e6644),
	.w5(32'hba3841c5),
	.w6(32'hb9ce1cfb),
	.w7(32'hba641a3a),
	.w8(32'h376fc5c4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36dde4f4),
	.w1(32'hba3d4490),
	.w2(32'hba1e1d5f),
	.w3(32'h39e27ebd),
	.w4(32'hba26271c),
	.w5(32'hbae046bb),
	.w6(32'h39a4da09),
	.w7(32'hbab4d9ea),
	.w8(32'hba96c584),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0adb11),
	.w1(32'h3ae1b172),
	.w2(32'h3901f29e),
	.w3(32'hbb2d85a0),
	.w4(32'h3ac04405),
	.w5(32'h3a4c6bb1),
	.w6(32'hba79083d),
	.w7(32'h3b66c9e2),
	.w8(32'h3a7d5400),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e0e84),
	.w1(32'h3a91f055),
	.w2(32'h3a7bc54b),
	.w3(32'h3a017f2a),
	.w4(32'hb9f44b2a),
	.w5(32'h3a5d4ff3),
	.w6(32'h39be7c4e),
	.w7(32'hba0f5efc),
	.w8(32'hba772665),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c46b0b),
	.w1(32'hba0a0239),
	.w2(32'hbad4965e),
	.w3(32'h3ab66f96),
	.w4(32'h394e11c9),
	.w5(32'hba0991c8),
	.w6(32'h3ab0a4db),
	.w7(32'h3b22b6e5),
	.w8(32'h3a82b77f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb428ce9),
	.w1(32'hbb18572c),
	.w2(32'hbb66a7bc),
	.w3(32'hbb18195b),
	.w4(32'hba6979d1),
	.w5(32'hbab1fedf),
	.w6(32'hb96a87c6),
	.w7(32'hb99189a8),
	.w8(32'hba9a2212),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3ba4e),
	.w1(32'h3aa78053),
	.w2(32'h3981e310),
	.w3(32'hbb409460),
	.w4(32'hb92e5e9a),
	.w5(32'hba5e1ff1),
	.w6(32'hbb0daa1c),
	.w7(32'h38d520b4),
	.w8(32'h3a011c58),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb476449),
	.w1(32'hbb1c7f4a),
	.w2(32'hbb4133b3),
	.w3(32'hba94ba23),
	.w4(32'hba2cae27),
	.w5(32'hbb1b1f22),
	.w6(32'h398e265b),
	.w7(32'h3b38ca47),
	.w8(32'hba938119),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b1a8a0),
	.w1(32'h3aa27127),
	.w2(32'hba967d68),
	.w3(32'h39d8c3f5),
	.w4(32'h3abf11f6),
	.w5(32'hba7eecf8),
	.w6(32'h3ad5fd92),
	.w7(32'h3aed60ff),
	.w8(32'hba3e49e6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63c1c5),
	.w1(32'hbb4dd2b3),
	.w2(32'hbb962134),
	.w3(32'hbaa8e861),
	.w4(32'h39b8e6af),
	.w5(32'hba4937b7),
	.w6(32'h39587bb2),
	.w7(32'h39354702),
	.w8(32'hba34d1d7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ac83a),
	.w1(32'hba2aee54),
	.w2(32'hbb109f3f),
	.w3(32'h3ab2dfa2),
	.w4(32'hba1191fb),
	.w5(32'hbb2496c0),
	.w6(32'h3afeb144),
	.w7(32'h3b376b8f),
	.w8(32'h3a48ce27),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada8ec8),
	.w1(32'h3aa0f1a4),
	.w2(32'hba04872b),
	.w3(32'hbacba8da),
	.w4(32'h3ac4a9e9),
	.w5(32'hbad46d1a),
	.w6(32'h39b94ead),
	.w7(32'h3a96308a),
	.w8(32'h398b8ed1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e96a35),
	.w1(32'hb9b7ae9d),
	.w2(32'hb7a13f03),
	.w3(32'h39b55ac9),
	.w4(32'hb965b895),
	.w5(32'hba1052f8),
	.w6(32'hb9414086),
	.w7(32'hba818b70),
	.w8(32'hba21b42e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa8397),
	.w1(32'hbb1048be),
	.w2(32'hbb996321),
	.w3(32'hb9ac8596),
	.w4(32'hba387244),
	.w5(32'hbb264eed),
	.w6(32'h39903519),
	.w7(32'hba216b0d),
	.w8(32'hbb319e44),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee539),
	.w1(32'hbaac9d6d),
	.w2(32'hbb027ad2),
	.w3(32'hbab58d28),
	.w4(32'h3a13f2f2),
	.w5(32'hb9b11737),
	.w6(32'h3a8ed192),
	.w7(32'h3ab290d0),
	.w8(32'h3a05f8a5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba45b82),
	.w1(32'h39612966),
	.w2(32'hbb15f67b),
	.w3(32'hb9eba5bc),
	.w4(32'h3a4f8d8f),
	.w5(32'hbb4abd36),
	.w6(32'hba41656e),
	.w7(32'h3ab01e10),
	.w8(32'hbb420387),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad67307),
	.w1(32'h3ba45bf8),
	.w2(32'h3b62a655),
	.w3(32'hbb255e7a),
	.w4(32'h3b97bbd3),
	.w5(32'h3b14683a),
	.w6(32'h3a8d6f78),
	.w7(32'h3bfea4a2),
	.w8(32'h3b8ddd97),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb299b28),
	.w1(32'hbb808cc6),
	.w2(32'hbbb97a7f),
	.w3(32'hbabe07d9),
	.w4(32'hbb0faf75),
	.w5(32'hbb88346e),
	.w6(32'hbaa4b00e),
	.w7(32'hba6b9549),
	.w8(32'hbb328a3d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b53b5),
	.w1(32'h39f4c317),
	.w2(32'hbb00d637),
	.w3(32'h38bdd2e2),
	.w4(32'hb9242b8b),
	.w5(32'hbb433437),
	.w6(32'h3af0b3b3),
	.w7(32'h3b33bfba),
	.w8(32'hbaa16644),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38cf49),
	.w1(32'hba1d8e7d),
	.w2(32'h38cfa217),
	.w3(32'h3a076659),
	.w4(32'hb94c566d),
	.w5(32'hbaa3e6f7),
	.w6(32'h39b2dabf),
	.w7(32'h3a031669),
	.w8(32'h39b615ad),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb426ca0),
	.w1(32'hbab9f826),
	.w2(32'hbb01f960),
	.w3(32'hbab66ea1),
	.w4(32'h3b2ff4f7),
	.w5(32'hba3498c0),
	.w6(32'hba33d2f2),
	.w7(32'h3aedf765),
	.w8(32'hbb0a3a1b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7d6eb),
	.w1(32'hb99ad7b2),
	.w2(32'hbb078d63),
	.w3(32'hba98d2bf),
	.w4(32'hba597446),
	.w5(32'hbb122175),
	.w6(32'hba5df33f),
	.w7(32'hb99287b1),
	.w8(32'hbb03a412),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba808cd0),
	.w1(32'h38cf1c03),
	.w2(32'h398c1b4a),
	.w3(32'hba285985),
	.w4(32'h361810e1),
	.w5(32'hb9ed8335),
	.w6(32'hb98dc35d),
	.w7(32'hb8135d5f),
	.w8(32'hb96a5c4b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f3e6b),
	.w1(32'hba38d57e),
	.w2(32'hba622bf4),
	.w3(32'hba1ec83d),
	.w4(32'h39d898f7),
	.w5(32'h3920c6ce),
	.w6(32'hb9cf4a4f),
	.w7(32'h38ee6479),
	.w8(32'h3960f51f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb144929),
	.w1(32'hbb50f586),
	.w2(32'hbb828ff9),
	.w3(32'hb88a98fb),
	.w4(32'hbb08a34a),
	.w5(32'hbb38a1fa),
	.w6(32'hba9c8966),
	.w7(32'hbb0630c2),
	.w8(32'hbb4b618b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93cc53),
	.w1(32'hba8f2c57),
	.w2(32'hbb38c15e),
	.w3(32'h3a1b2645),
	.w4(32'hba0be3a7),
	.w5(32'hbb1a2105),
	.w6(32'hb9292849),
	.w7(32'hba56dd06),
	.w8(32'hbb4f4a6e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c0037),
	.w1(32'hba82df90),
	.w2(32'hbafcb5d1),
	.w3(32'hbabf9f41),
	.w4(32'h39adb019),
	.w5(32'hb8362fe4),
	.w6(32'hbb1b09ef),
	.w7(32'hb96da3cd),
	.w8(32'hba52cdcd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f84a8),
	.w1(32'hbaa0c5c6),
	.w2(32'hbb123c6e),
	.w3(32'hb9e34222),
	.w4(32'hba272ca9),
	.w5(32'hbb16dfc4),
	.w6(32'hba991e04),
	.w7(32'h38525bed),
	.w8(32'hba70683c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7fe4c),
	.w1(32'h3a511043),
	.w2(32'h39259600),
	.w3(32'hbb0ed582),
	.w4(32'hb9a802b6),
	.w5(32'hba28242f),
	.w6(32'hbb16b791),
	.w7(32'h3a42857d),
	.w8(32'h3a46e972),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ad438),
	.w1(32'hbb36172d),
	.w2(32'hbb3b0a98),
	.w3(32'hb9a67ee3),
	.w4(32'hba81204f),
	.w5(32'hbb0d684b),
	.w6(32'h39039e17),
	.w7(32'hb98d2049),
	.w8(32'hba743979),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73ca6c),
	.w1(32'hb9740715),
	.w2(32'hbaa60b96),
	.w3(32'hba95b052),
	.w4(32'h3a970118),
	.w5(32'h39af23be),
	.w6(32'hba420fcb),
	.w7(32'h3ac1d731),
	.w8(32'h39651ca3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6027c),
	.w1(32'hba4bafce),
	.w2(32'hba6362f0),
	.w3(32'h3a0f80da),
	.w4(32'hb98fb77e),
	.w5(32'hba14278b),
	.w6(32'h3a89a7ae),
	.w7(32'hb9edc0d5),
	.w8(32'hba07b292),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe4d46),
	.w1(32'hba2b6445),
	.w2(32'hba0d9885),
	.w3(32'hbadf810f),
	.w4(32'hb9cb68b9),
	.w5(32'hb9db6219),
	.w6(32'hba9caa0f),
	.w7(32'hba8eaa71),
	.w8(32'hb915ed68),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd54cb),
	.w1(32'hb90cf0df),
	.w2(32'hba36c50c),
	.w3(32'h39ce27b5),
	.w4(32'h3a7c73dc),
	.w5(32'h39d6be48),
	.w6(32'h39dd77d2),
	.w7(32'h3970486b),
	.w8(32'hba0ed36b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a12d37),
	.w1(32'h39db65d0),
	.w2(32'h3a196af7),
	.w3(32'h39787d8c),
	.w4(32'hba47f488),
	.w5(32'h3a38e0f7),
	.w6(32'h38259a6c),
	.w7(32'hb9e09bf8),
	.w8(32'hba17d8ed),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02c65c),
	.w1(32'hba681ce9),
	.w2(32'hbaebda09),
	.w3(32'h39327b77),
	.w4(32'h3a1742ec),
	.w5(32'hbac1e86d),
	.w6(32'hb9dd8004),
	.w7(32'h3ace2abc),
	.w8(32'h39e45205),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb879b606),
	.w1(32'hb9dd0aa6),
	.w2(32'hb87a2d3d),
	.w3(32'h3a665291),
	.w4(32'hba0f3786),
	.w5(32'hb95c16b1),
	.w6(32'h3ad7cc0b),
	.w7(32'hb9abfeb2),
	.w8(32'h393690ec),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a1837),
	.w1(32'hb8a64190),
	.w2(32'hbadbe867),
	.w3(32'hba27599d),
	.w4(32'hb9f7197c),
	.w5(32'hbab4192d),
	.w6(32'h3a725872),
	.w7(32'h392d4164),
	.w8(32'hb882239c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29595b),
	.w1(32'hba526759),
	.w2(32'hba7f98b6),
	.w3(32'hbac3b1dc),
	.w4(32'hb99226fa),
	.w5(32'hba96a1c9),
	.w6(32'hba02347d),
	.w7(32'h3914d253),
	.w8(32'hbab64c62),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377b8ecc),
	.w1(32'hb733f654),
	.w2(32'hba269c4f),
	.w3(32'hba051477),
	.w4(32'hb97dfaac),
	.w5(32'hbae6e216),
	.w6(32'h3967ecb2),
	.w7(32'h39fe0130),
	.w8(32'hb90f3f4f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a7c6c),
	.w1(32'hba31f859),
	.w2(32'hba526236),
	.w3(32'hba2c09cc),
	.w4(32'hbaa62d15),
	.w5(32'hba9caa44),
	.w6(32'hb9d303d1),
	.w7(32'hbabce8ca),
	.w8(32'hba578902),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a34e23),
	.w1(32'h392cb91d),
	.w2(32'hb8986f54),
	.w3(32'hb9a93b1a),
	.w4(32'h3953dc90),
	.w5(32'h399806c0),
	.w6(32'hb9465b85),
	.w7(32'hb9abdca5),
	.w8(32'hbab31f0b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b6263),
	.w1(32'hbac83eb1),
	.w2(32'hbad38a8e),
	.w3(32'hb8cfc1ae),
	.w4(32'h393d54db),
	.w5(32'hb9bd7ddb),
	.w6(32'hbacfbf4b),
	.w7(32'h3a3e1d62),
	.w8(32'h39f650eb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c3d4d),
	.w1(32'hbb0023be),
	.w2(32'hbaea2efc),
	.w3(32'h3a9a5de0),
	.w4(32'hba5f01e3),
	.w5(32'hbb05891c),
	.w6(32'h393ec2e6),
	.w7(32'h3975897f),
	.w8(32'hbb1533e0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba925e12),
	.w1(32'hbb073ed6),
	.w2(32'hbb81dad3),
	.w3(32'hbaa3b144),
	.w4(32'hb9a3019c),
	.w5(32'hbb0e6378),
	.w6(32'hba3503dd),
	.w7(32'h3a7e38d4),
	.w8(32'hbaf3bbc2),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0559d2),
	.w1(32'hb9e900db),
	.w2(32'hba092d1f),
	.w3(32'h3991ea87),
	.w4(32'hb978c63f),
	.w5(32'hbaadeab8),
	.w6(32'h39cc7d5c),
	.w7(32'hba28219b),
	.w8(32'hbaa04686),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb6b34),
	.w1(32'hbab4f45d),
	.w2(32'hba8bba15),
	.w3(32'hbb1cc1c2),
	.w4(32'hbaed29bb),
	.w5(32'hba8d1b69),
	.w6(32'hbb1885c3),
	.w7(32'hba7bc3be),
	.w8(32'hb910626a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909fd0e),
	.w1(32'h38c7b791),
	.w2(32'hb9ef8f7f),
	.w3(32'hb62b81cc),
	.w4(32'hb8d5c918),
	.w5(32'hb9d47b39),
	.w6(32'h39e0a273),
	.w7(32'h38a09091),
	.w8(32'hb8aa6bab),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcc87b),
	.w1(32'hba64c39a),
	.w2(32'hbae0d523),
	.w3(32'hba5d0659),
	.w4(32'hba054159),
	.w5(32'hba7abfc1),
	.w6(32'hba0cacef),
	.w7(32'hb9d90e7c),
	.w8(32'hba10eb52),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafb580),
	.w1(32'hbaed2439),
	.w2(32'hbb3df4e1),
	.w3(32'hba1de7ed),
	.w4(32'hba32f4f0),
	.w5(32'hbaeb102d),
	.w6(32'h3a2d4ab9),
	.w7(32'hb9a4216a),
	.w8(32'hb7a554c0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4e25e),
	.w1(32'hb9c3e5c3),
	.w2(32'hbb3a3feb),
	.w3(32'hb9c72838),
	.w4(32'hb9de872c),
	.w5(32'hbb112111),
	.w6(32'h399d3626),
	.w7(32'hba454287),
	.w8(32'hbb5d933b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39064529),
	.w1(32'hb9686577),
	.w2(32'hbacd84bf),
	.w3(32'hb92814c5),
	.w4(32'h3a3baa2f),
	.w5(32'hb9ab980c),
	.w6(32'hba9b771b),
	.w7(32'hb8849c63),
	.w8(32'hbaa3ee7e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39260c75),
	.w1(32'hba3ddd6e),
	.w2(32'hbb2324c1),
	.w3(32'h3a8ac095),
	.w4(32'h3ad348dd),
	.w5(32'hba7c3638),
	.w6(32'h3a44231e),
	.w7(32'h3b2e444a),
	.w8(32'h3904e356),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5d1a8),
	.w1(32'hba844ade),
	.w2(32'hbb4fc158),
	.w3(32'hb9c4f82d),
	.w4(32'h39d838c4),
	.w5(32'hbad3fbe9),
	.w6(32'h3a33b360),
	.w7(32'hb9876105),
	.w8(32'hbb08a990),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ae996),
	.w1(32'hbaa2e6c5),
	.w2(32'hbaf05731),
	.w3(32'hba6cb1d8),
	.w4(32'hb9ec8f71),
	.w5(32'hbac5b530),
	.w6(32'hba9566c5),
	.w7(32'h37e56b5f),
	.w8(32'hba900d1e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba775e1d),
	.w1(32'hbad3e8bc),
	.w2(32'hbb4fbab7),
	.w3(32'hb89c56c1),
	.w4(32'hba9003af),
	.w5(32'hbaef34a5),
	.w6(32'h3a8345cc),
	.w7(32'h398a8158),
	.w8(32'hba37f68a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba491de1),
	.w1(32'hb80db257),
	.w2(32'h378b2f63),
	.w3(32'hba54808e),
	.w4(32'h3a35a4c8),
	.w5(32'h371f022f),
	.w6(32'h3a0496bf),
	.w7(32'h3a19fb49),
	.w8(32'hb7ea3f51),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93fe0f4),
	.w1(32'h3b32e883),
	.w2(32'h3858077f),
	.w3(32'hbad7f54f),
	.w4(32'h3ab080da),
	.w5(32'hbb003a43),
	.w6(32'hba7cc802),
	.w7(32'h3b5e0210),
	.w8(32'h3aba0ff1),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4dd208),
	.w1(32'h382505e3),
	.w2(32'hb98a5692),
	.w3(32'h3a9a9f96),
	.w4(32'h3a5f6c9b),
	.w5(32'hb9c9b14f),
	.w6(32'h3af39c93),
	.w7(32'h39ceb1f2),
	.w8(32'h39a67ed0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d469e2),
	.w1(32'hb9c208ff),
	.w2(32'h3691848c),
	.w3(32'h39bcf214),
	.w4(32'hb9681222),
	.w5(32'h395a2f94),
	.w6(32'h387cd50e),
	.w7(32'h3969f331),
	.w8(32'h3a4e6d07),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a072db9),
	.w1(32'hb9d7a7af),
	.w2(32'hb9c10a35),
	.w3(32'h37d29aac),
	.w4(32'hb9e7f941),
	.w5(32'hb8c29aab),
	.w6(32'h3a36d087),
	.w7(32'hba8df891),
	.w8(32'hba2c0796),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba690f63),
	.w1(32'h39fe0f39),
	.w2(32'hb95275c3),
	.w3(32'hba289bf3),
	.w4(32'hb99e880c),
	.w5(32'hb9fc7c7f),
	.w6(32'hba6aeb4f),
	.w7(32'h3a514b41),
	.w8(32'hb91343ab),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadc7c8),
	.w1(32'hba7a1983),
	.w2(32'hbb1566ac),
	.w3(32'h39d6e4f3),
	.w4(32'h3abc852d),
	.w5(32'hbae6d770),
	.w6(32'h3abfc1ae),
	.w7(32'h3b09169f),
	.w8(32'hb9daa7fd),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f8934),
	.w1(32'hbb5ec04c),
	.w2(32'hbb693459),
	.w3(32'hbb6551de),
	.w4(32'hbb3e8f16),
	.w5(32'hbb40b63b),
	.w6(32'hbb4f06fa),
	.w7(32'hbb60c409),
	.w8(32'hbb3a8e10),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d21c71),
	.w1(32'h3916a61e),
	.w2(32'hb9b04663),
	.w3(32'hbad95f48),
	.w4(32'h39b7ad76),
	.w5(32'hb97a7a5b),
	.w6(32'hb9a7e185),
	.w7(32'h3926b045),
	.w8(32'hb9aaa134),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91c2a0),
	.w1(32'hbb350075),
	.w2(32'hbb3cbb1d),
	.w3(32'hba0a99fb),
	.w4(32'hba6acb79),
	.w5(32'hba91b09d),
	.w6(32'h39b43eb0),
	.w7(32'hbb048d79),
	.w8(32'hbb00ff44),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393068b2),
	.w1(32'hbacc67ec),
	.w2(32'hbb6280ba),
	.w3(32'h3a0c99ab),
	.w4(32'hb9f0e858),
	.w5(32'hba987ab2),
	.w6(32'h3a5d19f1),
	.w7(32'h38fbec77),
	.w8(32'hba975b4f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7257),
	.w1(32'hbaebc070),
	.w2(32'hbb86a2c1),
	.w3(32'hb9afb367),
	.w4(32'hbb377697),
	.w5(32'hbb9e9993),
	.w6(32'hb95676a2),
	.w7(32'hba9534e7),
	.w8(32'hbb373ba3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b0e29),
	.w1(32'h3ad0e12c),
	.w2(32'hbaeda3f5),
	.w3(32'hbb1005cb),
	.w4(32'h3af9526b),
	.w5(32'hbaaa2e10),
	.w6(32'hbada140c),
	.w7(32'h3ac38e19),
	.w8(32'h3a3fd32f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386f5b26),
	.w1(32'hb7c90569),
	.w2(32'hba8d55a9),
	.w3(32'hb92706a9),
	.w4(32'hb7495466),
	.w5(32'hbb0932b4),
	.w6(32'hb98269b8),
	.w7(32'h3a09bb31),
	.w8(32'hba3e57f6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e3a61),
	.w1(32'hba9c6bb1),
	.w2(32'hb958e622),
	.w3(32'hbac7365d),
	.w4(32'hbab4eb99),
	.w5(32'hba85ff49),
	.w6(32'h39193252),
	.w7(32'hba860e95),
	.w8(32'hba4b63fc),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee0b6e),
	.w1(32'h39cece11),
	.w2(32'hba332941),
	.w3(32'hb933ec58),
	.w4(32'h3a2c02a7),
	.w5(32'hba4ca80b),
	.w6(32'hba91bb8f),
	.w7(32'h3a9d174a),
	.w8(32'h3a3c6dd4),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e54065),
	.w1(32'h3a0375f1),
	.w2(32'hba279144),
	.w3(32'hba0f2c11),
	.w4(32'h3b1b68ca),
	.w5(32'h39d0fd32),
	.w6(32'h3a555fae),
	.w7(32'h3b774a97),
	.w8(32'h394f5e05),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bbbe8),
	.w1(32'h3a9f286e),
	.w2(32'h3a8debe4),
	.w3(32'hbaf89959),
	.w4(32'h3a9d50da),
	.w5(32'h3a1660c9),
	.w6(32'hbb02db73),
	.w7(32'h3ad7df90),
	.w8(32'h3a51440e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8210b7d),
	.w1(32'hb9b5191d),
	.w2(32'hbab6d66d),
	.w3(32'hba14cee0),
	.w4(32'hb99c633b),
	.w5(32'hb9408b6b),
	.w6(32'h39548fac),
	.w7(32'h39ba37d6),
	.w8(32'hb9f7c164),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e75180),
	.w1(32'hb9c50dc5),
	.w2(32'hba04d09c),
	.w3(32'h39d4e6e3),
	.w4(32'h382aec65),
	.w5(32'hba09a465),
	.w6(32'hba0815bc),
	.w7(32'hb97a4712),
	.w8(32'h39bf7805),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6acc15),
	.w1(32'hba8191c4),
	.w2(32'hbb03f7e5),
	.w3(32'h3a858948),
	.w4(32'h387140ee),
	.w5(32'hba802311),
	.w6(32'h3ab858e9),
	.w7(32'h385e7366),
	.w8(32'hba67be4b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394da77b),
	.w1(32'hb9d9a9c5),
	.w2(32'hba860782),
	.w3(32'h397cad46),
	.w4(32'hba81cb4e),
	.w5(32'hba3b0862),
	.w6(32'h395f2bcf),
	.w7(32'hb9a4e2bd),
	.w8(32'hba04b3bd),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22ba92),
	.w1(32'h3aa072c9),
	.w2(32'h38456c4f),
	.w3(32'h3aa0a30f),
	.w4(32'h3a929ff6),
	.w5(32'hb938a144),
	.w6(32'hb4d0e8dc),
	.w7(32'h3af3633a),
	.w8(32'h3ab081b3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acaf935),
	.w1(32'h398b7ab7),
	.w2(32'h391f3e1e),
	.w3(32'h3a6d3cde),
	.w4(32'h3a09a053),
	.w5(32'h39e9827d),
	.w6(32'h3a9174ef),
	.w7(32'h39378008),
	.w8(32'hb9a056b5),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab85812),
	.w1(32'hba50dafe),
	.w2(32'h39730918),
	.w3(32'hbae092e1),
	.w4(32'hbaca05a5),
	.w5(32'hba86bb33),
	.w6(32'hbab837e8),
	.w7(32'hba7f51e4),
	.w8(32'hb9167be8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0e0ba),
	.w1(32'h39a12325),
	.w2(32'h39fefe41),
	.w3(32'hb978acc9),
	.w4(32'h3a14a6d4),
	.w5(32'h397c6019),
	.w6(32'hb991bd4a),
	.w7(32'h39b9bb7e),
	.w8(32'h3a309256),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e51c1b),
	.w1(32'h38e6c6c7),
	.w2(32'hb9c86093),
	.w3(32'hb9878f5e),
	.w4(32'hba19daf9),
	.w5(32'hbad37b80),
	.w6(32'h3916ccd0),
	.w7(32'hb892b8a5),
	.w8(32'hb9b9eb70),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ba414),
	.w1(32'h39b97e2f),
	.w2(32'hba62dced),
	.w3(32'h39b3bfe4),
	.w4(32'h3a9dc59c),
	.w5(32'h37c6b4d3),
	.w6(32'h3a2b675b),
	.w7(32'h3acd0690),
	.w8(32'h3a444f08),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58683b),
	.w1(32'hbb4f1269),
	.w2(32'hbbad9e97),
	.w3(32'h3b09f957),
	.w4(32'hba9ad5a0),
	.w5(32'hbbb0d438),
	.w6(32'h3b351ead),
	.w7(32'h3b0650b8),
	.w8(32'hbb12f3be),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9ae8),
	.w1(32'hba42622a),
	.w2(32'hb9163970),
	.w3(32'hbb453ebc),
	.w4(32'hbad26bb0),
	.w5(32'hbab6adb4),
	.w6(32'hbad0a4ca),
	.w7(32'hbac2940b),
	.w8(32'hb9518634),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb237647),
	.w1(32'hbb1a55d4),
	.w2(32'hbb6606a5),
	.w3(32'hba8c3b11),
	.w4(32'hba422b66),
	.w5(32'hbb001b82),
	.w6(32'hba5e220b),
	.w7(32'h3956774d),
	.w8(32'hba883feb),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95c7d0),
	.w1(32'h3897f536),
	.w2(32'hba47b50d),
	.w3(32'hbab62b50),
	.w4(32'h396ce849),
	.w5(32'hba75a05b),
	.w6(32'hba7992c0),
	.w7(32'h398373ab),
	.w8(32'hb94d060f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ef41c),
	.w1(32'hbb4d2000),
	.w2(32'hbbbaadb8),
	.w3(32'hbb5e204a),
	.w4(32'hbab6c6b9),
	.w5(32'hbb940e41),
	.w6(32'hbb2267c8),
	.w7(32'hba0ba7b3),
	.w8(32'hbb1d5728),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139baf),
	.w1(32'hbabefaec),
	.w2(32'hbb321a1e),
	.w3(32'hba43da85),
	.w4(32'h38aeaf44),
	.w5(32'hba84e086),
	.w6(32'h3902de7c),
	.w7(32'h39c16bd1),
	.w8(32'hb9ad3afc),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81333f),
	.w1(32'hb9c1c568),
	.w2(32'hbb346c39),
	.w3(32'hb99384c4),
	.w4(32'h3955c7b4),
	.w5(32'hbb0a9f8f),
	.w6(32'h3a1f6e78),
	.w7(32'h395ebc13),
	.w8(32'hbb2ff4a3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f2540),
	.w1(32'hba6eca81),
	.w2(32'hba52efff),
	.w3(32'hba782f6d),
	.w4(32'hba39c35c),
	.w5(32'hba54242e),
	.w6(32'hba4dc50c),
	.w7(32'hba051a24),
	.w8(32'hba81c487),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9485490),
	.w1(32'h394b10c3),
	.w2(32'hbb1778ca),
	.w3(32'h3a654569),
	.w4(32'h3a876098),
	.w5(32'hbae7a0b9),
	.w6(32'h3ac66c2e),
	.w7(32'h3a4302ba),
	.w8(32'hba962b41),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cdeab),
	.w1(32'h390e0a7f),
	.w2(32'h3880cca7),
	.w3(32'hbac060d2),
	.w4(32'hb741eea5),
	.w5(32'hb9d6530e),
	.w6(32'hbaad6298),
	.w7(32'hb8ebacea),
	.w8(32'h389fe5eb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b79ad),
	.w1(32'hb9975c2c),
	.w2(32'hba628f6f),
	.w3(32'hba962585),
	.w4(32'hba4edf5a),
	.w5(32'hba1cd74e),
	.w6(32'h37979ce6),
	.w7(32'hb961fe92),
	.w8(32'hb97e19a4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ae8d7),
	.w1(32'hba8ec6f1),
	.w2(32'hba675faf),
	.w3(32'hb943ffe3),
	.w4(32'hba1995da),
	.w5(32'hba5ec37f),
	.w6(32'hb9024b39),
	.w7(32'hbaaed19a),
	.w8(32'hba9b4780),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dd79b),
	.w1(32'hbab45271),
	.w2(32'hbb3767da),
	.w3(32'hbb1da623),
	.w4(32'hbac2d05a),
	.w5(32'hbad24137),
	.w6(32'hbb1ae6b9),
	.w7(32'hba8e9be4),
	.w8(32'hbacf339b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a052bbb),
	.w1(32'h3ab59558),
	.w2(32'h3a4b40d5),
	.w3(32'h398f2a89),
	.w4(32'h3aa48243),
	.w5(32'h3a8e5dc7),
	.w6(32'h39f93da5),
	.w7(32'h3a425349),
	.w8(32'hb8b8d5c7),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac61932),
	.w1(32'hb8fe0e14),
	.w2(32'h39ee24e9),
	.w3(32'h3a835a65),
	.w4(32'hb9f84cfe),
	.w5(32'h39a171e4),
	.w6(32'h3a302fbc),
	.w7(32'hbab2d12a),
	.w8(32'hba04619e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917e8a1),
	.w1(32'h395d0e82),
	.w2(32'hb9a8685a),
	.w3(32'hb90d0235),
	.w4(32'h3aa3f141),
	.w5(32'h38806d2c),
	.w6(32'hbad61824),
	.w7(32'h3ad9b1e8),
	.w8(32'h38c0199e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb190860),
	.w1(32'hbab2275f),
	.w2(32'hbb19b99f),
	.w3(32'hbaf8c80e),
	.w4(32'hbaaacc0e),
	.w5(32'hbb03ab8f),
	.w6(32'hba8d4758),
	.w7(32'h3843c2e9),
	.w8(32'hba33968b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacccde3),
	.w1(32'hb993faa6),
	.w2(32'hb9532461),
	.w3(32'hb9c77ee2),
	.w4(32'h3a1af798),
	.w5(32'h38dd0d42),
	.w6(32'h3a00de87),
	.w7(32'h399b2455),
	.w8(32'hb9128a3b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96cf355),
	.w1(32'hba87a0a9),
	.w2(32'hbadd7377),
	.w3(32'h3a1fa94c),
	.w4(32'hbaaabac5),
	.w5(32'hbab13ad4),
	.w6(32'h39d2ba72),
	.w7(32'hbad10f61),
	.w8(32'hbadfcf66),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaffff1),
	.w1(32'hbb02e9fc),
	.w2(32'hbbf4686b),
	.w3(32'hbb9d03ce),
	.w4(32'hba9e8170),
	.w5(32'hbb9f4686),
	.w6(32'hbb255103),
	.w7(32'h39c2e271),
	.w8(32'hbb043831),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9440f),
	.w1(32'hb9da4f90),
	.w2(32'hbb7085e3),
	.w3(32'hba9b3430),
	.w4(32'h3b1d63b1),
	.w5(32'hba657183),
	.w6(32'h3af0b06f),
	.w7(32'h3b453142),
	.w8(32'h3a44d633),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba249afb),
	.w1(32'hb9c3f60f),
	.w2(32'hba1205d0),
	.w3(32'h394024d2),
	.w4(32'hb9ebab6c),
	.w5(32'hba9bb281),
	.w6(32'h3933b8b4),
	.w7(32'hb9bb8236),
	.w8(32'hb711c203),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389caf51),
	.w1(32'h394d57c4),
	.w2(32'h37ed447e),
	.w3(32'h3a510084),
	.w4(32'hb969fd5c),
	.w5(32'hba35d525),
	.w6(32'h39afe3d5),
	.w7(32'h37861187),
	.w8(32'h3983b708),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1971e),
	.w1(32'hba5e7b58),
	.w2(32'hbaa52f73),
	.w3(32'hb9ea0cb9),
	.w4(32'hba258394),
	.w5(32'hba1c29e3),
	.w6(32'h3965e68b),
	.w7(32'h39b5bd95),
	.w8(32'hb91df05c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b2ca9),
	.w1(32'h3ad9213f),
	.w2(32'h3a4bad04),
	.w3(32'hbaa39030),
	.w4(32'h3a34bbd5),
	.w5(32'hb9493034),
	.w6(32'hb915efc3),
	.w7(32'h3ac4e911),
	.w8(32'h39f40e9f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04ee12),
	.w1(32'hb9398838),
	.w2(32'hbac7fb33),
	.w3(32'h3ac7ffe6),
	.w4(32'hb974e8e1),
	.w5(32'hbb17eec7),
	.w6(32'h3b1d8ca8),
	.w7(32'h39f942b1),
	.w8(32'hba5abe22),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3d7fc),
	.w1(32'hba546e28),
	.w2(32'hbb25d5c4),
	.w3(32'hb9395f5b),
	.w4(32'h3a85f22d),
	.w5(32'hb9ff2320),
	.w6(32'h3a708513),
	.w7(32'h3aabf42e),
	.w8(32'hbab18942),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb882b46),
	.w1(32'hbb2ac89d),
	.w2(32'hbb5732a6),
	.w3(32'hbb2801a2),
	.w4(32'hb9d498f3),
	.w5(32'hbb136a37),
	.w6(32'hbb4af9bf),
	.w7(32'hba37712a),
	.w8(32'hbaf9f448),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c8180),
	.w1(32'h3812a65b),
	.w2(32'h3a7822a9),
	.w3(32'hba28807e),
	.w4(32'h38ffd430),
	.w5(32'h3a1ba550),
	.w6(32'hbaaaaf3a),
	.w7(32'h3927897c),
	.w8(32'h39b48f12),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02e4cb),
	.w1(32'hbb34951c),
	.w2(32'hbb752533),
	.w3(32'hba4574e3),
	.w4(32'hbac5bbb9),
	.w5(32'hbb251be3),
	.w6(32'hbaa73267),
	.w7(32'hba900e67),
	.w8(32'hbb055785),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801f74),
	.w1(32'hba0f0136),
	.w2(32'hba3ade94),
	.w3(32'hba3f3981),
	.w4(32'hba123905),
	.w5(32'hba54e77c),
	.w6(32'hba64f90e),
	.w7(32'hba2cc06c),
	.w8(32'hba58c595),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3801b557),
	.w1(32'h37744c95),
	.w2(32'h37b4bf1f),
	.w3(32'h379e2b4d),
	.w4(32'h3648a3bf),
	.w5(32'h3729228c),
	.w6(32'h376edb4b),
	.w7(32'h358558b9),
	.w8(32'h37213edb),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86668b),
	.w1(32'hba2ae46a),
	.w2(32'hb7cfc41e),
	.w3(32'hba4014ae),
	.w4(32'hba1b31bc),
	.w5(32'h3993a196),
	.w6(32'hba29b618),
	.w7(32'hb93301b8),
	.w8(32'h36f712d4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3866a17b),
	.w1(32'h379a52d3),
	.w2(32'h38396cc6),
	.w3(32'h3818335d),
	.w4(32'hb55c6614),
	.w5(32'h379b2df0),
	.w6(32'h37ea2c45),
	.w7(32'hb6e3613c),
	.w8(32'h37c0a454),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf0e78),
	.w1(32'hba0efedf),
	.w2(32'hba31c3ac),
	.w3(32'hb9030599),
	.w4(32'h3a0cd050),
	.w5(32'h38369e2c),
	.w6(32'hb9b3cc8a),
	.w7(32'hb778b762),
	.w8(32'hba7b4bdb),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6e0f4),
	.w1(32'h3a784164),
	.w2(32'h3a2805e0),
	.w3(32'hba834476),
	.w4(32'h3b0a6bdd),
	.w5(32'h3a81490b),
	.w6(32'hb9706bf3),
	.w7(32'h3b4c2d18),
	.w8(32'h3ace4798),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91fe06),
	.w1(32'hba5c2a12),
	.w2(32'hbb05628b),
	.w3(32'hb9c15180),
	.w4(32'h392b4549),
	.w5(32'hba8c420e),
	.w6(32'hb880acf6),
	.w7(32'h3a4ea740),
	.w8(32'hba31b876),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ddcc5),
	.w1(32'h39bebc0b),
	.w2(32'h3a33324e),
	.w3(32'hb9f7f61e),
	.w4(32'h37ac0c25),
	.w5(32'h39b18045),
	.w6(32'hba081aae),
	.w7(32'h35f8080b),
	.w8(32'h39d22477),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5d636),
	.w1(32'hbafdb818),
	.w2(32'hbb417e56),
	.w3(32'hba47bbc2),
	.w4(32'h37a1cda9),
	.w5(32'hbaa88e5f),
	.w6(32'hba391953),
	.w7(32'h3980287c),
	.w8(32'hba799465),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1c9a4),
	.w1(32'hba8b5131),
	.w2(32'hbacd8548),
	.w3(32'hba098854),
	.w4(32'hb9825dbb),
	.w5(32'hba4fdf86),
	.w6(32'hb8ef8991),
	.w7(32'hb8b81a75),
	.w8(32'hb9fef957),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb727588),
	.w1(32'hbb3a8d67),
	.w2(32'hbb580683),
	.w3(32'hbb948614),
	.w4(32'hbb242b8f),
	.w5(32'hbb27b884),
	.w6(32'hbb47b3f5),
	.w7(32'hbaa67cdb),
	.w8(32'hbb4542aa),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3635b138),
	.w1(32'hb6a9163b),
	.w2(32'h3467ddc4),
	.w3(32'h365a9577),
	.w4(32'hb694bed4),
	.w5(32'h368bcbe5),
	.w6(32'h36b1c24f),
	.w7(32'hb626fe93),
	.w8(32'h3717ecbe),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3818efcf),
	.w1(32'h37930634),
	.w2(32'h37dcbfde),
	.w3(32'h37cfb5b4),
	.w4(32'h36fe8eee),
	.w5(32'hb79e1491),
	.w6(32'hb80c42a9),
	.w7(32'h35b7e1ad),
	.w8(32'hb5eb4517),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2063cf),
	.w1(32'hba625b53),
	.w2(32'hbb02b324),
	.w3(32'hba0e0f7e),
	.w4(32'hb7d2ca46),
	.w5(32'hbabf5e92),
	.w6(32'hb96e1b28),
	.w7(32'h3a595d03),
	.w8(32'hba87d4c9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5a59b),
	.w1(32'hba834654),
	.w2(32'hbb3cf608),
	.w3(32'h3abf42f1),
	.w4(32'h3a95c757),
	.w5(32'hba9bb570),
	.w6(32'h3a863715),
	.w7(32'h3ac4689b),
	.w8(32'hba40e557),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeeba0),
	.w1(32'hbaad33ef),
	.w2(32'hbb432896),
	.w3(32'hb9d9b8cb),
	.w4(32'h3956a506),
	.w5(32'hbae765e0),
	.w6(32'hba3136eb),
	.w7(32'h39cafdf0),
	.w8(32'hbacbb17b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c1df0),
	.w1(32'hb8965f4e),
	.w2(32'hb84b9471),
	.w3(32'h36f0128e),
	.w4(32'hb9c79fd9),
	.w5(32'hba1f2990),
	.w6(32'h3ad9463d),
	.w7(32'h3a0b83ed),
	.w8(32'hba10d126),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba27e3),
	.w1(32'hb899ee52),
	.w2(32'h38298be8),
	.w3(32'hb782eaa1),
	.w4(32'h36bd555a),
	.w5(32'hb7c1afb5),
	.w6(32'hb7e1379a),
	.w7(32'hb852822c),
	.w8(32'h389c833b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d76fd3),
	.w1(32'hb99d5024),
	.w2(32'hb9099664),
	.w3(32'hb97c5408),
	.w4(32'hb93232eb),
	.w5(32'hb867d782),
	.w6(32'hb8a37a78),
	.w7(32'hb89a2c50),
	.w8(32'hb8edfa57),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9081ffa),
	.w1(32'h3aa3c965),
	.w2(32'hba36b6a5),
	.w3(32'h3aaf4883),
	.w4(32'h39f6aef9),
	.w5(32'hbb13f83f),
	.w6(32'h3ab9511e),
	.w7(32'h3b07c17e),
	.w8(32'hbb09c4f4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a980f),
	.w1(32'hbb54e3ba),
	.w2(32'hbb844eac),
	.w3(32'hbb4c8c3d),
	.w4(32'hbb36400a),
	.w5(32'hbb3dec28),
	.w6(32'hbb37bcd6),
	.w7(32'hbb0d9b5b),
	.w8(32'hbb01cdd5),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38037ae9),
	.w1(32'hb9d6c1e7),
	.w2(32'hbaf5844e),
	.w3(32'h3a2d75dd),
	.w4(32'h381bc862),
	.w5(32'hbae128ca),
	.w6(32'h3aa3b63b),
	.w7(32'h3a12dfae),
	.w8(32'hbac8d52e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956532c),
	.w1(32'h3b0532e3),
	.w2(32'h3aa393c0),
	.w3(32'hba24dcb5),
	.w4(32'h3ae00266),
	.w5(32'h39feb057),
	.w6(32'hb9953476),
	.w7(32'h3afbb5ca),
	.w8(32'h3a25aa8e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dbfdc),
	.w1(32'hbabc39ac),
	.w2(32'hbb0699e7),
	.w3(32'hbae133bc),
	.w4(32'h39226c65),
	.w5(32'hba632b30),
	.w6(32'hba7c01ec),
	.w7(32'h3a953bd9),
	.w8(32'h39cc153b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373de0b8),
	.w1(32'h36db8467),
	.w2(32'h370622dc),
	.w3(32'h36d72f3c),
	.w4(32'h35b97df3),
	.w5(32'h35359074),
	.w6(32'h366c1a92),
	.w7(32'h3558b087),
	.w8(32'h350142fd),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372ba052),
	.w1(32'h36a44469),
	.w2(32'h3742a25b),
	.w3(32'h364374c5),
	.w4(32'hb642130f),
	.w5(32'h36a44bb3),
	.w6(32'h368c08ad),
	.w7(32'h34890dbd),
	.w8(32'h37224ee8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7a9bc),
	.w1(32'h3933d5fb),
	.w2(32'h390a3d13),
	.w3(32'h39f5951a),
	.w4(32'hb8e9214c),
	.w5(32'hb989af17),
	.w6(32'h399d6ee3),
	.w7(32'h383d5c47),
	.w8(32'h394bc998),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c959d2),
	.w1(32'hb6bf717f),
	.w2(32'hb677260e),
	.w3(32'h37813895),
	.w4(32'hb75454b7),
	.w5(32'hb70e5713),
	.w6(32'h375548a9),
	.w7(32'hb731aca4),
	.w8(32'hb6e1b97b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bf0e5a),
	.w1(32'hb99d1147),
	.w2(32'hb9df4dae),
	.w3(32'h393f2ce7),
	.w4(32'hb9d316f0),
	.w5(32'hba334bac),
	.w6(32'h3a0ca8b6),
	.w7(32'hb8fa55f4),
	.w8(32'hb9eea6f1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf6878),
	.w1(32'hba8b92b7),
	.w2(32'hbb0c9e38),
	.w3(32'h3a88b06b),
	.w4(32'h39ed9d58),
	.w5(32'hba99105b),
	.w6(32'h3a11fdbf),
	.w7(32'h3a6352ac),
	.w8(32'hba01784b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6546f2),
	.w1(32'hba963eb0),
	.w2(32'hbb015513),
	.w3(32'hb9bbd491),
	.w4(32'hb98be5a7),
	.w5(32'hba654537),
	.w6(32'h3a0b0fa7),
	.w7(32'h3a1f3985),
	.w8(32'hba13d22c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3777996f),
	.w1(32'h3780c807),
	.w2(32'h3740e88a),
	.w3(32'h3759ed75),
	.w4(32'h374568eb),
	.w5(32'h36de8503),
	.w6(32'h370d4b0d),
	.w7(32'h375cb34b),
	.w8(32'h373583c6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac289e1),
	.w1(32'hb99b5c6f),
	.w2(32'hbb2bd00c),
	.w3(32'hb9c58df1),
	.w4(32'hb97e5ba8),
	.w5(32'hbafa8fe2),
	.w6(32'h3a451039),
	.w7(32'hb64151f6),
	.w8(32'hbb394e87),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9611877),
	.w1(32'hb962e52e),
	.w2(32'hba4ff81d),
	.w3(32'h3a01acba),
	.w4(32'h35925483),
	.w5(32'hba2ab4a4),
	.w6(32'h39b1df6e),
	.w7(32'hb9261f52),
	.w8(32'hba391ff1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb804c203),
	.w1(32'hb861270b),
	.w2(32'hb7c085a4),
	.w3(32'h374dc70e),
	.w4(32'hb82c56ab),
	.w5(32'h37fb6dbd),
	.w6(32'hb6f82e18),
	.w7(32'hb5ed6938),
	.w8(32'h3876805a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9850677),
	.w1(32'hb909c944),
	.w2(32'hba43bade),
	.w3(32'h39a01b29),
	.w4(32'hb6f2bc3f),
	.w5(32'hba4ad01e),
	.w6(32'h3a093885),
	.w7(32'h39489039),
	.w8(32'hb9f97c49),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d8afcf),
	.w1(32'hb75ea211),
	.w2(32'h377a997b),
	.w3(32'h37177a36),
	.w4(32'h3766135c),
	.w5(32'h36122d43),
	.w6(32'h35d9fc7c),
	.w7(32'h370b8d6b),
	.w8(32'hb6591174),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aea68e),
	.w1(32'h393fb946),
	.w2(32'h386f6c3b),
	.w3(32'h388a1839),
	.w4(32'h38710d38),
	.w5(32'hb82f9392),
	.w6(32'h3832217a),
	.w7(32'h375e0d96),
	.w8(32'hb80d64dd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e66972),
	.w1(32'hb507a42b),
	.w2(32'h36c575b8),
	.w3(32'h37504f44),
	.w4(32'h3759859f),
	.w5(32'h378dcd6d),
	.w6(32'h37e263b0),
	.w7(32'h370f3147),
	.w8(32'h37a5a25a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3772592e),
	.w1(32'h36914c43),
	.w2(32'h37460ee2),
	.w3(32'h36fd41fe),
	.w4(32'h3614f1cd),
	.w5(32'h368c7fd7),
	.w6(32'h369b4155),
	.w7(32'h363785ba),
	.w8(32'h368455e9),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c62a96),
	.w1(32'h39ab266a),
	.w2(32'hb812af70),
	.w3(32'hba38a5d2),
	.w4(32'h3967a6d8),
	.w5(32'hb9e994e4),
	.w6(32'hba24ffa2),
	.w7(32'h39b5bcf1),
	.w8(32'hb9b3c581),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabea3f),
	.w1(32'hbb1935a6),
	.w2(32'hbb880601),
	.w3(32'h3702e16b),
	.w4(32'hba1139b2),
	.w5(32'hbb3629bd),
	.w6(32'h3a1de3f0),
	.w7(32'hba20e400),
	.w8(32'hbae9e4f2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f8e6b),
	.w1(32'hba2eb53e),
	.w2(32'hbaf6c836),
	.w3(32'h3955420f),
	.w4(32'h3992d005),
	.w5(32'hba99859c),
	.w6(32'h3a8ad071),
	.w7(32'h3a1a054d),
	.w8(32'hba1e65fe),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae42f7f),
	.w1(32'hbb1552b3),
	.w2(32'hbb73cf66),
	.w3(32'hba4472ac),
	.w4(32'hba86a15b),
	.w5(32'hbb287d63),
	.w6(32'hb9aca7a6),
	.w7(32'hbaab75d4),
	.w8(32'hbb017812),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e72673),
	.w1(32'h386d32ef),
	.w2(32'h384d61f7),
	.w3(32'h3757632d),
	.w4(32'h38629224),
	.w5(32'h386c687f),
	.w6(32'hb74a9075),
	.w7(32'h37a7a3cd),
	.w8(32'h380cd484),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9422f36),
	.w1(32'hb9497df6),
	.w2(32'hb8c8b5d2),
	.w3(32'hb886a7f0),
	.w4(32'hb913e9c1),
	.w5(32'h372ca233),
	.w6(32'hb7ce9bae),
	.w7(32'hb8611047),
	.w8(32'h374f6826),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367f9e3d),
	.w1(32'h34529a91),
	.w2(32'h36c30f47),
	.w3(32'h36947232),
	.w4(32'h35f811d0),
	.w5(32'h35e7e68d),
	.w6(32'h3565b415),
	.w7(32'hb6b24560),
	.w8(32'hb4fb0ee6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374cdd84),
	.w1(32'h374d829f),
	.w2(32'h37cec46a),
	.w3(32'h363b28f7),
	.w4(32'hb6ed2867),
	.w5(32'h361208c9),
	.w6(32'h370ff950),
	.w7(32'hb68e73fd),
	.w8(32'hb6d8425a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4d305),
	.w1(32'hbab0cd28),
	.w2(32'hbb2f8f47),
	.w3(32'hb94c893c),
	.w4(32'hb98c523f),
	.w5(32'hba8e459a),
	.w6(32'h3937a8d0),
	.w7(32'hb9705ae0),
	.w8(32'hba84abe4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b2cca4),
	.w1(32'h37b31e31),
	.w2(32'h3822e5bd),
	.w3(32'h37917839),
	.w4(32'h38185826),
	.w5(32'h383d74eb),
	.w6(32'hb6a850be),
	.w7(32'h36b83165),
	.w8(32'h375bacfc),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c712f6),
	.w1(32'h38822447),
	.w2(32'h39ab423a),
	.w3(32'hba31696e),
	.w4(32'hb9af7dba),
	.w5(32'hb7b1a3d0),
	.w6(32'hba24ebb9),
	.w7(32'hb9775486),
	.w8(32'hb628d709),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47df93),
	.w1(32'hb9a5e068),
	.w2(32'h37be17bd),
	.w3(32'hba6d392c),
	.w4(32'hb95c673a),
	.w5(32'h38f44eae),
	.w6(32'hba307e44),
	.w7(32'hb94b0f9a),
	.w8(32'h388013e8),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c7102c),
	.w1(32'h3577a1ae),
	.w2(32'h37ab69e0),
	.w3(32'hb7489b00),
	.w4(32'h36848684),
	.w5(32'h37aa5fa6),
	.w6(32'hb794f243),
	.w7(32'hb6997686),
	.w8(32'h373b1246),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d9996),
	.w1(32'hba3341f9),
	.w2(32'hba586538),
	.w3(32'hba12fd5f),
	.w4(32'hba064114),
	.w5(32'hba39b77b),
	.w6(32'hb99a158b),
	.w7(32'hba037659),
	.w8(32'hba53ff52),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ebfda9),
	.w1(32'hb930e25a),
	.w2(32'hb8538fee),
	.w3(32'hb8e5c905),
	.w4(32'hb91175e9),
	.w5(32'hb80acea4),
	.w6(32'hb86868e9),
	.w7(32'hb92440b2),
	.w8(32'hb8a06aa8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ed913),
	.w1(32'hbb3241ef),
	.w2(32'hbb97fc6c),
	.w3(32'hbaccf45c),
	.w4(32'hba7c6ceb),
	.w5(32'hbb0df81a),
	.w6(32'hba6985ce),
	.w7(32'hb9bedcc7),
	.w8(32'hb9a3f38e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb700c836),
	.w1(32'hb7f819ed),
	.w2(32'hb6c78e90),
	.w3(32'h3807d138),
	.w4(32'hb7a50f4e),
	.w5(32'h3781ca51),
	.w6(32'h379d9ac0),
	.w7(32'hb79f7a5b),
	.w8(32'h371386bb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16f023),
	.w1(32'h3ac82b23),
	.w2(32'h3ab9376c),
	.w3(32'h3a0e339b),
	.w4(32'h3afddf60),
	.w5(32'h3adbd7ea),
	.w6(32'h393a20f8),
	.w7(32'h3b097e87),
	.w8(32'h3a9271d2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule