module layer_10_featuremap_357(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cd9f0),
	.w1(32'h3952abae),
	.w2(32'hba679208),
	.w3(32'hba6cc728),
	.w4(32'hb99d6d3f),
	.w5(32'hb9d890d7),
	.w6(32'h39ab0206),
	.w7(32'hba570a40),
	.w8(32'hb9cff844),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3bafc),
	.w1(32'hbaec0e97),
	.w2(32'hbb2537cc),
	.w3(32'hbb1d2dba),
	.w4(32'hbafc6c21),
	.w5(32'hbaeefd1d),
	.w6(32'hba4f72c7),
	.w7(32'hbaaafd61),
	.w8(32'hbb986752),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb246365),
	.w1(32'hbaf970f3),
	.w2(32'h3903f957),
	.w3(32'hbb1fa48f),
	.w4(32'hba6e0579),
	.w5(32'h3a9e5bf0),
	.w6(32'hbab8e298),
	.w7(32'hbaedbfd6),
	.w8(32'h3af1e137),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9cc36),
	.w1(32'h3b046931),
	.w2(32'h39f977b5),
	.w3(32'hb9d5f8d9),
	.w4(32'h38e6c4a7),
	.w5(32'hbaf9b59a),
	.w6(32'h3a76e43d),
	.w7(32'h3878ec7c),
	.w8(32'h3aad1e4c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1887ee),
	.w1(32'h3ab58981),
	.w2(32'h39a3cdb2),
	.w3(32'hbaafc0a7),
	.w4(32'hbaa824a8),
	.w5(32'h3a0499a8),
	.w6(32'h3a7f4677),
	.w7(32'h3ac6210f),
	.w8(32'h39e5c635),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb960ba81),
	.w1(32'hb97b626d),
	.w2(32'hba2fbc31),
	.w3(32'h391a72db),
	.w4(32'h3aa35f8c),
	.w5(32'h3796c2ee),
	.w6(32'h37faa9a7),
	.w7(32'h384c0bf2),
	.w8(32'hb8e9cafb),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c9ba5),
	.w1(32'h3a6a17d4),
	.w2(32'hb9d2b106),
	.w3(32'h3bb81b9f),
	.w4(32'h3b5e29c0),
	.w5(32'hbaf7533f),
	.w6(32'h3bb17504),
	.w7(32'h3b4faa88),
	.w8(32'hbb5966fb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17858d),
	.w1(32'hbb48d136),
	.w2(32'hba973bec),
	.w3(32'hbb1c4e51),
	.w4(32'hbb10c8bc),
	.w5(32'h390a15b4),
	.w6(32'h3993b1a0),
	.w7(32'hbba5bb48),
	.w8(32'hb833e4fc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8694e8),
	.w1(32'hb9adfedf),
	.w2(32'h394208dc),
	.w3(32'hb7e30acf),
	.w4(32'h3a8c648a),
	.w5(32'h39c4b444),
	.w6(32'hbabbcc4e),
	.w7(32'hb9b089c5),
	.w8(32'h3a954975),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac233ce),
	.w1(32'hbae7c1dc),
	.w2(32'hbade2e64),
	.w3(32'h3b6825be),
	.w4(32'h39b53921),
	.w5(32'hba68fce0),
	.w6(32'h3bc512a4),
	.w7(32'h39b4cc70),
	.w8(32'hbab8f523),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc9fcd),
	.w1(32'h371914e6),
	.w2(32'hb81bb419),
	.w3(32'h38f2d9e5),
	.w4(32'h3af0809c),
	.w5(32'h3ac56d31),
	.w6(32'h3a2f9237),
	.w7(32'h3a2a8654),
	.w8(32'hba819d06),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57f500),
	.w1(32'h39d0c497),
	.w2(32'h3adf6cb4),
	.w3(32'h3b7d1550),
	.w4(32'h3ba690e5),
	.w5(32'hbacb3839),
	.w6(32'h3bba265c),
	.w7(32'h3bb09dce),
	.w8(32'hbaca4596),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ab1d5),
	.w1(32'hbb2367c3),
	.w2(32'hba844f9b),
	.w3(32'h3b789413),
	.w4(32'hba889794),
	.w5(32'hbae29299),
	.w6(32'h3bc70428),
	.w7(32'h396fe606),
	.w8(32'hbb041672),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4940d0),
	.w1(32'hbacc43af),
	.w2(32'hba18ead3),
	.w3(32'h3ae26fc3),
	.w4(32'hbadabc91),
	.w5(32'hba55611c),
	.w6(32'h3ae8b233),
	.w7(32'hb9dcf7d6),
	.w8(32'h3a91b7fa),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77d3e6),
	.w1(32'h385d51eb),
	.w2(32'hba84664d),
	.w3(32'h3af5f92d),
	.w4(32'h3ab7e348),
	.w5(32'hba60bb69),
	.w6(32'h3b1b6a45),
	.w7(32'hb91f33c3),
	.w8(32'hbaf7b202),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25c66e),
	.w1(32'hbadc6625),
	.w2(32'hbb20feb8),
	.w3(32'hb994ece9),
	.w4(32'hbb680548),
	.w5(32'hbbab417c),
	.w6(32'h3b7dc5f7),
	.w7(32'hbaf9ef59),
	.w8(32'hbb6bb5a8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23cc27),
	.w1(32'h39781d4b),
	.w2(32'hb96afce0),
	.w3(32'hb996f30c),
	.w4(32'h3a3bac9c),
	.w5(32'hba8acd54),
	.w6(32'h381bbb52),
	.w7(32'h3a43dcfe),
	.w8(32'hbac85038),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391cc58e),
	.w1(32'hbb3a1512),
	.w2(32'hbaeff8a8),
	.w3(32'h3b8d2104),
	.w4(32'hb941c36d),
	.w5(32'hba9d8b40),
	.w6(32'h3ad301da),
	.w7(32'hbacc07de),
	.w8(32'hb98ddf73),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3eeda4),
	.w1(32'h39465663),
	.w2(32'h39ff601b),
	.w3(32'h3b32c10a),
	.w4(32'h3a7f9850),
	.w5(32'h39873a83),
	.w6(32'h3b7344f4),
	.w7(32'h3a8c2210),
	.w8(32'hba87add5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b203d1),
	.w1(32'h3a6437fa),
	.w2(32'h3a9aca1d),
	.w3(32'h3a85dfc3),
	.w4(32'h3a28cc65),
	.w5(32'h3985b31e),
	.w6(32'h3afb9b34),
	.w7(32'h3a923474),
	.w8(32'hb94ee5a3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90238f0),
	.w1(32'h3b16893b),
	.w2(32'h3a52db51),
	.w3(32'h3a86f2ef),
	.w4(32'hb9995de7),
	.w5(32'h3aee2d01),
	.w6(32'h3ad6705c),
	.w7(32'h3a60bca5),
	.w8(32'h3b2f75bb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecf7ed),
	.w1(32'h3b52d249),
	.w2(32'h3b261ffd),
	.w3(32'hba7b57e0),
	.w4(32'h39db1bb1),
	.w5(32'h3ad21410),
	.w6(32'h39041b04),
	.w7(32'h3b05e81b),
	.w8(32'h3a0cdc99),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad2038),
	.w1(32'hbb926780),
	.w2(32'hbb9b15bc),
	.w3(32'h3bc96c29),
	.w4(32'hba5597d5),
	.w5(32'hbbc073dc),
	.w6(32'h3b6097a5),
	.w7(32'h3a73cbfe),
	.w8(32'hbb8f7784),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941bb61),
	.w1(32'hbb10dd16),
	.w2(32'hbb3c7f65),
	.w3(32'hbae7d60f),
	.w4(32'hbadf8262),
	.w5(32'hbb48ff6f),
	.w6(32'h3b24edab),
	.w7(32'hba08101e),
	.w8(32'hbb88bbb9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb791543),
	.w1(32'hbb989a6b),
	.w2(32'hbb81521d),
	.w3(32'hbbaaa656),
	.w4(32'hbb74f131),
	.w5(32'hbb707aea),
	.w6(32'hb9a80034),
	.w7(32'hbab8ff70),
	.w8(32'hbb2545fe),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cb987),
	.w1(32'h3aa1305a),
	.w2(32'hba59ceb2),
	.w3(32'h3aeeebf0),
	.w4(32'h39eb367d),
	.w5(32'hbaffb674),
	.w6(32'h3b6cd4a1),
	.w7(32'h3a232e61),
	.w8(32'hba49a67f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a2013),
	.w1(32'h3a0c4a82),
	.w2(32'h3ad56c2d),
	.w3(32'hba963487),
	.w4(32'hba0f0d14),
	.w5(32'hba1ce8a3),
	.w6(32'hb93a8e3e),
	.w7(32'h3a53cc94),
	.w8(32'h399cf067),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ceb53),
	.w1(32'h3ab6f64b),
	.w2(32'h3aa30f7b),
	.w3(32'hbb307a56),
	.w4(32'hbaf9107c),
	.w5(32'hbaf1dae5),
	.w6(32'h3a0a21a4),
	.w7(32'h3a7b0323),
	.w8(32'h3b8a845b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acaf941),
	.w1(32'h3b0f4aac),
	.w2(32'h3963c8e5),
	.w3(32'hb96644a6),
	.w4(32'h3a8dc147),
	.w5(32'h3a4b64f2),
	.w6(32'h398761c6),
	.w7(32'h36ebb438),
	.w8(32'h3ab6f007),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08fcaf),
	.w1(32'hbb98a169),
	.w2(32'hbb49fe94),
	.w3(32'hbaca70bd),
	.w4(32'hbba1a7f4),
	.w5(32'hbbdd4fe6),
	.w6(32'h3b4da4c3),
	.w7(32'hbb3680d4),
	.w8(32'hbb7b5634),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f4fd9),
	.w1(32'h3a15fb0d),
	.w2(32'h3a8b38ab),
	.w3(32'h3abef67c),
	.w4(32'h3aad7e0a),
	.w5(32'hb998ee4d),
	.w6(32'h3ac8fe65),
	.w7(32'h3a1e2c10),
	.w8(32'hbb80c43e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb190264),
	.w1(32'hbb4af4b5),
	.w2(32'hba4931d8),
	.w3(32'hbaef6aa7),
	.w4(32'h3839e551),
	.w5(32'hbb477493),
	.w6(32'hbafde276),
	.w7(32'hbb10a061),
	.w8(32'h39c2695c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6c7f8),
	.w1(32'hb960c457),
	.w2(32'hbae14883),
	.w3(32'h3b871ac1),
	.w4(32'hbab492d0),
	.w5(32'hbaf74356),
	.w6(32'h3b8f6b51),
	.w7(32'hbaba1231),
	.w8(32'hbb02542b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1499c2),
	.w1(32'hbbbd7639),
	.w2(32'hbb6e3da3),
	.w3(32'h3a24ab9b),
	.w4(32'hba72a1d2),
	.w5(32'h3a2cd265),
	.w6(32'hb8a8c2bf),
	.w7(32'hbaa06684),
	.w8(32'h39aa1619),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fedd3),
	.w1(32'h3a499877),
	.w2(32'h387b4e68),
	.w3(32'h3a34d84f),
	.w4(32'hbaaebd1e),
	.w5(32'h3a056864),
	.w6(32'h3b2754cf),
	.w7(32'h39149a71),
	.w8(32'h3a66fe23),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a426060),
	.w1(32'hbb4b07f4),
	.w2(32'hbad5b439),
	.w3(32'h3bc7d188),
	.w4(32'h3a3dd5fd),
	.w5(32'h3a4280f9),
	.w6(32'h395f5b60),
	.w7(32'h3a951f1d),
	.w8(32'hba2c7db3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8abbcbb),
	.w1(32'hbc0ddf7c),
	.w2(32'hbc03f85e),
	.w3(32'hba90521e),
	.w4(32'hbbe671ac),
	.w5(32'hbc166f17),
	.w6(32'h3b47c35c),
	.w7(32'h3b106371),
	.w8(32'hbc1c230c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399daaf9),
	.w1(32'h3b604683),
	.w2(32'h3aca70c4),
	.w3(32'h388625e8),
	.w4(32'h3b11eacb),
	.w5(32'hbb3eddbc),
	.w6(32'hb9806a78),
	.w7(32'h3b1c806f),
	.w8(32'hbb2b37cf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fcad0),
	.w1(32'hb899e146),
	.w2(32'hba853e6d),
	.w3(32'hbb62d588),
	.w4(32'hb8a7def2),
	.w5(32'h3a512ce4),
	.w6(32'hbb1447c7),
	.w7(32'h39529b9a),
	.w8(32'h3b951504),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0651b),
	.w1(32'hba665bc4),
	.w2(32'hbb1964de),
	.w3(32'hbb5051d3),
	.w4(32'hbb9052ca),
	.w5(32'h3936c9f1),
	.w6(32'h3a046507),
	.w7(32'hbb3bcaab),
	.w8(32'h394c2027),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34ce68),
	.w1(32'h397f46ff),
	.w2(32'h3aa2e599),
	.w3(32'h37dfd499),
	.w4(32'h3a821ba7),
	.w5(32'hb9a00db6),
	.w6(32'hba0651f2),
	.w7(32'hb9285bc5),
	.w8(32'h3a0a205e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98772c0),
	.w1(32'h3aa2e54a),
	.w2(32'hb93a20a2),
	.w3(32'hba365bc7),
	.w4(32'h3a1155a7),
	.w5(32'h3aff521e),
	.w6(32'h3a6690f4),
	.w7(32'hb8ae64b1),
	.w8(32'h3a2872f0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61b96e),
	.w1(32'h3b0a610c),
	.w2(32'h3a2fa133),
	.w3(32'h3b8c45a2),
	.w4(32'h3b73feaa),
	.w5(32'h3a48f8ae),
	.w6(32'h3b214a72),
	.w7(32'h3b0f1c1e),
	.w8(32'hbaa0446b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35bff0),
	.w1(32'h39a0851b),
	.w2(32'h3a107ccc),
	.w3(32'h3b166741),
	.w4(32'h3ab95b0c),
	.w5(32'hba742809),
	.w6(32'h3b16d3b7),
	.w7(32'hbb4dc29e),
	.w8(32'h39188761),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0849ba),
	.w1(32'hba1f5374),
	.w2(32'hbb39e7f1),
	.w3(32'h3b1e3341),
	.w4(32'hba9fa321),
	.w5(32'hbb9461b0),
	.w6(32'h3b88dac0),
	.w7(32'h3a3b974f),
	.w8(32'hbb67ada6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b53864),
	.w1(32'hbb34e06f),
	.w2(32'hbb984d7b),
	.w3(32'h3a9953e8),
	.w4(32'hbacc6f1a),
	.w5(32'hbb43660e),
	.w6(32'h3b2c784f),
	.w7(32'hbaab6d30),
	.w8(32'hbb836a13),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad77f9),
	.w1(32'hb9ff79a7),
	.w2(32'hba341682),
	.w3(32'hba3366f3),
	.w4(32'hbab884f6),
	.w5(32'hbab6be40),
	.w6(32'h3ab46594),
	.w7(32'hb9ae8dc9),
	.w8(32'hb94e818f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd4885),
	.w1(32'h3b9fd390),
	.w2(32'h3b28ddd7),
	.w3(32'h3bbf747f),
	.w4(32'h3b230f53),
	.w5(32'hbb0fe82c),
	.w6(32'h3bfae0e3),
	.w7(32'h3b19e8ed),
	.w8(32'hbb486049),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53f26b),
	.w1(32'hbb173e27),
	.w2(32'hb9c43116),
	.w3(32'hba9651a3),
	.w4(32'h376461d6),
	.w5(32'h3ac98e2d),
	.w6(32'h394a0e3a),
	.w7(32'h3a4305a7),
	.w8(32'h3b385f89),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b081607),
	.w1(32'h3b272bd2),
	.w2(32'h3b0a6c16),
	.w3(32'hb9b43b4e),
	.w4(32'hba258ea1),
	.w5(32'hbb3de1d2),
	.w6(32'h3a32792d),
	.w7(32'h3a45efc3),
	.w8(32'hbabe79dd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1db876),
	.w1(32'hba9b2b33),
	.w2(32'h39854fbb),
	.w3(32'hbb56d875),
	.w4(32'hba7b47fe),
	.w5(32'h3a7af947),
	.w6(32'hba644de2),
	.w7(32'h3a832dab),
	.w8(32'h3a840e70),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea9e43),
	.w1(32'hba129a0f),
	.w2(32'hba422f27),
	.w3(32'h3af9a18e),
	.w4(32'h3977a403),
	.w5(32'hba00544f),
	.w6(32'h3b074de7),
	.w7(32'h3a9e75e3),
	.w8(32'hba9f3fa1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d230db),
	.w1(32'hba57aac8),
	.w2(32'hba13c793),
	.w3(32'hb95cf154),
	.w4(32'h3a5b57d6),
	.w5(32'hbae3d428),
	.w6(32'h39ce3eec),
	.w7(32'h3748a84f),
	.w8(32'hb96f0241),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04840a),
	.w1(32'h3ac37be4),
	.w2(32'hbafd44c5),
	.w3(32'h3b5b1077),
	.w4(32'h3b2eb79e),
	.w5(32'hba0ff924),
	.w6(32'h3bfcb02d),
	.w7(32'h3b07802c),
	.w8(32'hba464761),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9471c32),
	.w1(32'h39becf63),
	.w2(32'h390012aa),
	.w3(32'h3ab5fe89),
	.w4(32'h3adfeca9),
	.w5(32'h39e2fdc4),
	.w6(32'h3ae89736),
	.w7(32'h3a7dfa8e),
	.w8(32'h3a16b700),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962b7b9),
	.w1(32'hba326114),
	.w2(32'hba54c336),
	.w3(32'hbadc5aed),
	.w4(32'hbad19406),
	.w5(32'h3a96e421),
	.w6(32'h3a0e0a9c),
	.w7(32'hba70f27f),
	.w8(32'h3a940b31),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a751ab4),
	.w1(32'h399fe5f4),
	.w2(32'h3a6f7583),
	.w3(32'h3a01ee6a),
	.w4(32'h3a45a064),
	.w5(32'h3a013f2b),
	.w6(32'h39c5c302),
	.w7(32'h3a4ba2eb),
	.w8(32'h394dfc93),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72563f),
	.w1(32'h3adee23d),
	.w2(32'h3aef3d2f),
	.w3(32'h3aabd675),
	.w4(32'h3aa08c07),
	.w5(32'h3a21e0f4),
	.w6(32'h3b329900),
	.w7(32'h39e8bfcf),
	.w8(32'h3ad78e98),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17d48f),
	.w1(32'h3b32e65f),
	.w2(32'h3acbe411),
	.w3(32'h39d2e9d2),
	.w4(32'h3a8c8db0),
	.w5(32'h3992492c),
	.w6(32'h3aa656d7),
	.w7(32'h3ac060f5),
	.w8(32'hbb0bc2ab),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f026ad),
	.w1(32'h39d2f48d),
	.w2(32'h3a9029be),
	.w3(32'hba18dc85),
	.w4(32'h3b1e3761),
	.w5(32'hb9ee7ddb),
	.w6(32'hbb0573ea),
	.w7(32'h3b1f9dc7),
	.w8(32'h380a9649),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c445f),
	.w1(32'h3a4ad3f1),
	.w2(32'h39e245c5),
	.w3(32'h3aef4e4d),
	.w4(32'hb9acccd9),
	.w5(32'hba9c3134),
	.w6(32'h3abf2a8b),
	.w7(32'h39073a9c),
	.w8(32'h3a8e1471),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fc629),
	.w1(32'h3b5bc9d4),
	.w2(32'hba826638),
	.w3(32'hba614e1b),
	.w4(32'h3a19556b),
	.w5(32'hbaa94f08),
	.w6(32'h3b3421e2),
	.w7(32'h3a9e9f68),
	.w8(32'h3acf159d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad67e92),
	.w1(32'h38fc7a47),
	.w2(32'hb9d7aee7),
	.w3(32'hbb08642a),
	.w4(32'hbaced5cf),
	.w5(32'h3a0124be),
	.w6(32'h3ace06ba),
	.w7(32'h3a3089b3),
	.w8(32'h3a036438),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9520c4a),
	.w1(32'h37feb1b1),
	.w2(32'h37bc3cc8),
	.w3(32'hba944e40),
	.w4(32'hba8a270e),
	.w5(32'h38458ab9),
	.w6(32'hb9a9d5fb),
	.w7(32'hba4266e0),
	.w8(32'h3a32b8d1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2d91a),
	.w1(32'h398b842f),
	.w2(32'hb9066b83),
	.w3(32'hba36e54d),
	.w4(32'hb981c8d0),
	.w5(32'h3ac7d130),
	.w6(32'h3ae91ed5),
	.w7(32'h3738676c),
	.w8(32'hb9c9fc27),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392350e6),
	.w1(32'hba8f87c3),
	.w2(32'h398c5dec),
	.w3(32'h3a579636),
	.w4(32'h3aa38a8b),
	.w5(32'h390dfaa2),
	.w6(32'h37ccfcb8),
	.w7(32'h3a1ebaac),
	.w8(32'hba3173a5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54e6d),
	.w1(32'h3b5cb716),
	.w2(32'h3b434156),
	.w3(32'hbb42f7a8),
	.w4(32'hbacc0a1d),
	.w5(32'hbb474567),
	.w6(32'h3c01da0a),
	.w7(32'h3ac7f29f),
	.w8(32'h3badeddc),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc16af),
	.w1(32'hba99ea78),
	.w2(32'hbb5f488b),
	.w3(32'h3b61ed51),
	.w4(32'h3aa2d43e),
	.w5(32'hba97d3e6),
	.w6(32'h3b05f56c),
	.w7(32'hb8b97ec9),
	.w8(32'hbbb2aec0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb228d4d),
	.w1(32'hbade9e4b),
	.w2(32'hbad21770),
	.w3(32'h3b0c081d),
	.w4(32'h3a9abc1a),
	.w5(32'hb98fb2dc),
	.w6(32'hba8c8d2a),
	.w7(32'hb9e5b6dd),
	.w8(32'hba68a598),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87096c),
	.w1(32'hbbd1199a),
	.w2(32'hbb8df9a8),
	.w3(32'hb8b7cacb),
	.w4(32'hba17268b),
	.w5(32'hbb62c953),
	.w6(32'hbba6dfc8),
	.w7(32'hbafb8b8a),
	.w8(32'hbb686eed),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af46edc),
	.w1(32'h3a045c4e),
	.w2(32'h3a364aa8),
	.w3(32'h3b54857b),
	.w4(32'h3a986b31),
	.w5(32'hbb0bb627),
	.w6(32'h3afac99d),
	.w7(32'h3ac21a8e),
	.w8(32'h397dbe94),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba992026),
	.w1(32'hba8d778c),
	.w2(32'hba949c0f),
	.w3(32'hba2dcc69),
	.w4(32'hbb19026f),
	.w5(32'h3a1b1fd9),
	.w6(32'hbb05c1b8),
	.w7(32'hbacfe07d),
	.w8(32'hbb26cba2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5c81a),
	.w1(32'h3a3db413),
	.w2(32'h39178643),
	.w3(32'h3b31bff8),
	.w4(32'h3a85832a),
	.w5(32'hb9fae23d),
	.w6(32'hbab397d0),
	.w7(32'hba71b648),
	.w8(32'hb98fc019),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92d7c1),
	.w1(32'hba72d647),
	.w2(32'hbb022e18),
	.w3(32'h3b3e7013),
	.w4(32'h3aefe5d2),
	.w5(32'h3af83e6f),
	.w6(32'h3accd3d0),
	.w7(32'hba3bf30c),
	.w8(32'h39a22eb8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a92e1),
	.w1(32'h39293e82),
	.w2(32'hba22e3db),
	.w3(32'hba7200d1),
	.w4(32'h39c969f2),
	.w5(32'hbac57cfd),
	.w6(32'h39a5547b),
	.w7(32'hb9f07095),
	.w8(32'hbb2aeecf),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a434),
	.w1(32'hbb90adbb),
	.w2(32'hbb2933e2),
	.w3(32'h3aac7c78),
	.w4(32'h3a8a8319),
	.w5(32'h39e9dd6f),
	.w6(32'h3b6b156b),
	.w7(32'h3aefd90c),
	.w8(32'h39cd2357),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa8b70),
	.w1(32'h3b1e6f31),
	.w2(32'h3ae24844),
	.w3(32'h3b8ebdce),
	.w4(32'h3b302eae),
	.w5(32'hbaa5e545),
	.w6(32'h3b480cfa),
	.w7(32'hba80fdd7),
	.w8(32'hb8bc8b93),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af23e50),
	.w1(32'hbb13ab23),
	.w2(32'hbae7bf8d),
	.w3(32'h399dd5e4),
	.w4(32'hbb2c3c7a),
	.w5(32'hbbca2420),
	.w6(32'h3ae87d52),
	.w7(32'hbad1ea5f),
	.w8(32'hbbb4b2a9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53948f),
	.w1(32'hbad47ff2),
	.w2(32'hbb265a8d),
	.w3(32'hbabb086e),
	.w4(32'hbb380fe8),
	.w5(32'hbb1e7745),
	.w6(32'h3ab5f239),
	.w7(32'hbad4bdf1),
	.w8(32'hbadfdb12),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48b021),
	.w1(32'h3a921fb3),
	.w2(32'h37ddf4e0),
	.w3(32'h3aa1b27d),
	.w4(32'h3aaf69f3),
	.w5(32'hbb91d7ca),
	.w6(32'h3b9d7da2),
	.w7(32'h3aeac92c),
	.w8(32'hbaa468e6),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5ebc1),
	.w1(32'hba803f64),
	.w2(32'hbb2ee5d3),
	.w3(32'hbb6d0b9a),
	.w4(32'hbb6433ac),
	.w5(32'hbb24b137),
	.w6(32'h3a72fae9),
	.w7(32'hbaac708b),
	.w8(32'hbb711b2a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad16d5b),
	.w1(32'hbb30b052),
	.w2(32'hbb0770ea),
	.w3(32'h3baab715),
	.w4(32'h3b43edc9),
	.w5(32'h3a00a8eb),
	.w6(32'h3b02be41),
	.w7(32'h3a917cf4),
	.w8(32'hba330857),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2adfc6),
	.w1(32'hb9e5369a),
	.w2(32'h3aa1cc54),
	.w3(32'hb8b1501b),
	.w4(32'h39cbe5f1),
	.w5(32'hbaa22bb7),
	.w6(32'hb923374b),
	.w7(32'hb9d87ba8),
	.w8(32'h3a9df38e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96bccb7),
	.w1(32'hba028739),
	.w2(32'hbac8666c),
	.w3(32'hbba51c74),
	.w4(32'hbb58e26c),
	.w5(32'h3a173926),
	.w6(32'h39f386d9),
	.w7(32'hb9fb81d2),
	.w8(32'h395f60d4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ab62a),
	.w1(32'hbac577d3),
	.w2(32'hb9efa803),
	.w3(32'hb9921312),
	.w4(32'hb873c9c9),
	.w5(32'hb904ad36),
	.w6(32'hb81ae1cb),
	.w7(32'hb9ea2304),
	.w8(32'hbb0b6472),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2820f5),
	.w1(32'h39c65abb),
	.w2(32'h39f71382),
	.w3(32'hbaa5286b),
	.w4(32'h3abcacaf),
	.w5(32'hba29577e),
	.w6(32'hb8aaacfc),
	.w7(32'h3a574c3b),
	.w8(32'h39d06ac9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801e16),
	.w1(32'hbb5c38eb),
	.w2(32'hba9ab249),
	.w3(32'hbb88c17a),
	.w4(32'hbb277bce),
	.w5(32'hbb97101b),
	.w6(32'hbac36b38),
	.w7(32'hbaaa004f),
	.w8(32'hbb361df0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a621d),
	.w1(32'h3ad713bc),
	.w2(32'h3af1ba5e),
	.w3(32'h390d4b9f),
	.w4(32'h39ee0993),
	.w5(32'h39f99646),
	.w6(32'h37db5c93),
	.w7(32'h3af90009),
	.w8(32'h3a5aa5f9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae53e71),
	.w1(32'hbac41d35),
	.w2(32'hbaa04720),
	.w3(32'hba4a1203),
	.w4(32'hb9a3be15),
	.w5(32'hba620fff),
	.w6(32'hb9d9053a),
	.w7(32'hbaf1728a),
	.w8(32'hba5ec6e1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c6082),
	.w1(32'h3aae6a94),
	.w2(32'h3a84d371),
	.w3(32'h3baae750),
	.w4(32'h3b63c35d),
	.w5(32'h3a63eddf),
	.w6(32'h3bcd8ec5),
	.w7(32'h3b8d6182),
	.w8(32'h3a96d6b8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a9059),
	.w1(32'h39ea6ff0),
	.w2(32'hba9ca5f9),
	.w3(32'hbb5cdf5c),
	.w4(32'hba7d432b),
	.w5(32'hbae3ce7c),
	.w6(32'h3a445466),
	.w7(32'h3720ef73),
	.w8(32'h3adfda37),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc29853),
	.w1(32'h3b07ca1e),
	.w2(32'hbad4a0c3),
	.w3(32'h3bad7d8c),
	.w4(32'hbaf66652),
	.w5(32'hbbe5cc24),
	.w6(32'h3c00316c),
	.w7(32'h3b100a47),
	.w8(32'hba13ddad),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13d7c2),
	.w1(32'hba20f7a7),
	.w2(32'h3923ddad),
	.w3(32'hbae073ed),
	.w4(32'hba62d8e1),
	.w5(32'hba4950f2),
	.w6(32'hbace99e3),
	.w7(32'hbaedcc6a),
	.w8(32'h3a0018e0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8711ed),
	.w1(32'h3974a011),
	.w2(32'hbab0cafd),
	.w3(32'hb8e6745e),
	.w4(32'hbbbed1ee),
	.w5(32'hbc030247),
	.w6(32'h3ac09f80),
	.w7(32'hbb6a87fe),
	.w8(32'hbb6f1b1e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393cda55),
	.w1(32'hb99e8078),
	.w2(32'hbab92db0),
	.w3(32'hba36fd6f),
	.w4(32'hbb430443),
	.w5(32'hbb2b9112),
	.w6(32'h3b0d6534),
	.w7(32'hbaa6c441),
	.w8(32'hbb832b8a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21f75e),
	.w1(32'hbb217d02),
	.w2(32'hba8305d3),
	.w3(32'hbb032515),
	.w4(32'hbb74de78),
	.w5(32'hbbad8edf),
	.w6(32'hbafc512b),
	.w7(32'hbb1a0559),
	.w8(32'hbb3b73d0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43e1ab),
	.w1(32'hba877997),
	.w2(32'hbb2f1f5e),
	.w3(32'hbb5675ae),
	.w4(32'hbb339fe1),
	.w5(32'hbb0dd1e8),
	.w6(32'h3a8638dd),
	.w7(32'hbb0e1ff8),
	.w8(32'h3aa5894e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac43603),
	.w1(32'hba017830),
	.w2(32'hb8eb9968),
	.w3(32'h3baa9c95),
	.w4(32'h38a60e58),
	.w5(32'hbb4387bb),
	.w6(32'h3baafdb8),
	.w7(32'hba6f1b98),
	.w8(32'hbb9088ff),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4f2ae),
	.w1(32'hb8c6db2c),
	.w2(32'h3781baa6),
	.w3(32'hbb3e3449),
	.w4(32'hbb36dc63),
	.w5(32'hbb06ef31),
	.w6(32'h3b88a0b9),
	.w7(32'hbad77aa2),
	.w8(32'h3a449950),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b215396),
	.w1(32'hbae00d2a),
	.w2(32'hbb16d8d9),
	.w3(32'h3b2d5b99),
	.w4(32'hba9bcefe),
	.w5(32'hbbdef5c1),
	.w6(32'hb6f0dbc4),
	.w7(32'h3b358064),
	.w8(32'hbbfb655a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b7dd9),
	.w1(32'hba24bb6d),
	.w2(32'hb9d71624),
	.w3(32'hbae8299b),
	.w4(32'h3b453a51),
	.w5(32'h3b020a4d),
	.w6(32'hbb4763f9),
	.w7(32'h3a15e1f7),
	.w8(32'h3bae955d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8cf11),
	.w1(32'h3b9c91f8),
	.w2(32'h3b7656f6),
	.w3(32'h3b6c34e1),
	.w4(32'h39ac4aa1),
	.w5(32'hbb9fc05e),
	.w6(32'h3c3b0092),
	.w7(32'h3bdb58b1),
	.w8(32'hbbd53ec4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c667e6),
	.w1(32'hbb7c963a),
	.w2(32'hbb66212c),
	.w3(32'h3a8381de),
	.w4(32'hbb4ffdeb),
	.w5(32'hbbcc99e8),
	.w6(32'h3ba47b7b),
	.w7(32'h3a533610),
	.w8(32'hbb7e6730),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba76411b),
	.w1(32'hb9dbf512),
	.w2(32'h3978d5d9),
	.w3(32'hbadc932e),
	.w4(32'hbab2cd42),
	.w5(32'hb9d8e1dc),
	.w6(32'h38a5227f),
	.w7(32'hb92113e0),
	.w8(32'hb9931c2d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3df195),
	.w1(32'hbb742258),
	.w2(32'hbb73c1a9),
	.w3(32'hbb47f885),
	.w4(32'hbbbeb79e),
	.w5(32'hbba50f69),
	.w6(32'h3b5859bd),
	.w7(32'hbaff5047),
	.w8(32'hbbac3589),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab77d16),
	.w1(32'h3af242ef),
	.w2(32'hba4f677b),
	.w3(32'h3af8f21f),
	.w4(32'h3ac2da5e),
	.w5(32'hba93e3d1),
	.w6(32'h3b4c34f9),
	.w7(32'h3b0f4519),
	.w8(32'hb9b122d9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99504de),
	.w1(32'h3a6baccd),
	.w2(32'h3a74af54),
	.w3(32'h3a117241),
	.w4(32'hb98100a9),
	.w5(32'hb9ac572f),
	.w6(32'hba64f98f),
	.w7(32'h38d3a8a2),
	.w8(32'hb9a285d0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc3469),
	.w1(32'hba1bd4c5),
	.w2(32'hba795ba0),
	.w3(32'hb9d7bd90),
	.w4(32'hb8e9e0ba),
	.w5(32'hba8b2ee6),
	.w6(32'hba596642),
	.w7(32'hba22aa38),
	.w8(32'hbb3012bc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0f5ab),
	.w1(32'hba844e97),
	.w2(32'hbae9ff6b),
	.w3(32'h3b7a215a),
	.w4(32'hb9cd5812),
	.w5(32'hbb8e742e),
	.w6(32'h3b91a5f3),
	.w7(32'hbab39508),
	.w8(32'hbbadb7d2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37afe0),
	.w1(32'hbb42ea74),
	.w2(32'hbb6a6a4b),
	.w3(32'h38869df6),
	.w4(32'hbb104325),
	.w5(32'hbb541f9e),
	.w6(32'h39c5d259),
	.w7(32'hbb154b8a),
	.w8(32'hbb5d45fb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39691c0a),
	.w1(32'hba875dde),
	.w2(32'hb8b667ca),
	.w3(32'hbadfafc9),
	.w4(32'hbad23d32),
	.w5(32'hb9d9572d),
	.w6(32'h39d6ef32),
	.w7(32'hba40ed2b),
	.w8(32'h3ac72862),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a858fc),
	.w1(32'hba045f04),
	.w2(32'hb9803b84),
	.w3(32'hba222304),
	.w4(32'hba4f39b2),
	.w5(32'hbb079d51),
	.w6(32'h3a4b3f1f),
	.w7(32'h3a18d02d),
	.w8(32'hbb223c4f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0971dc),
	.w1(32'hb954028b),
	.w2(32'hba949815),
	.w3(32'h3b3c6638),
	.w4(32'h3ae43f01),
	.w5(32'h3b21c5b1),
	.w6(32'hbb2a575d),
	.w7(32'hba943816),
	.w8(32'hb9c58611),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c53a52),
	.w1(32'hba1ecef5),
	.w2(32'h39a6f0a0),
	.w3(32'h3b22ef9e),
	.w4(32'h3a43eaa2),
	.w5(32'hbb108ed1),
	.w6(32'h3b5888f7),
	.w7(32'h3afa8805),
	.w8(32'hb9070549),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf9f8d),
	.w1(32'hba9ea680),
	.w2(32'hbb120bee),
	.w3(32'h3ac15dcc),
	.w4(32'hba54cc8f),
	.w5(32'hba0a8d5c),
	.w6(32'h3acdf32a),
	.w7(32'hbad9b4fe),
	.w8(32'h3a09e792),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b908c2c),
	.w1(32'h3b8dc776),
	.w2(32'h3ac88806),
	.w3(32'h3a88adb7),
	.w4(32'h3a184134),
	.w5(32'h3b13b82f),
	.w6(32'h3b38b967),
	.w7(32'h3b428062),
	.w8(32'h3ab2e9d7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f5cab),
	.w1(32'hba2f5898),
	.w2(32'hba11f1b6),
	.w3(32'h3b0080f1),
	.w4(32'h3aa6ec7d),
	.w5(32'h3a96f4bc),
	.w6(32'h3aca9120),
	.w7(32'h3a2118f6),
	.w8(32'h3b079a19),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9bf30),
	.w1(32'h3b468029),
	.w2(32'h3b4e7fcd),
	.w3(32'h3acfa905),
	.w4(32'h39f39be4),
	.w5(32'hbb0cef9a),
	.w6(32'h3b65f833),
	.w7(32'h3b4b43a4),
	.w8(32'hbb1cd1c7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0723dc),
	.w1(32'hbaa71a7a),
	.w2(32'hba1e5b4e),
	.w3(32'hbb00109f),
	.w4(32'hba9cc4d6),
	.w5(32'hbb65354a),
	.w6(32'hbaafa5bc),
	.w7(32'hba627b64),
	.w8(32'hbb849ec6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8ffbc),
	.w1(32'hbbac5a5e),
	.w2(32'hbb8c5b88),
	.w3(32'hbb1832b8),
	.w4(32'hbb236f47),
	.w5(32'hbb8355a3),
	.w6(32'hbb04c960),
	.w7(32'hbb601e66),
	.w8(32'hbb710bde),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa944c9),
	.w1(32'hb9b19407),
	.w2(32'h39fb414c),
	.w3(32'hbaea314c),
	.w4(32'hbae8ea68),
	.w5(32'hba676edf),
	.w6(32'hbacd34d5),
	.w7(32'hba42d59e),
	.w8(32'hba38797a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64c994),
	.w1(32'h3a46c58d),
	.w2(32'hba0d937d),
	.w3(32'h3ab41300),
	.w4(32'h38e3a8b3),
	.w5(32'h3985d3f8),
	.w6(32'h3b13f62e),
	.w7(32'hb97e9f03),
	.w8(32'h3a19a649),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb908364a),
	.w1(32'hb9bef1f0),
	.w2(32'hba52f69c),
	.w3(32'hbaec8ff5),
	.w4(32'hbb37cca9),
	.w5(32'hbb743c27),
	.w6(32'hba4f30c8),
	.w7(32'hba30c7ea),
	.w8(32'hbb49c1c9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bbfb08),
	.w1(32'hb9d9679c),
	.w2(32'hba20935a),
	.w3(32'hba7b41f8),
	.w4(32'hba29afcc),
	.w5(32'hb9dec41d),
	.w6(32'hba617934),
	.w7(32'hba5d86aa),
	.w8(32'hba131870),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f65d8),
	.w1(32'h3ad582c4),
	.w2(32'h3a8e661d),
	.w3(32'h38b2889b),
	.w4(32'h39f3e266),
	.w5(32'h3af6c9c3),
	.w6(32'hba9a1cdf),
	.w7(32'hb9cd2f3d),
	.w8(32'h3a5dea58),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9b506),
	.w1(32'h3ad635fe),
	.w2(32'h3afc5f16),
	.w3(32'h3aa7a307),
	.w4(32'h3aa3813e),
	.w5(32'h3a27ee34),
	.w6(32'h3a43e054),
	.w7(32'h3a9c2ca9),
	.w8(32'h39a1081a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b3c2af),
	.w1(32'hb805818c),
	.w2(32'hb9678b14),
	.w3(32'h3a8ae631),
	.w4(32'h3a02fcfb),
	.w5(32'h3a7681d7),
	.w6(32'h3a492ca2),
	.w7(32'hb96bfbdd),
	.w8(32'h3af7c2d1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0338ad),
	.w1(32'h39b66ae0),
	.w2(32'hbac8619b),
	.w3(32'h3c39a259),
	.w4(32'h3b25f3e6),
	.w5(32'hba946aa6),
	.w6(32'h3b67dd34),
	.w7(32'hbb04cd83),
	.w8(32'hbc080f99),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa670b1),
	.w1(32'h39527fe5),
	.w2(32'hb9827ad0),
	.w3(32'h3b646524),
	.w4(32'h3a218832),
	.w5(32'hbacaa94c),
	.w6(32'h3b4be946),
	.w7(32'hb9da0053),
	.w8(32'hbaffa57a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397f8bee),
	.w1(32'h3746636a),
	.w2(32'h3930b56b),
	.w3(32'h394111e9),
	.w4(32'hba3a1fbd),
	.w5(32'hb9c9e5cc),
	.w6(32'hb9a01547),
	.w7(32'hba660ff3),
	.w8(32'hb967890d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b279666),
	.w1(32'h3b5a42ee),
	.w2(32'h3a81258f),
	.w3(32'hba80659d),
	.w4(32'hba67703c),
	.w5(32'h393a79be),
	.w6(32'hba13f4f0),
	.w7(32'hb96abb02),
	.w8(32'hba2fd606),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b9fd2),
	.w1(32'h39abf5db),
	.w2(32'hb924dab7),
	.w3(32'h365c6ac9),
	.w4(32'hb94a5deb),
	.w5(32'hbaf64f82),
	.w6(32'h3a1e3661),
	.w7(32'h38ecdcbd),
	.w8(32'hbaefe9c1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c16b62),
	.w1(32'hba8bb8a5),
	.w2(32'hb9182c5f),
	.w3(32'hbab0969f),
	.w4(32'hbaf28d32),
	.w5(32'hbae1c26d),
	.w6(32'hba7561a9),
	.w7(32'hbabc486a),
	.w8(32'hbafd6612),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed2d4c),
	.w1(32'hba651146),
	.w2(32'hbb0a9fa1),
	.w3(32'hb9b6a01b),
	.w4(32'hbacdf4f2),
	.w5(32'hba926450),
	.w6(32'h3a266cd2),
	.w7(32'hba80fc00),
	.w8(32'hba3ab375),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88b296),
	.w1(32'h3ae4d014),
	.w2(32'h39e808d8),
	.w3(32'h3bae7a64),
	.w4(32'h3b0fdad6),
	.w5(32'hba935e79),
	.w6(32'h3bd39c05),
	.w7(32'h3b19f690),
	.w8(32'hba498aa6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7ac8),
	.w1(32'hbb254649),
	.w2(32'hbb1b1260),
	.w3(32'hba3a7018),
	.w4(32'hbaba1a65),
	.w5(32'hbb264855),
	.w6(32'h3a63dab1),
	.w7(32'hba677428),
	.w8(32'hbb448822),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386c11c4),
	.w1(32'hbb1f9319),
	.w2(32'hba9f0bfd),
	.w3(32'hb8a63a5e),
	.w4(32'hbae95e77),
	.w5(32'hbb0503cb),
	.w6(32'hb9c9678c),
	.w7(32'hbab90eef),
	.w8(32'hbaff591b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad98989),
	.w1(32'h3912446f),
	.w2(32'hba6f90de),
	.w3(32'h3b300add),
	.w4(32'hba335a69),
	.w5(32'hbae0825d),
	.w6(32'h3b6595cf),
	.w7(32'h3948407b),
	.w8(32'hbaf8863f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95be5a),
	.w1(32'hba769eed),
	.w2(32'hbae4a57c),
	.w3(32'hb9bb66ed),
	.w4(32'hba6e82b3),
	.w5(32'hbb59d4bf),
	.w6(32'hba5abec4),
	.w7(32'hba8c8163),
	.w8(32'hbb7d3b3a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac82b4e),
	.w1(32'hbad4eccc),
	.w2(32'hba98e0fc),
	.w3(32'h3aad762f),
	.w4(32'hba183f44),
	.w5(32'hbae890c8),
	.w6(32'h3b361a77),
	.w7(32'h39b4bee5),
	.w8(32'hba932c26),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5210b0),
	.w1(32'hb982b261),
	.w2(32'hba124d74),
	.w3(32'hb8aa1a09),
	.w4(32'hba861fd7),
	.w5(32'h39034b5e),
	.w6(32'h393b36f1),
	.w7(32'hba11847d),
	.w8(32'hba6e8e1e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac7965),
	.w1(32'hbb8cf494),
	.w2(32'hbadf3c0f),
	.w3(32'hbb278028),
	.w4(32'hbbd57056),
	.w5(32'hbb85a15f),
	.w6(32'hb791f895),
	.w7(32'hbb6ab41f),
	.w8(32'hbb1fc03b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafb06d),
	.w1(32'hbac64988),
	.w2(32'hbadd4000),
	.w3(32'hba59720f),
	.w4(32'hbae5dfd2),
	.w5(32'hba8fae5d),
	.w6(32'hba6a5264),
	.w7(32'hbaf8cdd2),
	.w8(32'hba8b2c3f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a453af9),
	.w1(32'h3ac5ccef),
	.w2(32'h3adabd01),
	.w3(32'h3ac5628e),
	.w4(32'h3aa0171a),
	.w5(32'h37874ca9),
	.w6(32'h3a09a7ef),
	.w7(32'h39a328d8),
	.w8(32'hbab9362f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1c088),
	.w1(32'hba872f63),
	.w2(32'hbaa2637d),
	.w3(32'h3923f01b),
	.w4(32'h388debcf),
	.w5(32'hba0dcff9),
	.w6(32'hbadf056d),
	.w7(32'hbad4a252),
	.w8(32'hba5bacb3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d4668),
	.w1(32'h3a0dce56),
	.w2(32'hba0fc79a),
	.w3(32'hba6c09fb),
	.w4(32'hba8e3fe7),
	.w5(32'hba2ff1fd),
	.w6(32'hba6cd7ba),
	.w7(32'hba7c43a7),
	.w8(32'h3ada14a8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d8614),
	.w1(32'hbad30f59),
	.w2(32'hbada8610),
	.w3(32'hbb70d8d7),
	.w4(32'hbb904b68),
	.w5(32'hbb0abe26),
	.w6(32'h3a6598d1),
	.w7(32'hba863bb0),
	.w8(32'hbb066b9b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d956c),
	.w1(32'h3aec752a),
	.w2(32'hba888810),
	.w3(32'h3ba3d4da),
	.w4(32'h3afee30a),
	.w5(32'hba94d157),
	.w6(32'h3b86b262),
	.w7(32'h39f3c5b6),
	.w8(32'hbb023a32),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be625c),
	.w1(32'h39c3e590),
	.w2(32'hb88abd5c),
	.w3(32'hb8f40c9e),
	.w4(32'hb8ab0c4e),
	.w5(32'h3af87ee3),
	.w6(32'hb9d9f11b),
	.w7(32'hba6114de),
	.w8(32'h398ea2d5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b633a5),
	.w1(32'hbabf2b1d),
	.w2(32'hbacc52e3),
	.w3(32'h3b7d4c3c),
	.w4(32'h3aa16682),
	.w5(32'hba995f29),
	.w6(32'h3b957e6e),
	.w7(32'hb9c53818),
	.w8(32'hba96da9c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a057b83),
	.w1(32'hb997687f),
	.w2(32'hb89aaeff),
	.w3(32'h3b25cd55),
	.w4(32'h3a8611ae),
	.w5(32'hbb52334a),
	.w6(32'h3b2e120b),
	.w7(32'h393f089d),
	.w8(32'hbb4028f4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4376db),
	.w1(32'h3a6cd96e),
	.w2(32'hb99e92d8),
	.w3(32'h3b177242),
	.w4(32'hbae84fcb),
	.w5(32'hbaa80f7e),
	.w6(32'h3b84eb71),
	.w7(32'hba671e36),
	.w8(32'h3b33aa51),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd5108),
	.w1(32'h3bd02fe2),
	.w2(32'h3b6a237f),
	.w3(32'hbb1e3db5),
	.w4(32'hb917689e),
	.w5(32'hbac5970f),
	.w6(32'h3c0459a9),
	.w7(32'h3b93979a),
	.w8(32'hba0a818d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1578fa),
	.w1(32'hbacfb345),
	.w2(32'hbadb3d30),
	.w3(32'h3a66dddb),
	.w4(32'h3a6d0a39),
	.w5(32'hbac38ce7),
	.w6(32'h3a6826d5),
	.w7(32'h39680591),
	.w8(32'hbac2f115),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d79c87),
	.w1(32'hb9c4fca7),
	.w2(32'h37f49e93),
	.w3(32'hb8bcd63b),
	.w4(32'h39a9ce9f),
	.w5(32'hbb0bbe13),
	.w6(32'hba2bca39),
	.w7(32'hb7f5736d),
	.w8(32'hbb2992d3),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb077d3a),
	.w1(32'hbac13b6c),
	.w2(32'hbac397fb),
	.w3(32'hbab6808f),
	.w4(32'hbacf1c2e),
	.w5(32'hbac22c3f),
	.w6(32'hbac726a7),
	.w7(32'hbb08d44c),
	.w8(32'hbad3feb0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74e4ac3),
	.w1(32'h3b40ae26),
	.w2(32'h3b35e37d),
	.w3(32'hbb17415a),
	.w4(32'hba78b440),
	.w5(32'hbae08973),
	.w6(32'h3a383aa0),
	.w7(32'h3b1d4e8c),
	.w8(32'hb9d3dfc4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab4078),
	.w1(32'hb962f4ad),
	.w2(32'hbaab8171),
	.w3(32'hbae038f1),
	.w4(32'hb78b4ddb),
	.w5(32'h3b1ed437),
	.w6(32'hbb182f8c),
	.w7(32'hb9c4db02),
	.w8(32'h3b56ae48),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10e488),
	.w1(32'h3a779ad3),
	.w2(32'h39334d13),
	.w3(32'h3b1efb97),
	.w4(32'h3ae7b96a),
	.w5(32'hba7a4e47),
	.w6(32'h3b8c70b2),
	.w7(32'h3b35e06e),
	.w8(32'hba5c1202),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63ff99),
	.w1(32'h3a9d1f1a),
	.w2(32'h39d7b5ac),
	.w3(32'hba0aee28),
	.w4(32'hba26cee8),
	.w5(32'h3ad018bf),
	.w6(32'hba673dd3),
	.w7(32'hba6c1a31),
	.w8(32'h3b658b5c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd11b4),
	.w1(32'h3b08ec09),
	.w2(32'hb9bef090),
	.w3(32'h3b861522),
	.w4(32'h3b36316c),
	.w5(32'hba1e1da0),
	.w6(32'h3bed16e8),
	.w7(32'h3b603f56),
	.w8(32'hbace16e7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1db003),
	.w1(32'h3aba23ee),
	.w2(32'h3a1aa6ce),
	.w3(32'h3a1b6217),
	.w4(32'h389d716b),
	.w5(32'hb971692e),
	.w6(32'h3a060710),
	.w7(32'h39b888cd),
	.w8(32'h3a21cb9b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9967084),
	.w1(32'hb9bb04fa),
	.w2(32'hb897949e),
	.w3(32'h3a25e04d),
	.w4(32'hba4d6306),
	.w5(32'hb9c1589f),
	.w6(32'h3a8230a8),
	.w7(32'hba829a73),
	.w8(32'hba84a74f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0e25f),
	.w1(32'h3a510f4d),
	.w2(32'hbab884f0),
	.w3(32'hb98aad34),
	.w4(32'hbac99592),
	.w5(32'h3ae258d6),
	.w6(32'hb9b850c2),
	.w7(32'hbacd5426),
	.w8(32'h3b6bd25e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee4ef4),
	.w1(32'h3b4ab9a2),
	.w2(32'h3b56a2a4),
	.w3(32'h3b8baeaf),
	.w4(32'h3b91816f),
	.w5(32'h3b34b201),
	.w6(32'h3bacfad3),
	.w7(32'h3b9ef248),
	.w8(32'h3a520d98),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3fafc),
	.w1(32'h3a52d284),
	.w2(32'h3ac5aca2),
	.w3(32'h38adde07),
	.w4(32'h39cff9ea),
	.w5(32'hba6fe1ee),
	.w6(32'hb7252dd5),
	.w7(32'h3a2d982e),
	.w8(32'hba16a3f5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97430b5),
	.w1(32'h38a1b8a9),
	.w2(32'hb8ddc264),
	.w3(32'hba8cddbb),
	.w4(32'hbac97563),
	.w5(32'hba329102),
	.w6(32'hba6fb93c),
	.w7(32'hba63855c),
	.w8(32'hbb12202b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb507a1c),
	.w1(32'hbb8ad004),
	.w2(32'hbb8e87a1),
	.w3(32'h3a6a66ba),
	.w4(32'hb928bed1),
	.w5(32'hbb0403d2),
	.w6(32'h3a3a1cd2),
	.w7(32'hbad1e709),
	.w8(32'hbb217282),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a162a81),
	.w1(32'hbab1caa6),
	.w2(32'h373e13e2),
	.w3(32'h3bab42dd),
	.w4(32'h3b2131fb),
	.w5(32'hb99d0b34),
	.w6(32'h3b800f2a),
	.w7(32'h3aabab05),
	.w8(32'hbb827d35),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12b06a),
	.w1(32'h3a0b229e),
	.w2(32'h3922bfb8),
	.w3(32'h3ac1eba5),
	.w4(32'h3b32920f),
	.w5(32'h3ad6fbc7),
	.w6(32'hb917388b),
	.w7(32'h3a61c160),
	.w8(32'h3b015131),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff5b8c),
	.w1(32'hbac0dc1c),
	.w2(32'hbb0ec6b5),
	.w3(32'h3b03e39b),
	.w4(32'hbb0cfad5),
	.w5(32'hbbaabd2f),
	.w6(32'h3b5e1c56),
	.w7(32'hba0cffb9),
	.w8(32'hbbb9011a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04c82a),
	.w1(32'h3945120d),
	.w2(32'hba95273f),
	.w3(32'hbafbcbc8),
	.w4(32'hba9b58b4),
	.w5(32'hba102f05),
	.w6(32'hba92a2b4),
	.w7(32'hba1bdbeb),
	.w8(32'h362b7d99),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafacc13),
	.w1(32'hbae5bfc5),
	.w2(32'hbb2aa778),
	.w3(32'h3a6e10de),
	.w4(32'h3a887a5c),
	.w5(32'h3994cdce),
	.w6(32'h3a07e27e),
	.w7(32'hbae4a8bb),
	.w8(32'h3a84d088),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ba743),
	.w1(32'hb9ca28b7),
	.w2(32'hba5a4cad),
	.w3(32'h3ae41ea3),
	.w4(32'h3ae8e8b3),
	.w5(32'hbab2818e),
	.w6(32'h3b762f16),
	.w7(32'h3b0a4721),
	.w8(32'hba913eee),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe14e8),
	.w1(32'hbb4a6023),
	.w2(32'hbb1b99cb),
	.w3(32'h3b1c951e),
	.w4(32'hb9b38508),
	.w5(32'hba18f922),
	.w6(32'h3b308c10),
	.w7(32'hba9b5ee0),
	.w8(32'hbadf9544),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2037c4),
	.w1(32'h39ea9e88),
	.w2(32'h3a4ef3cf),
	.w3(32'h3ab46d8c),
	.w4(32'h3a9eedf1),
	.w5(32'hb9959f80),
	.w6(32'h3986c05d),
	.w7(32'h396ea58d),
	.w8(32'hba0df49a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bf930),
	.w1(32'hbb1e2222),
	.w2(32'hbb3162b1),
	.w3(32'hbb36a41f),
	.w4(32'hbb7dffdc),
	.w5(32'hbb0609a2),
	.w6(32'hbaac1c94),
	.w7(32'hbb415f18),
	.w8(32'hbaed71dc),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba601a79),
	.w1(32'hba796570),
	.w2(32'hb9641392),
	.w3(32'h3aa78de0),
	.w4(32'h3ada5ce6),
	.w5(32'h3a0c4b4d),
	.w6(32'hb9071b8d),
	.w7(32'h38c0ca1e),
	.w8(32'h39ec8b66),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d49b73),
	.w1(32'hb97f5c98),
	.w2(32'hbb22d8e8),
	.w3(32'h3ab2d87a),
	.w4(32'hba2d48dd),
	.w5(32'hb937d706),
	.w6(32'hb9295a7d),
	.w7(32'hbadfcf69),
	.w8(32'hb9e8c774),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb07f8),
	.w1(32'h3a24db8e),
	.w2(32'hb80e8043),
	.w3(32'hba01a6b4),
	.w4(32'hbae3c817),
	.w5(32'hba9c1cd1),
	.w6(32'h397ab31e),
	.w7(32'hb9ad6850),
	.w8(32'hb9e67a21),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43a264),
	.w1(32'hb9d12eb2),
	.w2(32'hbab91d03),
	.w3(32'hb9861c1b),
	.w4(32'hbb1c79b9),
	.w5(32'hbb4559ce),
	.w6(32'h3ad8607e),
	.w7(32'hba93f411),
	.w8(32'hbb15bbd1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4959d6),
	.w1(32'hbafb961b),
	.w2(32'hbb017377),
	.w3(32'hb95bfd25),
	.w4(32'hba40d9bd),
	.w5(32'h3b4a4c90),
	.w6(32'hba15880f),
	.w7(32'hba922b42),
	.w8(32'h3b4bfe13),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdf082),
	.w1(32'h3ab737b1),
	.w2(32'h397fe1d0),
	.w3(32'h3b26ad08),
	.w4(32'h3a5d7cce),
	.w5(32'hbb1c67fb),
	.w6(32'h3b3c9d73),
	.w7(32'h3aba7f29),
	.w8(32'hbb2f12bc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bf92b),
	.w1(32'hb9eb77b9),
	.w2(32'h3a71c141),
	.w3(32'hbb0934f2),
	.w4(32'hbaf6572f),
	.w5(32'hb9b15cc4),
	.w6(32'hbb052d42),
	.w7(32'hbb25eee6),
	.w8(32'hba69d1ef),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f0c60),
	.w1(32'hbaf6ec6b),
	.w2(32'hbb853472),
	.w3(32'hba2a3313),
	.w4(32'hba6dfcd4),
	.w5(32'hbbbd2f31),
	.w6(32'h3b194d70),
	.w7(32'h3902bace),
	.w8(32'hbbcab958),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fd2a6),
	.w1(32'hba8bf1dc),
	.w2(32'hba017639),
	.w3(32'hbad6cdb3),
	.w4(32'hbb1a9ff9),
	.w5(32'h3a701624),
	.w6(32'h399a710b),
	.w7(32'h3a7f82f1),
	.w8(32'hba8ac6e5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7c632),
	.w1(32'hba064228),
	.w2(32'hb606ce0e),
	.w3(32'h3aeb69c5),
	.w4(32'h3b0640f7),
	.w5(32'h3ad33ec8),
	.w6(32'h37ee3866),
	.w7(32'h398794de),
	.w8(32'h3a889644),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0cb20),
	.w1(32'h3b32810f),
	.w2(32'h3b4bb491),
	.w3(32'h3c2b0c69),
	.w4(32'h3ba56d43),
	.w5(32'h3a7266b1),
	.w6(32'h3c08abf2),
	.w7(32'h3b33f1c4),
	.w8(32'hbb0b9507),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16f7c7),
	.w1(32'h3b18d4d3),
	.w2(32'hba86d39e),
	.w3(32'hbacf04d7),
	.w4(32'hb7723c14),
	.w5(32'hbb0775f1),
	.w6(32'h3b15101f),
	.w7(32'hbb197cef),
	.w8(32'h3a8e45b4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b707e7a),
	.w1(32'h3ae255f1),
	.w2(32'h3a52ae02),
	.w3(32'h3b39b7e5),
	.w4(32'h3aea9152),
	.w5(32'hb9b9db07),
	.w6(32'h3b9090a1),
	.w7(32'h3b18b001),
	.w8(32'hb86edbfb),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39484700),
	.w1(32'h399bb458),
	.w2(32'h39dceb15),
	.w3(32'hba18246e),
	.w4(32'hba3b2f68),
	.w5(32'hb9792120),
	.w6(32'hb91c008a),
	.w7(32'h39e75b86),
	.w8(32'hb9547984),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f4d42),
	.w1(32'hb92bdec7),
	.w2(32'h3a8e77ea),
	.w3(32'hb9022fe0),
	.w4(32'h3937daa3),
	.w5(32'hba98ab91),
	.w6(32'hb9a278e6),
	.w7(32'h3a02d409),
	.w8(32'hba17d9e4),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85c2b2a),
	.w1(32'hba471d71),
	.w2(32'hbb1ce923),
	.w3(32'hbaac5013),
	.w4(32'hbb5158b8),
	.w5(32'h3a87a6af),
	.w6(32'hbab35369),
	.w7(32'hbb3f4735),
	.w8(32'h3afddc6b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8599cc),
	.w1(32'h3617bcb4),
	.w2(32'hba8e9c19),
	.w3(32'h3b9a54e7),
	.w4(32'h3b14feba),
	.w5(32'hb99adbae),
	.w6(32'h3bb99598),
	.w7(32'h3b488ee0),
	.w8(32'hbab3b4e8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fe32c),
	.w1(32'hba500f78),
	.w2(32'hb8c90d7d),
	.w3(32'h3b16283c),
	.w4(32'hb996df70),
	.w5(32'hbb298c36),
	.w6(32'h39cf4b58),
	.w7(32'hbae278fe),
	.w8(32'hbb39b6e2),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb643946),
	.w1(32'hbba0ab1d),
	.w2(32'hbbcbe4c7),
	.w3(32'hbb19f644),
	.w4(32'hbb9ebc32),
	.w5(32'hba94ade4),
	.w6(32'hba9f3725),
	.w7(32'hbb850f09),
	.w8(32'hb9814804),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a0586),
	.w1(32'h3b3a8dfe),
	.w2(32'h39dba8cc),
	.w3(32'h3b2b31d2),
	.w4(32'h3a550489),
	.w5(32'hb94e9f09),
	.w6(32'h3b730bfb),
	.w7(32'h3a3513c1),
	.w8(32'hba0ea3ad),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78e0f2),
	.w1(32'h39266b46),
	.w2(32'hbab7a604),
	.w3(32'h3b8d7ce8),
	.w4(32'h3a0a6038),
	.w5(32'hba97fc48),
	.w6(32'h3b793f4a),
	.w7(32'h39ad08a4),
	.w8(32'hbaeb2348),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa66e05),
	.w1(32'hba59df73),
	.w2(32'hb995cbe3),
	.w3(32'h38c500e3),
	.w4(32'h3a3c0cc2),
	.w5(32'hbae874af),
	.w6(32'h379b34cc),
	.w7(32'h398e1b0a),
	.w8(32'hbb215156),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae4d58),
	.w1(32'hba8449d1),
	.w2(32'hba5b6ace),
	.w3(32'hba84f942),
	.w4(32'hba2c609f),
	.w5(32'hba35491f),
	.w6(32'hba8c9bdb),
	.w7(32'hba6ae77d),
	.w8(32'hba81ea54),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fa640),
	.w1(32'hbb1f9b53),
	.w2(32'hb99da867),
	.w3(32'hbb4c426b),
	.w4(32'hbb4ad0df),
	.w5(32'hba726882),
	.w6(32'hba9a44ab),
	.w7(32'hbaac062f),
	.w8(32'h39827687),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983441f),
	.w1(32'h399ff5d4),
	.w2(32'h3a505a80),
	.w3(32'h3a3f9efc),
	.w4(32'h389a3259),
	.w5(32'h3a1ca052),
	.w6(32'h39d638e6),
	.w7(32'h3a82ed23),
	.w8(32'hb9857067),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cb285),
	.w1(32'h3a97a50c),
	.w2(32'hba90f1c4),
	.w3(32'h3b7097b1),
	.w4(32'h3aaeefa1),
	.w5(32'hbb136878),
	.w6(32'h3b17e052),
	.w7(32'h3a065b53),
	.w8(32'hbb1a45b7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567efc),
	.w1(32'hbaa0ad94),
	.w2(32'hba8fec21),
	.w3(32'hbbce7694),
	.w4(32'hbb548474),
	.w5(32'hbabde335),
	.w6(32'hbba0a696),
	.w7(32'hbb218c63),
	.w8(32'hbae56eb2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9911e6),
	.w1(32'hbac13d0a),
	.w2(32'hbaec7d2a),
	.w3(32'h3af0a491),
	.w4(32'h3a6e50a1),
	.w5(32'hbacba073),
	.w6(32'h3af2190a),
	.w7(32'h398ad01a),
	.w8(32'hbb0582b9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84d2a5),
	.w1(32'h3a849480),
	.w2(32'hb97bc0ee),
	.w3(32'h3a32b47e),
	.w4(32'h3987cc10),
	.w5(32'hba6a2414),
	.w6(32'h3a06c9e5),
	.w7(32'hb7fa0228),
	.w8(32'hba6ba80c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63f445),
	.w1(32'hbb0c9ee4),
	.w2(32'hbb549238),
	.w3(32'hb9cda4c7),
	.w4(32'hbacd8578),
	.w5(32'hbb23aeda),
	.w6(32'h3ab44718),
	.w7(32'hbaa13970),
	.w8(32'hbb357275),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94ffd9),
	.w1(32'hb906ce28),
	.w2(32'hba458665),
	.w3(32'h3b5bf6d3),
	.w4(32'h3a15b99c),
	.w5(32'hbb06261b),
	.w6(32'h3b4e7a7c),
	.w7(32'hb764061b),
	.w8(32'hbae13d14),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2201bf),
	.w1(32'hb99a15d3),
	.w2(32'h3a80f3f3),
	.w3(32'h3ab53a3e),
	.w4(32'h3a66c0b0),
	.w5(32'h3a2ce2f7),
	.w6(32'h3b35c4f9),
	.w7(32'h3aaee3d9),
	.w8(32'h39be1dd9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a849972),
	.w1(32'h3a553f25),
	.w2(32'hb8a5fbe9),
	.w3(32'h395bffc9),
	.w4(32'hb9d7947b),
	.w5(32'h39c67190),
	.w6(32'h39f0e842),
	.w7(32'h39e9fa15),
	.w8(32'h3af3b0da),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9188fb),
	.w1(32'h3b6d93bb),
	.w2(32'h3a467f3c),
	.w3(32'hba317822),
	.w4(32'hba869cc4),
	.w5(32'hb9e1c41a),
	.w6(32'h3b0ed315),
	.w7(32'h3a255fd6),
	.w8(32'hb8cbb2c7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109989),
	.w1(32'hb9d33b09),
	.w2(32'hbade590c),
	.w3(32'h3b15ea92),
	.w4(32'h373148df),
	.w5(32'h39e1d041),
	.w6(32'h3a811158),
	.w7(32'hba647122),
	.w8(32'hbb7102da),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cc9e3),
	.w1(32'h3a1aded9),
	.w2(32'hb95dd14c),
	.w3(32'h3b2767b4),
	.w4(32'hbab07be8),
	.w5(32'hbabc2102),
	.w6(32'h3b3d9dd3),
	.w7(32'hba235614),
	.w8(32'hbb2eae96),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e0f34),
	.w1(32'h39996604),
	.w2(32'hbabc5d10),
	.w3(32'h3a5cc577),
	.w4(32'hb9f713bc),
	.w5(32'hbb43052d),
	.w6(32'h3b10a2a7),
	.w7(32'h39abf999),
	.w8(32'hbbb79ef6),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b277a7e),
	.w1(32'hb9cbe525),
	.w2(32'hba97d087),
	.w3(32'hb9ba6da1),
	.w4(32'hbb635b9a),
	.w5(32'hbac16c27),
	.w6(32'h3baaab2e),
	.w7(32'hb9c975e0),
	.w8(32'h39ee5b5a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba901062),
	.w1(32'hba73b3b2),
	.w2(32'hbab7a093),
	.w3(32'h3ac1793c),
	.w4(32'h39f81482),
	.w5(32'h3a2cedbe),
	.w6(32'hbaa80fb6),
	.w7(32'hbac115bf),
	.w8(32'hb956be98),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab8ba9),
	.w1(32'hba624440),
	.w2(32'hba909902),
	.w3(32'h3a014e7e),
	.w4(32'hba16cb4e),
	.w5(32'h39f68344),
	.w6(32'h39a0ef14),
	.w7(32'hba782c4e),
	.w8(32'h3a0c6165),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91450f),
	.w1(32'h3b312922),
	.w2(32'hba84f43e),
	.w3(32'h3bcc334f),
	.w4(32'h3bd1c1d9),
	.w5(32'h3710ef70),
	.w6(32'h3a36f858),
	.w7(32'h3b93f7f3),
	.w8(32'hbb4ba420),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aaef1),
	.w1(32'h3b432fba),
	.w2(32'h3a2e6448),
	.w3(32'h3bb8332e),
	.w4(32'h3abe1df4),
	.w5(32'h39d3b7cc),
	.w6(32'h3b364a0c),
	.w7(32'hba39afcc),
	.w8(32'hba191233),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b453a21),
	.w1(32'h37e54778),
	.w2(32'hba98581e),
	.w3(32'h3b026a60),
	.w4(32'h3872a809),
	.w5(32'hbb9572d9),
	.w6(32'h3b539ffd),
	.w7(32'h3a52be5f),
	.w8(32'hbb9cc730),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d4e9),
	.w1(32'hbb71f8f4),
	.w2(32'hbb1e611f),
	.w3(32'hbb951940),
	.w4(32'hbb4143fa),
	.w5(32'hbb001f77),
	.w6(32'hbba3a4d1),
	.w7(32'hbb583b9c),
	.w8(32'hba085066),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb105525),
	.w1(32'hbb46de83),
	.w2(32'hbb770b15),
	.w3(32'hbb1b9608),
	.w4(32'hbb214bdd),
	.w5(32'hbb5ea0ad),
	.w6(32'h397a53ac),
	.w7(32'hbad14e08),
	.w8(32'hbb2bb44e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56166c),
	.w1(32'h3a8b96a4),
	.w2(32'h3a8219fd),
	.w3(32'hb901a7b4),
	.w4(32'h37195dff),
	.w5(32'h398b3b94),
	.w6(32'h3a4898fd),
	.w7(32'h3a5416b2),
	.w8(32'h3934d537),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5e886),
	.w1(32'h3b2140b4),
	.w2(32'h3b21cfd9),
	.w3(32'h398ecb69),
	.w4(32'h3a16345c),
	.w5(32'hbb1682ab),
	.w6(32'hb9748e53),
	.w7(32'h39f45fd9),
	.w8(32'hbb197024),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cc49b),
	.w1(32'hbabec0d1),
	.w2(32'hba92510e),
	.w3(32'hba94b584),
	.w4(32'hbb1b5e13),
	.w5(32'hbaf3282a),
	.w6(32'hb9b77037),
	.w7(32'hbb01de20),
	.w8(32'hbb084355),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c020d),
	.w1(32'hbb5aa37f),
	.w2(32'hbac3cfe1),
	.w3(32'hba4cdba5),
	.w4(32'h39d38b37),
	.w5(32'h3ad72869),
	.w6(32'hbb1ccd9f),
	.w7(32'hbb0de647),
	.w8(32'h3a8b67f9),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7ac44),
	.w1(32'hb99621ed),
	.w2(32'h3b84c505),
	.w3(32'h3bd59d71),
	.w4(32'h3abe88eb),
	.w5(32'h3c624c48),
	.w6(32'hbb8814e7),
	.w7(32'h3b0afc6d),
	.w8(32'h3be193d7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c190f25),
	.w1(32'h3bdba673),
	.w2(32'h3b5bfa56),
	.w3(32'h3b4b929f),
	.w4(32'h3ad747de),
	.w5(32'hbb7580d8),
	.w6(32'h3cd3ec67),
	.w7(32'h3ac7ab59),
	.w8(32'hbbda04cb),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1de02d),
	.w1(32'hba4f395d),
	.w2(32'h3bc14da0),
	.w3(32'hb91d6e80),
	.w4(32'h3bd5d5ca),
	.w5(32'hbb646ead),
	.w6(32'h3abe387d),
	.w7(32'h3c198faf),
	.w8(32'h3bb34cfc),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfcb0e),
	.w1(32'hbc37acc7),
	.w2(32'hbad4f4d3),
	.w3(32'h3a3a2586),
	.w4(32'h3bc83484),
	.w5(32'h3afbc18d),
	.w6(32'h3c447256),
	.w7(32'hbbc4efb4),
	.w8(32'hbae709e0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa9e1e),
	.w1(32'hbb73af7e),
	.w2(32'hba185264),
	.w3(32'h3b3121a7),
	.w4(32'h3b538d99),
	.w5(32'h3c1ead73),
	.w6(32'hba527463),
	.w7(32'h3ba43cb7),
	.w8(32'h3c4ebcc0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2777e),
	.w1(32'h3c029124),
	.w2(32'h3c994568),
	.w3(32'h3ce6690e),
	.w4(32'h3c34d129),
	.w5(32'h3b8e3edd),
	.w6(32'h3c2bde94),
	.w7(32'h3c8519df),
	.w8(32'hbb345f28),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a8192),
	.w1(32'hbc048b24),
	.w2(32'hb9adf6b2),
	.w3(32'hbc31fe5d),
	.w4(32'h3b842d7d),
	.w5(32'hbc031754),
	.w6(32'h3bfeb6ba),
	.w7(32'h3a134807),
	.w8(32'hbbea8d92),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81cfde),
	.w1(32'hbc147c19),
	.w2(32'h3b17e55d),
	.w3(32'hbc11721d),
	.w4(32'hbc1bfcd5),
	.w5(32'hba4c90b3),
	.w6(32'hbc04941c),
	.w7(32'hbc3844ef),
	.w8(32'hbac61a65),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bb963),
	.w1(32'h3c808b0b),
	.w2(32'h3c38ba82),
	.w3(32'hbb8ce53d),
	.w4(32'hbb0a946a),
	.w5(32'hbb4efb07),
	.w6(32'h3bcd327f),
	.w7(32'h3c2dcafa),
	.w8(32'hbc07ac0f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e502),
	.w1(32'h3b52c657),
	.w2(32'hbad5fbb2),
	.w3(32'hbb4dc459),
	.w4(32'h3a904ec1),
	.w5(32'hbc71493d),
	.w6(32'h3b9587c7),
	.w7(32'hb9a03c8e),
	.w8(32'hbc96aecd),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc477290),
	.w1(32'hbc699cb2),
	.w2(32'hbba278e4),
	.w3(32'hbbcf782f),
	.w4(32'hbc578e97),
	.w5(32'h3b1f28ba),
	.w6(32'hbca0aff6),
	.w7(32'hbc55d2a9),
	.w8(32'hba4a0b7c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98da59b),
	.w1(32'hba104a4f),
	.w2(32'hbae83177),
	.w3(32'hbb19074d),
	.w4(32'hbaf8083a),
	.w5(32'h3c62eeb5),
	.w6(32'h3b90233a),
	.w7(32'hba0983d1),
	.w8(32'h3c8861d8),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e7ca9),
	.w1(32'h3cdc6250),
	.w2(32'h3c681b6b),
	.w3(32'h3ca07810),
	.w4(32'h3cc1e5a8),
	.w5(32'hbb8d4ef7),
	.w6(32'h3d09e2a7),
	.w7(32'h3d0ac22a),
	.w8(32'h3a993b3d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbc9ff),
	.w1(32'hbbbd65a3),
	.w2(32'hbb910dcc),
	.w3(32'h3b175122),
	.w4(32'h3a39e0dc),
	.w5(32'hbc25b6c1),
	.w6(32'h3b8d2eb0),
	.w7(32'hbbbb7159),
	.w8(32'hbc3358d0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9684a0),
	.w1(32'hbbb4824b),
	.w2(32'hbbd31b33),
	.w3(32'hbbc4ffa2),
	.w4(32'hbb73d700),
	.w5(32'h3a9d88b5),
	.w6(32'h39f1f74a),
	.w7(32'hbb6c7f6e),
	.w8(32'h3ad6511b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bd2eb),
	.w1(32'h3c0352f5),
	.w2(32'h3bfeca5b),
	.w3(32'h3a09eef6),
	.w4(32'hbbbf61a3),
	.w5(32'hbc1dabc3),
	.w6(32'hbb9daa70),
	.w7(32'hbb2150a0),
	.w8(32'hbc164765),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d1484),
	.w1(32'hbb9d4f79),
	.w2(32'hbc3e65b4),
	.w3(32'hbc48a797),
	.w4(32'hbbb523a4),
	.w5(32'h3b739783),
	.w6(32'hbc80093a),
	.w7(32'hbbcffed3),
	.w8(32'h3be04ab3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ef518),
	.w1(32'hbbf89248),
	.w2(32'hbb9682e9),
	.w3(32'h3be821f5),
	.w4(32'h3b52f6ea),
	.w5(32'hbb695b9e),
	.w6(32'h3c277358),
	.w7(32'hbc0cee46),
	.w8(32'hbac35094),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46b1c9),
	.w1(32'hbbc4054c),
	.w2(32'hbb429c9e),
	.w3(32'hba85d574),
	.w4(32'hbbb4ba8c),
	.w5(32'h3aff058e),
	.w6(32'hbbd48405),
	.w7(32'hbb933244),
	.w8(32'hbbcae9b1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a7072),
	.w1(32'hbbb31fd0),
	.w2(32'h3a4a949c),
	.w3(32'h3b48e42f),
	.w4(32'hba9d5d84),
	.w5(32'h3c7e58fb),
	.w6(32'hbc16e348),
	.w7(32'h3c061f9b),
	.w8(32'h3bd43aba),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2c033),
	.w1(32'hbc0734b1),
	.w2(32'h3b0b1e92),
	.w3(32'h3b72342d),
	.w4(32'hba815964),
	.w5(32'h3c7ae8de),
	.w6(32'hbb8a032c),
	.w7(32'hbc057568),
	.w8(32'h3cf6e8ff),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac1bf4),
	.w1(32'h3c7a5814),
	.w2(32'h3ce2c950),
	.w3(32'h3d07572a),
	.w4(32'h3c6819b3),
	.w5(32'h39ad310e),
	.w6(32'hbbed226b),
	.w7(32'h3c4d1ca6),
	.w8(32'hba9910fc),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b844b),
	.w1(32'h36994834),
	.w2(32'h3bc22fce),
	.w3(32'h3acf5ab6),
	.w4(32'h3b8f1b54),
	.w5(32'h3b20d388),
	.w6(32'hba1339df),
	.w7(32'h3bc6df0c),
	.w8(32'h3b71019a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47bdeb),
	.w1(32'h3be58d1c),
	.w2(32'h3b01af0a),
	.w3(32'hbb4eddbc),
	.w4(32'h3b072444),
	.w5(32'hba94392b),
	.w6(32'hbbba6eab),
	.w7(32'h3bd6f776),
	.w8(32'hbc070e28),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dedb9),
	.w1(32'hbb11ea42),
	.w2(32'h3b726cd8),
	.w3(32'hbb87b3bb),
	.w4(32'h3a9c659a),
	.w5(32'h3b80bb75),
	.w6(32'hbbcd246e),
	.w7(32'hbba373ad),
	.w8(32'hbae50db2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4c44a),
	.w1(32'hbb32a3c2),
	.w2(32'h3b522c66),
	.w3(32'hb9e4a739),
	.w4(32'hbb676d15),
	.w5(32'h3b85bc53),
	.w6(32'hbb2be2e1),
	.w7(32'hbbc7b20e),
	.w8(32'hbc318a2e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f328f),
	.w1(32'hbb5fb0c1),
	.w2(32'hbc1e125e),
	.w3(32'hbabe64c0),
	.w4(32'h3aefd21d),
	.w5(32'hbb8d7317),
	.w6(32'hbac7f83f),
	.w7(32'h3ba30901),
	.w8(32'h3ba8d674),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905872a),
	.w1(32'h3c17e389),
	.w2(32'h3b92c6e8),
	.w3(32'h3badb5e9),
	.w4(32'h3b60c605),
	.w5(32'hba69386e),
	.w6(32'h3bf9048d),
	.w7(32'h3a36b6fb),
	.w8(32'hba2312ec),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b826c14),
	.w1(32'h39c5a94c),
	.w2(32'hbb7c3f71),
	.w3(32'hbb7e1663),
	.w4(32'hbb580cdf),
	.w5(32'hbb5b1ab3),
	.w6(32'hbb6b7898),
	.w7(32'h3af12243),
	.w8(32'h3be19257),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa7db5),
	.w1(32'h3c14531b),
	.w2(32'h3b71b61f),
	.w3(32'h3bc9b056),
	.w4(32'hb9505fc6),
	.w5(32'hbb8efd07),
	.w6(32'h3c0bada7),
	.w7(32'h3a923a18),
	.w8(32'hbc026ce7),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule