module layer_10_featuremap_35(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00f8e6),
	.w1(32'hbbd23fb1),
	.w2(32'h3c58f8ce),
	.w3(32'h3a8fb3e4),
	.w4(32'hba2ddb0b),
	.w5(32'h3b780ad7),
	.w6(32'hb16dd351),
	.w7(32'hbaa2f2b5),
	.w8(32'h3c506dab),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adafa9b),
	.w1(32'hbc1a22d9),
	.w2(32'h3bc8faef),
	.w3(32'h3bff5e4a),
	.w4(32'hbc025abd),
	.w5(32'hbb1d886d),
	.w6(32'h3b97b2cd),
	.w7(32'hb911bd21),
	.w8(32'hbc10aa3f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0c92),
	.w1(32'h3b116998),
	.w2(32'hbb7c600b),
	.w3(32'hbc2fc4af),
	.w4(32'hbac80f1a),
	.w5(32'hbaa34bbd),
	.w6(32'hbc094183),
	.w7(32'hbb8597c9),
	.w8(32'h3a1e29f6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a6cd3),
	.w1(32'hbabdd0b5),
	.w2(32'h3b694747),
	.w3(32'hbbb84327),
	.w4(32'hb90f9244),
	.w5(32'h3b0e4ccc),
	.w6(32'hba9fe22a),
	.w7(32'hbb419f32),
	.w8(32'hbbbf1932),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a2b6a),
	.w1(32'hbbe3edce),
	.w2(32'hbb873c9f),
	.w3(32'h3a148d5f),
	.w4(32'hbb223165),
	.w5(32'hbb41e676),
	.w6(32'hbb2ce627),
	.w7(32'hbc4ec3b7),
	.w8(32'hbbc5adb0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06ea28),
	.w1(32'hbc0d6eb7),
	.w2(32'hbbdaaf49),
	.w3(32'hbc1722f3),
	.w4(32'hbc66d64c),
	.w5(32'hbbbc164a),
	.w6(32'hbc420896),
	.w7(32'hbc59b885),
	.w8(32'hbb6140c5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eaebc),
	.w1(32'hbbb4e551),
	.w2(32'hbb2fe488),
	.w3(32'hbbb0a117),
	.w4(32'hbb93c2c1),
	.w5(32'hbc24def9),
	.w6(32'hbba8271c),
	.w7(32'hbb9fcad5),
	.w8(32'hbc0a0cf4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe263f3),
	.w1(32'hbba18758),
	.w2(32'hbb192cf9),
	.w3(32'hbba0f35f),
	.w4(32'hbb82a3b5),
	.w5(32'h3b168074),
	.w6(32'hbc21a8a9),
	.w7(32'hbc56d722),
	.w8(32'hbbda023c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3727fa00),
	.w1(32'hbbe72441),
	.w2(32'hbb497730),
	.w3(32'h3b36ce46),
	.w4(32'hbb527a17),
	.w5(32'hbc636e08),
	.w6(32'hbbd9f535),
	.w7(32'hbb8efa92),
	.w8(32'hbc2368e8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4f8dd),
	.w1(32'hbc328e4f),
	.w2(32'hbb29a6cf),
	.w3(32'hbd1a107b),
	.w4(32'hbcb0e055),
	.w5(32'hbc23b1fb),
	.w6(32'hbcf1d949),
	.w7(32'hbc0e3e7d),
	.w8(32'hbb489512),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39775dbb),
	.w1(32'h3ac4bb96),
	.w2(32'hbb88bf82),
	.w3(32'hba9d1dc5),
	.w4(32'h3a4070af),
	.w5(32'hb9f8bd6f),
	.w6(32'h3a650a83),
	.w7(32'h3b024e35),
	.w8(32'hb98f898b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cd179),
	.w1(32'hbb728bad),
	.w2(32'hbbb605ef),
	.w3(32'h385d78dd),
	.w4(32'hbad59cf6),
	.w5(32'hbbb85f28),
	.w6(32'h3b4a9dfa),
	.w7(32'h3b1db39b),
	.w8(32'hbbd128aa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd657db),
	.w1(32'hbc33f957),
	.w2(32'hbc23e511),
	.w3(32'hbceb6169),
	.w4(32'hbc48e682),
	.w5(32'hbc3ca845),
	.w6(32'hbc9e7ffc),
	.w7(32'hbb671b69),
	.w8(32'h3b0af23c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bdffc),
	.w1(32'hbb6bde19),
	.w2(32'h3c5e0f2f),
	.w3(32'hbb6e2e91),
	.w4(32'h3b3604fb),
	.w5(32'h3a22bf74),
	.w6(32'hba547dd0),
	.w7(32'hbbce378b),
	.w8(32'h3a2ab29a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ee94f),
	.w1(32'h3c943f5c),
	.w2(32'hbbbf702c),
	.w3(32'h39fb9be8),
	.w4(32'h3ba9a015),
	.w5(32'hbc13cf48),
	.w6(32'hbb7c8da9),
	.w7(32'h3b066420),
	.w8(32'hbc013649),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8910a2),
	.w1(32'hbb11bf78),
	.w2(32'h3995b6f8),
	.w3(32'hbc09b456),
	.w4(32'hbb5467ea),
	.w5(32'hbb0b839a),
	.w6(32'hbc5404c6),
	.w7(32'hbbdc3427),
	.w8(32'hb8447c0d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9870d),
	.w1(32'hb982f2fd),
	.w2(32'hba9e92ac),
	.w3(32'hba813a2f),
	.w4(32'h3a858bcc),
	.w5(32'hbb18e0c5),
	.w6(32'h3a3ed5f2),
	.w7(32'h3b5b1b11),
	.w8(32'hb97b9f44),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77055d),
	.w1(32'h3805c12b),
	.w2(32'hbb5e06e8),
	.w3(32'hbb3c0990),
	.w4(32'hbb2905db),
	.w5(32'hbc3345b6),
	.w6(32'hbaef079c),
	.w7(32'h3bbc332d),
	.w8(32'hb9c58a48),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12361a),
	.w1(32'hbb094886),
	.w2(32'h3c124d1e),
	.w3(32'hbb8bdae0),
	.w4(32'hba3812d0),
	.w5(32'hba78e739),
	.w6(32'hbbef1dcf),
	.w7(32'hbb44260b),
	.w8(32'h3b3f2fc0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b8131),
	.w1(32'h3bb0e913),
	.w2(32'h3aa385ba),
	.w3(32'h3c287b71),
	.w4(32'h3c103b0e),
	.w5(32'h3ac753c9),
	.w6(32'hbc4768bc),
	.w7(32'h3b307301),
	.w8(32'hba835322),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b805d5b),
	.w1(32'hb971efe7),
	.w2(32'h3bc61ead),
	.w3(32'h3b4ca787),
	.w4(32'hbb5ce2cf),
	.w5(32'h3af2cf69),
	.w6(32'hbb8985e6),
	.w7(32'hbbcb23da),
	.w8(32'h39c32fcb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc2ccc),
	.w1(32'h3b2d2e79),
	.w2(32'h3b4021d1),
	.w3(32'h3c0e2a0e),
	.w4(32'h3bbd3930),
	.w5(32'h3bf2b5c5),
	.w6(32'h3b4d5f67),
	.w7(32'h3baf0147),
	.w8(32'h3bf5a0c0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6923de),
	.w1(32'hba721d1e),
	.w2(32'hbc234dee),
	.w3(32'h3cc05896),
	.w4(32'h3c54f914),
	.w5(32'hbbac6d37),
	.w6(32'hbbccafad),
	.w7(32'hbba8d57f),
	.w8(32'hbc82b575),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1be358),
	.w1(32'hbb81fb00),
	.w2(32'hbc14bb0d),
	.w3(32'hbb35728c),
	.w4(32'hbba87f46),
	.w5(32'hbbe5c06b),
	.w6(32'hbc0337bf),
	.w7(32'hbba1048e),
	.w8(32'hbc054bd2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0c4b5),
	.w1(32'hba7a518b),
	.w2(32'h3a2e6cc8),
	.w3(32'h3b07dff7),
	.w4(32'h3b99b398),
	.w5(32'hbb03f0ba),
	.w6(32'hbc0841db),
	.w7(32'hbb812ab9),
	.w8(32'hb9893f13),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23ed5f),
	.w1(32'h3a72e17e),
	.w2(32'hbc35e811),
	.w3(32'h3c3ac366),
	.w4(32'h3b5edfcf),
	.w5(32'hba952fb7),
	.w6(32'hba0223aa),
	.w7(32'h3bb12d41),
	.w8(32'hb9e268f5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ffd57),
	.w1(32'hbab5d70f),
	.w2(32'h394d3824),
	.w3(32'h3ba18d90),
	.w4(32'h3bf5adda),
	.w5(32'h3ae591ed),
	.w6(32'hb9e73c58),
	.w7(32'h3c0ee03d),
	.w8(32'h3ac93001),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39b999),
	.w1(32'h3b4c32c6),
	.w2(32'h3c034103),
	.w3(32'h39bea6c1),
	.w4(32'h3ba8df1a),
	.w5(32'h39f6dba5),
	.w6(32'hbb0ac9e1),
	.w7(32'h3b2f12c0),
	.w8(32'h3c0434c5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cc585),
	.w1(32'h3c10dc5c),
	.w2(32'h3be1f1ae),
	.w3(32'hbc61d53d),
	.w4(32'h3b2e35ff),
	.w5(32'h3c1b0441),
	.w6(32'hbbbbb9c7),
	.w7(32'hb9c5fd93),
	.w8(32'h3a786230),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b32a7),
	.w1(32'h3b4ea396),
	.w2(32'hbbc9a70d),
	.w3(32'h3ceb4bdc),
	.w4(32'h3d07087c),
	.w5(32'hbbf36e7c),
	.w6(32'hbc45612b),
	.w7(32'h3c18dac5),
	.w8(32'hbc11088c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b00df),
	.w1(32'h3a7b398a),
	.w2(32'h3c01e93d),
	.w3(32'hbb269998),
	.w4(32'hbb27c0dc),
	.w5(32'h3ad8cf40),
	.w6(32'hbad48134),
	.w7(32'hba1e56ed),
	.w8(32'hba1db1e5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95bf250),
	.w1(32'hb89379f0),
	.w2(32'hbba10d68),
	.w3(32'h3b514d0d),
	.w4(32'hbaeb1f9c),
	.w5(32'hbbf5b0a7),
	.w6(32'hba560654),
	.w7(32'h3b8e679f),
	.w8(32'hbcebb2eb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03e552),
	.w1(32'hba7ec15d),
	.w2(32'hbb734d18),
	.w3(32'hba166d8e),
	.w4(32'hbb4307ae),
	.w5(32'hbb9773db),
	.w6(32'hbcf0cb5c),
	.w7(32'hbc876e85),
	.w8(32'h39f98a53),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19504d),
	.w1(32'hb8c2aaf2),
	.w2(32'hbbd59abc),
	.w3(32'hbb66601d),
	.w4(32'h39bd0082),
	.w5(32'h3bc71cfe),
	.w6(32'hbb39aba3),
	.w7(32'hbb03d094),
	.w8(32'h3c0c9daf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b6ab6),
	.w1(32'hbb5f2dc9),
	.w2(32'h3b9bbac8),
	.w3(32'hbb85724f),
	.w4(32'h3a8ad5ba),
	.w5(32'h3b5cf319),
	.w6(32'h3b089012),
	.w7(32'hb97e18b0),
	.w8(32'h3ac12a3d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4736c8),
	.w1(32'h3b77ee11),
	.w2(32'hba4e5e11),
	.w3(32'hba8d4e62),
	.w4(32'h3b59d3e8),
	.w5(32'hbbb21a42),
	.w6(32'h3af9c3fa),
	.w7(32'h3a62a8ac),
	.w8(32'hba84c2f9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81392a),
	.w1(32'hbbb8b5f0),
	.w2(32'hbb78f07f),
	.w3(32'hbb77d0e9),
	.w4(32'h3c2afce5),
	.w5(32'hbc3aba08),
	.w6(32'hbc5487c5),
	.w7(32'hbbf22991),
	.w8(32'hbac2960a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5ea9c),
	.w1(32'hba3824b3),
	.w2(32'h3c7dad44),
	.w3(32'hbc2f38fb),
	.w4(32'h3c233dcc),
	.w5(32'h3afc1105),
	.w6(32'hbc46a871),
	.w7(32'hbb68d27e),
	.w8(32'h3b5925f7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3a706b),
	.w1(32'h3c4074cc),
	.w2(32'h3c3699a3),
	.w3(32'h3bed0aee),
	.w4(32'h3cd9f49b),
	.w5(32'h3d4c9247),
	.w6(32'hbca73444),
	.w7(32'hbc46633c),
	.w8(32'hbadfd66f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6e301),
	.w1(32'hbc448b8f),
	.w2(32'hbad1600f),
	.w3(32'h3d14bcad),
	.w4(32'hbc365150),
	.w5(32'h3b4962c4),
	.w6(32'h3d1e241e),
	.w7(32'h3d159475),
	.w8(32'hba75a0d9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb326f2),
	.w1(32'h3a8ad0bb),
	.w2(32'hbbad529c),
	.w3(32'hbb00a6e6),
	.w4(32'hbbb8e94d),
	.w5(32'hbad7e04f),
	.w6(32'hbb2356d4),
	.w7(32'h3b1bcb3a),
	.w8(32'h3a9767ab),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18c2b8),
	.w1(32'hbbf9f12f),
	.w2(32'h3ca0cfe6),
	.w3(32'h3b8fdbfd),
	.w4(32'hbaa3fa0f),
	.w5(32'h3c406acc),
	.w6(32'hbbc94e87),
	.w7(32'hbb85b784),
	.w8(32'h3c1d4ebd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafdf77),
	.w1(32'h3c264e3f),
	.w2(32'h3a9d879e),
	.w3(32'h3d179f6e),
	.w4(32'h3d037c89),
	.w5(32'h3b00e363),
	.w6(32'h3c8452f5),
	.w7(32'h3c936109),
	.w8(32'h3aa02cf0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7e96d),
	.w1(32'hbbc33121),
	.w2(32'hbbcbfbf0),
	.w3(32'hbb992b95),
	.w4(32'h3951ee02),
	.w5(32'hbc4613a8),
	.w6(32'hbbeaf86f),
	.w7(32'hba90a9e6),
	.w8(32'hbb177f1d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e3c7),
	.w1(32'hbc48e4ae),
	.w2(32'hbbd41f4e),
	.w3(32'hbc132fb0),
	.w4(32'hbc3a25e2),
	.w5(32'h3b296c14),
	.w6(32'hbcafed00),
	.w7(32'hbc4af924),
	.w8(32'h39cdf1ed),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba86f92),
	.w1(32'hbbc18885),
	.w2(32'hbb9f936f),
	.w3(32'h3ab45636),
	.w4(32'hbc5af416),
	.w5(32'hbc258a4e),
	.w6(32'h3c1fabda),
	.w7(32'h3c270a96),
	.w8(32'hbb4110c9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8173d),
	.w1(32'h3bd57b54),
	.w2(32'hbbe98c51),
	.w3(32'h3c0f7333),
	.w4(32'h3c62c8c3),
	.w5(32'hbc3f6d7b),
	.w6(32'hbc76767f),
	.w7(32'h3bb3ca7e),
	.w8(32'hbc81031c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a7e5f),
	.w1(32'hbbf9dfb4),
	.w2(32'hbbacae19),
	.w3(32'hbc4ab7ad),
	.w4(32'hbc4f6173),
	.w5(32'hbc4ce4df),
	.w6(32'hbd18669d),
	.w7(32'hbc8d63a4),
	.w8(32'hb998c7a4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2a2bc),
	.w1(32'hbc38f494),
	.w2(32'h3be3f844),
	.w3(32'hbb9b9f5a),
	.w4(32'hbc050bc2),
	.w5(32'h3cdc1c2f),
	.w6(32'hbbebb7c6),
	.w7(32'hbc179a86),
	.w8(32'h3bfe9c67),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eeb2d),
	.w1(32'hbccc07d6),
	.w2(32'h39234a7d),
	.w3(32'h3c713de5),
	.w4(32'hbbd3670e),
	.w5(32'h3bca5f76),
	.w6(32'h3cca3920),
	.w7(32'h3ccc6f22),
	.w8(32'h3b16bb3d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa6ec3),
	.w1(32'hbbbc0e66),
	.w2(32'hbc04258e),
	.w3(32'h3c013e6c),
	.w4(32'hbb0839fb),
	.w5(32'hbc9e7f12),
	.w6(32'hba305c9e),
	.w7(32'h398b888c),
	.w8(32'hbc4dbe03),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d633e),
	.w1(32'hbca9f423),
	.w2(32'hbba41e56),
	.w3(32'hbc36baf6),
	.w4(32'hbb406cd7),
	.w5(32'hbb6b9bdd),
	.w6(32'hbc96e756),
	.w7(32'h3b21c04b),
	.w8(32'h3b286984),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb7c54),
	.w1(32'h3afed7bd),
	.w2(32'hbc5aa1a1),
	.w3(32'h3c1aed8b),
	.w4(32'h3ba74757),
	.w5(32'hbc116774),
	.w6(32'h3b7aa619),
	.w7(32'hb9cbb678),
	.w8(32'h3b99df50),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c0984),
	.w1(32'hbc322a95),
	.w2(32'hbc2511ec),
	.w3(32'hbcd29fb0),
	.w4(32'hbc9f1af7),
	.w5(32'hbc2d1e83),
	.w6(32'hbaa328b4),
	.w7(32'hbc325419),
	.w8(32'h3c6f7186),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5602f),
	.w1(32'hbca3604d),
	.w2(32'h3b2979b9),
	.w3(32'hbcc64047),
	.w4(32'hbc9176ea),
	.w5(32'h3c8b96fe),
	.w6(32'h3c621c52),
	.w7(32'hbc25da51),
	.w8(32'hbbec7e48),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82888a),
	.w1(32'hbb4b05fa),
	.w2(32'hbc30ffed),
	.w3(32'h3c64fdd8),
	.w4(32'h3b0a6e32),
	.w5(32'hbc488d69),
	.w6(32'h3c9e3b4b),
	.w7(32'h3c827503),
	.w8(32'h39e9c286),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74ed00),
	.w1(32'hbb699d25),
	.w2(32'hbb0b8b75),
	.w3(32'hbc1ceb80),
	.w4(32'hbbe8ea09),
	.w5(32'hbb8b45e4),
	.w6(32'hbcad38c7),
	.w7(32'hbc49e371),
	.w8(32'h3b37e0b1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba10af3),
	.w1(32'h3bff9cdb),
	.w2(32'h38e0d1fc),
	.w3(32'hbb0ae86e),
	.w4(32'hbb0513a5),
	.w5(32'hbafe649b),
	.w6(32'h3b9fea55),
	.w7(32'h3bb4d7e7),
	.w8(32'h389f7b58),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5169d9),
	.w1(32'h3b7d994c),
	.w2(32'hbbc71147),
	.w3(32'hbae7a747),
	.w4(32'h3ad116df),
	.w5(32'hbba50ede),
	.w6(32'hbb35e3ca),
	.w7(32'h3a49ea91),
	.w8(32'hbc33f332),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f47b1),
	.w1(32'hbcbd4aec),
	.w2(32'h3be986d0),
	.w3(32'hbc1c5857),
	.w4(32'hbcc6c21d),
	.w5(32'h3bf3d55e),
	.w6(32'hbb896dce),
	.w7(32'hbb916f19),
	.w8(32'hbbd8cfa5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c055441),
	.w1(32'h3bd0c634),
	.w2(32'h3c7f38ad),
	.w3(32'h3c972283),
	.w4(32'h3c4c4ce3),
	.w5(32'h3cd3f526),
	.w6(32'h3bd47fa9),
	.w7(32'h3c885e97),
	.w8(32'hbae0aba7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7344e8),
	.w1(32'hbae14ab8),
	.w2(32'h3b918358),
	.w3(32'h3d0d6391),
	.w4(32'h392a0512),
	.w5(32'hbbd94ed3),
	.w6(32'h3c6d60d0),
	.w7(32'h3c4dc993),
	.w8(32'hbb78f21b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb239619),
	.w1(32'h3b6dabcf),
	.w2(32'hba7037c0),
	.w3(32'h3a5a8bcd),
	.w4(32'hba7ddb7e),
	.w5(32'h3c356b85),
	.w6(32'hbc7e7407),
	.w7(32'hbc03defa),
	.w8(32'hbb5e0f97),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb052711),
	.w1(32'hbaff65de),
	.w2(32'h3a1b582d),
	.w3(32'h3c85f58d),
	.w4(32'h3caa4875),
	.w5(32'h3c4701b8),
	.w6(32'hbbd97f0f),
	.w7(32'hbbd3b4b6),
	.w8(32'hbb727786),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88ef19),
	.w1(32'h3c533f37),
	.w2(32'hbc2d4fa0),
	.w3(32'h3b1fe603),
	.w4(32'h3bb55eba),
	.w5(32'hbc13aaee),
	.w6(32'h3b3b2835),
	.w7(32'h3bb06578),
	.w8(32'h3a05888a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45991b),
	.w1(32'hbb5902ef),
	.w2(32'hb94e9010),
	.w3(32'hbca4a1a0),
	.w4(32'hbc4b9fb7),
	.w5(32'h3904a723),
	.w6(32'hbc099da7),
	.w7(32'hbc399149),
	.w8(32'h3bf21737),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba884ef3),
	.w1(32'hb994f265),
	.w2(32'h3c26e698),
	.w3(32'hba71df0a),
	.w4(32'h3bdefc06),
	.w5(32'h3a9d8e1b),
	.w6(32'hb802cdb3),
	.w7(32'h3b6ad3f7),
	.w8(32'h3c077aa4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaf9dd),
	.w1(32'h3a33e73e),
	.w2(32'hbb089676),
	.w3(32'h3c4eea7a),
	.w4(32'h3bff2d7d),
	.w5(32'hbb95aa17),
	.w6(32'h3bfb59cc),
	.w7(32'h3bc848d2),
	.w8(32'hbb563a21),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c338e34),
	.w1(32'h3b977b7a),
	.w2(32'hbb9d14bf),
	.w3(32'h3bdd9bbc),
	.w4(32'h3c5b1623),
	.w5(32'hbba8f26c),
	.w6(32'h3bf62d35),
	.w7(32'h3c202557),
	.w8(32'hbb6eb2f0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa66be1),
	.w1(32'hbb44f96d),
	.w2(32'hbb1b4615),
	.w3(32'h3b64b310),
	.w4(32'h3a9307cd),
	.w5(32'h3c2826d5),
	.w6(32'h3bbd807b),
	.w7(32'h3a8466bc),
	.w8(32'hbc0968e6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8038eb),
	.w1(32'hbcdee7d0),
	.w2(32'hbc4fea4a),
	.w3(32'hba538794),
	.w4(32'hbcbf7913),
	.w5(32'h3bc0dc39),
	.w6(32'h3a4f3631),
	.w7(32'hbc0990d8),
	.w8(32'h3ca8ef1e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e992a),
	.w1(32'h3c92441a),
	.w2(32'h3abbcaf8),
	.w3(32'hbc743bfa),
	.w4(32'hbc0c7db6),
	.w5(32'h3b704ca7),
	.w6(32'h3bc39ece),
	.w7(32'hbbdcee03),
	.w8(32'h3a038a1e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ace11),
	.w1(32'h3b7b6172),
	.w2(32'hbbbd5a52),
	.w3(32'h399d6201),
	.w4(32'h3b5b66db),
	.w5(32'h3ba8fd55),
	.w6(32'hbb3b4a91),
	.w7(32'hb935afb9),
	.w8(32'h3a0767e6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c56d7),
	.w1(32'hbc22a59c),
	.w2(32'h3b81eab6),
	.w3(32'h3b905d56),
	.w4(32'hbbbb1184),
	.w5(32'h3bfbf76a),
	.w6(32'hba223de4),
	.w7(32'h372d8496),
	.w8(32'h3b555daf),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3324a8),
	.w1(32'hbbeee1ed),
	.w2(32'h3ba29ba4),
	.w3(32'h3a81866f),
	.w4(32'hba8a42cc),
	.w5(32'h3bbd0713),
	.w6(32'hba89983c),
	.w7(32'hbac01b00),
	.w8(32'h3aba9153),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0086bb),
	.w1(32'hbb19e9e3),
	.w2(32'h3bb6543a),
	.w3(32'h3c40f541),
	.w4(32'h3be0edfa),
	.w5(32'h3c16dec3),
	.w6(32'hb95f35d4),
	.w7(32'hba23e90f),
	.w8(32'h3be7098b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff9c40),
	.w1(32'hbb25e400),
	.w2(32'h3b608360),
	.w3(32'h3ba41e98),
	.w4(32'h3bd3b00a),
	.w5(32'h3b0c256b),
	.w6(32'h3b80163e),
	.w7(32'h3bfb6593),
	.w8(32'h3bbbcd9c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2219),
	.w1(32'hbbe817a0),
	.w2(32'hbce21ac5),
	.w3(32'hbc3cd71b),
	.w4(32'hbb3410f3),
	.w5(32'hbc58bd4f),
	.w6(32'hbc820a1b),
	.w7(32'h3b31b2c3),
	.w8(32'h3c2ad8d5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb69c8d),
	.w1(32'hbc0fd7ca),
	.w2(32'hbb760712),
	.w3(32'hbccf54f7),
	.w4(32'hbca73314),
	.w5(32'hbc1273f4),
	.w6(32'hbc66d4fc),
	.w7(32'hbcadca21),
	.w8(32'h39bb2864),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da23a),
	.w1(32'h3ab60255),
	.w2(32'h3a698b59),
	.w3(32'hbc1f25c7),
	.w4(32'hbbe95c3b),
	.w5(32'h3b2eaead),
	.w6(32'hbb40b442),
	.w7(32'h3b1b15aa),
	.w8(32'hbbe65dee),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb217e1c),
	.w1(32'hbb813101),
	.w2(32'hbc3396a7),
	.w3(32'h3bb77e6a),
	.w4(32'h3b4e98bf),
	.w5(32'hbc1efe89),
	.w6(32'hbb7c4b4e),
	.w7(32'h3b5d1d46),
	.w8(32'hbbf0407d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d7d0d),
	.w1(32'h3b826a7d),
	.w2(32'hbb944ce3),
	.w3(32'hbc2db796),
	.w4(32'hbb2e67db),
	.w5(32'hbb470104),
	.w6(32'hbc2797b9),
	.w7(32'hbad4438f),
	.w8(32'hbbd13b28),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b447ff),
	.w1(32'hbc13aee9),
	.w2(32'h3cd394d2),
	.w3(32'hbba5a344),
	.w4(32'hbc4513e8),
	.w5(32'h3cc16e9e),
	.w6(32'hbaa34cfb),
	.w7(32'hbc15be66),
	.w8(32'h3c1546bc),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce65513),
	.w1(32'hbbc39213),
	.w2(32'h3c3f756b),
	.w3(32'h3d4bc6f8),
	.w4(32'h3d14a437),
	.w5(32'hba357e73),
	.w6(32'h3c8648dc),
	.w7(32'h3ca594ff),
	.w8(32'hbab1c620),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7c2b4),
	.w1(32'hb9fe98ae),
	.w2(32'hbbcce458),
	.w3(32'h3baea7de),
	.w4(32'h3c0e39d0),
	.w5(32'hbb214f5b),
	.w6(32'hbc57b0c7),
	.w7(32'hbb393b15),
	.w8(32'hbc0b1d20),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba369cb5),
	.w1(32'h3c6626db),
	.w2(32'hbc587b12),
	.w3(32'hba620633),
	.w4(32'h3b3fd776),
	.w5(32'hbc020d91),
	.w6(32'hb925a257),
	.w7(32'h3b93673c),
	.w8(32'hbac42229),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c6276),
	.w1(32'h3b9aea73),
	.w2(32'hbb24b23e),
	.w3(32'hbc643534),
	.w4(32'h3a6c2101),
	.w5(32'h3b4b0017),
	.w6(32'hbbdc654d),
	.w7(32'hbba63814),
	.w8(32'hbbccb8b1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c1848),
	.w1(32'hba951afd),
	.w2(32'hbb86db30),
	.w3(32'hba4109d5),
	.w4(32'hbb30d014),
	.w5(32'hba8e8563),
	.w6(32'hbba4feba),
	.w7(32'hbb47512e),
	.w8(32'h3aa68741),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b086a52),
	.w1(32'h3b47e4b5),
	.w2(32'h3baec142),
	.w3(32'h3c75a894),
	.w4(32'h3b067858),
	.w5(32'h3c9eecbf),
	.w6(32'h3ac761be),
	.w7(32'h3bbb24dc),
	.w8(32'h3c3db98d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b362c4e),
	.w1(32'hbc4773ed),
	.w2(32'hbc47ea41),
	.w3(32'h3c975a0b),
	.w4(32'h3c8316c0),
	.w5(32'h3ba7ce1f),
	.w6(32'h3c8b731b),
	.w7(32'h3c24f850),
	.w8(32'h3c83ef1c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb497a71),
	.w1(32'hba41e61e),
	.w2(32'h3b5ab845),
	.w3(32'hbba7ca64),
	.w4(32'hbb9234c5),
	.w5(32'h3be1dcc9),
	.w6(32'h3c7217c4),
	.w7(32'h3ad4ad84),
	.w8(32'h3b55928d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93c591),
	.w1(32'h3bbd3e81),
	.w2(32'hbc2caaa2),
	.w3(32'hbc28694b),
	.w4(32'hbc0187ea),
	.w5(32'hbc7afd82),
	.w6(32'hbb58e204),
	.w7(32'h39d27a77),
	.w8(32'hbc283d3f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ed96d),
	.w1(32'hbb8f7f81),
	.w2(32'hbb8172d4),
	.w3(32'hbc243d29),
	.w4(32'hbbfda71d),
	.w5(32'hbbc60e15),
	.w6(32'hbc4c3e57),
	.w7(32'hbbf43283),
	.w8(32'hbc08c888),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba735195),
	.w1(32'hbb8771fd),
	.w2(32'hbc18cb3c),
	.w3(32'h3c4d2145),
	.w4(32'h3c03930c),
	.w5(32'h3b16375b),
	.w6(32'h3c522c3a),
	.w7(32'h3c3acba0),
	.w8(32'h3c0bd5f4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d0af0),
	.w1(32'h3c05ab74),
	.w2(32'hbaa8d7ba),
	.w3(32'h3c424c46),
	.w4(32'h3c2bb3af),
	.w5(32'hbc0a0d5e),
	.w6(32'h3c38be4d),
	.w7(32'h3b517a50),
	.w8(32'hbbf45f03),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8262c2),
	.w1(32'hba5be2fc),
	.w2(32'h3b166e7e),
	.w3(32'hbc834cb9),
	.w4(32'h3af1f4cd),
	.w5(32'h3c487e53),
	.w6(32'hbc6dbd60),
	.w7(32'h3b651b3e),
	.w8(32'h3c5d5c2e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19e650),
	.w1(32'hbc401082),
	.w2(32'hba49f235),
	.w3(32'h3c39e0f2),
	.w4(32'h3be030ac),
	.w5(32'hbbda594f),
	.w6(32'h3c124d1a),
	.w7(32'h3b8c0c77),
	.w8(32'hbab63b58),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7477e0),
	.w1(32'h3c1013ab),
	.w2(32'hbc2be297),
	.w3(32'h3ae801ff),
	.w4(32'h3c162c13),
	.w5(32'hbb9ad0e9),
	.w6(32'hbc82e364),
	.w7(32'hbb90c1bc),
	.w8(32'hbb996493),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b4deb),
	.w1(32'hbc350ad5),
	.w2(32'hbb8b14ff),
	.w3(32'hb8e0a5dc),
	.w4(32'hb9051631),
	.w5(32'hbc641276),
	.w6(32'h3bba4e2f),
	.w7(32'h3c179834),
	.w8(32'hbc8f5d23),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb888fc8),
	.w1(32'hbbb2323a),
	.w2(32'h399ac43c),
	.w3(32'hbc01e31d),
	.w4(32'hbad8d884),
	.w5(32'hbcae6ef2),
	.w6(32'hbc65aadc),
	.w7(32'hbc49fbd9),
	.w8(32'hbc1872ca),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbdd18),
	.w1(32'h3bc2a961),
	.w2(32'h3bde524d),
	.w3(32'h3ca647ef),
	.w4(32'h3ce18841),
	.w5(32'h3c3a4506),
	.w6(32'h3c399e3f),
	.w7(32'h3cc368b2),
	.w8(32'hbb91fa2e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5df3ce),
	.w1(32'h3b125e2d),
	.w2(32'hbb921054),
	.w3(32'h3b5d414b),
	.w4(32'h3bd2e630),
	.w5(32'hbc190b88),
	.w6(32'hbc0cd2c7),
	.w7(32'hbbbcc52d),
	.w8(32'hbc3e3753),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb323087),
	.w1(32'hbb45112e),
	.w2(32'hbc2ff384),
	.w3(32'h3b8e1160),
	.w4(32'h3c426b03),
	.w5(32'hbb7c7733),
	.w6(32'hbaba7808),
	.w7(32'h3c6f5ebe),
	.w8(32'hbc28fac4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ec0d3),
	.w1(32'h3af4c139),
	.w2(32'hbbbe54e8),
	.w3(32'hbb99cc57),
	.w4(32'hbbc173dc),
	.w5(32'hbc24e71b),
	.w6(32'h39d6efad),
	.w7(32'hba8d1b76),
	.w8(32'hbc268673),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37b34d),
	.w1(32'hba380c4d),
	.w2(32'hbcae6bea),
	.w3(32'hbc8a0ace),
	.w4(32'hbbb778a0),
	.w5(32'hbc0513db),
	.w6(32'hbca2f840),
	.w7(32'hbc3fe215),
	.w8(32'h3b5a6baf),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1dd92),
	.w1(32'hbc001186),
	.w2(32'hbc5f16b6),
	.w3(32'hbc4fb7e2),
	.w4(32'hbc39eba2),
	.w5(32'hbbb479a8),
	.w6(32'h39fc876d),
	.w7(32'h3a5e8c9d),
	.w8(32'h3a25f00a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f01de),
	.w1(32'hbb3c3d6e),
	.w2(32'hbb8e2ee3),
	.w3(32'hbc84ed5a),
	.w4(32'hbc05e299),
	.w5(32'hbc83ee7c),
	.w6(32'hbbc54acd),
	.w7(32'hbbf78192),
	.w8(32'hbc77487c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbd6a0),
	.w1(32'hbc46cf49),
	.w2(32'h3b80708a),
	.w3(32'hbbe67da5),
	.w4(32'hbb50d698),
	.w5(32'hbc2e42c4),
	.w6(32'hbc79e631),
	.w7(32'hbc368b57),
	.w8(32'hbc38da10),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62278c),
	.w1(32'hbbcbe498),
	.w2(32'h3af5bfa8),
	.w3(32'h3ba9fe99),
	.w4(32'hbbd27c69),
	.w5(32'h3b671f77),
	.w6(32'hbc85b0b5),
	.w7(32'h3b924a88),
	.w8(32'h3b394dca),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f75f),
	.w1(32'hbc4e17bf),
	.w2(32'h3c86e56d),
	.w3(32'h3c617c2c),
	.w4(32'hba475469),
	.w5(32'hbbe73e22),
	.w6(32'h3bca8097),
	.w7(32'h3bd2916b),
	.w8(32'h3ad4627b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca09ff9),
	.w1(32'h38e4d6f3),
	.w2(32'hbc17e633),
	.w3(32'h3cfe22e6),
	.w4(32'h3c97542f),
	.w5(32'hbbe63052),
	.w6(32'hbbab16ae),
	.w7(32'h3c3a13cd),
	.w8(32'hbc0b4dc9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6c777),
	.w1(32'hbb30c1f6),
	.w2(32'h3c3c9426),
	.w3(32'h3a970ed3),
	.w4(32'h39ecd36b),
	.w5(32'hba4d385f),
	.w6(32'hbc5dde16),
	.w7(32'hbbf131c4),
	.w8(32'hbc8dff6a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1062ad),
	.w1(32'hbb9aeaa6),
	.w2(32'h3bb0dba5),
	.w3(32'h3b846342),
	.w4(32'hbc448855),
	.w5(32'h3cbc25f6),
	.w6(32'h3b7436f5),
	.w7(32'h3ac83811),
	.w8(32'h3c374b85),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a21cd),
	.w1(32'hbabb1380),
	.w2(32'h3c56d2be),
	.w3(32'h3cd13afc),
	.w4(32'h3be40ad3),
	.w5(32'h3c568427),
	.w6(32'h3c3275d1),
	.w7(32'h3cb3e917),
	.w8(32'hbc81534d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78d407),
	.w1(32'hba08d401),
	.w2(32'h37958e50),
	.w3(32'h3d1937d6),
	.w4(32'h3d1a5c2b),
	.w5(32'hbbfffa01),
	.w6(32'h3ba0f071),
	.w7(32'h3ce0447a),
	.w8(32'hbc39d6cf),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae3efe),
	.w1(32'hbb8d2411),
	.w2(32'h3c102015),
	.w3(32'h3b019c85),
	.w4(32'hbb5b23bf),
	.w5(32'h3c42729e),
	.w6(32'hbbda7de0),
	.w7(32'hbbc5a249),
	.w8(32'h3c64cebc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c640f19),
	.w1(32'h3c9379d3),
	.w2(32'hbb87e574),
	.w3(32'hb71acbcf),
	.w4(32'h3ba8d018),
	.w5(32'hbba98cbf),
	.w6(32'h3ae1b742),
	.w7(32'hbbc7eb60),
	.w8(32'hbc5427ce),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb017694),
	.w1(32'hbbb2740d),
	.w2(32'h3bc04312),
	.w3(32'h3b474ebe),
	.w4(32'h3b128e01),
	.w5(32'hbb06a3a4),
	.w6(32'hbc386242),
	.w7(32'hbbceaa01),
	.w8(32'hbb4b1e40),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a37c22),
	.w1(32'hbb1fbd32),
	.w2(32'h3b2f495a),
	.w3(32'h3ba3ae96),
	.w4(32'h39c969ef),
	.w5(32'h3a40406f),
	.w6(32'hbba6ab69),
	.w7(32'hba30188d),
	.w8(32'hbc4bc6a5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2daaa),
	.w1(32'h3b2e6a85),
	.w2(32'h3af8e2ad),
	.w3(32'h3a5b52f2),
	.w4(32'h3ba3df6a),
	.w5(32'h39a39122),
	.w6(32'hbc59ca5e),
	.w7(32'h3b078e5e),
	.w8(32'hbb686b88),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cd3d0),
	.w1(32'h3c0b3fa6),
	.w2(32'hbb5d05b1),
	.w3(32'h3be09571),
	.w4(32'h3bcd2df9),
	.w5(32'hbb63fc84),
	.w6(32'hbb74ab09),
	.w7(32'h3bb8fb66),
	.w8(32'hbb7cd2ca),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc370bdb),
	.w1(32'hbbae2b02),
	.w2(32'h39e49af4),
	.w3(32'hbc0835a1),
	.w4(32'hbb95f8a3),
	.w5(32'h3a89e385),
	.w6(32'hbbb3b1c8),
	.w7(32'hbbe9636d),
	.w8(32'h3b1292f6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadb34e),
	.w1(32'h3b6ea5d6),
	.w2(32'hbc3508e5),
	.w3(32'h39e83289),
	.w4(32'hbb579d36),
	.w5(32'h3b7c7e26),
	.w6(32'hbb1af221),
	.w7(32'hbbe1928c),
	.w8(32'h3bcb95cc),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b4ee6),
	.w1(32'h3b7be101),
	.w2(32'h395edfd4),
	.w3(32'hbc60e6a8),
	.w4(32'hbabda669),
	.w5(32'hbaa9a6aa),
	.w6(32'hbb07f9f8),
	.w7(32'hbc8e8a9f),
	.w8(32'hbb804ed2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bf813),
	.w1(32'h3aaf40e4),
	.w2(32'h3bfc1460),
	.w3(32'hbb561e65),
	.w4(32'hbba16985),
	.w5(32'h3962fcf5),
	.w6(32'hbab9f50d),
	.w7(32'hba4802b5),
	.w8(32'hbb7b7c38),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf46c7),
	.w1(32'hba8a2cde),
	.w2(32'h3c098a13),
	.w3(32'h3c12c430),
	.w4(32'hbbb9fdf1),
	.w5(32'h3bdbf21a),
	.w6(32'h3c0552d9),
	.w7(32'h3bd756d1),
	.w8(32'h3bab23e7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24843a),
	.w1(32'hbbc3449b),
	.w2(32'h3b94dd17),
	.w3(32'h3bdda73c),
	.w4(32'h3a419ac0),
	.w5(32'hba3bd8b0),
	.w6(32'h3985f487),
	.w7(32'h3c059c8b),
	.w8(32'h398fb96d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54a4dc),
	.w1(32'hbbb8d99c),
	.w2(32'hbb90e090),
	.w3(32'h3a846cc6),
	.w4(32'hbb13e658),
	.w5(32'h3b3f2f0e),
	.w6(32'hbbbe2c82),
	.w7(32'h3c21b6ba),
	.w8(32'hbbf1e53e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc092fbf),
	.w1(32'h3bcbe70e),
	.w2(32'h3bb0f389),
	.w3(32'h3c0913fd),
	.w4(32'h3a92cdce),
	.w5(32'h3ac72f57),
	.w6(32'h3b86fc6b),
	.w7(32'h3c47b93c),
	.w8(32'hbc7d1a9d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcea6e4),
	.w1(32'hbbb39eed),
	.w2(32'h3a321351),
	.w3(32'h3d04e74c),
	.w4(32'h3bf50150),
	.w5(32'h3c22485b),
	.w6(32'h3be89d48),
	.w7(32'h3c2c5788),
	.w8(32'h3c36bc9e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba8a21),
	.w1(32'h3c420b99),
	.w2(32'hbad68558),
	.w3(32'hbc2c0113),
	.w4(32'hbb7121e0),
	.w5(32'hbbbabc9b),
	.w6(32'h3c0b384b),
	.w7(32'hbb09f27c),
	.w8(32'h3b4a0f78),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6657e2),
	.w1(32'h3b884235),
	.w2(32'h3bc92d33),
	.w3(32'h3b5d19ae),
	.w4(32'h3b77330f),
	.w5(32'h3c3bce8d),
	.w6(32'hbc2e96b6),
	.w7(32'hbba3a5a3),
	.w8(32'hbc21daae),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbef212),
	.w1(32'hbb491dd1),
	.w2(32'h3bc1ec76),
	.w3(32'h3cab1413),
	.w4(32'h3c9a4932),
	.w5(32'h3c4374bc),
	.w6(32'h3a45bf2e),
	.w7(32'h3c1dacc7),
	.w8(32'h3bc61686),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5642c),
	.w1(32'hbc39e816),
	.w2(32'hbbaf11c5),
	.w3(32'h3d17614d),
	.w4(32'hbb56f896),
	.w5(32'hbae19749),
	.w6(32'h3d04f229),
	.w7(32'h3cd08fae),
	.w8(32'hbc110ede),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2319),
	.w1(32'hbacfaa30),
	.w2(32'h3c2d4290),
	.w3(32'hbbf3be72),
	.w4(32'h3b025bca),
	.w5(32'hbc3e28a3),
	.w6(32'hbc12bdff),
	.w7(32'h3b59e342),
	.w8(32'hbbb8ce3e),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b823091),
	.w1(32'hbb99dc69),
	.w2(32'hbcb4cbb2),
	.w3(32'h3b8ab926),
	.w4(32'h3b724fa3),
	.w5(32'hbc6f40b7),
	.w6(32'hbc3baa66),
	.w7(32'hbb11af27),
	.w8(32'h3c772c99),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc998201),
	.w1(32'h3b50d646),
	.w2(32'h3c30520d),
	.w3(32'hbd2586cb),
	.w4(32'hbbc56c1e),
	.w5(32'h3bf47196),
	.w6(32'hbc1b19af),
	.w7(32'hbc9f9e53),
	.w8(32'h3c4011cf),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6609d),
	.w1(32'h3cb0b2af),
	.w2(32'hbb21ab8e),
	.w3(32'h3b0f2742),
	.w4(32'h3cb1d8b4),
	.w5(32'hbb5d1a19),
	.w6(32'h3b1613c7),
	.w7(32'h3c751514),
	.w8(32'hbb339abb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6745be),
	.w1(32'h3c17bedd),
	.w2(32'hbad78ca0),
	.w3(32'h3b8e49fa),
	.w4(32'h3ba136b8),
	.w5(32'h3c1cd935),
	.w6(32'h3b369388),
	.w7(32'h3bc4ec9d),
	.w8(32'hbaec6cf0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac836c),
	.w1(32'h3c11e43d),
	.w2(32'h3b16dfcf),
	.w3(32'h3cabbd10),
	.w4(32'h3c4f081b),
	.w5(32'hba995165),
	.w6(32'hbae1ce91),
	.w7(32'h3c1a3c99),
	.w8(32'hbbcfe2cd),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa15b09),
	.w1(32'hbaa30780),
	.w2(32'h3bafc843),
	.w3(32'hb90619bf),
	.w4(32'hbb4b00c1),
	.w5(32'h3c07418f),
	.w6(32'hbb8e4208),
	.w7(32'hbb364e34),
	.w8(32'h3c12be85),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c90c7),
	.w1(32'h3b95fbc9),
	.w2(32'hbc354d5b),
	.w3(32'h3b3078f6),
	.w4(32'hb888233d),
	.w5(32'hbc2eb2f2),
	.w6(32'h3bbe7400),
	.w7(32'h3b967f9c),
	.w8(32'h3b4e796d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc822874),
	.w1(32'h3ba35fbb),
	.w2(32'hbbe6db6e),
	.w3(32'hbc9990f6),
	.w4(32'hbc96acc5),
	.w5(32'hbb6d9a3a),
	.w6(32'h3bfd9a41),
	.w7(32'hbb259986),
	.w8(32'hbc4a6099),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36cfde),
	.w1(32'hbc9211ee),
	.w2(32'hbaad4d08),
	.w3(32'hb8fc63d8),
	.w4(32'hbbb42f87),
	.w5(32'hbabcb415),
	.w6(32'hbb7b64ff),
	.w7(32'h3b800ef2),
	.w8(32'hbb4dae9f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae2bc0),
	.w1(32'h3bf65328),
	.w2(32'hbb7239df),
	.w3(32'h3a94e20d),
	.w4(32'h394bd5d2),
	.w5(32'hbb174f35),
	.w6(32'h3a3bbd0b),
	.w7(32'h3b296c66),
	.w8(32'h3bac7610),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bb1c8),
	.w1(32'hbb8ac586),
	.w2(32'hbaf14e1f),
	.w3(32'hbbc3e54d),
	.w4(32'hbb933306),
	.w5(32'h3ad1ae20),
	.w6(32'h3c2b2fd9),
	.w7(32'hbb25f249),
	.w8(32'hbab562b8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39838d3d),
	.w1(32'h3b1b5660),
	.w2(32'hbb38e7ee),
	.w3(32'h3af7692a),
	.w4(32'h3ac0637b),
	.w5(32'hbc528190),
	.w6(32'hbb0968f2),
	.w7(32'h3b9fea5a),
	.w8(32'h3c1bb2e4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd04b3b1),
	.w1(32'hbc5780fe),
	.w2(32'hbc1ca855),
	.w3(32'hbd18f3d1),
	.w4(32'hbd015d65),
	.w5(32'hbc2eb884),
	.w6(32'hbcdd6f53),
	.w7(32'hbcc6cad6),
	.w8(32'hbb832d0d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa4f0d),
	.w1(32'hba860308),
	.w2(32'hba94ac4f),
	.w3(32'hba013775),
	.w4(32'hbb89b504),
	.w5(32'hbab5962e),
	.w6(32'hbb597992),
	.w7(32'hbbc5c712),
	.w8(32'h3a0769b0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fd9ec),
	.w1(32'hbb241c90),
	.w2(32'h3c021ace),
	.w3(32'hbb0910a4),
	.w4(32'h3b508ba9),
	.w5(32'h3b287697),
	.w6(32'hbc8e148f),
	.w7(32'hbc02a806),
	.w8(32'hbcad5ae5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89a34a),
	.w1(32'hb9304458),
	.w2(32'h3aee9909),
	.w3(32'h3cb970dd),
	.w4(32'h3c8c814f),
	.w5(32'hbbe125c1),
	.w6(32'hbb877d12),
	.w7(32'h3b124c96),
	.w8(32'hbb918f7f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc135d14),
	.w1(32'hbb2943e7),
	.w2(32'hba9db0a9),
	.w3(32'hbc1d3b3c),
	.w4(32'hbb8bab0e),
	.w5(32'h3be4ec48),
	.w6(32'hbb89abb8),
	.w7(32'h3b0c7d62),
	.w8(32'h3c48ca95),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39929a),
	.w1(32'h3ab2a864),
	.w2(32'hbbd1242b),
	.w3(32'h3bf26231),
	.w4(32'h3b95fb5f),
	.w5(32'hbc8f65c8),
	.w6(32'h3bb4462f),
	.w7(32'hb8ae0f12),
	.w8(32'hbb4df807),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdba19e),
	.w1(32'h3c90fbe6),
	.w2(32'h3c05931b),
	.w3(32'h3a3e0190),
	.w4(32'h3c3c1e26),
	.w5(32'h3bdfaee1),
	.w6(32'h3b3224e1),
	.w7(32'hbc11b63d),
	.w8(32'h3bf55d1e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c286f96),
	.w1(32'h3c282357),
	.w2(32'h3b475881),
	.w3(32'h3c42f5bf),
	.w4(32'h3be7d57f),
	.w5(32'h3b417a12),
	.w6(32'h3c2389bf),
	.w7(32'h3c50b483),
	.w8(32'h3b2690b0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b676c7c),
	.w1(32'h3b2e3cd9),
	.w2(32'h3b78302d),
	.w3(32'h3bc47f6b),
	.w4(32'h3be6544d),
	.w5(32'h3c496aee),
	.w6(32'h3b5deae2),
	.w7(32'h3bea4ca6),
	.w8(32'h3c1186f8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29d1b0),
	.w1(32'hba453079),
	.w2(32'hbb53ea8e),
	.w3(32'h3c0c71d2),
	.w4(32'hbb18ab6f),
	.w5(32'h3bd500cd),
	.w6(32'h3bf69364),
	.w7(32'h3b84bba5),
	.w8(32'h3bd4d612),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc6ea3),
	.w1(32'h3c6a4918),
	.w2(32'h3b714347),
	.w3(32'h3b013af1),
	.w4(32'hb6f21fa4),
	.w5(32'h3bc1407a),
	.w6(32'h39b9435c),
	.w7(32'hbbb621e1),
	.w8(32'h3b2830e9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a6916),
	.w1(32'hbb6f6ed6),
	.w2(32'hbbb1b6bf),
	.w3(32'hbb02b1d5),
	.w4(32'hbbd37e8d),
	.w5(32'h3b82b3bb),
	.w6(32'hba78de15),
	.w7(32'hbbc2a9c2),
	.w8(32'h3c4dea29),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba849f7a),
	.w1(32'hbaff0b43),
	.w2(32'h3c6f32fa),
	.w3(32'h3c94b990),
	.w4(32'h3c0299f3),
	.w5(32'h3bb7602a),
	.w6(32'h3c57f74b),
	.w7(32'hbb3de4a4),
	.w8(32'h39a3a848),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ab78a),
	.w1(32'h3ba98533),
	.w2(32'hbbf37791),
	.w3(32'h3c041b73),
	.w4(32'h3c5900c7),
	.w5(32'hbb9b1df9),
	.w6(32'h3c4868e4),
	.w7(32'h3c54885f),
	.w8(32'hbc0fb3fe),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8787c),
	.w1(32'hbb251019),
	.w2(32'hbc028684),
	.w3(32'hba9a3fc6),
	.w4(32'h3b585e48),
	.w5(32'hbc989526),
	.w6(32'hbb062e55),
	.w7(32'h3a889de6),
	.w8(32'hbcffa2a8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc584c0e),
	.w1(32'hbc820c81),
	.w2(32'hbbb9d618),
	.w3(32'hbd475252),
	.w4(32'hbc680e96),
	.w5(32'hbbcd8d4b),
	.w6(32'hbcf6fa02),
	.w7(32'hba81e971),
	.w8(32'hbbaa7496),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bb4c0),
	.w1(32'h3b701e46),
	.w2(32'hbb15b490),
	.w3(32'h3a9b8cff),
	.w4(32'h3c237438),
	.w5(32'hbbb26dc5),
	.w6(32'h3b887ec8),
	.w7(32'h3c19bc9d),
	.w8(32'hbbdb1112),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf64d8),
	.w1(32'hbabb635a),
	.w2(32'h3a52a417),
	.w3(32'h3c5013f6),
	.w4(32'h3960e365),
	.w5(32'h3bfbb26a),
	.w6(32'hbb98b949),
	.w7(32'hbc3b8dd2),
	.w8(32'h3ba2c3d9),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1734fb),
	.w1(32'h3af15138),
	.w2(32'hb8b46f19),
	.w3(32'h3bc22edf),
	.w4(32'h3c45aaaf),
	.w5(32'h3b93bfcf),
	.w6(32'h3bbd1484),
	.w7(32'h3c1788e3),
	.w8(32'hb9ca6094),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d56cc),
	.w1(32'h3b38c554),
	.w2(32'hbc75b1a6),
	.w3(32'h3cccbcb8),
	.w4(32'h3c940530),
	.w5(32'hbbc7a156),
	.w6(32'h3baa3530),
	.w7(32'h3b98bd51),
	.w8(32'h3ae860e4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44c8e8),
	.w1(32'hbc15bbee),
	.w2(32'hbba4fe2c),
	.w3(32'h3c8543c1),
	.w4(32'hbbccffcf),
	.w5(32'hbbadf2eb),
	.w6(32'h3cb3f036),
	.w7(32'h3c40eee8),
	.w8(32'hbb66aaad),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1cc29),
	.w1(32'hbc3397e4),
	.w2(32'h3b81637f),
	.w3(32'hbbaee7c4),
	.w4(32'hbc8113e2),
	.w5(32'hbbc4bc85),
	.w6(32'hbbce430d),
	.w7(32'hbc711a51),
	.w8(32'hbc0e32ad),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bb052),
	.w1(32'h3b97b257),
	.w2(32'hba49d300),
	.w3(32'h3bb547c7),
	.w4(32'h3bf1cc37),
	.w5(32'hbae1407c),
	.w6(32'hbb94f6f6),
	.w7(32'h3c0a4dc6),
	.w8(32'hbaade87f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb318de0),
	.w1(32'h3ab0db54),
	.w2(32'hbc1c1749),
	.w3(32'h3ba0357b),
	.w4(32'h3b9b930d),
	.w5(32'hbc60dcf2),
	.w6(32'h3c0e07fd),
	.w7(32'h3c342d32),
	.w8(32'hbc0716da),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402beb),
	.w1(32'h3a191a5c),
	.w2(32'hbc988a07),
	.w3(32'hbb1b8f1a),
	.w4(32'h3bd94ddc),
	.w5(32'hbcc7858a),
	.w6(32'hbab5dd7b),
	.w7(32'h3b82c564),
	.w8(32'hbc1b77b3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2528f1),
	.w1(32'hbc887f57),
	.w2(32'hbc0bf667),
	.w3(32'hbcff5286),
	.w4(32'hbc5b2bac),
	.w5(32'hbadfb73b),
	.w6(32'hbc3c00ba),
	.w7(32'h3b35bfec),
	.w8(32'h3bbdd35f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab1b3d),
	.w1(32'h3be1686c),
	.w2(32'hbcefbe8c),
	.w3(32'hbc825b9c),
	.w4(32'hbb455c14),
	.w5(32'hbce2294b),
	.w6(32'hbc255c40),
	.w7(32'hbc26bf1c),
	.w8(32'hbc332413),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab630f),
	.w1(32'h3b2f0bef),
	.w2(32'hbd0ab07c),
	.w3(32'hbc7c9ef8),
	.w4(32'h3c3d70d2),
	.w5(32'hbd271553),
	.w6(32'hbb827b64),
	.w7(32'h3cad1b3b),
	.w8(32'hbc941be8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccabc7a),
	.w1(32'h3b43d363),
	.w2(32'hba58c353),
	.w3(32'hbd16c0d6),
	.w4(32'h3c790972),
	.w5(32'hba3e2cb8),
	.w6(32'hbc160b99),
	.w7(32'h3c3123e6),
	.w8(32'h3b001b43),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0bdd4),
	.w1(32'h3b3a7460),
	.w2(32'h3c55ccf8),
	.w3(32'h3ba00422),
	.w4(32'h3c3018ef),
	.w5(32'h3bf08628),
	.w6(32'h3bf24b86),
	.w7(32'h3c554d5f),
	.w8(32'hbbda9213),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5c029),
	.w1(32'hbc4f7965),
	.w2(32'hbb83b219),
	.w3(32'h3b11b947),
	.w4(32'hbc44da8d),
	.w5(32'hbc123118),
	.w6(32'hbc08cfe9),
	.w7(32'hbbf88ce9),
	.w8(32'h3947b9b9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe68e03),
	.w1(32'h3a1da644),
	.w2(32'hbc9785ac),
	.w3(32'h3c0e3091),
	.w4(32'h3c4a183a),
	.w5(32'hbbb6fb03),
	.w6(32'h3c791813),
	.w7(32'h3c0f94bb),
	.w8(32'h3c258722),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeceec8),
	.w1(32'h3c7b2051),
	.w2(32'h3bb2b13f),
	.w3(32'h3cd5588f),
	.w4(32'h3cb190e7),
	.w5(32'h3a3e7ddb),
	.w6(32'h3cba1809),
	.w7(32'h3c1c3b30),
	.w8(32'h3bbfa7a0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2f9a6),
	.w1(32'h3a114776),
	.w2(32'hbbf76f26),
	.w3(32'h3c3c81b9),
	.w4(32'h3bba9a0e),
	.w5(32'hbbf20a05),
	.w6(32'h3c732410),
	.w7(32'h3bf63987),
	.w8(32'h38746298),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52de5f),
	.w1(32'h3c9195bc),
	.w2(32'h3a33250e),
	.w3(32'h3b8b4be6),
	.w4(32'h3c397fa0),
	.w5(32'h3c266adf),
	.w6(32'hbad033fa),
	.w7(32'hbbcfbc1e),
	.w8(32'h3c2bfcd8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59c02c),
	.w1(32'h3ca1e9fb),
	.w2(32'hbb96e61b),
	.w3(32'h3ccb9cdc),
	.w4(32'h3c37c9cf),
	.w5(32'hbbfdee21),
	.w6(32'h3b011461),
	.w7(32'hbb7ed176),
	.w8(32'h39941077),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1109ef),
	.w1(32'h3a6772f3),
	.w2(32'hbc429bde),
	.w3(32'hbc213b18),
	.w4(32'hbb84abb6),
	.w5(32'hbc9677fa),
	.w6(32'h3b67e5e2),
	.w7(32'hbb05a654),
	.w8(32'hbb8e53b7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c016b1d),
	.w1(32'h3bac1e4c),
	.w2(32'h3c3d533f),
	.w3(32'h3ba3a0a9),
	.w4(32'h3c9de579),
	.w5(32'h3b9986ca),
	.w6(32'h3c4104b2),
	.w7(32'h3cd12ce0),
	.w8(32'hbba8d3cd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5477),
	.w1(32'hbb8025ad),
	.w2(32'h3b84bf10),
	.w3(32'hbcb49524),
	.w4(32'hbc8287e1),
	.w5(32'h3ba96f4a),
	.w6(32'hbc59ac99),
	.w7(32'hbbcfcbf3),
	.w8(32'h3b6e49d1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bf008),
	.w1(32'h3a00885c),
	.w2(32'h3b2c46e2),
	.w3(32'h3ba8bf36),
	.w4(32'h3b3598d4),
	.w5(32'h3b0b2d43),
	.w6(32'h3b2eaf5b),
	.w7(32'hbb84d256),
	.w8(32'hbbf38e78),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced7909),
	.w1(32'hbc8ba40b),
	.w2(32'hbb6adea4),
	.w3(32'hbc14c101),
	.w4(32'hbaba678b),
	.w5(32'h3c4dabcb),
	.w6(32'h3c01da1e),
	.w7(32'h3d09eac1),
	.w8(32'h3cdbe461),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fa1b8),
	.w1(32'h3b78986f),
	.w2(32'hbc363073),
	.w3(32'h3c78d6b6),
	.w4(32'h3a29c963),
	.w5(32'hbc52c39b),
	.w6(32'h3c61d2ce),
	.w7(32'hbbc16c60),
	.w8(32'hbc00f296),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2cf986),
	.w1(32'hbc059451),
	.w2(32'h3b8ba305),
	.w3(32'hbc7a9ff4),
	.w4(32'hbbc8480e),
	.w5(32'h3bd43fd2),
	.w6(32'h3bbfddc8),
	.w7(32'h3c12d9c0),
	.w8(32'h3bfcd6b8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15e08a),
	.w1(32'hba90fbaa),
	.w2(32'hbaeb096d),
	.w3(32'h3c7aeb87),
	.w4(32'h3bb52e6b),
	.w5(32'hbb508983),
	.w6(32'h3c85e7df),
	.w7(32'h3c2e7469),
	.w8(32'hba90685d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb928e0f),
	.w1(32'hbc79e5db),
	.w2(32'h3b47a4e1),
	.w3(32'hbc0189eb),
	.w4(32'hbc68fda7),
	.w5(32'h3c06c6d5),
	.w6(32'hbc3ffe58),
	.w7(32'hbc860700),
	.w8(32'h3bb4e887),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3300a),
	.w1(32'h3b8fb03b),
	.w2(32'h3c14fa98),
	.w3(32'h3b560a33),
	.w4(32'hbb75da4e),
	.w5(32'h3c2eb7ec),
	.w6(32'hbb2e69e8),
	.w7(32'hbbab84b2),
	.w8(32'h3c0ccde0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5464cd),
	.w1(32'h3a585d7c),
	.w2(32'hbbb1d2cb),
	.w3(32'h3a771dcc),
	.w4(32'hbb278725),
	.w5(32'hbb92d954),
	.w6(32'hbb86b414),
	.w7(32'hbba2865a),
	.w8(32'hbb3f0229),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3a799),
	.w1(32'hbc03e0f3),
	.w2(32'hbc20f4dd),
	.w3(32'hba299087),
	.w4(32'h3ad348d5),
	.w5(32'hbc2a6ee5),
	.w6(32'hbb1f37f6),
	.w7(32'hbbbc1000),
	.w8(32'hbca6b9fc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75c9cc),
	.w1(32'hbbb2f038),
	.w2(32'hbbe4f4a0),
	.w3(32'hbc9c832b),
	.w4(32'h3b273e1b),
	.w5(32'hba15d372),
	.w6(32'hbc220f71),
	.w7(32'h3bb4543d),
	.w8(32'hbb5fe81f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3077ef),
	.w1(32'hbb98223d),
	.w2(32'h3bd2dbab),
	.w3(32'h3b96d152),
	.w4(32'h3b20d7d6),
	.w5(32'h3bf98867),
	.w6(32'h3b8440d3),
	.w7(32'h3a680a28),
	.w8(32'h3ba1cefa),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b72fb),
	.w1(32'hbbadea89),
	.w2(32'hbcd687bd),
	.w3(32'hbbba87ff),
	.w4(32'hbc45d82a),
	.w5(32'hbccd13a3),
	.w6(32'hbc055d84),
	.w7(32'hbc17321f),
	.w8(32'hbc527a7d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2064d),
	.w1(32'h39db715d),
	.w2(32'hbaf8ced7),
	.w3(32'h3c302dfd),
	.w4(32'h3ab18459),
	.w5(32'hbba569ef),
	.w6(32'h3c12ae02),
	.w7(32'h3af85616),
	.w8(32'hb909f198),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90eed4),
	.w1(32'hbbafe072),
	.w2(32'hbc5c2676),
	.w3(32'hbc111d8c),
	.w4(32'hbc41604c),
	.w5(32'hbccbb5b0),
	.w6(32'hbab42d51),
	.w7(32'hbb95c030),
	.w8(32'hbc089771),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbee8b0),
	.w1(32'hbb0a22c7),
	.w2(32'h3b40870b),
	.w3(32'hbc02901d),
	.w4(32'h3c231daa),
	.w5(32'hbb3ca397),
	.w6(32'h39c07db1),
	.w7(32'h3c9eaa98),
	.w8(32'h3badebb9),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5945),
	.w1(32'hbc2293f0),
	.w2(32'h3a0ec8d6),
	.w3(32'hbb8972df),
	.w4(32'hbcada80c),
	.w5(32'h3b68a5fc),
	.w6(32'hbc38fd7f),
	.w7(32'hbca56400),
	.w8(32'h3b2e6f55),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cf486),
	.w1(32'hbb0bc43c),
	.w2(32'hbc851fff),
	.w3(32'h3b0524e6),
	.w4(32'h3b9773b7),
	.w5(32'hbcec7a96),
	.w6(32'hbb11b448),
	.w7(32'hbb0cbf0e),
	.w8(32'hbce296d6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf7264),
	.w1(32'h3c140b17),
	.w2(32'hbb3eefda),
	.w3(32'hbaa2568b),
	.w4(32'h3c9dae09),
	.w5(32'h3c4c9bde),
	.w6(32'hba929fd7),
	.w7(32'h3c2b9f51),
	.w8(32'h3bddb075),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0ebf0),
	.w1(32'h3c358910),
	.w2(32'hbc4d86c4),
	.w3(32'h3c71d262),
	.w4(32'h3c94a37b),
	.w5(32'hbc49021d),
	.w6(32'h3c810d7a),
	.w7(32'h3c267211),
	.w8(32'h3a5f73b6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03df38),
	.w1(32'h3b5b690d),
	.w2(32'hbc32bd62),
	.w3(32'hbb6bb5c3),
	.w4(32'h3c3c27ff),
	.w5(32'hbc55a245),
	.w6(32'h3b895b28),
	.w7(32'h3afe4aa8),
	.w8(32'hba0c890a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b5129),
	.w1(32'hb98a0ab1),
	.w2(32'h3a84337d),
	.w3(32'hbca429b1),
	.w4(32'h3c842b7f),
	.w5(32'h3b4d26dd),
	.w6(32'hbbab4567),
	.w7(32'h3c8f456b),
	.w8(32'hbb063815),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8c4c8),
	.w1(32'hba2dd72e),
	.w2(32'hbbd5c8d1),
	.w3(32'hbb74b574),
	.w4(32'hb987e371),
	.w5(32'hbc73b7f3),
	.w6(32'hbbeb0e55),
	.w7(32'hb9513278),
	.w8(32'hba8dec6a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd9471f),
	.w1(32'hbbdc63ec),
	.w2(32'hbb9d4c0a),
	.w3(32'hbcb0c8b3),
	.w4(32'hbb0e4028),
	.w5(32'h3ada3328),
	.w6(32'hbbf672bb),
	.w7(32'h3c4aed10),
	.w8(32'h3c1ca033),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c350054),
	.w1(32'h3acd5455),
	.w2(32'hbc49af66),
	.w3(32'h3c23ce07),
	.w4(32'h3acc4e30),
	.w5(32'hbc9d842e),
	.w6(32'h3b9db4a9),
	.w7(32'hbb9ad675),
	.w8(32'hbcae288b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c95c4),
	.w1(32'hbc31a1d6),
	.w2(32'hbcb8825b),
	.w3(32'hbc779060),
	.w4(32'hbc8be51b),
	.w5(32'hbca98b95),
	.w6(32'hbcba542a),
	.w7(32'hbc7e931a),
	.w8(32'hba9355a8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb2226),
	.w1(32'hbb939a38),
	.w2(32'hbc210cbe),
	.w3(32'hbccde522),
	.w4(32'h3c57788b),
	.w5(32'hbbe7f8d4),
	.w6(32'hbc0e9ba8),
	.w7(32'h3c3985b3),
	.w8(32'h3b1df3be),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39fae8),
	.w1(32'h3c5734ad),
	.w2(32'hbcca6e1c),
	.w3(32'h3c6647e3),
	.w4(32'h3d0de290),
	.w5(32'hbd283317),
	.w6(32'h3ca234b7),
	.w7(32'h3d0e1fc6),
	.w8(32'hbcb14289),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbdce28),
	.w1(32'h3b385921),
	.w2(32'h3bb70613),
	.w3(32'hbc0e7d5a),
	.w4(32'h3c36a486),
	.w5(32'h3b2f5d7a),
	.w6(32'hbb689d54),
	.w7(32'h3c8def46),
	.w8(32'h3b9e6c3c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23e139),
	.w1(32'hbc2c211c),
	.w2(32'hbbb6209a),
	.w3(32'hbc83b9c2),
	.w4(32'hbc7328cd),
	.w5(32'hbbf70cb8),
	.w6(32'hbc634dc2),
	.w7(32'hbc48f615),
	.w8(32'hbc0d79ae),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc05a27),
	.w1(32'hbb60636b),
	.w2(32'h3b6a42f8),
	.w3(32'hbbe49b24),
	.w4(32'hbbaae773),
	.w5(32'hb953af12),
	.w6(32'hbc0099aa),
	.w7(32'hbbaf4843),
	.w8(32'h3c199110),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d00e3),
	.w1(32'h3b0bfd90),
	.w2(32'h3aec0f3b),
	.w3(32'h3c0cfcc0),
	.w4(32'h3c9fa1e2),
	.w5(32'hbb9c65df),
	.w6(32'h3c99215d),
	.w7(32'h3c7c3536),
	.w8(32'hbc537bc1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1e470),
	.w1(32'h3c1330fc),
	.w2(32'hbc345c0c),
	.w3(32'hb94848aa),
	.w4(32'h3c70822b),
	.w5(32'h3b79316b),
	.w6(32'hbc546196),
	.w7(32'hbc2ff026),
	.w8(32'h3b9155c9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcefc5a9),
	.w1(32'hbc47ded7),
	.w2(32'h3b1b77ba),
	.w3(32'hbc2c1d66),
	.w4(32'h3afc8459),
	.w5(32'h3ccd57ff),
	.w6(32'hbbc04442),
	.w7(32'hbb8763eb),
	.w8(32'h3ca54396),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8aba1),
	.w1(32'hbc0e5fbf),
	.w2(32'h3af4fce3),
	.w3(32'h3be94577),
	.w4(32'hbcabfd21),
	.w5(32'hbbb543a4),
	.w6(32'hbb8f48b3),
	.w7(32'hbcb37831),
	.w8(32'hbb9a2387),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952a8a6),
	.w1(32'h3b0bcee0),
	.w2(32'h3a66ff30),
	.w3(32'hbbb9933c),
	.w4(32'h39a80ff5),
	.w5(32'h3a9065f0),
	.w6(32'hbb8fef21),
	.w7(32'hba537579),
	.w8(32'hbadb299c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e2b81b),
	.w1(32'hbb0b2d9c),
	.w2(32'hba32a41c),
	.w3(32'hb9ad4b32),
	.w4(32'hba84673a),
	.w5(32'h3bd0eb17),
	.w6(32'hbac1dad3),
	.w7(32'hbb4f5e9e),
	.w8(32'h3baad241),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b815c5d),
	.w1(32'h3b5c0f66),
	.w2(32'h3ca4b093),
	.w3(32'h3bf3c09e),
	.w4(32'h3c229e2c),
	.w5(32'h3c9b4f83),
	.w6(32'h3c15ee78),
	.w7(32'h3c009663),
	.w8(32'h3ba74526),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c304a9a),
	.w1(32'hbb104f6f),
	.w2(32'h3a9b264f),
	.w3(32'h3a95ffb4),
	.w4(32'h3ab3c839),
	.w5(32'hbc089c02),
	.w6(32'hbc412d76),
	.w7(32'hbc268b7e),
	.w8(32'hbc16e501),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf86416),
	.w1(32'h3bea2aa4),
	.w2(32'hb935d7c0),
	.w3(32'hbb1d718c),
	.w4(32'h3bdd69e4),
	.w5(32'hbb1d352e),
	.w6(32'hbb818703),
	.w7(32'hb9a012d0),
	.w8(32'h3c029456),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81807e),
	.w1(32'h3b82a27e),
	.w2(32'hbbdc82e4),
	.w3(32'h3c85e5ea),
	.w4(32'h3ca05468),
	.w5(32'hbc5f94e8),
	.w6(32'h3ca70bd6),
	.w7(32'h3cbb368d),
	.w8(32'hbae8ca1a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8c23a),
	.w1(32'hbb7e4672),
	.w2(32'hbcd32779),
	.w3(32'hbc92f2c7),
	.w4(32'h3a95d221),
	.w5(32'hbcb57bc7),
	.w6(32'hbb4a56c0),
	.w7(32'h3b926dea),
	.w8(32'hbc6d8421),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb581133),
	.w1(32'hbc4b4d81),
	.w2(32'h3b4ec51f),
	.w3(32'h3b6ae98a),
	.w4(32'h3b31ccab),
	.w5(32'h3c239abe),
	.w6(32'h3b7c71fa),
	.w7(32'hbbaed5d0),
	.w8(32'h3ba5948d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29e509),
	.w1(32'h3bbec871),
	.w2(32'hbb32de28),
	.w3(32'h3c465f4e),
	.w4(32'h3c189a4f),
	.w5(32'h3bea64f1),
	.w6(32'h3bec037d),
	.w7(32'hbb154ca7),
	.w8(32'h3bfaea06),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c436efe),
	.w1(32'h3c82458c),
	.w2(32'h3a65e3fd),
	.w3(32'h3c730553),
	.w4(32'h3c5778fa),
	.w5(32'hbbe83bf4),
	.w6(32'h3c1909be),
	.w7(32'h3b95352f),
	.w8(32'hbb3bfc78),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb957617),
	.w1(32'hbc114b2b),
	.w2(32'hbc952dde),
	.w3(32'hbc976ad4),
	.w4(32'hbc751826),
	.w5(32'hbcedcf4d),
	.w6(32'hbba8f935),
	.w7(32'hbb678de2),
	.w8(32'hbc6bda80),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c759c),
	.w1(32'hbb89c936),
	.w2(32'hbceefa46),
	.w3(32'hbb63c476),
	.w4(32'hbb3972da),
	.w5(32'hbce05462),
	.w6(32'hbba360a5),
	.w7(32'hbbde5d2c),
	.w8(32'hbc2ec8a2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc910a80),
	.w1(32'h3ab04fb9),
	.w2(32'h3a3e9a34),
	.w3(32'hbc2a1bb6),
	.w4(32'h3c6cc147),
	.w5(32'hb9ce452f),
	.w6(32'h3c102b50),
	.w7(32'h3cdf1f84),
	.w8(32'h3be085f4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d2b40),
	.w1(32'h39c82e5f),
	.w2(32'hbb80b8d7),
	.w3(32'hbbca8077),
	.w4(32'h3acd2937),
	.w5(32'hbb87a0ba),
	.w6(32'h3bac0759),
	.w7(32'h3bd327b0),
	.w8(32'h3b7bfcf7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea698b),
	.w1(32'h3c208c53),
	.w2(32'hbb9de65a),
	.w3(32'hbacd9b83),
	.w4(32'h3c5ed5bc),
	.w5(32'hbbd7e323),
	.w6(32'h3bfcd5a1),
	.w7(32'h3c64cbc6),
	.w8(32'h3ae2c191),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4be69),
	.w1(32'hbb1388d4),
	.w2(32'hbbc0bf53),
	.w3(32'h3baef360),
	.w4(32'h3bdd56f0),
	.w5(32'hbc264630),
	.w6(32'h3c0b0832),
	.w7(32'h3b4a061f),
	.w8(32'h3b69e8f3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22941e),
	.w1(32'h3bc90804),
	.w2(32'h3ae7f31c),
	.w3(32'h3c8904c5),
	.w4(32'h3ce7039f),
	.w5(32'h3ae11204),
	.w6(32'h3ccd818b),
	.w7(32'h3cd60c4d),
	.w8(32'h38fb8070),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999bab6),
	.w1(32'h3ae29919),
	.w2(32'h3b0cb8d7),
	.w3(32'hbb8fced8),
	.w4(32'h3b790cec),
	.w5(32'h3c388c31),
	.w6(32'h3a97b688),
	.w7(32'hbbe938e2),
	.w8(32'h3bff64cd),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd06976),
	.w1(32'h3c3b0dd9),
	.w2(32'hbc93d9f8),
	.w3(32'h3bfdde0a),
	.w4(32'h3c1c2858),
	.w5(32'hbcc3547c),
	.w6(32'h3ca83985),
	.w7(32'h3c499429),
	.w8(32'hbc1fa1aa),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0857ee),
	.w1(32'hbc410222),
	.w2(32'hbbb19099),
	.w3(32'hbbf5117a),
	.w4(32'hbb4fcf12),
	.w5(32'hbcc9a6fe),
	.w6(32'h3b099dc3),
	.w7(32'h3b6a76c9),
	.w8(32'hbc70ab35),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae80fb),
	.w1(32'hbca39260),
	.w2(32'hbb839b57),
	.w3(32'hbd24a834),
	.w4(32'hbc988cc2),
	.w5(32'hbc338a13),
	.w6(32'hbc9a4fa8),
	.w7(32'hbc490d39),
	.w8(32'hbaa7b2cd),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb1c0b),
	.w1(32'hbb9cfabd),
	.w2(32'h3b8a8496),
	.w3(32'hbbd7d486),
	.w4(32'hbb4f03a6),
	.w5(32'hbc1d284e),
	.w6(32'h3b758cf6),
	.w7(32'h3b5b3d6a),
	.w8(32'hba3703a7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf394d),
	.w1(32'hbb534e65),
	.w2(32'h3b2e5b79),
	.w3(32'hbcacf319),
	.w4(32'hbca69e97),
	.w5(32'h3b869fdc),
	.w6(32'hbc35c5d2),
	.w7(32'hbbb47948),
	.w8(32'hb9867b58),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d552),
	.w1(32'h3b65ec6b),
	.w2(32'hbc179d87),
	.w3(32'h3bb3633b),
	.w4(32'h3b9a4677),
	.w5(32'h3abbb5b6),
	.w6(32'hba0f9051),
	.w7(32'h3b87fe12),
	.w8(32'h3c171ef3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9684ea),
	.w1(32'h3c36c90f),
	.w2(32'h3ba69ede),
	.w3(32'h3c2b71b0),
	.w4(32'h3b85d4d4),
	.w5(32'h3ac7a4a0),
	.w6(32'h3bfee239),
	.w7(32'hbbb9941a),
	.w8(32'h3b1ee2ea),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6e1b0),
	.w1(32'h3b9b85a6),
	.w2(32'hbbe95c32),
	.w3(32'hbabf5749),
	.w4(32'h3bec1872),
	.w5(32'h3b5cb573),
	.w6(32'hba6507c2),
	.w7(32'h3bba0a8a),
	.w8(32'h3c0ac7da),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacafd5c),
	.w1(32'h3a523d97),
	.w2(32'h3bf91832),
	.w3(32'h3c6a37fb),
	.w4(32'h3c775223),
	.w5(32'h3c596093),
	.w6(32'h3c3bd2af),
	.w7(32'h3bf5ccac),
	.w8(32'h3bc4e81c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2364cb),
	.w1(32'h3bc86a67),
	.w2(32'h3be02b8c),
	.w3(32'h3c3ec679),
	.w4(32'h3be5a8c1),
	.w5(32'h3c34a2a5),
	.w6(32'h3c31cc87),
	.w7(32'h3aa87853),
	.w8(32'h3bc78a00),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76eca6),
	.w1(32'h3b0d31dc),
	.w2(32'h3b518a08),
	.w3(32'h3c50797a),
	.w4(32'h3b6922c5),
	.w5(32'h3b5aa2fc),
	.w6(32'h3c458c88),
	.w7(32'h3c1697f9),
	.w8(32'h3b071605),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27f509),
	.w1(32'hb89b0429),
	.w2(32'hbb394439),
	.w3(32'h3a906378),
	.w4(32'hb958d876),
	.w5(32'hbaab4ccb),
	.w6(32'h39423a55),
	.w7(32'h3b1995ab),
	.w8(32'hba9d1cc9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba125317),
	.w1(32'h3b661908),
	.w2(32'h3bab840f),
	.w3(32'h390e5a4c),
	.w4(32'h3bc5d8ba),
	.w5(32'h3bfc4fd0),
	.w6(32'h3b70e1a3),
	.w7(32'h3bae6514),
	.w8(32'h3c848616),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccff21e),
	.w1(32'hbce03736),
	.w2(32'h3c496cf0),
	.w3(32'hbd41d0a3),
	.w4(32'hbd25bb15),
	.w5(32'h3c2a93f1),
	.w6(32'hbc14daea),
	.w7(32'hbcba3af3),
	.w8(32'h3c38452b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e846c),
	.w1(32'hba52aa5e),
	.w2(32'hbcf4e5f4),
	.w3(32'hbb286005),
	.w4(32'hbb7f07af),
	.w5(32'hbd09e126),
	.w6(32'hb96b6657),
	.w7(32'hba7253a9),
	.w8(32'h3857b582),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06850d),
	.w1(32'hbc85c274),
	.w2(32'hbcccd8b1),
	.w3(32'hbc81dea5),
	.w4(32'hb95a6399),
	.w5(32'hbd110993),
	.w6(32'h3c0b463b),
	.w7(32'h3c15c3ce),
	.w8(32'hbcf34337),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99734b),
	.w1(32'hbc428828),
	.w2(32'hbc9ece69),
	.w3(32'hbcb0b316),
	.w4(32'hbb6e9599),
	.w5(32'hbd110b3e),
	.w6(32'hbc0064e7),
	.w7(32'h3bd419d3),
	.w8(32'hbcd252a9),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc633d0b),
	.w1(32'hbbe72e91),
	.w2(32'hbbb39106),
	.w3(32'hbc641113),
	.w4(32'h3c76a896),
	.w5(32'hbc18b944),
	.w6(32'h3b1ec99b),
	.w7(32'h3c4c2533),
	.w8(32'h3b61c688),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule