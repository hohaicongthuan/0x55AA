module layer_10_featuremap_261(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac73fa),
	.w1(32'h3c1b1644),
	.w2(32'hbbbcb3d1),
	.w3(32'hbb385b53),
	.w4(32'h3b74fb91),
	.w5(32'h39a4943f),
	.w6(32'h3c336ad4),
	.w7(32'h3b9cf0ad),
	.w8(32'hb93bb261),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6749dd),
	.w1(32'h3a20de38),
	.w2(32'h3a9c5048),
	.w3(32'h3bab8fa0),
	.w4(32'h39ebb652),
	.w5(32'h3b267565),
	.w6(32'hba1154eb),
	.w7(32'hbb40e874),
	.w8(32'hba740a4d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14721c),
	.w1(32'h3b9f0adf),
	.w2(32'hb8b1171e),
	.w3(32'hbb647f27),
	.w4(32'h3accbf55),
	.w5(32'hba8ce243),
	.w6(32'h3b79a9fa),
	.w7(32'h3b85afad),
	.w8(32'h3a07fa15),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9dfc),
	.w1(32'h3c285668),
	.w2(32'h3bd8a157),
	.w3(32'h3b81d00a),
	.w4(32'h3b8d2c32),
	.w5(32'h3c0333dd),
	.w6(32'h3bd657b5),
	.w7(32'h3b6cd5d4),
	.w8(32'h3bcf947b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3d01b),
	.w1(32'hbc37b96a),
	.w2(32'hbb96f5ef),
	.w3(32'hbb4e119c),
	.w4(32'h3b1d32bf),
	.w5(32'hbb6cf89e),
	.w6(32'hbbcf3c55),
	.w7(32'h3a1bf7b6),
	.w8(32'hbab0f9f1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28ee5b),
	.w1(32'h3baa48d3),
	.w2(32'h3af96f93),
	.w3(32'h3b45bd28),
	.w4(32'h3b43ea9e),
	.w5(32'h37d810d8),
	.w6(32'h3c22ee2b),
	.w7(32'h3b00d14c),
	.w8(32'hbb2c7fe7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb25b7a),
	.w1(32'h3b6359fa),
	.w2(32'hbb17cc41),
	.w3(32'h3b824b94),
	.w4(32'hba0aef57),
	.w5(32'hbbde46d0),
	.w6(32'h377584dc),
	.w7(32'hbbb37d3d),
	.w8(32'hbbcb1964),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27e0dc),
	.w1(32'hba0fb615),
	.w2(32'hbc50112e),
	.w3(32'hbc99df4f),
	.w4(32'hbc110537),
	.w5(32'h3bb80ad6),
	.w6(32'h3b8a2d08),
	.w7(32'hbc6c2830),
	.w8(32'hbbd2371a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb82bc),
	.w1(32'h3b59c189),
	.w2(32'h39596e3a),
	.w3(32'h3b2b216b),
	.w4(32'h3b377305),
	.w5(32'hbb779a5d),
	.w6(32'h3bcbb484),
	.w7(32'h3b1b1513),
	.w8(32'hba1a91cf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69b2fd),
	.w1(32'h3baa7c56),
	.w2(32'h3b05fd51),
	.w3(32'h3aa017fa),
	.w4(32'h3ae7a0aa),
	.w5(32'hbc00449a),
	.w6(32'h3bac623c),
	.w7(32'hbb6b0507),
	.w8(32'hbc266c63),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63bf8c),
	.w1(32'h3bca3a70),
	.w2(32'h3bede635),
	.w3(32'hba343c25),
	.w4(32'h3b911df5),
	.w5(32'h398b99ad),
	.w6(32'h3bec7c82),
	.w7(32'h3baa0381),
	.w8(32'h3b64b60c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2c42c),
	.w1(32'h3c0d3cba),
	.w2(32'hbc1a2a7d),
	.w3(32'h3c32d069),
	.w4(32'h3c329d4d),
	.w5(32'hbc142119),
	.w6(32'h3c8ece00),
	.w7(32'h3ba80d3f),
	.w8(32'hbc00ce10),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaa1fd),
	.w1(32'h3bdd4ab5),
	.w2(32'hbbdf44ea),
	.w3(32'hbbc6bd62),
	.w4(32'hbba84142),
	.w5(32'hbb5fa7f6),
	.w6(32'h3c3b1cb7),
	.w7(32'hbbf6cdd8),
	.w8(32'hbbca0bf7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb948fdc),
	.w1(32'hbbfbe403),
	.w2(32'hbc12d820),
	.w3(32'hbb1eb8f4),
	.w4(32'hbb8f8241),
	.w5(32'hbc04a15d),
	.w6(32'h3a813f16),
	.w7(32'hbb87d57c),
	.w8(32'hbba8d95d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec9a86),
	.w1(32'hbb2d1589),
	.w2(32'hbb01c80d),
	.w3(32'hbb10e34e),
	.w4(32'hba3ccb19),
	.w5(32'h3bd780bf),
	.w6(32'h3af825e2),
	.w7(32'hbb6b298c),
	.w8(32'h3c45aab0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18125a),
	.w1(32'hbbfe2102),
	.w2(32'hbc0309ba),
	.w3(32'hbc40241c),
	.w4(32'hbb7ec278),
	.w5(32'h3ab08182),
	.w6(32'hbc8b1e61),
	.w7(32'hbc0b028d),
	.w8(32'h3bb67eed),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba44cc5),
	.w1(32'h3b43b5ea),
	.w2(32'h3a32bca9),
	.w3(32'h3b4ec19d),
	.w4(32'hba70912e),
	.w5(32'h3b0f604e),
	.w6(32'h3b3d3f36),
	.w7(32'h3b30597d),
	.w8(32'h3967b966),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4d77a),
	.w1(32'hbc6bd812),
	.w2(32'hbc70eaa7),
	.w3(32'hbc72c4f6),
	.w4(32'hbcab2c1b),
	.w5(32'hbc42d94d),
	.w6(32'hbc69be4e),
	.w7(32'hbce3ad2d),
	.w8(32'hbc7e7e44),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69d79),
	.w1(32'hbbbb9f20),
	.w2(32'hbba7c2d5),
	.w3(32'hbc0654bc),
	.w4(32'hbbc86672),
	.w5(32'hbbc6f99d),
	.w6(32'hbbf8e5e8),
	.w7(32'hbc2503fc),
	.w8(32'hbbf1aded),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2b524),
	.w1(32'hbaa1ee90),
	.w2(32'h3b669ec2),
	.w3(32'h3b62de01),
	.w4(32'h3b2cf700),
	.w5(32'h3b5f266b),
	.w6(32'hbb851fb0),
	.w7(32'h3a832051),
	.w8(32'h3c05d688),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb574fdb),
	.w1(32'hbc4371bd),
	.w2(32'h39a0d352),
	.w3(32'hbc1c5240),
	.w4(32'h3b67eb4f),
	.w5(32'h3b4aebc7),
	.w6(32'hbc3cc541),
	.w7(32'h3ba2e630),
	.w8(32'h3b52d81b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be587ae),
	.w1(32'h3adcd6e8),
	.w2(32'h3b6c1487),
	.w3(32'hbab9af71),
	.w4(32'hbafc2a5b),
	.w5(32'h3ba1d278),
	.w6(32'hbb4f1e97),
	.w7(32'h3b0ef1d2),
	.w8(32'h3b0f0f9c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5578e9),
	.w1(32'hbc503b1f),
	.w2(32'hbc96113e),
	.w3(32'hbc757e03),
	.w4(32'hbc062d46),
	.w5(32'hbcd387cb),
	.w6(32'hbcc3792f),
	.w7(32'hbc95480a),
	.w8(32'hbd0e1e74),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc553724),
	.w1(32'hbbb130b4),
	.w2(32'hb8b455a2),
	.w3(32'hbbc9f7f8),
	.w4(32'hbb1581b5),
	.w5(32'h3bc816ce),
	.w6(32'hbb649678),
	.w7(32'h39873587),
	.w8(32'hb9ffdf4e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380e9886),
	.w1(32'h3a5ae0f3),
	.w2(32'h3c177435),
	.w3(32'hbb25f5a7),
	.w4(32'h3b990240),
	.w5(32'h3b99e23f),
	.w6(32'hbb06e792),
	.w7(32'h3bb430de),
	.w8(32'h3ba660dc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a4fc39),
	.w1(32'hbb4d06bd),
	.w2(32'h3b2575e9),
	.w3(32'hbb6837eb),
	.w4(32'hbb610da8),
	.w5(32'hbb088800),
	.w6(32'hbb7f6ebb),
	.w7(32'hbba47286),
	.w8(32'hbae26a30),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4746ac),
	.w1(32'h3b783f36),
	.w2(32'h3ae358b5),
	.w3(32'h39a88be7),
	.w4(32'h391e6e68),
	.w5(32'h3b861d87),
	.w6(32'h3891b330),
	.w7(32'hb8c3431d),
	.w8(32'h3bd6045c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c172a62),
	.w1(32'h3b07b104),
	.w2(32'hbb48bb1e),
	.w3(32'h3badec86),
	.w4(32'h3c0abcde),
	.w5(32'hba5d2ccc),
	.w6(32'h3c6919f0),
	.w7(32'h3c02dd79),
	.w8(32'h3b21f391),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0905d9),
	.w1(32'h3b70cf3b),
	.w2(32'h3aefa790),
	.w3(32'h3b120490),
	.w4(32'hbb6c6d7a),
	.w5(32'hbc17b89f),
	.w6(32'h3b461a7b),
	.w7(32'h389e81b7),
	.w8(32'hbc09e2b5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaaa86),
	.w1(32'h3c55e62a),
	.w2(32'h3ab71e7e),
	.w3(32'h3bdd6f31),
	.w4(32'h3c091727),
	.w5(32'hb9097529),
	.w6(32'h3ce5dd96),
	.w7(32'h3bef2584),
	.w8(32'h3b9dd94b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39925fb9),
	.w1(32'hbbc73467),
	.w2(32'hb961308d),
	.w3(32'h3b88f3b7),
	.w4(32'h3b3a59ba),
	.w5(32'h3b356991),
	.w6(32'hbb9c9867),
	.w7(32'hbb7624e6),
	.w8(32'h3b904933),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb551be),
	.w1(32'hba3ce885),
	.w2(32'h38349462),
	.w3(32'hbbe01c2d),
	.w4(32'hbbc1056a),
	.w5(32'h398fe6c5),
	.w6(32'hbaf84520),
	.w7(32'h3a701a46),
	.w8(32'h3b1602af),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa20435),
	.w1(32'hba5abdfe),
	.w2(32'hba9d1d00),
	.w3(32'h3a40aca2),
	.w4(32'hbbc3bd52),
	.w5(32'hba229229),
	.w6(32'hbb506292),
	.w7(32'hbb852cb0),
	.w8(32'hbbb0e843),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3595b),
	.w1(32'h3a476ab5),
	.w2(32'h39913349),
	.w3(32'h3badaa01),
	.w4(32'hba0ada69),
	.w5(32'hbb42abe2),
	.w6(32'h3bdbfdaa),
	.w7(32'h3aa44ae5),
	.w8(32'h3a12fdd1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9defaa5),
	.w1(32'h3a684dca),
	.w2(32'h3b41e469),
	.w3(32'hbae784ef),
	.w4(32'h3a792645),
	.w5(32'h3bc33502),
	.w6(32'hbb173a4d),
	.w7(32'h3a7c0e79),
	.w8(32'hba588cfd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b137e78),
	.w1(32'h3b56f22b),
	.w2(32'h3b011e25),
	.w3(32'h39a17960),
	.w4(32'h3a14557d),
	.w5(32'hbaef0921),
	.w6(32'h3a35dd86),
	.w7(32'h3b51c978),
	.w8(32'hbbc86b88),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd8917),
	.w1(32'h3ba51bcf),
	.w2(32'hbc38ec7d),
	.w3(32'h3b80d3c4),
	.w4(32'h3bc9e492),
	.w5(32'hbc362f4c),
	.w6(32'h3b0e48ff),
	.w7(32'h3bd36e8a),
	.w8(32'hbcafd03f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51f822),
	.w1(32'h3bc5a35c),
	.w2(32'h3c30746a),
	.w3(32'h3c2179fc),
	.w4(32'h3c858edc),
	.w5(32'h3ca56377),
	.w6(32'h3b8b284c),
	.w7(32'h3c43fb2c),
	.w8(32'h3bbac338),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb05e80),
	.w1(32'h3c1c044a),
	.w2(32'h3c308756),
	.w3(32'h3c5354ca),
	.w4(32'h3c3749d5),
	.w5(32'h3c5e0dba),
	.w6(32'h3b5b66a4),
	.w7(32'h3c2db545),
	.w8(32'h3c6fb701),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bd38a),
	.w1(32'h3b8a44b0),
	.w2(32'hba66efbc),
	.w3(32'h3b9ac213),
	.w4(32'hba8afcba),
	.w5(32'h3b4b6885),
	.w6(32'h3af0f417),
	.w7(32'hbae934da),
	.w8(32'h3af51b70),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad28f14),
	.w1(32'h3bfb29f5),
	.w2(32'hbb2b5b63),
	.w3(32'h3bf7b406),
	.w4(32'h3ae0aefc),
	.w5(32'h3b00bc74),
	.w6(32'h3c5eccf2),
	.w7(32'hba03e893),
	.w8(32'h3ab7dc58),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33fe61),
	.w1(32'h3aeedf70),
	.w2(32'h3b9b63fe),
	.w3(32'hbaab309f),
	.w4(32'hbaa00a79),
	.w5(32'h3ab3ae96),
	.w6(32'h39ea8caf),
	.w7(32'h3a6cf62b),
	.w8(32'hba8140d8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0eb512),
	.w1(32'h3a69ab2f),
	.w2(32'hbaa5222d),
	.w3(32'h3a9706a6),
	.w4(32'hbaa4e8cc),
	.w5(32'h39b8317f),
	.w6(32'h3b318cff),
	.w7(32'h3926707f),
	.w8(32'hba996a57),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3a69d),
	.w1(32'hbac3e24d),
	.w2(32'hbb067255),
	.w3(32'hbb8cf00c),
	.w4(32'hbbb453a5),
	.w5(32'hbbee5cf5),
	.w6(32'hbc44617c),
	.w7(32'hbbe89e29),
	.w8(32'hbbf1156c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f03d3d),
	.w1(32'h3bb6909b),
	.w2(32'h3b866846),
	.w3(32'h368e0a22),
	.w4(32'h3b909f78),
	.w5(32'h3a827ea6),
	.w6(32'h3bc8979e),
	.w7(32'h3c03aa4a),
	.w8(32'h3b1568b9),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bfa88),
	.w1(32'h3bc64098),
	.w2(32'h3b8cc7de),
	.w3(32'h3b401054),
	.w4(32'h3b6421c2),
	.w5(32'hba18bec1),
	.w6(32'h3b9c80f2),
	.w7(32'h3ab7b4fe),
	.w8(32'hba8e4c84),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6cf85),
	.w1(32'h3b1a9c30),
	.w2(32'h3ba1753c),
	.w3(32'h3b4eaebf),
	.w4(32'h3b68766b),
	.w5(32'h3b937439),
	.w6(32'hbad3d33f),
	.w7(32'h3b005c4d),
	.w8(32'h3b9b3634),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd002a9),
	.w1(32'hbb993544),
	.w2(32'hbc47730e),
	.w3(32'hbca7978d),
	.w4(32'hbc9f524a),
	.w5(32'hbca39cd2),
	.w6(32'hbcc441d6),
	.w7(32'hbcca1bc1),
	.w8(32'hbccdcb87),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addb7cf),
	.w1(32'hbabe09c9),
	.w2(32'hbbd3800a),
	.w3(32'h3ac4d261),
	.w4(32'hbacb8a83),
	.w5(32'hb89b6221),
	.w6(32'h3bc574e3),
	.w7(32'hbac60183),
	.w8(32'hb98da7a9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c8044),
	.w1(32'hbb627dd4),
	.w2(32'h3aae9326),
	.w3(32'hbc102f88),
	.w4(32'hbb039c02),
	.w5(32'h3b5d7259),
	.w6(32'hbc0ffd31),
	.w7(32'h3ab5f442),
	.w8(32'hbb246868),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e5a61),
	.w1(32'hbc37b02a),
	.w2(32'hbb089aa7),
	.w3(32'hb96e746e),
	.w4(32'h3b8ce7d9),
	.w5(32'h3ab12558),
	.w6(32'hbb99efc3),
	.w7(32'h399f0487),
	.w8(32'h3ab63620),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee1474),
	.w1(32'hbb5fbdf1),
	.w2(32'hbad51e7e),
	.w3(32'hbba1872c),
	.w4(32'hb99d56f4),
	.w5(32'hbb50e7d5),
	.w6(32'hbb5f0f3c),
	.w7(32'hbb80a90a),
	.w8(32'hbc341c6e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb258e28),
	.w1(32'h3bb3fd64),
	.w2(32'hbb90895f),
	.w3(32'hba8ac16c),
	.w4(32'hb9d9d806),
	.w5(32'hb943cf1a),
	.w6(32'h3b41d7ad),
	.w7(32'hbb8fba08),
	.w8(32'h3abcd4af),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb488255),
	.w1(32'h3ac7dcaf),
	.w2(32'hbc7cdfad),
	.w3(32'hbb9e4874),
	.w4(32'hbbda4dcc),
	.w5(32'hbb29224d),
	.w6(32'h39fee4fa),
	.w7(32'hbc9b3930),
	.w8(32'hbbd84ca3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31044d),
	.w1(32'h3a37f863),
	.w2(32'h3b4c0087),
	.w3(32'h3acfbaec),
	.w4(32'h38a2c6c4),
	.w5(32'h3a4038e7),
	.w6(32'hbae668ba),
	.w7(32'hb9f827bc),
	.w8(32'h3b082a28),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ad42a),
	.w1(32'hbb7b6d8b),
	.w2(32'hba5568ff),
	.w3(32'hba143155),
	.w4(32'h3a79a2af),
	.w5(32'h3a9ed4b2),
	.w6(32'hbb9e5267),
	.w7(32'h39d3160a),
	.w8(32'h3b1a30c2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafa545),
	.w1(32'h3afa1e44),
	.w2(32'hbab80763),
	.w3(32'h3bad097f),
	.w4(32'hbadd476c),
	.w5(32'hba63928c),
	.w6(32'h3b6b307a),
	.w7(32'hbb291eea),
	.w8(32'hbaf4dd37),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34e683),
	.w1(32'hbb43ccd3),
	.w2(32'hbb12a1e1),
	.w3(32'h3b40e0de),
	.w4(32'hba36d26c),
	.w5(32'h3b1b17ee),
	.w6(32'hba64627c),
	.w7(32'hbb80a290),
	.w8(32'h3a85bb6a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b454790),
	.w1(32'hbb151a80),
	.w2(32'h3b33d907),
	.w3(32'hbc19c164),
	.w4(32'hba9b3d42),
	.w5(32'h3c3cd4df),
	.w6(32'hbbe9056e),
	.w7(32'h3b6062b6),
	.w8(32'h3ad3ea29),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b927ee0),
	.w1(32'hbbbec49b),
	.w2(32'h3beaa5ae),
	.w3(32'hb9f2e1e6),
	.w4(32'hbac8b1d4),
	.w5(32'hbbcb9934),
	.w6(32'hbc7aba42),
	.w7(32'hbb4db707),
	.w8(32'hbbfc1bdd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae3911),
	.w1(32'hbb962eb3),
	.w2(32'hbba934ac),
	.w3(32'hbc0b44b3),
	.w4(32'hbbe9343a),
	.w5(32'hbbf0664a),
	.w6(32'hbc6ee4f0),
	.w7(32'hbbf2d044),
	.w8(32'hbb0027ad),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe18aa3),
	.w1(32'hbc06bd75),
	.w2(32'hbb7b1667),
	.w3(32'hbc13484a),
	.w4(32'hbc0288a9),
	.w5(32'hb995e705),
	.w6(32'hbbd9b3b4),
	.w7(32'hbc193541),
	.w8(32'h3b3b9450),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f6e777),
	.w1(32'hbae082c5),
	.w2(32'hb9a5e0ed),
	.w3(32'hba84b130),
	.w4(32'hbae22da1),
	.w5(32'hba280ec8),
	.w6(32'hbb796e62),
	.w7(32'hbb01f407),
	.w8(32'hb9594acb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53f5f1),
	.w1(32'hbab99bb3),
	.w2(32'hb8963d88),
	.w3(32'h3a6fca03),
	.w4(32'h3aacda4e),
	.w5(32'hbb163d6d),
	.w6(32'hba13c96a),
	.w7(32'hba712460),
	.w8(32'h398ea145),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f26174),
	.w1(32'h3b98d4bb),
	.w2(32'h3b853328),
	.w3(32'h3bd3c913),
	.w4(32'h3b253625),
	.w5(32'h3b5c0a93),
	.w6(32'h3a2aa375),
	.w7(32'h3acb5be5),
	.w8(32'h3b762f69),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e083b3),
	.w1(32'hba844a9f),
	.w2(32'h3a3a3e85),
	.w3(32'h39e50a6f),
	.w4(32'h3b14dfea),
	.w5(32'hbc1c1480),
	.w6(32'hbb0bfe61),
	.w7(32'h3a236716),
	.w8(32'hbc234704),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a0109),
	.w1(32'h3bf43db1),
	.w2(32'hbb67ff28),
	.w3(32'hbbc9336d),
	.w4(32'h3bd29e2d),
	.w5(32'h3bfda40a),
	.w6(32'h3c598415),
	.w7(32'hbb67ca60),
	.w8(32'h3c32fe18),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1445c),
	.w1(32'h3bb6e32c),
	.w2(32'h3c05b4ba),
	.w3(32'h3c387b5c),
	.w4(32'h3b99f64e),
	.w5(32'hbc022094),
	.w6(32'h3beb333c),
	.w7(32'h39e56c50),
	.w8(32'hbc4f7f5a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b7415),
	.w1(32'hbb9621d8),
	.w2(32'hbbbb57f6),
	.w3(32'hbbba6b23),
	.w4(32'hbb83fbff),
	.w5(32'hbc253d87),
	.w6(32'hbbb2a73e),
	.w7(32'hbc3f3562),
	.w8(32'hbc017a88),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba3263),
	.w1(32'h3bc4ff8a),
	.w2(32'h3b9d09a3),
	.w3(32'h3beeef3d),
	.w4(32'h3c2318b9),
	.w5(32'h3bde9ce4),
	.w6(32'h3c2fedce),
	.w7(32'h3c27a243),
	.w8(32'h3bcbf2c9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965df20),
	.w1(32'hba5ee8b2),
	.w2(32'h3a33e1f2),
	.w3(32'h3ae597a6),
	.w4(32'h39dec571),
	.w5(32'h3bf91066),
	.w6(32'hba8b82b9),
	.w7(32'hb8b42f89),
	.w8(32'h3b923342),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b3b3d),
	.w1(32'hbc160dfa),
	.w2(32'hbb75f66c),
	.w3(32'hbb2e95e9),
	.w4(32'hbb8fd383),
	.w5(32'h3c0917e9),
	.w6(32'hbc4f1fc2),
	.w7(32'h3a7f1f02),
	.w8(32'h3b235c6f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b2802),
	.w1(32'h3b240990),
	.w2(32'h3bbf8fb7),
	.w3(32'h3b293344),
	.w4(32'hbada52a2),
	.w5(32'h39d6afd4),
	.w6(32'hbbf10a90),
	.w7(32'hbb1366a6),
	.w8(32'hbaf368f9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb176952),
	.w1(32'h3a0aab53),
	.w2(32'hb9992e95),
	.w3(32'hba445cf8),
	.w4(32'hbbc3fc65),
	.w5(32'hbc04f256),
	.w6(32'hbb7490d3),
	.w7(32'hbc0e61d1),
	.w8(32'hbc4395f1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ec74a),
	.w1(32'h3c71a59b),
	.w2(32'h3a84750a),
	.w3(32'hb81b3b5c),
	.w4(32'h3bbb70d3),
	.w5(32'h39c50968),
	.w6(32'h3ca4687e),
	.w7(32'h3b4ee5b5),
	.w8(32'hbb2257c7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fb26f),
	.w1(32'hbbffbc67),
	.w2(32'hbc2ff0b1),
	.w3(32'hbb70bf69),
	.w4(32'hbbb2fe8d),
	.w5(32'h3a85bd00),
	.w6(32'h3911b522),
	.w7(32'hbc07bdd9),
	.w8(32'hbc05fa99),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb485a3b),
	.w1(32'hbb9f2095),
	.w2(32'hbc31250b),
	.w3(32'hbbfe7908),
	.w4(32'hbc1574aa),
	.w5(32'hbc01c2c7),
	.w6(32'hbba62b41),
	.w7(32'hbc7a4a10),
	.w8(32'hbc6aa984),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f4e44),
	.w1(32'hba1abd8c),
	.w2(32'h3b3a2f75),
	.w3(32'hbbe96b26),
	.w4(32'h388f8709),
	.w5(32'hbb85afbd),
	.w6(32'hbb51764b),
	.w7(32'h3a4cf363),
	.w8(32'hb910a394),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4274c0),
	.w1(32'h3a4f93f5),
	.w2(32'hbbb068ab),
	.w3(32'hba0ac2d9),
	.w4(32'h3b475a9d),
	.w5(32'hbb3cb2bf),
	.w6(32'h3c229c66),
	.w7(32'hbbaec7f9),
	.w8(32'hbade27ca),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b5baa),
	.w1(32'h3adac119),
	.w2(32'hbb81a283),
	.w3(32'h3badc035),
	.w4(32'h3aa8a7c5),
	.w5(32'hbc033a30),
	.w6(32'h3c2744e4),
	.w7(32'hbbca9e37),
	.w8(32'hbbb5773d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75bd8f),
	.w1(32'hbabc7f3e),
	.w2(32'hbbe54d95),
	.w3(32'hbb7647ad),
	.w4(32'hbb883dd9),
	.w5(32'h399c5bd3),
	.w6(32'h3bdae7f3),
	.w7(32'hbb3249bb),
	.w8(32'hbb057b20),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb562ff4),
	.w1(32'hbbe0fa7e),
	.w2(32'hbc158a28),
	.w3(32'hbbbec426),
	.w4(32'hbbd4243d),
	.w5(32'hbb4bec42),
	.w6(32'hbb8e544a),
	.w7(32'hbc274a7a),
	.w8(32'hbc443ea6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95cce4),
	.w1(32'h3bad042b),
	.w2(32'h3aaf7090),
	.w3(32'h3a18003a),
	.w4(32'h3ae1b594),
	.w5(32'hbbc7ef1b),
	.w6(32'h3baae1bc),
	.w7(32'h39a3fde5),
	.w8(32'hbaa0e7f4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989bd39),
	.w1(32'h3c935cef),
	.w2(32'h3c6fceae),
	.w3(32'h3b8a5c4e),
	.w4(32'h3bc11502),
	.w5(32'h3b830cb1),
	.w6(32'h3c64f78d),
	.w7(32'h3c2aadf1),
	.w8(32'hba701b06),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7496c6),
	.w1(32'h3b2ae41e),
	.w2(32'h39b9d969),
	.w3(32'hbb4352b7),
	.w4(32'h38d21fb5),
	.w5(32'hbbc91283),
	.w6(32'hbb19819d),
	.w7(32'hba9a160f),
	.w8(32'hbb855f40),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a467a),
	.w1(32'hb980ebd3),
	.w2(32'h3af212ff),
	.w3(32'hbad96647),
	.w4(32'h3b2cb63a),
	.w5(32'h3b7e57a9),
	.w6(32'h3bb678b0),
	.w7(32'h3b44019e),
	.w8(32'h3a1e8650),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b023f),
	.w1(32'h3a9006b8),
	.w2(32'h3b296c88),
	.w3(32'h3b567f11),
	.w4(32'h3bb94b4b),
	.w5(32'h3c12f644),
	.w6(32'h3b751004),
	.w7(32'h3bc6cd7f),
	.w8(32'h3b9875ff),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22f670),
	.w1(32'hbaabf48f),
	.w2(32'h398be176),
	.w3(32'h3b6768fc),
	.w4(32'h3b72c81d),
	.w5(32'h39f3fcc0),
	.w6(32'hbb14e2ee),
	.w7(32'h3af787fc),
	.w8(32'h3b7b76c2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e04ff6),
	.w1(32'hbb2538da),
	.w2(32'hbacb651a),
	.w3(32'hbc1521aa),
	.w4(32'hbbc240b0),
	.w5(32'hbc154276),
	.w6(32'hbb993545),
	.w7(32'hbae79376),
	.w8(32'hba51f98b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5502f8),
	.w1(32'hba89b1ac),
	.w2(32'hbc97e196),
	.w3(32'hbbaf4f11),
	.w4(32'hbc927486),
	.w5(32'hbc96f68f),
	.w6(32'h3c9b5485),
	.w7(32'hbcbe328c),
	.w8(32'hbcc02e38),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c8773),
	.w1(32'h3bb06dc1),
	.w2(32'h3bb882fb),
	.w3(32'h3c4d0c02),
	.w4(32'h3c040472),
	.w5(32'h3b2c1734),
	.w6(32'h3bcfa478),
	.w7(32'h3c1202f3),
	.w8(32'hba4e18de),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba40f47),
	.w1(32'h3b63d3e8),
	.w2(32'h3a423dad),
	.w3(32'h3a92edb3),
	.w4(32'h3c1de814),
	.w5(32'h3b30e44b),
	.w6(32'hbb97395a),
	.w7(32'h3c0e75f8),
	.w8(32'hbb638ead),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ad03),
	.w1(32'hbb7bf3f9),
	.w2(32'h3b595c61),
	.w3(32'hbb9410d6),
	.w4(32'h3aa09c95),
	.w5(32'h3c0da0d3),
	.w6(32'hbadf0202),
	.w7(32'h3bcc560c),
	.w8(32'h3b6d9226),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b5572),
	.w1(32'hbb4a03f7),
	.w2(32'hbb23aad0),
	.w3(32'hbaf3a7f7),
	.w4(32'h3b74b3d8),
	.w5(32'h3b68b59b),
	.w6(32'hbaf412d0),
	.w7(32'hbadf1b90),
	.w8(32'h3bf8e882),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2939c),
	.w1(32'hbb1ca2af),
	.w2(32'hbb0ef15c),
	.w3(32'h3bfc506b),
	.w4(32'h3ac0c4b6),
	.w5(32'h3acc9c65),
	.w6(32'h3a2b371f),
	.w7(32'hbaa26303),
	.w8(32'h3b127e8e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafa981),
	.w1(32'h3b1c2ff1),
	.w2(32'h3a9038db),
	.w3(32'h39803ee5),
	.w4(32'h3b94dd75),
	.w5(32'h3c31481b),
	.w6(32'h3afd19c7),
	.w7(32'h3befe9ad),
	.w8(32'h3c14b7a6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe009e),
	.w1(32'h3af8db2a),
	.w2(32'h3b529b6e),
	.w3(32'h3b24d028),
	.w4(32'h3b939845),
	.w5(32'h3aed5a0e),
	.w6(32'hbaeee8e2),
	.w7(32'h3b20b91c),
	.w8(32'h3b8dd016),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2bd98),
	.w1(32'hbc25d4dc),
	.w2(32'hbbf7b5c3),
	.w3(32'h3b08e1c1),
	.w4(32'hbbe3e687),
	.w5(32'h394d191d),
	.w6(32'hbb6008ca),
	.w7(32'hbc66e0c2),
	.w8(32'hbbe19519),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeeafa4),
	.w1(32'hbb458c6a),
	.w2(32'hbb380737),
	.w3(32'h3b8add2f),
	.w4(32'h3c3b0f39),
	.w5(32'h3a305af3),
	.w6(32'h3ab4d502),
	.w7(32'hba46bc84),
	.w8(32'hbc8c62a7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b402d24),
	.w1(32'h3ad2bbc9),
	.w2(32'hbc2301cd),
	.w3(32'hbc8f666c),
	.w4(32'hbc27f630),
	.w5(32'hbb473d4d),
	.w6(32'hbb46d9d4),
	.w7(32'hbc663bba),
	.w8(32'hbc559ff4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb03e0),
	.w1(32'h3cbd562b),
	.w2(32'h3c9df0bd),
	.w3(32'h3ccf2f34),
	.w4(32'h3cd27e23),
	.w5(32'h3c35058e),
	.w6(32'hb9a14fe3),
	.w7(32'h3cb22910),
	.w8(32'hba8c85e4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bfb03),
	.w1(32'hbb66403d),
	.w2(32'h3b9be9a8),
	.w3(32'hbbd265f1),
	.w4(32'h3bc4ce53),
	.w5(32'hba171a7e),
	.w6(32'hb986b88c),
	.w7(32'hbb8f3e0d),
	.w8(32'hba020f9f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8b149),
	.w1(32'h3bb0969e),
	.w2(32'hbc07f226),
	.w3(32'h3c11848e),
	.w4(32'h3bf7c4a9),
	.w5(32'h3c4feba1),
	.w6(32'hb9199937),
	.w7(32'h3a03971f),
	.w8(32'h3ad16d98),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88a8fb),
	.w1(32'h3c7664f3),
	.w2(32'h3c73fb6b),
	.w3(32'h3c7c7d33),
	.w4(32'h3c1905c1),
	.w5(32'hbbadae8c),
	.w6(32'h3c014fd8),
	.w7(32'h3ba8acf6),
	.w8(32'hbb16830b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f7a7a),
	.w1(32'hbbc4f69b),
	.w2(32'hbcc9cdc4),
	.w3(32'hbcd8a86b),
	.w4(32'hbc58f756),
	.w5(32'hbc93a415),
	.w6(32'hbab66e6c),
	.w7(32'hbc10a8f0),
	.w8(32'hbcd302f6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb809585f),
	.w1(32'hbb8c6167),
	.w2(32'hbbe5a11b),
	.w3(32'hb9db2781),
	.w4(32'h3bb9483c),
	.w5(32'hbbd1beea),
	.w6(32'hbab9bd39),
	.w7(32'h3bbf26c4),
	.w8(32'hbcaa4fb4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39474dac),
	.w1(32'hbb627fec),
	.w2(32'hbac0e7e4),
	.w3(32'hbc1cfd76),
	.w4(32'hbaffc50c),
	.w5(32'h3b27dacb),
	.w6(32'hbc069a1a),
	.w7(32'hbb1c04ee),
	.w8(32'h3b0d7869),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3fa14),
	.w1(32'hb9c76dc7),
	.w2(32'h3b25c92e),
	.w3(32'h3ade0a3e),
	.w4(32'h3b47fa29),
	.w5(32'hbaefee32),
	.w6(32'hbb885ea2),
	.w7(32'h3b5ccae5),
	.w8(32'hbbafd916),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98fd48),
	.w1(32'hbbaa9d19),
	.w2(32'hbb7ba724),
	.w3(32'hbbe43c3c),
	.w4(32'hbb1e4bd0),
	.w5(32'hb84a936f),
	.w6(32'hbc00463a),
	.w7(32'hbc57e184),
	.w8(32'hbb4949ef),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b350b25),
	.w1(32'hbae956f8),
	.w2(32'h3ac770eb),
	.w3(32'hbb111a2c),
	.w4(32'h3b0f17a9),
	.w5(32'hbb8db258),
	.w6(32'hbad1266a),
	.w7(32'hb9ce388d),
	.w8(32'hbb6f563a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb854218),
	.w1(32'hbc64fb5f),
	.w2(32'hbbd61862),
	.w3(32'hbc5ac6ff),
	.w4(32'hbc0ba340),
	.w5(32'h3abc35a4),
	.w6(32'h3bb14b86),
	.w7(32'hbb565b32),
	.w8(32'hbab1fe5f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb029171),
	.w1(32'h3bb9f55b),
	.w2(32'h3bb79423),
	.w3(32'h3bbec7e7),
	.w4(32'h3b864bfb),
	.w5(32'hbbbc7d65),
	.w6(32'h3b8ccb79),
	.w7(32'h3b889bb9),
	.w8(32'hbc2924e3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab747b9),
	.w1(32'h3b26fffe),
	.w2(32'h3aacf4af),
	.w3(32'hbc1021f6),
	.w4(32'hba51f586),
	.w5(32'hb9eb5f20),
	.w6(32'hbc20185e),
	.w7(32'h3b0a0146),
	.w8(32'h3b2a0602),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1f695),
	.w1(32'hbb1e48a2),
	.w2(32'hbc0a8add),
	.w3(32'hbbb1da4e),
	.w4(32'hbb222312),
	.w5(32'hbb95d3b4),
	.w6(32'hbc4af94d),
	.w7(32'hbc4eacbd),
	.w8(32'hbbb56d1b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06d9c0),
	.w1(32'h3b32d726),
	.w2(32'h3bbbb4bb),
	.w3(32'hbb09f74c),
	.w4(32'h3b768893),
	.w5(32'h3b784f67),
	.w6(32'hb8f7edbe),
	.w7(32'hbb938f3b),
	.w8(32'hbb842e46),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ddd4c),
	.w1(32'hbb96bf9f),
	.w2(32'h3954b46a),
	.w3(32'h3aac09a9),
	.w4(32'h3a83eef9),
	.w5(32'hbbdd728e),
	.w6(32'h3b477bb2),
	.w7(32'hbb20a8c5),
	.w8(32'hbc1beb37),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94151b),
	.w1(32'hbbeac3dc),
	.w2(32'hbb8f4694),
	.w3(32'hbbe8b10c),
	.w4(32'hbb0bffb0),
	.w5(32'h3a58c64c),
	.w6(32'hbc567c89),
	.w7(32'hbbe27a20),
	.w8(32'hbb4ee701),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc044214),
	.w1(32'hbb5896ba),
	.w2(32'hbbfb7172),
	.w3(32'hbbeb501d),
	.w4(32'hbb89a08f),
	.w5(32'h3bd49157),
	.w6(32'h3c9ff83c),
	.w7(32'h3bbe7b24),
	.w8(32'h3b36baf8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e1932),
	.w1(32'h3bc7d81b),
	.w2(32'h3bda3402),
	.w3(32'h38d56d81),
	.w4(32'h3bd2513d),
	.w5(32'h3b8c1b38),
	.w6(32'hbc0124af),
	.w7(32'h398f5fa8),
	.w8(32'hba49042f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d306ec),
	.w1(32'h3c8d73ab),
	.w2(32'h3c21fc2d),
	.w3(32'h3c9eca21),
	.w4(32'h3c1d5e83),
	.w5(32'h3baae184),
	.w6(32'h3cb15717),
	.w7(32'h3bf12a70),
	.w8(32'hba4f69c7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9747),
	.w1(32'h3a57aa73),
	.w2(32'h3b9c8d29),
	.w3(32'hba42eacb),
	.w4(32'h3b61901f),
	.w5(32'hbbb3b346),
	.w6(32'hbbe92469),
	.w7(32'h3a1e8776),
	.w8(32'hbb9ec5e2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffe0cb),
	.w1(32'hba79431c),
	.w2(32'hb8ae8d11),
	.w3(32'hbb69a881),
	.w4(32'hbb8d08c6),
	.w5(32'hbc4d40a8),
	.w6(32'hbba19060),
	.w7(32'h3a4da9ba),
	.w8(32'hbc52d83c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb550cfd),
	.w1(32'h3b8ca9f8),
	.w2(32'hbaa46ab0),
	.w3(32'hbc1b434e),
	.w4(32'hbb0f076a),
	.w5(32'hbb8a8c8b),
	.w6(32'h3a4347d5),
	.w7(32'hbbb90b3a),
	.w8(32'hbc200b33),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6bcea),
	.w1(32'hbb3b804e),
	.w2(32'h3a9ecb89),
	.w3(32'h3936db29),
	.w4(32'hba57462f),
	.w5(32'hbbd89109),
	.w6(32'hba47a6cb),
	.w7(32'hbb90bc41),
	.w8(32'hbb821ee1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe68b90),
	.w1(32'h3b62419f),
	.w2(32'hba7fb185),
	.w3(32'hbbf77d80),
	.w4(32'hbb4824ce),
	.w5(32'h3bc2afcc),
	.w6(32'hbaca052c),
	.w7(32'hbb261959),
	.w8(32'h3b9f3f00),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ac549),
	.w1(32'hbb0b3415),
	.w2(32'h3a896c6e),
	.w3(32'h3ae1864d),
	.w4(32'hb93bd88f),
	.w5(32'hbb093f65),
	.w6(32'h3ba18714),
	.w7(32'h3b544487),
	.w8(32'hbbc0049c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64e16e),
	.w1(32'hbb0a07b2),
	.w2(32'h3a0abab8),
	.w3(32'hbb603e37),
	.w4(32'hba9d53c1),
	.w5(32'h3b84a38b),
	.w6(32'hbaeef87e),
	.w7(32'hbae7a43d),
	.w8(32'h3b844e03),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3633d9),
	.w1(32'h3bc659d0),
	.w2(32'h3b4f9ed4),
	.w3(32'h3c1c6fee),
	.w4(32'h3b240f06),
	.w5(32'hbad08a7d),
	.w6(32'hba8349fc),
	.w7(32'hba0da527),
	.w8(32'hbbb747e1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01542e),
	.w1(32'hbab43b2b),
	.w2(32'hb9b43e4e),
	.w3(32'hbb7ced3d),
	.w4(32'hba60fa57),
	.w5(32'hbb910c37),
	.w6(32'hbc3c5030),
	.w7(32'hbc05058e),
	.w8(32'hbc0ba3c9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88230e),
	.w1(32'hba7c81da),
	.w2(32'hbab007c9),
	.w3(32'hbb793f5a),
	.w4(32'hbbc17159),
	.w5(32'hbb113986),
	.w6(32'hbb7d7e7b),
	.w7(32'hbb2696e4),
	.w8(32'hbc08b698),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9e2b9),
	.w1(32'hbb6904e6),
	.w2(32'hbc2afabf),
	.w3(32'hbc1bc701),
	.w4(32'hbb5ee6d8),
	.w5(32'h3b93d650),
	.w6(32'h3a83477a),
	.w7(32'hba7cfbba),
	.w8(32'h3a8309df),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89c208),
	.w1(32'h3baa58ea),
	.w2(32'h3c084b17),
	.w3(32'h3aa91154),
	.w4(32'h3bb2ec0b),
	.w5(32'hbb031087),
	.w6(32'h3c177eeb),
	.w7(32'h3bf5585a),
	.w8(32'hbc19754b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248337),
	.w1(32'hbb8d1c0d),
	.w2(32'hba69aec0),
	.w3(32'h3a371f0f),
	.w4(32'h3ba50ad2),
	.w5(32'hbad24e4a),
	.w6(32'hbbfec6e8),
	.w7(32'hbb407f65),
	.w8(32'hbb4c197e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba617a5),
	.w1(32'hbaf9debb),
	.w2(32'h3b05f46c),
	.w3(32'hbb402eca),
	.w4(32'h3b731024),
	.w5(32'hbb667810),
	.w6(32'hbb8867bf),
	.w7(32'h39921c6a),
	.w8(32'hbba5ab6b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb53fd4),
	.w1(32'hbc435997),
	.w2(32'hbc47b738),
	.w3(32'hbc4a7076),
	.w4(32'hbc4871d1),
	.w5(32'hbbd58c41),
	.w6(32'hbc71978e),
	.w7(32'hbc7a85c2),
	.w8(32'hbc41b190),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03fd59),
	.w1(32'h397c5b41),
	.w2(32'h396faf4d),
	.w3(32'h392e573a),
	.w4(32'h3b80e585),
	.w5(32'hbb311dbf),
	.w6(32'hbb58c8d5),
	.w7(32'h3a61e383),
	.w8(32'hbac4ddf5),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4184),
	.w1(32'hbb7dae1a),
	.w2(32'hbbb4e30a),
	.w3(32'hbab6cd31),
	.w4(32'h38fd1d0e),
	.w5(32'hba06ae58),
	.w6(32'hbc04bbf2),
	.w7(32'hbbdd7578),
	.w8(32'hbb475b4b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399757d5),
	.w1(32'hbbca719a),
	.w2(32'hbbd98abb),
	.w3(32'hbb889480),
	.w4(32'hbb461e02),
	.w5(32'hbbee53e1),
	.w6(32'hbbac78de),
	.w7(32'hbbe3f9c6),
	.w8(32'hbc2dc8c2),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0309d0),
	.w1(32'hbad3c803),
	.w2(32'h3b9ce75a),
	.w3(32'hbbeaab5e),
	.w4(32'hbac491da),
	.w5(32'h39fe7b2d),
	.w6(32'hbb84bd31),
	.w7(32'h3b405adc),
	.w8(32'hbb825fa6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b31f9),
	.w1(32'hba4fedc4),
	.w2(32'hbbf53b66),
	.w3(32'hbbaa5a25),
	.w4(32'hbb9f9feb),
	.w5(32'hbc473fad),
	.w6(32'hbc327c8b),
	.w7(32'hbc43d123),
	.w8(32'hbc610694),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb507894),
	.w1(32'h3c11daab),
	.w2(32'hbc1077b3),
	.w3(32'hb988a337),
	.w4(32'hbc3fd89b),
	.w5(32'hbbbc877a),
	.w6(32'h3c859ff4),
	.w7(32'hbc6038fc),
	.w8(32'hbb8bc0c6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb790aca),
	.w1(32'h3b9bd65b),
	.w2(32'h3c322c10),
	.w3(32'h3c047b45),
	.w4(32'h3bc6a641),
	.w5(32'hbabe0348),
	.w6(32'h3c9713a2),
	.w7(32'h3c6c694e),
	.w8(32'h3aa5ecfc),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc73a9),
	.w1(32'hbb5eaa37),
	.w2(32'hbb321032),
	.w3(32'hbc08b79b),
	.w4(32'hbb312d91),
	.w5(32'h3b869c46),
	.w6(32'h3b78cde3),
	.w7(32'hbb7c5d8d),
	.w8(32'h3a3dc1c7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986b1de),
	.w1(32'hba960814),
	.w2(32'hbad1f7fe),
	.w3(32'hbba8ffea),
	.w4(32'hba2983d9),
	.w5(32'hbb8d311b),
	.w6(32'hbc0426fd),
	.w7(32'hbb5ae577),
	.w8(32'hbbf7883e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1835ca),
	.w1(32'hbadafb30),
	.w2(32'hba8aeafd),
	.w3(32'hbbbba015),
	.w4(32'hbb53604f),
	.w5(32'hbb361a18),
	.w6(32'hbbece34b),
	.w7(32'hbbb8b013),
	.w8(32'hbc32b23a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac62444),
	.w1(32'hbad25f0b),
	.w2(32'h3a689857),
	.w3(32'hbbd310f0),
	.w4(32'hbacb37f5),
	.w5(32'hbc086a9a),
	.w6(32'hbb67b680),
	.w7(32'hbbc82833),
	.w8(32'h3b839f58),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0db18),
	.w1(32'hbb1020da),
	.w2(32'hbb574fd9),
	.w3(32'hbbc270bd),
	.w4(32'h3a9b8c0d),
	.w5(32'h3b0f858f),
	.w6(32'h3c50ee4c),
	.w7(32'h3a0dbace),
	.w8(32'hbb94241b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb686a75),
	.w1(32'h3c27ed91),
	.w2(32'h3bc6f0ec),
	.w3(32'hbc182f8c),
	.w4(32'hbc08d2c2),
	.w5(32'h3c5e15b9),
	.w6(32'hbc21131c),
	.w7(32'hbbbc9e33),
	.w8(32'h3c828cbf),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3f325),
	.w1(32'h3c127b70),
	.w2(32'h3af124c6),
	.w3(32'h3c008184),
	.w4(32'h3b7fe0a0),
	.w5(32'hbbeb020f),
	.w6(32'h3b28447c),
	.w7(32'h3b1ac3e6),
	.w8(32'hbc44ae4e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf60386),
	.w1(32'hbc18cbb5),
	.w2(32'hbbe15c0b),
	.w3(32'hbc1a0c3f),
	.w4(32'hbbd1517f),
	.w5(32'hbb3324bb),
	.w6(32'hbc96c253),
	.w7(32'hbc706a33),
	.w8(32'hbbac7fc9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb690a45),
	.w1(32'h3b017696),
	.w2(32'hba7bedca),
	.w3(32'h3b11e33b),
	.w4(32'h3b0d18b8),
	.w5(32'h3b6f2a9b),
	.w6(32'hbb980b98),
	.w7(32'hbb78f3ec),
	.w8(32'h3be61ff6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e7fd0),
	.w1(32'hbb89e1aa),
	.w2(32'hbb66e9e5),
	.w3(32'h3badf766),
	.w4(32'hbaaff9c5),
	.w5(32'hba58d669),
	.w6(32'hbc1d8352),
	.w7(32'hbbb91a66),
	.w8(32'hbc641df2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48cc72),
	.w1(32'hbb2a727b),
	.w2(32'h3b55cc6c),
	.w3(32'h3c30c922),
	.w4(32'h3c6ab310),
	.w5(32'h3b0cbabc),
	.w6(32'h3c488c84),
	.w7(32'hbb0c666e),
	.w8(32'h3a5128f7),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace9bd6),
	.w1(32'h3b19313a),
	.w2(32'h3b105b30),
	.w3(32'hbb329a13),
	.w4(32'h3b4320fc),
	.w5(32'hb98f75a7),
	.w6(32'h3b1c6d10),
	.w7(32'h3af15341),
	.w8(32'h3bc64e2a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49edf6),
	.w1(32'h3b343c1b),
	.w2(32'h3b5fb7eb),
	.w3(32'hba46040b),
	.w4(32'hb9863924),
	.w5(32'h3ae20561),
	.w6(32'h3bf1c5b9),
	.w7(32'h3bcc604a),
	.w8(32'h3a8d9fc2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f19d54),
	.w1(32'hbb787175),
	.w2(32'hbb05eb7e),
	.w3(32'hbb35ed23),
	.w4(32'h3aa96987),
	.w5(32'h3b8d9c9a),
	.w6(32'hbb9b6536),
	.w7(32'h38bf5afd),
	.w8(32'h3a4dd81a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94cb92),
	.w1(32'hba34dcf4),
	.w2(32'hb985229d),
	.w3(32'h3bb889ec),
	.w4(32'hbb1d4bbf),
	.w5(32'hbb31294e),
	.w6(32'h3aef3a56),
	.w7(32'h3b0b813e),
	.w8(32'hbbb2f98b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba813e7d),
	.w1(32'h3b64dac2),
	.w2(32'h3b9c1882),
	.w3(32'h3a891e65),
	.w4(32'h3bf8cb91),
	.w5(32'hbbef0f67),
	.w6(32'hbb23d7c2),
	.w7(32'h3c133934),
	.w8(32'h3bb84825),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45673c),
	.w1(32'hbc916769),
	.w2(32'hbc8a7718),
	.w3(32'hbc17d0b3),
	.w4(32'hbc1e71ce),
	.w5(32'hbc0fa58a),
	.w6(32'hbafa89fc),
	.w7(32'hbc381552),
	.w8(32'hbb8d93ad),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82e458),
	.w1(32'hba3fd9b1),
	.w2(32'hbc04b042),
	.w3(32'hbbb7232e),
	.w4(32'hbb1343a6),
	.w5(32'hbb95e3d0),
	.w6(32'hbbd17716),
	.w7(32'hbc530314),
	.w8(32'h3b915ccb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab6b1d),
	.w1(32'hbb122fa3),
	.w2(32'hbc0652fb),
	.w3(32'h3aae6d35),
	.w4(32'h3bb2aed2),
	.w5(32'hbc0de041),
	.w6(32'hbb83b09c),
	.w7(32'hbbf921e6),
	.w8(32'hbca8cc21),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99341d7),
	.w1(32'h3ab1c67a),
	.w2(32'h3bd45491),
	.w3(32'hbbc0b702),
	.w4(32'h3b4b0452),
	.w5(32'h3be5129d),
	.w6(32'hbbf36e75),
	.w7(32'hbb091b09),
	.w8(32'hbbb74afd),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ada05),
	.w1(32'h3a75c84f),
	.w2(32'h3be7d42e),
	.w3(32'h3aa91e97),
	.w4(32'h3b22df63),
	.w5(32'h3ba8e8a5),
	.w6(32'hbbfde1ec),
	.w7(32'hbb27fc5e),
	.w8(32'hbaa10cd3),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08c283),
	.w1(32'hbb482443),
	.w2(32'hb9352068),
	.w3(32'hbb4084ff),
	.w4(32'hbbbadbdf),
	.w5(32'hbad04b1c),
	.w6(32'hbbca4022),
	.w7(32'hbc0ddcbc),
	.w8(32'hbc375466),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2033df),
	.w1(32'hbb3d3419),
	.w2(32'hbbcdd5e7),
	.w3(32'h3c74ee5b),
	.w4(32'h3b163e25),
	.w5(32'hba63f95b),
	.w6(32'hbb0b87c8),
	.w7(32'hbc267e8c),
	.w8(32'h3bc40dfb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5aaaea),
	.w1(32'h3b4a83de),
	.w2(32'h3a8b91db),
	.w3(32'h3baeca0b),
	.w4(32'h38243493),
	.w5(32'hbb8b2385),
	.w6(32'h3c170338),
	.w7(32'h3c2cc37a),
	.w8(32'hbbfcc343),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00ac4c),
	.w1(32'hbb0eed57),
	.w2(32'h3a4420d1),
	.w3(32'hb9b47079),
	.w4(32'hbb84ad9c),
	.w5(32'h3c9d03b8),
	.w6(32'hbb810230),
	.w7(32'hbb6f2b22),
	.w8(32'h3b04f336),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dbd50),
	.w1(32'h3c13cfc6),
	.w2(32'h3ca2bcf2),
	.w3(32'h3c5dc837),
	.w4(32'h3ccdd3ea),
	.w5(32'h3b3d6424),
	.w6(32'hbc46550b),
	.w7(32'h3c5f1b74),
	.w8(32'h3b9ecb61),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f29b4),
	.w1(32'h3bd717cb),
	.w2(32'hbbbea3b7),
	.w3(32'h3a856b63),
	.w4(32'hbba7f899),
	.w5(32'hbbc3cb2b),
	.w6(32'hbb0a6d46),
	.w7(32'hbc06f8de),
	.w8(32'hbc82b05d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a202b16),
	.w1(32'h3b33319c),
	.w2(32'h3bab339c),
	.w3(32'h3b287ddf),
	.w4(32'h3b9db0a5),
	.w5(32'h3ca9acf5),
	.w6(32'hb926d9a6),
	.w7(32'h3b46a996),
	.w8(32'h3cb7eddc),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9caa30),
	.w1(32'h3c571a75),
	.w2(32'h3c10c6cd),
	.w3(32'h3c458fb5),
	.w4(32'h3c464a2b),
	.w5(32'hbc1a305b),
	.w6(32'h3cc7457f),
	.w7(32'h3c9df45d),
	.w8(32'hbb6bd872),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7219b9),
	.w1(32'hbb4538e6),
	.w2(32'hbafe9b40),
	.w3(32'hbc1def31),
	.w4(32'hbc23c950),
	.w5(32'h3c337e8e),
	.w6(32'h3b7e410b),
	.w7(32'h3a86ac88),
	.w8(32'h3b637ccf),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac6f6a),
	.w1(32'h3c04546b),
	.w2(32'h3c8b8b07),
	.w3(32'h3b85941a),
	.w4(32'h3c3833e4),
	.w5(32'hbc79040b),
	.w6(32'hbc238e4e),
	.w7(32'h3b483ad4),
	.w8(32'hbc855589),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2d357),
	.w1(32'hbc5af8dc),
	.w2(32'hbc388cb3),
	.w3(32'hbc5fd057),
	.w4(32'hbc5fe764),
	.w5(32'hbc539069),
	.w6(32'hbbf7baa2),
	.w7(32'hbc363e0f),
	.w8(32'hbc643cf0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60980b),
	.w1(32'hbc376b60),
	.w2(32'hbc6f5220),
	.w3(32'hbc78ccba),
	.w4(32'hbca51ec4),
	.w5(32'hbc61a899),
	.w6(32'hbbe2b6b9),
	.w7(32'hbcad4735),
	.w8(32'hbc8851d3),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85f65d),
	.w1(32'hbc1ba9ed),
	.w2(32'hbc057fc7),
	.w3(32'hbc35e6c6),
	.w4(32'hbc0b0972),
	.w5(32'hbb9d5605),
	.w6(32'hbc7e676b),
	.w7(32'hbc6b98de),
	.w8(32'h3b1a3c00),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02dc51),
	.w1(32'h3abb2a10),
	.w2(32'hbbc63ba4),
	.w3(32'hba92e1ca),
	.w4(32'hbb43f362),
	.w5(32'hbbb94b78),
	.w6(32'h3bdcf929),
	.w7(32'hbb270d4b),
	.w8(32'hbc44640e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc9d52),
	.w1(32'hbb6843ae),
	.w2(32'hbb1f3768),
	.w3(32'hbb7f451c),
	.w4(32'hbb3a7885),
	.w5(32'h3be0e2b0),
	.w6(32'hbc79c936),
	.w7(32'hbc1d67d7),
	.w8(32'hba449a5b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb78637),
	.w1(32'h3c02bf71),
	.w2(32'h3bbdc925),
	.w3(32'h3c2c1198),
	.w4(32'hbb4a2ebc),
	.w5(32'h394a7ff0),
	.w6(32'h3bcd193e),
	.w7(32'hbb810145),
	.w8(32'h3c0b9f0e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23ac5f),
	.w1(32'h3abb244b),
	.w2(32'h39bf01c5),
	.w3(32'hbb15cbf9),
	.w4(32'hba7e10d3),
	.w5(32'hbb3f8308),
	.w6(32'h3cc9ecf6),
	.w7(32'h3be6a705),
	.w8(32'hb805fd10),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e2bd4),
	.w1(32'hbb974b84),
	.w2(32'h3af71196),
	.w3(32'hbc1ba7b3),
	.w4(32'hbb2767fa),
	.w5(32'hbc3b21a2),
	.w6(32'hbc3a9761),
	.w7(32'hbb137052),
	.w8(32'hbbfc5e3a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8423e7),
	.w1(32'hbc1aa7be),
	.w2(32'h3b82d034),
	.w3(32'hbc5b42cf),
	.w4(32'hba7f99cc),
	.w5(32'h3b1da50c),
	.w6(32'hbcc7b194),
	.w7(32'hbadb3b40),
	.w8(32'hba5b4025),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ad374),
	.w1(32'h3b343660),
	.w2(32'hba1286e7),
	.w3(32'h3ae45e11),
	.w4(32'h3a013942),
	.w5(32'hbb773cc1),
	.w6(32'hbbc45943),
	.w7(32'hba19ad18),
	.w8(32'hbb9d1276),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a237),
	.w1(32'h3aa14bee),
	.w2(32'h3b9893f2),
	.w3(32'hbb28cd4d),
	.w4(32'hbaf32ab3),
	.w5(32'hb8f31edb),
	.w6(32'hbabdc095),
	.w7(32'hbb47048c),
	.w8(32'hbbb8dd23),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d14440),
	.w1(32'hba59dde1),
	.w2(32'hba111d1f),
	.w3(32'h3bfbdf13),
	.w4(32'hbb2c0af0),
	.w5(32'hbb365ef4),
	.w6(32'h3aa778b0),
	.w7(32'hbb8f0b9f),
	.w8(32'hbc6b2b21),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad2508),
	.w1(32'h3be4b895),
	.w2(32'h3be4a894),
	.w3(32'hbbc3a220),
	.w4(32'h3c33ea06),
	.w5(32'hbb8d2fc0),
	.w6(32'hbc63e6f7),
	.w7(32'h3c57a8c8),
	.w8(32'hbc72856d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e3ae3),
	.w1(32'hbb75cb24),
	.w2(32'hba3b1719),
	.w3(32'hbb8150fe),
	.w4(32'hba418e35),
	.w5(32'hbc2bc3cd),
	.w6(32'hbc889432),
	.w7(32'hbc17a635),
	.w8(32'hbb15be5e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f744b),
	.w1(32'hbb8a3ef1),
	.w2(32'hbba70121),
	.w3(32'hbba4d13a),
	.w4(32'hbc0da871),
	.w5(32'hbbd1e617),
	.w6(32'h3c1225a6),
	.w7(32'h3af0d6ac),
	.w8(32'hbbb5a209),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c5b84),
	.w1(32'h3b8db775),
	.w2(32'h3bcb024a),
	.w3(32'h3c00ae02),
	.w4(32'h3c6ab5ba),
	.w5(32'h3aab96f8),
	.w6(32'h3bc8ca0a),
	.w7(32'h3c23c999),
	.w8(32'h3b8b1fc7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba4a8f),
	.w1(32'hbb80f097),
	.w2(32'hbc00e061),
	.w3(32'hbc126276),
	.w4(32'hbbc620c9),
	.w5(32'hbaa5faab),
	.w6(32'h3b8edb92),
	.w7(32'hbbd670fa),
	.w8(32'hbbeadfe1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0786c5),
	.w1(32'h3b81001e),
	.w2(32'h3c1e32ae),
	.w3(32'hbb896cd5),
	.w4(32'hba783cdf),
	.w5(32'h3b83d287),
	.w6(32'hbc0f48e7),
	.w7(32'hbbc58abd),
	.w8(32'hbb2558b9),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ffa49),
	.w1(32'h3c178616),
	.w2(32'h3b8e78a1),
	.w3(32'h3c20b96a),
	.w4(32'h3ada3a1d),
	.w5(32'h3afbef02),
	.w6(32'h3bda04bd),
	.w7(32'hba8e0123),
	.w8(32'h3a8947af),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc84250),
	.w1(32'h3bb21404),
	.w2(32'h3a325bbd),
	.w3(32'h3bc59390),
	.w4(32'hb9ee309f),
	.w5(32'hba2864ed),
	.w6(32'h3ba9081c),
	.w7(32'hba728928),
	.w8(32'hbb5756ac),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0421e3),
	.w1(32'h393cf59d),
	.w2(32'hbb54993c),
	.w3(32'h3a5b8359),
	.w4(32'h3b47dbcf),
	.w5(32'hbbd6c950),
	.w6(32'hbc20f6cc),
	.w7(32'hbb986a65),
	.w8(32'hbc410535),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53a29c),
	.w1(32'hbb53f0e9),
	.w2(32'hba01c230),
	.w3(32'hbb1f7dff),
	.w4(32'hbb01a9e5),
	.w5(32'hbbe4af6a),
	.w6(32'hbbb72a7e),
	.w7(32'hbb83bbc0),
	.w8(32'h3881598f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c568c),
	.w1(32'h3bee7211),
	.w2(32'h3b79204a),
	.w3(32'hba457c56),
	.w4(32'h3a889f80),
	.w5(32'h3bca4d3d),
	.w6(32'h3ca0aab1),
	.w7(32'h3c0dca9c),
	.w8(32'h3c48eca0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7b309),
	.w1(32'hbb022b09),
	.w2(32'hbad1d770),
	.w3(32'hbac5132f),
	.w4(32'h39f22317),
	.w5(32'h3a8455d9),
	.w6(32'hbb6af105),
	.w7(32'h3ae8deaa),
	.w8(32'h3abd67aa),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4628e7),
	.w1(32'hbaa8c98a),
	.w2(32'hbb38a0c8),
	.w3(32'hbc0ffca6),
	.w4(32'hbafd44ff),
	.w5(32'h3bd0f11d),
	.w6(32'h3beee602),
	.w7(32'hbbc31019),
	.w8(32'h3c4ec208),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad58b4),
	.w1(32'h3c57c2de),
	.w2(32'h3ba4d8fa),
	.w3(32'h3c90afbf),
	.w4(32'h3c1a01f7),
	.w5(32'h3ba55887),
	.w6(32'h3cb1f92f),
	.w7(32'h3c81bbd0),
	.w8(32'h3912bf8a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b445a09),
	.w1(32'hbb469a0d),
	.w2(32'h3aeabc45),
	.w3(32'h3b625f9b),
	.w4(32'h3a94c698),
	.w5(32'hbc1715f6),
	.w6(32'hbb897da4),
	.w7(32'hba24139e),
	.w8(32'hbb157465),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb46f9),
	.w1(32'hbc28f861),
	.w2(32'hbc1c5f81),
	.w3(32'hbc568f21),
	.w4(32'hbc550bc1),
	.w5(32'hba937586),
	.w6(32'hbb078a0e),
	.w7(32'hbbd9831a),
	.w8(32'hbbd2128b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb729345),
	.w1(32'h3a4bc67b),
	.w2(32'hbb9a40ee),
	.w3(32'h39ea2b24),
	.w4(32'h39c4f38a),
	.w5(32'hbaf3ce2e),
	.w6(32'h3b96c960),
	.w7(32'h3a56e78f),
	.w8(32'hbb828177),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba099460),
	.w1(32'h3b006e32),
	.w2(32'hbba8bf87),
	.w3(32'hbbfcd2e9),
	.w4(32'hbb94a9eb),
	.w5(32'hbb2fd373),
	.w6(32'hbbd0012c),
	.w7(32'hbb8d1903),
	.w8(32'h3a9cf44e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b518ff0),
	.w1(32'h3c0698a8),
	.w2(32'h3b92c50c),
	.w3(32'h3bfcb3dd),
	.w4(32'h3bc6d81b),
	.w5(32'h3b76a76d),
	.w6(32'h3cb7e28c),
	.w7(32'h3c02e0a9),
	.w8(32'h3beddd89),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb851a0a),
	.w1(32'h3b27994d),
	.w2(32'hbb1c0c6a),
	.w3(32'h3ac20dda),
	.w4(32'hb8c7723b),
	.w5(32'h3a10723a),
	.w6(32'hbb0be5a4),
	.w7(32'hbb41456e),
	.w8(32'hbbde4c95),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b802264),
	.w1(32'hb9807907),
	.w2(32'h3c3a2532),
	.w3(32'hbb5f08ae),
	.w4(32'h3c07ac29),
	.w5(32'hbb9ebb62),
	.w6(32'hbbb4a912),
	.w7(32'hb9e7ec40),
	.w8(32'h3b36b5fe),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81a2fa),
	.w1(32'h3aba7986),
	.w2(32'hbb9d96a9),
	.w3(32'hbb528fe9),
	.w4(32'hbb4bd9a5),
	.w5(32'hbbaa5249),
	.w6(32'h3c6f1b25),
	.w7(32'h3bbcf45e),
	.w8(32'hbb93a231),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf37fac),
	.w1(32'hbb696c11),
	.w2(32'hbba323fd),
	.w3(32'hbc29619d),
	.w4(32'hbc15496b),
	.w5(32'h3c99fe80),
	.w6(32'hbc019303),
	.w7(32'hbc3ae901),
	.w8(32'h3cae5b19),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafe803),
	.w1(32'h3c29944e),
	.w2(32'h3bb5a934),
	.w3(32'h3c1ccd35),
	.w4(32'h3c3d3a2b),
	.w5(32'hbb92764a),
	.w6(32'hb953d8bb),
	.w7(32'h3bb3fa5a),
	.w8(32'hbbe2062d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3df06),
	.w1(32'hbc035551),
	.w2(32'hbc076084),
	.w3(32'hbbe463d8),
	.w4(32'hbba4ab56),
	.w5(32'h39958f1e),
	.w6(32'hbb56304e),
	.w7(32'hbc20ab59),
	.w8(32'h39d8cbd9),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77ad8d),
	.w1(32'hb9705289),
	.w2(32'hbc192bf4),
	.w3(32'h3b389b9b),
	.w4(32'hb9ae031e),
	.w5(32'h3b2f9789),
	.w6(32'h3bcdb158),
	.w7(32'h3b68a707),
	.w8(32'h3c6a6c7d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b993180),
	.w1(32'h3c030e52),
	.w2(32'h3c1b795a),
	.w3(32'h3bb2ac11),
	.w4(32'h3c2ad716),
	.w5(32'h3b248bee),
	.w6(32'h3cbb02ce),
	.w7(32'h3c9be5dd),
	.w8(32'h3a54e118),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ba7cd),
	.w1(32'hbb173945),
	.w2(32'hbc220f83),
	.w3(32'hb9bc6d32),
	.w4(32'h3b12a023),
	.w5(32'hbc8cf3d2),
	.w6(32'hbb7382ea),
	.w7(32'hba609bd6),
	.w8(32'hbc9515ae),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c2b2c),
	.w1(32'hbb818cb1),
	.w2(32'h3b11dadb),
	.w3(32'hbba98c59),
	.w4(32'hbb8fdca0),
	.w5(32'h3bc92b46),
	.w6(32'h3a92ec0d),
	.w7(32'h3b9be8a6),
	.w8(32'hbbdbd179),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b099486),
	.w1(32'hbad75602),
	.w2(32'hbb27d2ea),
	.w3(32'hb989e212),
	.w4(32'h3ab5d20e),
	.w5(32'h3b28b283),
	.w6(32'hbc046762),
	.w7(32'hbb7945dc),
	.w8(32'h39c742bb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d5c0e),
	.w1(32'hb9daa94a),
	.w2(32'hb8ad1e6a),
	.w3(32'hba9f099d),
	.w4(32'hbabca3f0),
	.w5(32'hbbaa3716),
	.w6(32'hbbb00761),
	.w7(32'hbb02ae9e),
	.w8(32'hbc161cc2),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ac32a),
	.w1(32'hbb7de914),
	.w2(32'hbb496895),
	.w3(32'hbbf1b439),
	.w4(32'hbb919f97),
	.w5(32'hbaa501bd),
	.w6(32'hbbe05d00),
	.w7(32'hbbf885b0),
	.w8(32'hbc0d913e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b865ab9),
	.w1(32'h3c291005),
	.w2(32'hbbc3b66e),
	.w3(32'h3c21cedd),
	.w4(32'h3c6fe3df),
	.w5(32'hbacbacbc),
	.w6(32'h39a84b53),
	.w7(32'h3b88db0a),
	.w8(32'hbb956381),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e59fd),
	.w1(32'hbc0c658d),
	.w2(32'hbab687a9),
	.w3(32'hbbb83310),
	.w4(32'hbb06b0fb),
	.w5(32'hbbc53649),
	.w6(32'hbc076b75),
	.w7(32'hbbe940ea),
	.w8(32'hbc257c5e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cf0f3),
	.w1(32'h3be20f37),
	.w2(32'hbb6cd206),
	.w3(32'hbb16302c),
	.w4(32'hbb652a47),
	.w5(32'hbb8b1dda),
	.w6(32'hbc3ddcad),
	.w7(32'hbc318671),
	.w8(32'hbc78eb60),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc097035),
	.w1(32'h3bb0ab9e),
	.w2(32'h3c1564b2),
	.w3(32'hbba5d20d),
	.w4(32'h3a3e1952),
	.w5(32'h3c23f9ef),
	.w6(32'hbb2d0598),
	.w7(32'h3b2b1338),
	.w8(32'h3c43df8d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd6afa),
	.w1(32'h3c00de72),
	.w2(32'h3a12526c),
	.w3(32'h3bc76ce0),
	.w4(32'h3b7c1b2e),
	.w5(32'h3c75cbb8),
	.w6(32'h3c82535c),
	.w7(32'h3c02d232),
	.w8(32'h3c79c458),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62e444),
	.w1(32'h3c0f1e08),
	.w2(32'h3b9cd09b),
	.w3(32'h3c2b65ca),
	.w4(32'h3bd65932),
	.w5(32'h3bde9d1a),
	.w6(32'h3b16b3be),
	.w7(32'h3b4edcb8),
	.w8(32'h3c8826f5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ea611),
	.w1(32'h3c61f9d2),
	.w2(32'h3b062b25),
	.w3(32'hbb4fa222),
	.w4(32'hb985cee1),
	.w5(32'h3b26198f),
	.w6(32'h3c8acb34),
	.w7(32'h3bed9301),
	.w8(32'h3c2798fb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9d62a),
	.w1(32'h39e08ac2),
	.w2(32'hbbb9169d),
	.w3(32'h3c0ab2b0),
	.w4(32'hbba4c85e),
	.w5(32'hba4e0b89),
	.w6(32'h3c8288ee),
	.w7(32'h399c1f35),
	.w8(32'h3c13e733),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53a2d0),
	.w1(32'hbbc23333),
	.w2(32'hbbf5134b),
	.w3(32'hbb4e81d1),
	.w4(32'hbbdf3228),
	.w5(32'h3a62e996),
	.w6(32'hbc06e852),
	.w7(32'hbc634683),
	.w8(32'h39e989ec),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3296c2),
	.w1(32'hbb01174a),
	.w2(32'hbb4d23e5),
	.w3(32'h38de5f27),
	.w4(32'h38b79a48),
	.w5(32'hbb93606a),
	.w6(32'hbaa928bf),
	.w7(32'hba9f6000),
	.w8(32'hbc1d13c4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d16b3),
	.w1(32'h3ba91caf),
	.w2(32'hbb8e5347),
	.w3(32'hbb5e8a45),
	.w4(32'hba9348ca),
	.w5(32'hb97df4c0),
	.w6(32'hba8613cb),
	.w7(32'hbbac84b2),
	.w8(32'hbbee5f82),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba116362),
	.w1(32'hbb476df8),
	.w2(32'h3af29312),
	.w3(32'h3a9a57fc),
	.w4(32'h3be24cff),
	.w5(32'hbad54a91),
	.w6(32'hba97cd82),
	.w7(32'h3bf7e160),
	.w8(32'h3b03dc80),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0602df),
	.w1(32'hbb9090a5),
	.w2(32'h3b855585),
	.w3(32'hbb74606b),
	.w4(32'hbbc11f77),
	.w5(32'hbb122af0),
	.w6(32'hbb4e7383),
	.w7(32'hbbe3a5da),
	.w8(32'hba12cafb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5be7d8),
	.w1(32'h3b9bb0de),
	.w2(32'hbbfecbfb),
	.w3(32'hbbcaded7),
	.w4(32'hbba595fe),
	.w5(32'hbbf14b20),
	.w6(32'hbbeaa19d),
	.w7(32'hbc3e1a57),
	.w8(32'hbc75a8ac),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f26eb),
	.w1(32'h3a91f264),
	.w2(32'hbadf9ae4),
	.w3(32'hba4a9032),
	.w4(32'hbb25d950),
	.w5(32'hbaabe97f),
	.w6(32'hbb4c67ab),
	.w7(32'hbbc077e8),
	.w8(32'hbb55ac24),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80e2fa),
	.w1(32'hbbd124ee),
	.w2(32'hbb53a46f),
	.w3(32'h3af5af33),
	.w4(32'h3bbe56e8),
	.w5(32'hbaa7c2a8),
	.w6(32'h3b710ce0),
	.w7(32'h3aab4607),
	.w8(32'hbb34eaed),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab683a),
	.w1(32'hba225f07),
	.w2(32'hbc1e39f6),
	.w3(32'h3a2fcf7a),
	.w4(32'h3ac73f8e),
	.w5(32'hbb4948e0),
	.w6(32'hbbca1845),
	.w7(32'hbbfe1b89),
	.w8(32'hbbbd7a71),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb915a),
	.w1(32'h3c0b3ba6),
	.w2(32'hba93bb09),
	.w3(32'h398627f2),
	.w4(32'h3b96f8d3),
	.w5(32'hb9cf5d89),
	.w6(32'hbac4198a),
	.w7(32'h3b6c81c4),
	.w8(32'hba1304ea),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac19d77),
	.w1(32'h3b375736),
	.w2(32'hbb21af3e),
	.w3(32'h3abd9e0a),
	.w4(32'h3a028a43),
	.w5(32'h3b6380c8),
	.w6(32'h39e7b05f),
	.w7(32'hbae4b010),
	.w8(32'h3b218298),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b810272),
	.w1(32'h39069fb4),
	.w2(32'hbae6b8dd),
	.w3(32'h3a12dc39),
	.w4(32'h3a9f72d2),
	.w5(32'h3a1783ba),
	.w6(32'hbaa57cea),
	.w7(32'hb896e83d),
	.w8(32'h3bd9cd3e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2a4e1),
	.w1(32'h3bcbd5b1),
	.w2(32'h3b03c036),
	.w3(32'hbb46528e),
	.w4(32'hbb512bfd),
	.w5(32'h3b26571b),
	.w6(32'h3a13eab3),
	.w7(32'hbb47706c),
	.w8(32'hbb506c97),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b768215),
	.w1(32'h3c256be9),
	.w2(32'h3b5b2d79),
	.w3(32'h3b86cc66),
	.w4(32'h3bca125e),
	.w5(32'h3a1d7638),
	.w6(32'h3c1721da),
	.w7(32'h3c193d93),
	.w8(32'hbb65a71f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98c0e0),
	.w1(32'h3b4a602b),
	.w2(32'hba6e0a41),
	.w3(32'hbbc3a0f4),
	.w4(32'hba37477a),
	.w5(32'hbb811ddd),
	.w6(32'hbb9e853a),
	.w7(32'hbb957b59),
	.w8(32'hbb46993f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a8d6e),
	.w1(32'h3b43efe4),
	.w2(32'h3b72adfe),
	.w3(32'hbb5608a5),
	.w4(32'hb9cead1f),
	.w5(32'hbb00fed6),
	.w6(32'hba74f166),
	.w7(32'hba162c1b),
	.w8(32'hbb903241),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6ea5c),
	.w1(32'h3949ad73),
	.w2(32'h3b340ced),
	.w3(32'h39f574fd),
	.w4(32'hb9a52a12),
	.w5(32'h39d3f1e5),
	.w6(32'hbb7e3f88),
	.w7(32'hbb8d8533),
	.w8(32'hbbdac855),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aad09),
	.w1(32'hbb30e34d),
	.w2(32'hbaf47995),
	.w3(32'h3b9b5de2),
	.w4(32'h3b02b3c3),
	.w5(32'hbb073dcb),
	.w6(32'h3aa40753),
	.w7(32'hbaa26d27),
	.w8(32'hbb4f24b5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8210a5),
	.w1(32'h3b71cac5),
	.w2(32'h3b8851c5),
	.w3(32'hbb8d9ca9),
	.w4(32'hba808f0e),
	.w5(32'h3b0eba19),
	.w6(32'hbb42dd8b),
	.w7(32'hbabd8968),
	.w8(32'hbae34d36),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8154a),
	.w1(32'hbacfef7f),
	.w2(32'h3a95a22f),
	.w3(32'h3a98c8d0),
	.w4(32'hbb2bf010),
	.w5(32'hbb6ae0f1),
	.w6(32'hbabdb501),
	.w7(32'h3a1b2f44),
	.w8(32'hbb73c63d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914fc88),
	.w1(32'hbbcf30ff),
	.w2(32'hbb7d462e),
	.w3(32'h3b0bb641),
	.w4(32'h3b1919ff),
	.w5(32'h3b27753b),
	.w6(32'hbbe8d931),
	.w7(32'hbb8da093),
	.w8(32'h3a962608),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ba350),
	.w1(32'hba91de81),
	.w2(32'hbad72783),
	.w3(32'hbbb7e8f7),
	.w4(32'hbbaa05d6),
	.w5(32'hbbd7f1d0),
	.w6(32'hbbc2aea0),
	.w7(32'hbbf41be5),
	.w8(32'hbc1a748c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde294f),
	.w1(32'hbbdc5017),
	.w2(32'hbbbbbf28),
	.w3(32'hbc0f3b46),
	.w4(32'hbba6ade5),
	.w5(32'hbb8feadc),
	.w6(32'hbc2016a2),
	.w7(32'hbbc6031f),
	.w8(32'hbb816d88),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb931174),
	.w1(32'h3ae88446),
	.w2(32'h393b7182),
	.w3(32'hbb82917c),
	.w4(32'hbaca780d),
	.w5(32'h3a4902a4),
	.w6(32'hbb4556cc),
	.w7(32'hbadacb48),
	.w8(32'h3a2bcd52),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf747ff),
	.w1(32'h3be434f6),
	.w2(32'h3aa90fc2),
	.w3(32'hbbf30813),
	.w4(32'hbae47433),
	.w5(32'h3b401b99),
	.w6(32'h3a9dd023),
	.w7(32'h3b4f1284),
	.w8(32'hbc1107fa),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05780f),
	.w1(32'h3a84cd25),
	.w2(32'hbc17cdd4),
	.w3(32'h3b9bbdc5),
	.w4(32'h3ad1971a),
	.w5(32'hbb7ed95b),
	.w6(32'hbbb81f7f),
	.w7(32'hbbed5702),
	.w8(32'h3c6523db),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb383e9),
	.w1(32'hba7609fd),
	.w2(32'hbaa54543),
	.w3(32'hbc12316a),
	.w4(32'hbbac3bed),
	.w5(32'h3ae4b11c),
	.w6(32'h3be8df69),
	.w7(32'hbb24edb2),
	.w8(32'h39a7a4b2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1486f4),
	.w1(32'hbbd33bdc),
	.w2(32'hbafe49b8),
	.w3(32'h3aa1be09),
	.w4(32'hbb1cb28c),
	.w5(32'h3a9db8f9),
	.w6(32'h3bdbedad),
	.w7(32'hba9294e0),
	.w8(32'h3b404ace),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e340b),
	.w1(32'hbb0baff1),
	.w2(32'h3af0256a),
	.w3(32'hbb090df0),
	.w4(32'h39bf6450),
	.w5(32'h3a805357),
	.w6(32'hbbd5879f),
	.w7(32'hbbaa30e6),
	.w8(32'h3afe7d88),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeca191),
	.w1(32'hbb341c61),
	.w2(32'hba7953c3),
	.w3(32'hb92e197a),
	.w4(32'hbb6f75e4),
	.w5(32'hbb240b93),
	.w6(32'h3b2bfbb2),
	.w7(32'hbb4306cd),
	.w8(32'hb9d3e2b7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15d27a),
	.w1(32'h3a37be2e),
	.w2(32'h3bd7a3c3),
	.w3(32'hbb165ee3),
	.w4(32'h3b7f988d),
	.w5(32'h3b3821c6),
	.w6(32'hbbd9935c),
	.w7(32'h3b5422b4),
	.w8(32'h3c173620),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule