module layer_10_featuremap_292(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacb7de),
	.w1(32'hb9a360ac),
	.w2(32'hb977b54a),
	.w3(32'h3b41fb4c),
	.w4(32'h3a2acc9b),
	.w5(32'hba69bd4b),
	.w6(32'h3b1083dd),
	.w7(32'hb8be1611),
	.w8(32'hbabf5602),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15db0a),
	.w1(32'h3aa3b13d),
	.w2(32'h3a6100be),
	.w3(32'hba9b908e),
	.w4(32'hbae0290a),
	.w5(32'h3a8acfac),
	.w6(32'h37914148),
	.w7(32'hb9c01a0b),
	.w8(32'h39694ded),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb265bda),
	.w1(32'hbb2052af),
	.w2(32'hbaf3ea31),
	.w3(32'h390e4753),
	.w4(32'hbaff7966),
	.w5(32'hba9ed109),
	.w6(32'h398e58d9),
	.w7(32'h39f8f72e),
	.w8(32'hba6d4668),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9828f2f),
	.w1(32'hb9b5e1b4),
	.w2(32'h39517119),
	.w3(32'hba87b176),
	.w4(32'hba9579cf),
	.w5(32'hbb75bbb5),
	.w6(32'hbab29088),
	.w7(32'hba646981),
	.w8(32'hbb839b84),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dc936),
	.w1(32'hbbc7beac),
	.w2(32'hbbb3fff5),
	.w3(32'hbbbd8bf6),
	.w4(32'hbb8daa88),
	.w5(32'h3b67e2dd),
	.w6(32'hbbe37929),
	.w7(32'hbb92e900),
	.w8(32'h3b816876),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dc8be),
	.w1(32'h3af9fdab),
	.w2(32'h38cc0975),
	.w3(32'h3b310f39),
	.w4(32'h3a913a85),
	.w5(32'hb94acbd0),
	.w6(32'h3b5bb7d1),
	.w7(32'h3a5a9baa),
	.w8(32'h3a52a3c6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad68e26),
	.w1(32'h3aa8c146),
	.w2(32'h3a1cf5be),
	.w3(32'h39271a57),
	.w4(32'h3968ca04),
	.w5(32'h3a1ad5e2),
	.w6(32'h3ab3eddf),
	.w7(32'h3aa31a1c),
	.w8(32'h3980b6fd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba353f63),
	.w1(32'hbad89bf6),
	.w2(32'hb9fc49d6),
	.w3(32'h39ace8ee),
	.w4(32'hba267a6c),
	.w5(32'h3b85a59b),
	.w6(32'hba950e09),
	.w7(32'hba573520),
	.w8(32'h3b98290f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77d455),
	.w1(32'h3b384bc2),
	.w2(32'h3af5c68b),
	.w3(32'h3b38dbe1),
	.w4(32'h3b5471e1),
	.w5(32'h3ac6521f),
	.w6(32'h3b37ed26),
	.w7(32'h3b09caa7),
	.w8(32'h3afaef27),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f2c5a),
	.w1(32'h3a53f8c3),
	.w2(32'hb96053e2),
	.w3(32'h3a37ca81),
	.w4(32'hb92f5ac5),
	.w5(32'hb9afc23a),
	.w6(32'h3aa469a0),
	.w7(32'h39f2a969),
	.w8(32'h388877d0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa178d0),
	.w1(32'hbaba02d5),
	.w2(32'hba9f9a47),
	.w3(32'hb99519eb),
	.w4(32'hba96c256),
	.w5(32'h398221bd),
	.w6(32'hb8a02edf),
	.w7(32'hba4cda45),
	.w8(32'hb8597da8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a115b72),
	.w1(32'hb9c79bf7),
	.w2(32'hbb11cb26),
	.w3(32'h3adc6113),
	.w4(32'hb98ec712),
	.w5(32'hbb29f0ec),
	.w6(32'h3ad1e1c5),
	.w7(32'hb9f80fa6),
	.w8(32'hbb69dc0d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40f5af),
	.w1(32'hbb7ce594),
	.w2(32'hbb594f42),
	.w3(32'hbb630b4f),
	.w4(32'hbb5e8fa5),
	.w5(32'hbaf0a480),
	.w6(32'hbb9440a3),
	.w7(32'hbb9ffa5c),
	.w8(32'hbb2fe718),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c4371),
	.w1(32'hbba47295),
	.w2(32'hba7882ef),
	.w3(32'hbb7a31d9),
	.w4(32'hba97db61),
	.w5(32'h38c0630c),
	.w6(32'hbbb4ea37),
	.w7(32'hbb151146),
	.w8(32'hb827f2f6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f2afe),
	.w1(32'hb9d1d896),
	.w2(32'h39a65c91),
	.w3(32'h38f2e52a),
	.w4(32'hb8216f38),
	.w5(32'hbabd6b85),
	.w6(32'h397219cc),
	.w7(32'h39e051cb),
	.w8(32'hbb599c01),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d8034),
	.w1(32'hbb4dd9f3),
	.w2(32'hbb462f45),
	.w3(32'hbb0158ec),
	.w4(32'hbb36d82a),
	.w5(32'h3b9b3330),
	.w6(32'hbb112de4),
	.w7(32'hbb614d3b),
	.w8(32'h3b89ce1f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8937d1),
	.w1(32'h3b15789e),
	.w2(32'h39b4af6b),
	.w3(32'h3b810483),
	.w4(32'h3b003111),
	.w5(32'hbae3d1a0),
	.w6(32'h3b94ee17),
	.w7(32'h3a82c4a8),
	.w8(32'hbb0c157a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004503),
	.w1(32'hbae1864f),
	.w2(32'hbad9ff8f),
	.w3(32'hbb1b0128),
	.w4(32'hbb4fc84e),
	.w5(32'hb9c685dd),
	.w6(32'hbafc75f6),
	.w7(32'hbb2a0bc1),
	.w8(32'hbaf29096),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba027465),
	.w1(32'h3873777c),
	.w2(32'hb9699ed7),
	.w3(32'h3995f3ef),
	.w4(32'h3a100bd0),
	.w5(32'hbb346913),
	.w6(32'h3abf3218),
	.w7(32'h39f3d60e),
	.w8(32'hba872cbe),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad66a3a),
	.w1(32'hb9934bac),
	.w2(32'hb86a043e),
	.w3(32'hbabc9e35),
	.w4(32'hb9aa5b67),
	.w5(32'hb8657ad2),
	.w6(32'hba709d9e),
	.w7(32'hb9b22b6d),
	.w8(32'hbabe3f3f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b90e3),
	.w1(32'h3a146307),
	.w2(32'h3aa8d077),
	.w3(32'h3b00f730),
	.w4(32'h3925c2bd),
	.w5(32'h3b4adae7),
	.w6(32'h3ab651cd),
	.w7(32'h3a7447c2),
	.w8(32'h3b79006e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73df1f),
	.w1(32'h3b830b22),
	.w2(32'h3b45aeae),
	.w3(32'h3ae1be00),
	.w4(32'h3aae640b),
	.w5(32'hb9e361a6),
	.w6(32'h3b0bdbfa),
	.w7(32'h3ab84bb2),
	.w8(32'hb9c7b450),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95205d),
	.w1(32'hba9bcb38),
	.w2(32'hbb0944da),
	.w3(32'hba400a3b),
	.w4(32'hbaf414b3),
	.w5(32'hbaf4210d),
	.w6(32'hba0e6bfd),
	.w7(32'hbadb4bc9),
	.w8(32'hbb0cc910),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084ffd),
	.w1(32'hbab89656),
	.w2(32'hbb253bf5),
	.w3(32'hbab15023),
	.w4(32'hbb4087ce),
	.w5(32'hbab2c71d),
	.w6(32'hbb09d7ca),
	.w7(32'hbae8b008),
	.w8(32'hbb038ee8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa957b),
	.w1(32'hbb140d57),
	.w2(32'hbb3606dc),
	.w3(32'hbb512eeb),
	.w4(32'hbb0ee030),
	.w5(32'h3a46159e),
	.w6(32'hb980214e),
	.w7(32'h38402810),
	.w8(32'hb9ad1468),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fca6ab),
	.w1(32'h38dec76a),
	.w2(32'h3a7b5ca6),
	.w3(32'h3ad7dc89),
	.w4(32'h3adcb7ea),
	.w5(32'h3a0a9f37),
	.w6(32'h3b02be69),
	.w7(32'h3ac5c136),
	.w8(32'h3a3b19f1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12c091),
	.w1(32'hbab86183),
	.w2(32'hb8bd9457),
	.w3(32'h3982502c),
	.w4(32'h3a9b813b),
	.w5(32'h3bb3caf0),
	.w6(32'hb914932b),
	.w7(32'hb98a047c),
	.w8(32'h3bd1403a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a1b6f),
	.w1(32'h3b57d9cc),
	.w2(32'h3b255ca8),
	.w3(32'h3b871557),
	.w4(32'h3b290e46),
	.w5(32'hbb4397c6),
	.w6(32'h3b62c29c),
	.w7(32'h3b33e4a0),
	.w8(32'hbb3a3363),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba892c56),
	.w1(32'hb85e5f5b),
	.w2(32'hbaae1835),
	.w3(32'hbb07f99e),
	.w4(32'hba651b49),
	.w5(32'hbadf27c5),
	.w6(32'hba9bc720),
	.w7(32'hbaa65f54),
	.w8(32'hbb25d7f9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb021a88),
	.w1(32'hba924e7e),
	.w2(32'h399a5ed4),
	.w3(32'hba5d10f9),
	.w4(32'hba9038cf),
	.w5(32'hbb1e6ec0),
	.w6(32'hbb193ba3),
	.w7(32'hbab05118),
	.w8(32'hbac7d5cf),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3a933),
	.w1(32'hba95a45e),
	.w2(32'hba105a92),
	.w3(32'hbb9b17db),
	.w4(32'hbade9017),
	.w5(32'h3b1816bc),
	.w6(32'hba9537fc),
	.w7(32'hba136a52),
	.w8(32'hbb14d6c1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82d750),
	.w1(32'hbaeb0016),
	.w2(32'hbb71b819),
	.w3(32'h3b6db4d6),
	.w4(32'h3ad69415),
	.w5(32'hbb43cb9d),
	.w6(32'hba18d133),
	.w7(32'hb841217f),
	.w8(32'hbba4ed96),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98c6c3),
	.w1(32'hbb1986de),
	.w2(32'hba8aaf06),
	.w3(32'hbb7550e4),
	.w4(32'h398fe537),
	.w5(32'hbb0be2e0),
	.w6(32'hbaf5cfb8),
	.w7(32'hbb069ef4),
	.w8(32'hbb2c6566),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15852a),
	.w1(32'hbb20962c),
	.w2(32'hbb311e61),
	.w3(32'hbb1e700b),
	.w4(32'hbb4fcd46),
	.w5(32'hba8fa5fe),
	.w6(32'hbae12608),
	.w7(32'hbb99f528),
	.w8(32'h3a83b6c4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71e979),
	.w1(32'hba5a08bd),
	.w2(32'hbb330ba7),
	.w3(32'hbae0e855),
	.w4(32'hba7d49f7),
	.w5(32'hbb4660c3),
	.w6(32'hba790f0d),
	.w7(32'hbb0aaa6f),
	.w8(32'hbac68bb2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3be48c),
	.w1(32'hbb3f4f5f),
	.w2(32'hbb62bb98),
	.w3(32'hbb148121),
	.w4(32'hbb2b4943),
	.w5(32'hba880605),
	.w6(32'h38dea179),
	.w7(32'hbacb332a),
	.w8(32'hba84ffa7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb50f58be),
	.w1(32'h393e9ffa),
	.w2(32'hba84568f),
	.w3(32'hb93151dd),
	.w4(32'h3ab98832),
	.w5(32'h3a4c06bd),
	.w6(32'hb81afbe4),
	.w7(32'hba846044),
	.w8(32'hba7cd1ca),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb751f21d),
	.w1(32'h3924bc98),
	.w2(32'hb8e67208),
	.w3(32'h3adea624),
	.w4(32'h3b6e06a8),
	.w5(32'hbb4ebee6),
	.w6(32'h396235a4),
	.w7(32'hb95ee11a),
	.w8(32'h3b240dd2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2584f2),
	.w1(32'h3b23b8a6),
	.w2(32'h3af5bbca),
	.w3(32'hbb3a253b),
	.w4(32'hba054ffa),
	.w5(32'h3b0a8c2e),
	.w6(32'h3b343773),
	.w7(32'h3aadea62),
	.w8(32'h3b62e33b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b596e16),
	.w1(32'h3b9d5e7a),
	.w2(32'h3a8d2464),
	.w3(32'h3a74c153),
	.w4(32'hb9648255),
	.w5(32'hb6fe96e8),
	.w6(32'h3ae0ca3e),
	.w7(32'hba89a12f),
	.w8(32'hb9f30031),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a938e),
	.w1(32'hb9e28fca),
	.w2(32'h3a331bfb),
	.w3(32'hb9bc55fe),
	.w4(32'h38e39901),
	.w5(32'hba8a600c),
	.w6(32'hb9d3866c),
	.w7(32'hba282a21),
	.w8(32'hb9bfa0fd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1aad9d),
	.w1(32'h39458ee3),
	.w2(32'hba8ed1a0),
	.w3(32'h395a2ee5),
	.w4(32'hbadb42ab),
	.w5(32'h3a236eb0),
	.w6(32'h3b13898a),
	.w7(32'hba037da5),
	.w8(32'h3a2f70a2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c5e4),
	.w1(32'h3a413bd8),
	.w2(32'h3a96c036),
	.w3(32'h3aa78d73),
	.w4(32'h3a393c47),
	.w5(32'hbb26e6a6),
	.w6(32'h3a971f38),
	.w7(32'h3b1eb748),
	.w8(32'hbb2838d8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f7fbb),
	.w1(32'hbbe77f57),
	.w2(32'hbbd33c1f),
	.w3(32'hbb98f326),
	.w4(32'hbbb0b800),
	.w5(32'hbacee80d),
	.w6(32'hbb568583),
	.w7(32'hbbc3da0f),
	.w8(32'hba805428),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfd197),
	.w1(32'h3ad789f3),
	.w2(32'h3a75a65e),
	.w3(32'h3aa53d3f),
	.w4(32'h3adcbcd2),
	.w5(32'h3a8ebd38),
	.w6(32'h3af202c6),
	.w7(32'h3a7d1802),
	.w8(32'h3b332473),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b310457),
	.w1(32'h3ab786ac),
	.w2(32'h39027189),
	.w3(32'h3a4aaeeb),
	.w4(32'hbb0cc449),
	.w5(32'hba5c65db),
	.w6(32'h3b996e8c),
	.w7(32'h3abfdb72),
	.w8(32'hba0cfdd7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24086d),
	.w1(32'hba8af1e1),
	.w2(32'hbafb45c8),
	.w3(32'hb8836ff3),
	.w4(32'hbab0b2e8),
	.w5(32'h3bcca640),
	.w6(32'h39f68ecb),
	.w7(32'hbb00d3f5),
	.w8(32'h3bb795d6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd6256),
	.w1(32'h3bb4d1f1),
	.w2(32'h3b99305e),
	.w3(32'h3b9ce72c),
	.w4(32'h3bad81c1),
	.w5(32'hbb592037),
	.w6(32'h3b7bf326),
	.w7(32'h3b6f0e5d),
	.w8(32'hbb57f509),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c3160),
	.w1(32'hbb5fc866),
	.w2(32'hbb4e906e),
	.w3(32'hbb79c61a),
	.w4(32'hbb2c47b7),
	.w5(32'h3b2bb957),
	.w6(32'hbb841d9e),
	.w7(32'hbb58ced8),
	.w8(32'h3b08d565),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b45df),
	.w1(32'h3b1f9f32),
	.w2(32'h3aae63ad),
	.w3(32'h3af323a9),
	.w4(32'h3a5db36c),
	.w5(32'h3a560769),
	.w6(32'h3a9a162d),
	.w7(32'hb92a99d8),
	.w8(32'h3abe11d0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a970b),
	.w1(32'hbb81dd87),
	.w2(32'hba4e1f19),
	.w3(32'hbb836455),
	.w4(32'hbad777ee),
	.w5(32'hbaa3607d),
	.w6(32'hbb2fbecc),
	.w7(32'hb995740d),
	.w8(32'hba8acede),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b3a96),
	.w1(32'h38e87620),
	.w2(32'hb890e0e5),
	.w3(32'hb8863bc6),
	.w4(32'hba4c2044),
	.w5(32'h3a4f4e04),
	.w6(32'h3b17e7ec),
	.w7(32'h3ac07c74),
	.w8(32'hb98c7473),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42c12b),
	.w1(32'hbb0f5540),
	.w2(32'hbaf1087c),
	.w3(32'h3b094757),
	.w4(32'hba00ab0e),
	.w5(32'hbb863296),
	.w6(32'h3a003c74),
	.w7(32'hba3c8e26),
	.w8(32'hbb7fe491),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402311),
	.w1(32'hbb18cf65),
	.w2(32'hbbb5aca8),
	.w3(32'hbb158c53),
	.w4(32'hbb6120ff),
	.w5(32'hbb4a0ed9),
	.w6(32'hbad87ba8),
	.w7(32'hbba53179),
	.w8(32'hbae631a1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fff9e),
	.w1(32'h39d078b7),
	.w2(32'h39256468),
	.w3(32'hba0b757a),
	.w4(32'hb9b8d9ee),
	.w5(32'hbae7850c),
	.w6(32'h39ec8e0a),
	.w7(32'hb979e1e6),
	.w8(32'hba464623),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7cfd3),
	.w1(32'hbb1aae6b),
	.w2(32'hbb4ec8bc),
	.w3(32'hbb624411),
	.w4(32'hbb03211a),
	.w5(32'hb9e1eae8),
	.w6(32'hbb07750b),
	.w7(32'hbb19251d),
	.w8(32'hb93dfbab),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0022c4),
	.w1(32'hb9b8e640),
	.w2(32'h39edceab),
	.w3(32'hb9f1b912),
	.w4(32'h3a999c6a),
	.w5(32'hbab01e08),
	.w6(32'hb93660db),
	.w7(32'h3a9808a6),
	.w8(32'hba8e72e6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18a1ae),
	.w1(32'hbaed3bd7),
	.w2(32'hbabace50),
	.w3(32'hbb03a5cc),
	.w4(32'hbaba6cb4),
	.w5(32'h3b1d1b1f),
	.w6(32'hbb23ac27),
	.w7(32'hbb237fd7),
	.w8(32'h3af9eeab),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46425b),
	.w1(32'h3b21e14b),
	.w2(32'h3b051ec0),
	.w3(32'h3b3734ea),
	.w4(32'h3b17acc0),
	.w5(32'h3a650323),
	.w6(32'h3af6d8a5),
	.w7(32'h3ae7db4c),
	.w8(32'h3adf9c5f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d2524),
	.w1(32'h3b61863e),
	.w2(32'h3b12ae7f),
	.w3(32'h3a5a64e6),
	.w4(32'h3b3ff65b),
	.w5(32'hba076092),
	.w6(32'h3adbfd70),
	.w7(32'h3b603a7d),
	.w8(32'h3b73687e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4585ea),
	.w1(32'h3b07005b),
	.w2(32'h3ac7dff7),
	.w3(32'hb9bd7304),
	.w4(32'h3a1ffaf0),
	.w5(32'hbab02dbc),
	.w6(32'h3b3390e6),
	.w7(32'h3acad3ae),
	.w8(32'hbab4716e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3821ee7f),
	.w1(32'h383bc2c2),
	.w2(32'hbaa362db),
	.w3(32'hbacc00e7),
	.w4(32'hbb8912da),
	.w5(32'hbb1d47cb),
	.w6(32'h3a36ca19),
	.w7(32'hbaefeb30),
	.w8(32'hbaacedc1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fd927e),
	.w1(32'hbb06334c),
	.w2(32'hbb1524b9),
	.w3(32'hbb2f5f0d),
	.w4(32'hbab8cf58),
	.w5(32'hbb06e8dc),
	.w6(32'hba85451d),
	.w7(32'hb9bfcda3),
	.w8(32'hba8116a9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2581b5),
	.w1(32'hbad2e59e),
	.w2(32'hba6633d5),
	.w3(32'hbb1369f4),
	.w4(32'hbaa62bb0),
	.w5(32'hbb5dfc75),
	.w6(32'hbaf41bbd),
	.w7(32'hbb02a468),
	.w8(32'hbaa34dce),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c0a9e),
	.w1(32'hba61322b),
	.w2(32'hba46caef),
	.w3(32'hbb6d7cbd),
	.w4(32'hbb15ea84),
	.w5(32'hbb2c1e32),
	.w6(32'hbb4fd62d),
	.w7(32'hbacfed71),
	.w8(32'hbafd7e23),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf2f8f),
	.w1(32'hbac3b1be),
	.w2(32'hbae6213f),
	.w3(32'hba3400bb),
	.w4(32'h39a88c0d),
	.w5(32'h3a368c0b),
	.w6(32'hba28289c),
	.w7(32'hba41e2a9),
	.w8(32'h399b4497),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bb1a4),
	.w1(32'hbb299d13),
	.w2(32'hbb2ef509),
	.w3(32'h3a551f77),
	.w4(32'hbb1628b4),
	.w5(32'hbb1d646f),
	.w6(32'h380225c3),
	.w7(32'hbb51f408),
	.w8(32'hbad0bfcc),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68228c),
	.w1(32'hb9a7a4f3),
	.w2(32'h3a92b524),
	.w3(32'hbb0ae1e9),
	.w4(32'h38435b12),
	.w5(32'hbb0bbac6),
	.w6(32'hbaf47ee0),
	.w7(32'h39bac0c3),
	.w8(32'hbb437cad),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb018a10),
	.w1(32'hbb77e415),
	.w2(32'hbae97397),
	.w3(32'hbb6efd57),
	.w4(32'hbb390d6e),
	.w5(32'hba3d389d),
	.w6(32'hbb88761b),
	.w7(32'hbb209b88),
	.w8(32'h37f0b89a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3c38d),
	.w1(32'hbb3c1317),
	.w2(32'hbb6b21a8),
	.w3(32'hbb0fc036),
	.w4(32'hbaf394bd),
	.w5(32'hb9fa1e18),
	.w6(32'h3a40a3a7),
	.w7(32'hbb6965c0),
	.w8(32'hba365aac),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af3b90),
	.w1(32'h38f9a7a5),
	.w2(32'h3a23bfaf),
	.w3(32'h3a5cec52),
	.w4(32'h3b01f6f2),
	.w5(32'hbaf04389),
	.w6(32'hb9a17695),
	.w7(32'hb7f5c4aa),
	.w8(32'hbae05540),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bce6ef),
	.w1(32'hb827f2e6),
	.w2(32'h3a7b20cd),
	.w3(32'hbb25b34d),
	.w4(32'hba6d6b4f),
	.w5(32'h3a021431),
	.w6(32'h3a432252),
	.w7(32'h3acf45cd),
	.w8(32'h388bdebe),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96352a),
	.w1(32'h3b926369),
	.w2(32'h3b30f8f8),
	.w3(32'h39ceef12),
	.w4(32'h3a9d7adb),
	.w5(32'hbb12b64d),
	.w6(32'h3aaade3f),
	.w7(32'h3a22e33d),
	.w8(32'hbb0e6eb2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba536cd9),
	.w1(32'hba0ed6f3),
	.w2(32'hba6e3b68),
	.w3(32'hbb18461b),
	.w4(32'hbb2529d3),
	.w5(32'h3b11b58a),
	.w6(32'hba454fa8),
	.w7(32'hbb3d334a),
	.w8(32'h3abd7642),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9894d1),
	.w1(32'hba7dcdd0),
	.w2(32'hbb278820),
	.w3(32'h3b31b17d),
	.w4(32'h39b26322),
	.w5(32'hbb2f8874),
	.w6(32'h3b2317e9),
	.w7(32'hbb8e2835),
	.w8(32'hbb22dcfa),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143346),
	.w1(32'hbb1ac6e1),
	.w2(32'hbade876d),
	.w3(32'hbb0a2686),
	.w4(32'hbade7177),
	.w5(32'hbab1fd59),
	.w6(32'hbafc26be),
	.w7(32'hbadfbaf9),
	.w8(32'hbad4ef77),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafadd8d),
	.w1(32'hbb038cf3),
	.w2(32'hba91d346),
	.w3(32'hba91ad24),
	.w4(32'hba9a51ee),
	.w5(32'hbb03ff88),
	.w6(32'hbafff7e6),
	.w7(32'hbab103bd),
	.w8(32'hbb20cc90),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab914c4),
	.w1(32'hbae1cb3e),
	.w2(32'hba870d0a),
	.w3(32'hba512de8),
	.w4(32'hbaf35c24),
	.w5(32'hb932b94b),
	.w6(32'hba82f206),
	.w7(32'hbaccc2c5),
	.w8(32'hba79cc32),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba237e),
	.w1(32'hba880822),
	.w2(32'h398e5dd8),
	.w3(32'hbadc8e92),
	.w4(32'hbb0dd3c0),
	.w5(32'h3b117e81),
	.w6(32'hbb23c767),
	.w7(32'hbabe0a44),
	.w8(32'h3b41109b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebc59b),
	.w1(32'h3abaafbd),
	.w2(32'hba0572ff),
	.w3(32'h3a428842),
	.w4(32'hba5aeb0b),
	.w5(32'hbad37301),
	.w6(32'h3b26bb2c),
	.w7(32'hb9f1c8bf),
	.w8(32'hbb063175),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b36e5),
	.w1(32'hbaedd82e),
	.w2(32'h3a88af05),
	.w3(32'hba6e49b0),
	.w4(32'h393766f1),
	.w5(32'hbb32ae29),
	.w6(32'hbb6ffbe9),
	.w7(32'hba04b8c1),
	.w8(32'hbb01ac93),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade670c),
	.w1(32'hba8d119a),
	.w2(32'hba23e9fe),
	.w3(32'hbb1fc442),
	.w4(32'hbaee8008),
	.w5(32'hb9e5189a),
	.w6(32'hba585e7b),
	.w7(32'hba5a4f14),
	.w8(32'hbabb7c57),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277a94),
	.w1(32'hbb2525af),
	.w2(32'hbb178f88),
	.w3(32'hba95bbd0),
	.w4(32'hbaaa02f3),
	.w5(32'h3aa02e2b),
	.w6(32'hbb1859d4),
	.w7(32'hbb04631e),
	.w8(32'h3a6878d9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ace92d),
	.w1(32'h3a66b370),
	.w2(32'h3a1b80ac),
	.w3(32'h3b7015f7),
	.w4(32'h3a85264d),
	.w5(32'h3a0ea41c),
	.w6(32'h3b3f3a5f),
	.w7(32'h3a3b2b70),
	.w8(32'hba7d00b8),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f09b7),
	.w1(32'hbb19dd0b),
	.w2(32'hbb3432f1),
	.w3(32'hb8c99d5e),
	.w4(32'hba4029f4),
	.w5(32'h39dd23f8),
	.w6(32'hba47fdb1),
	.w7(32'hbacffb78),
	.w8(32'h3b18c8f8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06a6f8),
	.w1(32'hb99d1f2d),
	.w2(32'h39c0ebe2),
	.w3(32'h3b22b317),
	.w4(32'h3abc24e6),
	.w5(32'hbb41b7f5),
	.w6(32'h3b2239ff),
	.w7(32'h3b66b597),
	.w8(32'hbb1ced49),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10c70f),
	.w1(32'hbaa5f2dd),
	.w2(32'hbb46debf),
	.w3(32'hbb23d992),
	.w4(32'hbb0c40b8),
	.w5(32'hbaeb6c33),
	.w6(32'hba2d93c8),
	.w7(32'hbae26aa1),
	.w8(32'hba1849fd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0cc09),
	.w1(32'hb98a2d85),
	.w2(32'hbadfc128),
	.w3(32'hba8dd9dd),
	.w4(32'hba29e007),
	.w5(32'h3b378714),
	.w6(32'h384f7957),
	.w7(32'h387064fb),
	.w8(32'h3b3d64de),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f925e),
	.w1(32'h3aed6b03),
	.w2(32'h3980fc19),
	.w3(32'h3b15fe3e),
	.w4(32'h39a25b42),
	.w5(32'h39ebb46c),
	.w6(32'h3b349f9d),
	.w7(32'h39821eac),
	.w8(32'h3a0c425e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1f8c4),
	.w1(32'hba8720d8),
	.w2(32'h3a17345d),
	.w3(32'hba71ab8e),
	.w4(32'h393add51),
	.w5(32'h3b3d8b39),
	.w6(32'hbb06b52f),
	.w7(32'h3a2a2fb9),
	.w8(32'h3b1aa96d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12b523),
	.w1(32'h3b20c698),
	.w2(32'hba3e3584),
	.w3(32'h3a763e7c),
	.w4(32'hba178d89),
	.w5(32'hbb5d4bbe),
	.w6(32'h3af3a08f),
	.w7(32'hba1b5a11),
	.w8(32'hbb77a602),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62e64b),
	.w1(32'hbb8556c4),
	.w2(32'hba7be455),
	.w3(32'hbba358b9),
	.w4(32'hbaffba81),
	.w5(32'hbb4bf531),
	.w6(32'hbbd294fa),
	.w7(32'hbb0b6d5d),
	.w8(32'hbba967f2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba526a5),
	.w1(32'hbbe4e5de),
	.w2(32'hbbcf7707),
	.w3(32'hbb643f5c),
	.w4(32'hbb5adbf5),
	.w5(32'h39e6465e),
	.w6(32'hbb9eaa2a),
	.w7(32'hbb9f0e05),
	.w8(32'h38fb458c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3664f58c),
	.w1(32'hba915a23),
	.w2(32'hba4e8185),
	.w3(32'hba79431a),
	.w4(32'hba485de9),
	.w5(32'hbb0e2c4b),
	.w6(32'hbaa14546),
	.w7(32'hba547447),
	.w8(32'hbb7c52d7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd8d51),
	.w1(32'hba0053c1),
	.w2(32'h3a0a1664),
	.w3(32'hbaf39acb),
	.w4(32'h39edab50),
	.w5(32'h3ac04094),
	.w6(32'hbacfce69),
	.w7(32'h3a1289ad),
	.w8(32'hba387499),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4e749),
	.w1(32'hbb270cdb),
	.w2(32'hbb09dbbb),
	.w3(32'h3b07e4b3),
	.w4(32'h3a6b1c6a),
	.w5(32'hbaabdb6d),
	.w6(32'h3aed2d26),
	.w7(32'h3a713854),
	.w8(32'hb9cfe934),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942a686),
	.w1(32'h3afc2798),
	.w2(32'h3ae1ea9d),
	.w3(32'hbab7f7ff),
	.w4(32'hbade2d8a),
	.w5(32'hb955db27),
	.w6(32'hba2796a1),
	.w7(32'hb9ba9c4a),
	.w8(32'hbb2c8d52),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ec552),
	.w1(32'hba475473),
	.w2(32'hba47746a),
	.w3(32'hba9af249),
	.w4(32'h3a31bd2f),
	.w5(32'h3bcfcf16),
	.w6(32'hbaff9dc6),
	.w7(32'hbaaefea1),
	.w8(32'hb88781dd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdb713),
	.w1(32'hbb3e6000),
	.w2(32'h3ac485c8),
	.w3(32'h3b09e3a7),
	.w4(32'h3bc0d034),
	.w5(32'hbc1b26ee),
	.w6(32'hbb81aca7),
	.w7(32'h3b0a2515),
	.w8(32'h3b192b21),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3623d9),
	.w1(32'h3a7fac30),
	.w2(32'hbb5afc53),
	.w3(32'hbbda073e),
	.w4(32'hba8043b6),
	.w5(32'h3b96d22d),
	.w6(32'h3b84321f),
	.w7(32'h3a0bf1ab),
	.w8(32'hbbbf8ea5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcaa28),
	.w1(32'h3889cddb),
	.w2(32'hbabd8882),
	.w3(32'h3a54d80d),
	.w4(32'h3ae93983),
	.w5(32'h3ac7a8ad),
	.w6(32'hbc49db9a),
	.w7(32'hbb7b5227),
	.w8(32'h3c5d8f8c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30226a),
	.w1(32'h3b64dbbf),
	.w2(32'hbbc21625),
	.w3(32'h3b0ef4fd),
	.w4(32'hbb0d9f7f),
	.w5(32'h3a4f5deb),
	.w6(32'h3c894f0b),
	.w7(32'h3a6f31e9),
	.w8(32'hbb9d99ef),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bc0ae),
	.w1(32'hbbaaf23c),
	.w2(32'h3c1030de),
	.w3(32'hbc400e49),
	.w4(32'hbbfd7759),
	.w5(32'h3a03e401),
	.w6(32'hbc1fd99d),
	.w7(32'hbbf3217d),
	.w8(32'h3a855f82),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d653a),
	.w1(32'hbb6d54e6),
	.w2(32'hbb9063c3),
	.w3(32'h3aa39469),
	.w4(32'h3b6a9d3d),
	.w5(32'hba4a26c6),
	.w6(32'hba7c9b56),
	.w7(32'h3bb0a119),
	.w8(32'hbb878e6e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa92cd4),
	.w1(32'h3b3afd00),
	.w2(32'h3b8004c8),
	.w3(32'hbb9bb019),
	.w4(32'h3a885027),
	.w5(32'hbb013d22),
	.w6(32'hbba01bde),
	.w7(32'h3b245ae0),
	.w8(32'hbb43d0ba),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8b5f4),
	.w1(32'hbaaeb69a),
	.w2(32'hbb3cef13),
	.w3(32'hbb1e81f7),
	.w4(32'h39abeea1),
	.w5(32'hba83d5ec),
	.w6(32'hbbd45dd9),
	.w7(32'hbbb018c3),
	.w8(32'h398a04a8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c2e34),
	.w1(32'hbc3b9c47),
	.w2(32'hbadb56a1),
	.w3(32'hbb01266b),
	.w4(32'h3c01bc96),
	.w5(32'hbb124711),
	.w6(32'h3ba87da6),
	.w7(32'h3b83787f),
	.w8(32'hba840dec),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab80165),
	.w1(32'hbaeb1375),
	.w2(32'hbb1af6d0),
	.w3(32'hbbc278bf),
	.w4(32'hbb89323d),
	.w5(32'h3be099e6),
	.w6(32'hbb4e927f),
	.w7(32'hbbd12165),
	.w8(32'hbb344b21),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0c55e),
	.w1(32'hbb59a908),
	.w2(32'h3b8a4795),
	.w3(32'hba2683ce),
	.w4(32'h3bd36684),
	.w5(32'h3a42166b),
	.w6(32'hbc09fb89),
	.w7(32'h3b5c8bf9),
	.w8(32'hb9d84a35),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c2890),
	.w1(32'h3ae06b2c),
	.w2(32'h39c9d9b0),
	.w3(32'h3a28449b),
	.w4(32'hba4328be),
	.w5(32'hbb447eb3),
	.w6(32'hbb80c97c),
	.w7(32'hbb66627d),
	.w8(32'h3aae3095),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad317ee),
	.w1(32'hbac1d97c),
	.w2(32'h3b58fde2),
	.w3(32'hbbcc2632),
	.w4(32'hba17ae13),
	.w5(32'h3b8da4b0),
	.w6(32'hbb35e653),
	.w7(32'hba8d33b9),
	.w8(32'h3c8a58fd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca715e0),
	.w1(32'h3cbd6ee5),
	.w2(32'h3bb90af7),
	.w3(32'h3cdcffe4),
	.w4(32'h3c632b49),
	.w5(32'hbb10f057),
	.w6(32'h3cf5fc78),
	.w7(32'h3ae2b952),
	.w8(32'h3b07c404),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ee041),
	.w1(32'h3b646023),
	.w2(32'h3b3d12b7),
	.w3(32'hb9de1d5d),
	.w4(32'h3a1c6c1b),
	.w5(32'h3ca5e4c8),
	.w6(32'h3b6f6e9c),
	.w7(32'h3bf6fca7),
	.w8(32'h3ae7b29f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb68b8b),
	.w1(32'h3b9e2036),
	.w2(32'h3c2ae545),
	.w3(32'h3bc5035b),
	.w4(32'h3c19591f),
	.w5(32'hba634836),
	.w6(32'hba53305e),
	.w7(32'hba84a542),
	.w8(32'h3aac9440),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b538498),
	.w1(32'hbb2f1c97),
	.w2(32'hbb634886),
	.w3(32'h3aa1b53b),
	.w4(32'hbb709ba0),
	.w5(32'hba9875d7),
	.w6(32'hbaf5bda6),
	.w7(32'hbb053223),
	.w8(32'h3c330e8a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf2b5d),
	.w1(32'h3c4c51db),
	.w2(32'hbbd50bef),
	.w3(32'h3c9234d5),
	.w4(32'h3c6654da),
	.w5(32'h3ab738f9),
	.w6(32'h3cab843c),
	.w7(32'h3a2399bf),
	.w8(32'hb9fac2ec),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a007f1c),
	.w1(32'hb9e686b3),
	.w2(32'h3aa8ebcb),
	.w3(32'hbb55e185),
	.w4(32'hbb702d68),
	.w5(32'h3b8cbda0),
	.w6(32'hbb17fbf3),
	.w7(32'hbb7758d8),
	.w8(32'hbb4d037b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73e7ee),
	.w1(32'hbbf9ab48),
	.w2(32'hbb5d51b7),
	.w3(32'hbb4669a1),
	.w4(32'h3a2425d0),
	.w5(32'h3abff638),
	.w6(32'h3bab6391),
	.w7(32'h3b61f074),
	.w8(32'hbb32e615),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3fb29),
	.w1(32'hbb35dea8),
	.w2(32'h3ba492e3),
	.w3(32'hbb3c07e8),
	.w4(32'h3948a2ee),
	.w5(32'h39841488),
	.w6(32'hbba4e8f4),
	.w7(32'hbacff741),
	.w8(32'hb99cca75),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a277b),
	.w1(32'hbb3d72c5),
	.w2(32'hba88bf51),
	.w3(32'hbba5bab9),
	.w4(32'hbb920588),
	.w5(32'hbbec1b3c),
	.w6(32'hbba020fa),
	.w7(32'h3a1c69c9),
	.w8(32'h3b4b1f0c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f0eab),
	.w1(32'h3c8f4f52),
	.w2(32'h3beb70ad),
	.w3(32'h3ad0447d),
	.w4(32'hb9586427),
	.w5(32'hbaf54846),
	.w6(32'h3c2f8100),
	.w7(32'hbbc62aad),
	.w8(32'hbb17b501),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade4a66),
	.w1(32'h3b435f2f),
	.w2(32'hba733557),
	.w3(32'h3a1136d6),
	.w4(32'hbb902071),
	.w5(32'h3b71c4dd),
	.w6(32'hbb453444),
	.w7(32'hbabad178),
	.w8(32'h3bc12e2b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b473bfe),
	.w1(32'h3b8925a1),
	.w2(32'h3bfa4f5a),
	.w3(32'hba29cb85),
	.w4(32'hbb2b6702),
	.w5(32'hbba112c6),
	.w6(32'h3bcd9d0c),
	.w7(32'h3b3bdbf8),
	.w8(32'hbb49a913),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2609e4),
	.w1(32'hb9917c8b),
	.w2(32'hbac85f9d),
	.w3(32'hbaba9e6e),
	.w4(32'hbae73792),
	.w5(32'hbbaef4bb),
	.w6(32'hbb8da2f7),
	.w7(32'h3a66d775),
	.w8(32'h3b90f7e4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7f802),
	.w1(32'h3c1a51bf),
	.w2(32'h3b3ae8b3),
	.w3(32'hbc009d26),
	.w4(32'hbc00581a),
	.w5(32'hbb7c2300),
	.w6(32'h3ba6c806),
	.w7(32'h3b6a7f30),
	.w8(32'hbc588327),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33e27c),
	.w1(32'h3bbd1264),
	.w2(32'h3b78aca3),
	.w3(32'hbc553112),
	.w4(32'hbc4c69fe),
	.w5(32'hb9f4e57f),
	.w6(32'hbbcde809),
	.w7(32'hbc2dd72c),
	.w8(32'hba801c96),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb937ccd),
	.w1(32'hbb0de0f9),
	.w2(32'hba5137c0),
	.w3(32'hbb16892e),
	.w4(32'hbb7d79d3),
	.w5(32'h3c0a5aa7),
	.w6(32'hbabe3be1),
	.w7(32'hbaa56131),
	.w8(32'h3ae2e628),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a749012),
	.w1(32'hbb813aa9),
	.w2(32'hbb8c8685),
	.w3(32'h3c15741d),
	.w4(32'hba835d4d),
	.w5(32'hbb74bf10),
	.w6(32'hba066f24),
	.w7(32'hbb736951),
	.w8(32'h3af6bdf0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d81fc),
	.w1(32'hbab7075e),
	.w2(32'hbab77463),
	.w3(32'hbaced777),
	.w4(32'hbb5bab89),
	.w5(32'hbb045c3a),
	.w6(32'hbacfd286),
	.w7(32'hbb7b024a),
	.w8(32'hba40be1b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c40f2),
	.w1(32'hb995f4cd),
	.w2(32'hbb6f1044),
	.w3(32'hbb036761),
	.w4(32'hbb9b1d14),
	.w5(32'hbc216a66),
	.w6(32'hbab7e5de),
	.w7(32'hbaaad9ac),
	.w8(32'hba8d9f31),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dfc81),
	.w1(32'h3c8e28d2),
	.w2(32'h3b9ae6ff),
	.w3(32'hbbbb5a36),
	.w4(32'h3b033788),
	.w5(32'h3ac02d30),
	.w6(32'h3c3f1a2d),
	.w7(32'h3c13851d),
	.w8(32'hba940a72),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b3639),
	.w1(32'hbacc0e4e),
	.w2(32'h3a4b96f8),
	.w3(32'hbb48a0d4),
	.w4(32'hbb71903f),
	.w5(32'hbb82778e),
	.w6(32'hba3652a6),
	.w7(32'hb8d78dfd),
	.w8(32'h3c8903c1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02295d),
	.w1(32'hbc31434a),
	.w2(32'hbb405e86),
	.w3(32'hbc2b6499),
	.w4(32'h38856c2b),
	.w5(32'h3b7fbc72),
	.w6(32'h3c88cc16),
	.w7(32'h3c95fd70),
	.w8(32'h3b035400),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33fd07),
	.w1(32'h3b39a7b0),
	.w2(32'h3ac1586c),
	.w3(32'h3b002b4b),
	.w4(32'h3a6d297d),
	.w5(32'hbac069ca),
	.w6(32'h3aeeaf40),
	.w7(32'hba0bb4ad),
	.w8(32'h39104215),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cf7a0),
	.w1(32'h3902eb3c),
	.w2(32'hba179dc6),
	.w3(32'hbb066d8f),
	.w4(32'hbaf85e6b),
	.w5(32'hbb4d6dc9),
	.w6(32'hba4ced0c),
	.w7(32'hb80977b8),
	.w8(32'hba8bfa7a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d73b5),
	.w1(32'hbbaa718c),
	.w2(32'h3a4a48fd),
	.w3(32'hbbb6553e),
	.w4(32'hbb860309),
	.w5(32'h3a34eb98),
	.w6(32'hbb60808d),
	.w7(32'hbb759339),
	.w8(32'h3b0a45f4),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29e4fc),
	.w1(32'h3ac3c74f),
	.w2(32'h3ae99785),
	.w3(32'h393b5cf9),
	.w4(32'hb901129b),
	.w5(32'h3b7e8f1f),
	.w6(32'hb99033d4),
	.w7(32'h3a173681),
	.w8(32'h3ae44aae),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa617c9),
	.w1(32'h3abae175),
	.w2(32'h3ab01d3e),
	.w3(32'h3b05b277),
	.w4(32'h3a8451f9),
	.w5(32'h3b3f8611),
	.w6(32'h3aa951c5),
	.w7(32'hba74ae86),
	.w8(32'h3b716534),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a9cc7),
	.w1(32'h3b677f04),
	.w2(32'h3b2bc37c),
	.w3(32'hbac5fdb9),
	.w4(32'hbb256440),
	.w5(32'hba327eb9),
	.w6(32'h3bb8df10),
	.w7(32'h3ad2a87f),
	.w8(32'hba6e4752),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad4609),
	.w1(32'hbaba4ebf),
	.w2(32'h3ad0dbbd),
	.w3(32'hbb493392),
	.w4(32'hbb4c6bd5),
	.w5(32'hbbbf6e21),
	.w6(32'hbaea7505),
	.w7(32'hb9a1d2ee),
	.w8(32'h3b680174),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c6086),
	.w1(32'hba8a05a8),
	.w2(32'h39ee7eab),
	.w3(32'hba131c62),
	.w4(32'h3acf747a),
	.w5(32'hbc23c49f),
	.w6(32'h3b8ef295),
	.w7(32'h3b8f73f0),
	.w8(32'h3a6a757b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1a181),
	.w1(32'hbc7b2cc1),
	.w2(32'hbc0d9c99),
	.w3(32'hbb4b3ebc),
	.w4(32'h3ac99e54),
	.w5(32'h3a84de8a),
	.w6(32'h3a7ddf57),
	.w7(32'hb8fade5d),
	.w8(32'h39daf964),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c153e),
	.w1(32'h389794e8),
	.w2(32'h3b4505af),
	.w3(32'h398468d9),
	.w4(32'h3a5b2cca),
	.w5(32'h3ad000d4),
	.w6(32'hbb2c21cb),
	.w7(32'h3b228e49),
	.w8(32'hbae3a677),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe795d1),
	.w1(32'hbb806507),
	.w2(32'hbb1358d4),
	.w3(32'hbb49c279),
	.w4(32'hbb6cda4e),
	.w5(32'hba25fd61),
	.w6(32'h3a134430),
	.w7(32'hba86409e),
	.w8(32'h3b53c2ed),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31049d),
	.w1(32'h3b943c4f),
	.w2(32'h3b093189),
	.w3(32'hba5c9671),
	.w4(32'hb9a636a0),
	.w5(32'hbba65cef),
	.w6(32'h3ad811b0),
	.w7(32'h3b20f4d4),
	.w8(32'hba806bb7),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c925c),
	.w1(32'h3a3b9dee),
	.w2(32'h3aea9706),
	.w3(32'hbb5602c4),
	.w4(32'h39dd8e47),
	.w5(32'hbaa923fa),
	.w6(32'hba919995),
	.w7(32'h3ab2ec42),
	.w8(32'h3c113f26),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38efb5d3),
	.w1(32'h3b0ebfd5),
	.w2(32'hba13d50d),
	.w3(32'hba066539),
	.w4(32'h3aa19c44),
	.w5(32'h3b4b4f3e),
	.w6(32'h3b9a5888),
	.w7(32'h3bcb93e3),
	.w8(32'hbbe0d129),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5d334),
	.w1(32'h3be93891),
	.w2(32'hbacf47bc),
	.w3(32'h3b75d2da),
	.w4(32'hbad762b9),
	.w5(32'hbb0fb024),
	.w6(32'hbbd08819),
	.w7(32'hbc2f1bde),
	.w8(32'hbb34ff14),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48f5f3),
	.w1(32'hba1ff76a),
	.w2(32'h3a9457c7),
	.w3(32'hbb881c65),
	.w4(32'hbb0fb2a4),
	.w5(32'h3b46ed6a),
	.w6(32'hbb1283dd),
	.w7(32'h3abe1aca),
	.w8(32'hbb2ac166),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2e08a),
	.w1(32'hbb3e6c75),
	.w2(32'hba44f294),
	.w3(32'hbb0a4aa0),
	.w4(32'hba3c9820),
	.w5(32'h3c3ece66),
	.w6(32'hbbc5eab0),
	.w7(32'hbb46d9fc),
	.w8(32'hba8d43aa),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba947b),
	.w1(32'hbbc937f2),
	.w2(32'h3b42d6d1),
	.w3(32'h3b864b1a),
	.w4(32'h3c1f59da),
	.w5(32'hbb2b1a11),
	.w6(32'hbabf339f),
	.w7(32'hb9c144e1),
	.w8(32'h39694b87),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85c7bc),
	.w1(32'hbb824889),
	.w2(32'hb9b8f47b),
	.w3(32'hba29286e),
	.w4(32'h39ab5c61),
	.w5(32'h3b9857ae),
	.w6(32'h3c0084fd),
	.w7(32'hbbb8075b),
	.w8(32'h3bfe181c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb293c2c),
	.w1(32'h3bc548e3),
	.w2(32'hbb573255),
	.w3(32'h3a775847),
	.w4(32'h3b2a6c27),
	.w5(32'h3a2abde7),
	.w6(32'h3be4501e),
	.w7(32'h3ac50939),
	.w8(32'hbb7233e8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0886a),
	.w1(32'hbb12919c),
	.w2(32'hba229d9c),
	.w3(32'hbb18c3f7),
	.w4(32'hbb8ba496),
	.w5(32'h3ab73ecb),
	.w6(32'hbc22e0d1),
	.w7(32'hbb857afc),
	.w8(32'hb89d0eaa),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18f521),
	.w1(32'hbbb3eb68),
	.w2(32'hba761cf2),
	.w3(32'hbbba309e),
	.w4(32'hbad98114),
	.w5(32'hba42f2af),
	.w6(32'hbbf49315),
	.w7(32'h39393678),
	.w8(32'h3ad06da9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b4e98),
	.w1(32'h3abd1672),
	.w2(32'hb8c0e457),
	.w3(32'h3a6aa719),
	.w4(32'hb995654b),
	.w5(32'hbc02d718),
	.w6(32'hbb29668b),
	.w7(32'hbae0f624),
	.w8(32'hbc5ff5f3),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f8aef),
	.w1(32'hbc2aeb44),
	.w2(32'hbc0ff00b),
	.w3(32'hbc160ebb),
	.w4(32'hbbe78a8f),
	.w5(32'hbb43cea3),
	.w6(32'hbc08d43a),
	.w7(32'hbc1c3ab5),
	.w8(32'hbb9ecd21),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf6f9f),
	.w1(32'hbb164e20),
	.w2(32'hbbed746d),
	.w3(32'h3b0ac289),
	.w4(32'hb98fe089),
	.w5(32'h3acca11f),
	.w6(32'hbba7bbc4),
	.w7(32'hbaa2241f),
	.w8(32'h3b39b5ce),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2d7cf),
	.w1(32'hbace8ed2),
	.w2(32'hba8ab5fe),
	.w3(32'h3b9cdce9),
	.w4(32'h38d7b699),
	.w5(32'hbb93b14a),
	.w6(32'h3bd9d15f),
	.w7(32'hbacd8857),
	.w8(32'h3c195efa),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48047b),
	.w1(32'h3ca682e6),
	.w2(32'h3c1a7d1b),
	.w3(32'hbbb310fc),
	.w4(32'hbbaa44a1),
	.w5(32'h3affa9e1),
	.w6(32'h3c633aa4),
	.w7(32'h3bf99469),
	.w8(32'h3c690eb2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af930be),
	.w1(32'hb9be668d),
	.w2(32'hbc166564),
	.w3(32'h3cace22d),
	.w4(32'hbb21d1cb),
	.w5(32'hbb4ffb4c),
	.w6(32'hbac1e799),
	.w7(32'hbc1d9e46),
	.w8(32'hbb09b18c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec0574),
	.w1(32'hbc0d79b6),
	.w2(32'hbb3b3b73),
	.w3(32'hbba749bb),
	.w4(32'hbb147667),
	.w5(32'h3c86af89),
	.w6(32'hbb552dcf),
	.w7(32'h3a13da94),
	.w8(32'h3c003cb8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a7f22),
	.w1(32'h3c7a25f5),
	.w2(32'h3ca2ee0d),
	.w3(32'h3c055cbc),
	.w4(32'h3b12d340),
	.w5(32'hbbc8c6fe),
	.w6(32'h3c4e3e83),
	.w7(32'h3c6f0187),
	.w8(32'h3a25551e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac08eae),
	.w1(32'hbac00aeb),
	.w2(32'hbbea9fdb),
	.w3(32'hbae671c1),
	.w4(32'h3b6ee835),
	.w5(32'h3c156508),
	.w6(32'h3ab2b2c5),
	.w7(32'hbb8ee208),
	.w8(32'hbb013c02),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb29b1a),
	.w1(32'hbbf6cc7e),
	.w2(32'hbbc7c4d1),
	.w3(32'h3bdb877e),
	.w4(32'h3b2fb989),
	.w5(32'h3b71b329),
	.w6(32'hbb23f2ac),
	.w7(32'h3b5f4824),
	.w8(32'hbad29ca5),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd92974),
	.w1(32'h3a9cf33b),
	.w2(32'h3baccb77),
	.w3(32'hbba8e155),
	.w4(32'hbaf115b2),
	.w5(32'hbb7efb05),
	.w6(32'hbbfbcbdd),
	.w7(32'hba7e711a),
	.w8(32'hba02c154),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd9709),
	.w1(32'hbb0d414a),
	.w2(32'hbb57f778),
	.w3(32'hbb9494ef),
	.w4(32'h3b0a5ca1),
	.w5(32'h3aac35ae),
	.w6(32'h3ab48719),
	.w7(32'hbac3b8a6),
	.w8(32'h3a7c9dd7),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9389e0),
	.w1(32'hbbdb38ee),
	.w2(32'hbb342e4c),
	.w3(32'hbab1bf89),
	.w4(32'h3bdfe4b8),
	.w5(32'hbc0f0c0a),
	.w6(32'hbacb4676),
	.w7(32'h3b5f02dd),
	.w8(32'hbc1bc526),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1809e1),
	.w1(32'hbbf1be1d),
	.w2(32'hbb3a55b5),
	.w3(32'hbc26a49f),
	.w4(32'hbc333468),
	.w5(32'hbb58b75b),
	.w6(32'hbc1d1713),
	.w7(32'hbc228ed5),
	.w8(32'hbb90e189),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7efe0),
	.w1(32'hbb12e60a),
	.w2(32'hbaf9a7d4),
	.w3(32'hbbe1e550),
	.w4(32'hbbda2328),
	.w5(32'h3ad59176),
	.w6(32'hbbebc778),
	.w7(32'hbb62bff6),
	.w8(32'h3a212994),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd63fc2),
	.w1(32'h3bdcfff2),
	.w2(32'h3b8d0796),
	.w3(32'hbbb5cf37),
	.w4(32'h3b5c0e3d),
	.w5(32'hbb1176c5),
	.w6(32'h3b1de4d5),
	.w7(32'h3a803d6b),
	.w8(32'h3beb4902),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aa5ed),
	.w1(32'hbb8c8e3c),
	.w2(32'hbba22111),
	.w3(32'hbb5b0f1d),
	.w4(32'hbac55ff8),
	.w5(32'hbb81f229),
	.w6(32'h3babce72),
	.w7(32'h3b59f5bb),
	.w8(32'hbb4797fe),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31a5eb),
	.w1(32'h3b06c58c),
	.w2(32'h3b123be6),
	.w3(32'hba8de847),
	.w4(32'hbb29a69c),
	.w5(32'hb99d0f61),
	.w6(32'hbb429d2c),
	.w7(32'hba0b0a77),
	.w8(32'hbbceb88b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1270ce),
	.w1(32'hbb4e0a1e),
	.w2(32'h380cce7b),
	.w3(32'h3a0045a0),
	.w4(32'hba191d85),
	.w5(32'h3b918cb2),
	.w6(32'hbbaea375),
	.w7(32'hbb9df490),
	.w8(32'h3b16b6ee),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae477d),
	.w1(32'hbb1d1607),
	.w2(32'hba7bac91),
	.w3(32'h3b34a14d),
	.w4(32'h3b398eea),
	.w5(32'h3aec0382),
	.w6(32'hbb21de30),
	.w7(32'h3ab5cf3f),
	.w8(32'h3b884d28),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a306ad8),
	.w1(32'h3af1e765),
	.w2(32'h3a85c026),
	.w3(32'h38bd8624),
	.w4(32'hbb37ec96),
	.w5(32'hba3a989a),
	.w6(32'h3a1a1a9d),
	.w7(32'h3b06b62f),
	.w8(32'h3b3bbb8d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02e294),
	.w1(32'h3b8693b4),
	.w2(32'h3b55ef6d),
	.w3(32'h3b0546f1),
	.w4(32'h3989da05),
	.w5(32'hba40389b),
	.w6(32'hbaa70177),
	.w7(32'hba1b89ff),
	.w8(32'hb93a17d6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65a7df),
	.w1(32'hbb86828c),
	.w2(32'hbb1e36f0),
	.w3(32'hbbbb6e6b),
	.w4(32'hbb9a88ac),
	.w5(32'hbbda8340),
	.w6(32'hbbf807a6),
	.w7(32'hba2cc7a3),
	.w8(32'h3b7639d7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f953c),
	.w1(32'hbc0183ad),
	.w2(32'hbc3b9e5b),
	.w3(32'h3a8b7320),
	.w4(32'h3c2e324b),
	.w5(32'h39a686b8),
	.w6(32'h3bb6ddd6),
	.w7(32'hb968c93c),
	.w8(32'hba856b26),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac7cb9),
	.w1(32'h3aa75d45),
	.w2(32'hb88b3697),
	.w3(32'hbb2bb608),
	.w4(32'h3b072019),
	.w5(32'hbca04c39),
	.w6(32'hba11c2fe),
	.w7(32'hbb64aee4),
	.w8(32'hbac39ecc),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad035e8),
	.w1(32'h3b96d473),
	.w2(32'hbc16464d),
	.w3(32'hbc085bdc),
	.w4(32'hbbfe2302),
	.w5(32'hbb0e4397),
	.w6(32'h3c5ebfc6),
	.w7(32'hbb5f2016),
	.w8(32'hbbcc9054),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca8c8),
	.w1(32'hbc093fc7),
	.w2(32'hbb898008),
	.w3(32'h388b17bd),
	.w4(32'hbb587ed9),
	.w5(32'hbc6baba1),
	.w6(32'hbb602cce),
	.w7(32'hbb30293f),
	.w8(32'hbc68a15c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b6b90),
	.w1(32'hbc27904f),
	.w2(32'hbc305f2b),
	.w3(32'hbc59fb51),
	.w4(32'hbc82f4f8),
	.w5(32'h3b894a14),
	.w6(32'hbc4ec873),
	.w7(32'hbc81f72e),
	.w8(32'h3c1520c3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bf3e6),
	.w1(32'h3c7a0187),
	.w2(32'h3c5728c7),
	.w3(32'hbc0a63b4),
	.w4(32'hbc3245f4),
	.w5(32'h3b52c3fd),
	.w6(32'h3be0d037),
	.w7(32'h3a85d103),
	.w8(32'h3a25b333),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb191470),
	.w1(32'h3b675574),
	.w2(32'h3bf481d7),
	.w3(32'hba20fd54),
	.w4(32'hbbe0856b),
	.w5(32'hbc15ce81),
	.w6(32'hbb43313b),
	.w7(32'hbb964e25),
	.w8(32'hbbad8f7b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c7791),
	.w1(32'h3b73c8ec),
	.w2(32'hbb0fc2e0),
	.w3(32'hbb1cdaf4),
	.w4(32'hbba456e3),
	.w5(32'hba6173ce),
	.w6(32'h3b8d3bcf),
	.w7(32'h3a13e74d),
	.w8(32'hb9f02fd6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac38ec7),
	.w1(32'hbb6b857c),
	.w2(32'hbb147f46),
	.w3(32'hbbcbce3c),
	.w4(32'hbbbeb189),
	.w5(32'h3bfa9ace),
	.w6(32'hbc054661),
	.w7(32'hbaf9ee50),
	.w8(32'h3ac78aea),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb8a9d),
	.w1(32'hbaccaf4e),
	.w2(32'h383fba5f),
	.w3(32'hba47cdb9),
	.w4(32'hba84188b),
	.w5(32'hbb485b4c),
	.w6(32'hbb710ab4),
	.w7(32'hbaa4fe9f),
	.w8(32'hbb3caee5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb535e93),
	.w1(32'hbb0bca55),
	.w2(32'hbadfe74f),
	.w3(32'hbb59608d),
	.w4(32'hb8a75fff),
	.w5(32'hbb5452c4),
	.w6(32'hbb3f8cba),
	.w7(32'hbb00ee25),
	.w8(32'hbb9499f6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfd594),
	.w1(32'hbbb32e63),
	.w2(32'hbb459b42),
	.w3(32'hbb9a31cd),
	.w4(32'hbbd50aa5),
	.w5(32'h3abf8565),
	.w6(32'hbba11398),
	.w7(32'hbb6cfc9c),
	.w8(32'h3cbc77e4),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f9f4d),
	.w1(32'hb9b82083),
	.w2(32'hbb50454c),
	.w3(32'h3b6a56cf),
	.w4(32'hb9c83a70),
	.w5(32'h3bb936e4),
	.w6(32'h3d07af67),
	.w7(32'h3cb79b07),
	.w8(32'h3b4911bb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb864b68),
	.w1(32'h3b649bf2),
	.w2(32'h3c6463ad),
	.w3(32'h3b46f90e),
	.w4(32'h3b57dbe3),
	.w5(32'hbc1d0371),
	.w6(32'h3b1b18d9),
	.w7(32'h3c03e5d4),
	.w8(32'hbc16ba88),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fa2c8),
	.w1(32'hbb19d30e),
	.w2(32'hbb1e6050),
	.w3(32'hbc9581dc),
	.w4(32'hbc94ebf1),
	.w5(32'hbc812630),
	.w6(32'hbb3c8b92),
	.w7(32'hbbeea1f4),
	.w8(32'hbc51b2cb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e22fa),
	.w1(32'hbc1ed5b0),
	.w2(32'hbc5b7fcd),
	.w3(32'hbc3e918a),
	.w4(32'hbc6738fc),
	.w5(32'hbbadb0ab),
	.w6(32'hbaca580c),
	.w7(32'hbc59e7fa),
	.w8(32'hbaa6f893),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb423e98),
	.w1(32'h3b05d245),
	.w2(32'h3b23c929),
	.w3(32'hbb2c0dd1),
	.w4(32'hbb31661d),
	.w5(32'h3b7d1e66),
	.w6(32'h3b014eff),
	.w7(32'h3b9a3441),
	.w8(32'h3b5c336a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02e5e1),
	.w1(32'hb9aaf5a9),
	.w2(32'h3aa2bd21),
	.w3(32'hba3107c0),
	.w4(32'h3a800d8c),
	.w5(32'hbc591a0f),
	.w6(32'hba03bbdf),
	.w7(32'h3a4ae70d),
	.w8(32'hbb93e2f9),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc156844),
	.w1(32'hbc8aca37),
	.w2(32'hbc4f053b),
	.w3(32'hbbb51ab6),
	.w4(32'hbc340a2f),
	.w5(32'h3b32ec56),
	.w6(32'hbc41dcd7),
	.w7(32'hbc492475),
	.w8(32'hb9c67cc9),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad10786),
	.w1(32'h3a954c92),
	.w2(32'h3b583f34),
	.w3(32'h3a2f18ec),
	.w4(32'h3b87af5a),
	.w5(32'h3b4dc3ef),
	.w6(32'hbc25a2ad),
	.w7(32'hbb876401),
	.w8(32'h3a9546f5),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adccfb3),
	.w1(32'h3a2d9d83),
	.w2(32'h3b55c942),
	.w3(32'hbaf03f9b),
	.w4(32'h3a59dcdf),
	.w5(32'hb9ff0b4b),
	.w6(32'hbb842091),
	.w7(32'h3b55bba1),
	.w8(32'hbb71f605),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4620ee),
	.w1(32'h3b8bde76),
	.w2(32'hbac886fb),
	.w3(32'hbb5900e9),
	.w4(32'hbb0dc2db),
	.w5(32'hba888ecc),
	.w6(32'h3b4be2b3),
	.w7(32'h3b3f54e7),
	.w8(32'hbb51ec52),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeacbb0),
	.w1(32'h3b5474b5),
	.w2(32'hb8a244de),
	.w3(32'hbbb17d66),
	.w4(32'hbb429634),
	.w5(32'hbb008a0f),
	.w6(32'hba95a85d),
	.w7(32'hbb262aa8),
	.w8(32'hbb60372b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc47f6f),
	.w1(32'hbb84523b),
	.w2(32'hbbbaafa3),
	.w3(32'hbaf86ba6),
	.w4(32'hba9abce7),
	.w5(32'hbaa027fb),
	.w6(32'hbb90aa22),
	.w7(32'hbb807565),
	.w8(32'h3a101487),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b77c5),
	.w1(32'h3b911247),
	.w2(32'h3b3fecd8),
	.w3(32'hbaf57e80),
	.w4(32'hbb19b472),
	.w5(32'hbabb5365),
	.w6(32'h3b75bea9),
	.w7(32'h3b3d6589),
	.w8(32'h3bb64209),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c68ef),
	.w1(32'hb96166d9),
	.w2(32'h3a188f43),
	.w3(32'hb9f50d50),
	.w4(32'h3ae37b9d),
	.w5(32'hbaed4c2b),
	.w6(32'h3bb1cfbf),
	.w7(32'h3bb7b36f),
	.w8(32'hbba3a0cd),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee47dc),
	.w1(32'h39e34c7e),
	.w2(32'h3c347ba2),
	.w3(32'hbc3755dd),
	.w4(32'hbbd5badf),
	.w5(32'hba8a78a3),
	.w6(32'hbbed7811),
	.w7(32'hbbabe6f5),
	.w8(32'hbb46808e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe771a),
	.w1(32'hbba2ed19),
	.w2(32'h3a88dcf7),
	.w3(32'h3ac93cbc),
	.w4(32'h3b8ad0cf),
	.w5(32'h3afa89bb),
	.w6(32'hba268389),
	.w7(32'h3b2caf52),
	.w8(32'h38578c6d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d0b39),
	.w1(32'hbad82506),
	.w2(32'h397607ad),
	.w3(32'h3a476420),
	.w4(32'h3b8a7ca3),
	.w5(32'h39e405e4),
	.w6(32'hbaa63917),
	.w7(32'h3b5dc994),
	.w8(32'h3b613d85),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb122559),
	.w1(32'h3a939d5b),
	.w2(32'hba0d33f1),
	.w3(32'h3a6c56b7),
	.w4(32'hbafcdfbe),
	.w5(32'h3bb97e83),
	.w6(32'h3b59619f),
	.w7(32'h3b4535d3),
	.w8(32'h3afe0402),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adadac0),
	.w1(32'hba6f61d3),
	.w2(32'hbb25a343),
	.w3(32'hba2776f4),
	.w4(32'hb9fd2dce),
	.w5(32'hbb65bd62),
	.w6(32'hbb40bc15),
	.w7(32'hbb8564da),
	.w8(32'hbad0e887),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cafb3),
	.w1(32'h3bc3541c),
	.w2(32'h3ac11d6f),
	.w3(32'hbb734ff9),
	.w4(32'h3a266d03),
	.w5(32'hbbfd4d99),
	.w6(32'hbaed3b76),
	.w7(32'hbb1daac6),
	.w8(32'hbb84e1fa),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb36991),
	.w1(32'hbc21a39d),
	.w2(32'hbb82ff53),
	.w3(32'hbc75c95e),
	.w4(32'hbc51f692),
	.w5(32'h39b6da11),
	.w6(32'hbbc935e1),
	.w7(32'hbc64cc15),
	.w8(32'hbb3203b4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b281e19),
	.w1(32'h3b1c5ca3),
	.w2(32'h3baaf455),
	.w3(32'hbb2864d2),
	.w4(32'h3921841a),
	.w5(32'hbb3f609f),
	.w6(32'hbb6b8aff),
	.w7(32'h3b8512c9),
	.w8(32'hbb303dcc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7da7c1),
	.w1(32'h3a1ee9ba),
	.w2(32'hbad8b7fe),
	.w3(32'hbbbdf4ea),
	.w4(32'h3a3c28be),
	.w5(32'hbaa6194f),
	.w6(32'h3b0954af),
	.w7(32'hbaf55716),
	.w8(32'h3be55f8a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8be44c),
	.w1(32'h3a2502da),
	.w2(32'hbaab4e6d),
	.w3(32'hbb0a7c62),
	.w4(32'hbbaf82d0),
	.w5(32'hbbeb3c39),
	.w6(32'h3bc7a767),
	.w7(32'hbb95dd98),
	.w8(32'hbba75e3e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a527288),
	.w1(32'hba1deb9d),
	.w2(32'hbbca33df),
	.w3(32'hbbaeb2f4),
	.w4(32'hbb315a57),
	.w5(32'hbbd50f80),
	.w6(32'hbb279462),
	.w7(32'hba518607),
	.w8(32'hbc871e09),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed2feb),
	.w1(32'h3bd62a91),
	.w2(32'h3c32f46e),
	.w3(32'hbc35b5ac),
	.w4(32'hbbb7181e),
	.w5(32'h3935062f),
	.w6(32'hbc5ba625),
	.w7(32'hbc802429),
	.w8(32'h3a845bcb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1df560),
	.w1(32'h3b53471c),
	.w2(32'h3b1b09c0),
	.w3(32'h39b28d4b),
	.w4(32'h3a07769f),
	.w5(32'hbb0af8fe),
	.w6(32'hb9df6ae4),
	.w7(32'h3afc0d14),
	.w8(32'h3a9a1d52),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b098612),
	.w1(32'hbad46fad),
	.w2(32'hbbbd1936),
	.w3(32'hbb6a9a85),
	.w4(32'hbb86be41),
	.w5(32'hbb43c11a),
	.w6(32'hba9fc68b),
	.w7(32'h3b35012a),
	.w8(32'hbb474763),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c8912),
	.w1(32'h3a8bcd3d),
	.w2(32'hba2c5318),
	.w3(32'hbab3b760),
	.w4(32'hbb4b0e28),
	.w5(32'hbbfdd1bb),
	.w6(32'hbaa6fc2e),
	.w7(32'hbba28804),
	.w8(32'h3acf87bd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395058a1),
	.w1(32'hbb2a1ae5),
	.w2(32'hbc112db1),
	.w3(32'hbb46b153),
	.w4(32'hbbc4566e),
	.w5(32'hbb198938),
	.w6(32'h3a94e7d3),
	.w7(32'hbb487cb4),
	.w8(32'h3c05cfc4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6da711),
	.w1(32'h3b9da329),
	.w2(32'hbafa476e),
	.w3(32'hbbb1496c),
	.w4(32'hbbb73bf7),
	.w5(32'hbbb866de),
	.w6(32'h3b992934),
	.w7(32'h3b8c638e),
	.w8(32'h3b625499),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e6ea0),
	.w1(32'h3b557e3b),
	.w2(32'h3bde40d4),
	.w3(32'hbbac562c),
	.w4(32'hb9ac0850),
	.w5(32'h3b053895),
	.w6(32'h3beb233b),
	.w7(32'h3be27b14),
	.w8(32'h3a977b4b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afde20),
	.w1(32'hba5edb94),
	.w2(32'hba8b279d),
	.w3(32'h39f04cbf),
	.w4(32'hba922266),
	.w5(32'h3bcdc583),
	.w6(32'hbb216404),
	.w7(32'h39a45214),
	.w8(32'h3c09d214),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab59a8e),
	.w1(32'h3b1eada6),
	.w2(32'hb9aee31e),
	.w3(32'h3ac1dc60),
	.w4(32'h3c34c425),
	.w5(32'h3bc9a914),
	.w6(32'h3bb58208),
	.w7(32'h3b5d6b78),
	.w8(32'h3aa604ef),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0c9bd),
	.w1(32'hbb4d4655),
	.w2(32'hb9d72719),
	.w3(32'h3b77649a),
	.w4(32'h3ba28a11),
	.w5(32'h3a3ccbc5),
	.w6(32'hbb1052c7),
	.w7(32'h3b0ffef8),
	.w8(32'h3b4e43be),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf44124),
	.w1(32'hbb0871a3),
	.w2(32'hba298668),
	.w3(32'hbb951129),
	.w4(32'hbbadec86),
	.w5(32'h3af6f6fa),
	.w6(32'h3afe5229),
	.w7(32'hbb89ce30),
	.w8(32'h3a83ca69),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7a162),
	.w1(32'hbc091906),
	.w2(32'hbbf2408c),
	.w3(32'hbbf5ca13),
	.w4(32'hb9979490),
	.w5(32'h3c5a44cb),
	.w6(32'hbc468c01),
	.w7(32'hbc4b550e),
	.w8(32'h3d030fc6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e9c18),
	.w1(32'hbc5a756a),
	.w2(32'hbcbd671d),
	.w3(32'hbc3be04e),
	.w4(32'hbcbe6101),
	.w5(32'h3c382793),
	.w6(32'hbc0c8d64),
	.w7(32'hbcfa3873),
	.w8(32'h3c846fb7),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83b9b8),
	.w1(32'hbbbbaf79),
	.w2(32'hbcd26563),
	.w3(32'hbbc7c936),
	.w4(32'hbc419bf6),
	.w5(32'h3c340823),
	.w6(32'hbc1d1fc0),
	.w7(32'hbcd02565),
	.w8(32'hbb530609),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9417f2),
	.w1(32'hbbe2dc6c),
	.w2(32'h3ab6aef7),
	.w3(32'h3c6d51ee),
	.w4(32'h3c2b61f5),
	.w5(32'hbadab9ab),
	.w6(32'h3bb4f403),
	.w7(32'h3b95d7ff),
	.w8(32'hbb672214),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d338c),
	.w1(32'hbc278195),
	.w2(32'hbb1715a6),
	.w3(32'hbc00f531),
	.w4(32'hbb8552e5),
	.w5(32'h3d7823ab),
	.w6(32'hbc163f29),
	.w7(32'hbbcbb350),
	.w8(32'h3dda1f58),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8a2aba),
	.w1(32'hbc25e810),
	.w2(32'hbd99baac),
	.w3(32'hbc9f9e55),
	.w4(32'hbd72ba49),
	.w5(32'h3b93a918),
	.w6(32'hba8cd6dc),
	.w7(32'hbdc2a36c),
	.w8(32'hbb916986),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f0bea),
	.w1(32'h3b6ebbaa),
	.w2(32'h3bd83080),
	.w3(32'h3c4e5253),
	.w4(32'h3c038314),
	.w5(32'h3c83c2d1),
	.w6(32'hbbb2ff76),
	.w7(32'h3c5bdaa2),
	.w8(32'h3cc0fb69),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89eefb),
	.w1(32'h3bf95521),
	.w2(32'hbcc37732),
	.w3(32'hbb22c476),
	.w4(32'hbcef543f),
	.w5(32'h3c2e4ee6),
	.w6(32'h3be134d9),
	.w7(32'hbcfd0ee4),
	.w8(32'h3c2e4ff5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a4542),
	.w1(32'hbbc05abb),
	.w2(32'h3b4a9a4d),
	.w3(32'hbc2cb3c6),
	.w4(32'h3ba0000f),
	.w5(32'hbb029e3e),
	.w6(32'hbcce2433),
	.w7(32'hbc1f27b0),
	.w8(32'h39db303e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e3bd9),
	.w1(32'hb8e31b25),
	.w2(32'h3c24157c),
	.w3(32'h3b1e0cb1),
	.w4(32'h3c2d1bd0),
	.w5(32'h3c1ffc61),
	.w6(32'h3bc00253),
	.w7(32'h3c240f81),
	.w8(32'h3b38b2b2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7787),
	.w1(32'hbc490b65),
	.w2(32'hbbdc4f49),
	.w3(32'hbc16131a),
	.w4(32'h3b72467b),
	.w5(32'hbc4f34a0),
	.w6(32'hbc884bf2),
	.w7(32'hbc3843c7),
	.w8(32'hbcf8e6c6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8e9bd),
	.w1(32'hbb0ed644),
	.w2(32'h3ca0a044),
	.w3(32'h3c3e9817),
	.w4(32'h3d030ace),
	.w5(32'hb9c64205),
	.w6(32'h3a4cfbea),
	.w7(32'h3ce6a828),
	.w8(32'hbb02d635),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cc9cb),
	.w1(32'h3b928a2d),
	.w2(32'hbb97bf59),
	.w3(32'hbb7fbc67),
	.w4(32'hbbc4d517),
	.w5(32'h3b8518c0),
	.w6(32'h3a67dc6c),
	.w7(32'hbad92070),
	.w8(32'hbbb277b3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6ff93),
	.w1(32'hb99c7c34),
	.w2(32'hbb27ef17),
	.w3(32'h3bc911be),
	.w4(32'hbbfcdc63),
	.w5(32'hbd0782ba),
	.w6(32'h3be8996b),
	.w7(32'hbb8dbd4a),
	.w8(32'hbd38328d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd00df59),
	.w1(32'hbadc5089),
	.w2(32'h3cc944b3),
	.w3(32'h3a6ecc57),
	.w4(32'h3cb61ad4),
	.w5(32'h3a59dce3),
	.w6(32'h392e7b69),
	.w7(32'h3d277326),
	.w8(32'h3ba30413),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b957e45),
	.w1(32'h3a21609f),
	.w2(32'hbb0527d8),
	.w3(32'hb9f7d34d),
	.w4(32'hba9eede0),
	.w5(32'hbb4b8537),
	.w6(32'hbb4d25f6),
	.w7(32'hbacd70f5),
	.w8(32'h3c82c305),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ed6bb),
	.w1(32'hbbe140f2),
	.w2(32'hbd07e3c3),
	.w3(32'hbc982ebf),
	.w4(32'hbc6ee8ac),
	.w5(32'h3c3b1a63),
	.w6(32'hbbffe5e0),
	.w7(32'hbcf0a38b),
	.w8(32'hbadaf013),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41f1fd),
	.w1(32'hbbad794d),
	.w2(32'hbb2c009d),
	.w3(32'h3c1de62d),
	.w4(32'hbb85cba4),
	.w5(32'hbcca6e29),
	.w6(32'h3a93ec7c),
	.w7(32'hbbcb917a),
	.w8(32'hbcfbd1f2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdc3b9e),
	.w1(32'hba94f106),
	.w2(32'h3cb3ac6a),
	.w3(32'hbb1f3922),
	.w4(32'h3c683405),
	.w5(32'h3c692c9b),
	.w6(32'hbba28986),
	.w7(32'h3ca43ed3),
	.w8(32'h3c98ce50),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed0693),
	.w1(32'hbb70e903),
	.w2(32'hbc06ea16),
	.w3(32'h39dc4dd1),
	.w4(32'h3b8ed933),
	.w5(32'h3c51086f),
	.w6(32'hb81905d6),
	.w7(32'hbb6d6f9a),
	.w8(32'h3cae6e84),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3dc7d2),
	.w1(32'hbbb9b457),
	.w2(32'hbc90308a),
	.w3(32'hbbbbb694),
	.w4(32'hbc881808),
	.w5(32'h3d0aeec2),
	.w6(32'hbbbd3091),
	.w7(32'hbcc2fb9a),
	.w8(32'h3d69d08c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d240f6a),
	.w1(32'hbb3d7d59),
	.w2(32'hbd17f06b),
	.w3(32'hbc3578e9),
	.w4(32'hbd00a13a),
	.w5(32'h3c388df3),
	.w6(32'hbbad4855),
	.w7(32'hbd80b8b0),
	.w8(32'h3b20910d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea27a6),
	.w1(32'hbb7f0b7b),
	.w2(32'hbc1970a4),
	.w3(32'h3bcafcdf),
	.w4(32'h39a1acc9),
	.w5(32'hbbd87643),
	.w6(32'hba1617d7),
	.w7(32'hb9f3c321),
	.w8(32'hbb204bb5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb929e793),
	.w1(32'hbba148ad),
	.w2(32'h3be562cc),
	.w3(32'hbc08a58c),
	.w4(32'h3a22b716),
	.w5(32'hbb8340d6),
	.w6(32'hbc1de0b8),
	.w7(32'h3bae2761),
	.w8(32'hbc8f0067),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09b683),
	.w1(32'h3b8ce381),
	.w2(32'h3c84c155),
	.w3(32'h3be6f0a0),
	.w4(32'h3c4f772b),
	.w5(32'hbb6021a0),
	.w6(32'h3b1c9f01),
	.w7(32'h3cba4881),
	.w8(32'hbc8895ba),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48f5bd),
	.w1(32'hbad97c30),
	.w2(32'h3ba28152),
	.w3(32'h3bc4645a),
	.w4(32'h3aad17a6),
	.w5(32'hbb2e8c2d),
	.w6(32'h3ba1dbdb),
	.w7(32'h3c0ad130),
	.w8(32'hbc3e4218),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ed92f),
	.w1(32'h3bec4cd0),
	.w2(32'h3c98eec2),
	.w3(32'h3ac9f896),
	.w4(32'h3b93e340),
	.w5(32'h3c35eb96),
	.w6(32'h3baff0dd),
	.w7(32'h3c969efa),
	.w8(32'h3aa946c0),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e3f01),
	.w1(32'hbacb1c3b),
	.w2(32'hbbc701a1),
	.w3(32'h3c0205ec),
	.w4(32'h3bbc5275),
	.w5(32'hbb841837),
	.w6(32'h3c1ff64a),
	.w7(32'hbba39dc0),
	.w8(32'hbc75da78),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6eac4e),
	.w1(32'hbbfeaf00),
	.w2(32'h3c0f2a5b),
	.w3(32'h3c01e3fa),
	.w4(32'h3c49a293),
	.w5(32'h3b85bb4f),
	.w6(32'hbae1af5b),
	.w7(32'h3c7d7d81),
	.w8(32'h3bccae6c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc25834),
	.w1(32'hbc066873),
	.w2(32'hbc6cf82d),
	.w3(32'hbbc6c077),
	.w4(32'hbc3e88ea),
	.w5(32'hbc22af84),
	.w6(32'h3a398af2),
	.w7(32'hbc90610b),
	.w8(32'hbc451c8e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule