module layer_10_featuremap_427(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba110e),
	.w1(32'h3c20e8bc),
	.w2(32'h3b4269c7),
	.w3(32'hbc243f51),
	.w4(32'h3bf53fcb),
	.w5(32'h3b3dd8ca),
	.w6(32'h399bd56c),
	.w7(32'h3c1e535d),
	.w8(32'h3b63034e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc107e63),
	.w1(32'h3b3b955a),
	.w2(32'hbacf5118),
	.w3(32'hbbc1e405),
	.w4(32'hb9ced6a1),
	.w5(32'hbbab3599),
	.w6(32'hb8b08491),
	.w7(32'h3b5c05b8),
	.w8(32'hbc06b381),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad524),
	.w1(32'h392e20ed),
	.w2(32'h3abf9cb0),
	.w3(32'hb98f69d7),
	.w4(32'hb9d03053),
	.w5(32'hbc22dfe9),
	.w6(32'hb8e4a75d),
	.w7(32'h3ac7a014),
	.w8(32'hbb4d5f71),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c460b60),
	.w1(32'h3b280b49),
	.w2(32'h3c5bdfa7),
	.w3(32'h3bad6963),
	.w4(32'h3a8c992d),
	.w5(32'h3c2c9a2e),
	.w6(32'hbb8fab88),
	.w7(32'h3b990e5f),
	.w8(32'h3c7813c2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f2629),
	.w1(32'h3addbbfa),
	.w2(32'h3b02106d),
	.w3(32'h3c66d037),
	.w4(32'hbac54a50),
	.w5(32'hbb5d41aa),
	.w6(32'h3c402685),
	.w7(32'h3b842d21),
	.w8(32'h3b3ff10c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba1aa3),
	.w1(32'h36a9d3b0),
	.w2(32'hbbd1b923),
	.w3(32'h3b4f2c64),
	.w4(32'h3b3f1063),
	.w5(32'h3bf440f9),
	.w6(32'h3a8f3112),
	.w7(32'h3a12c251),
	.w8(32'h3a56f8b4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6435b),
	.w1(32'hbc5c079a),
	.w2(32'hbc65f26a),
	.w3(32'hbb123853),
	.w4(32'hbce620e0),
	.w5(32'hbd0fcfef),
	.w6(32'hb99d6f05),
	.w7(32'hbce188e8),
	.w8(32'hbce7f556),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b314a),
	.w1(32'hbc41daf2),
	.w2(32'hba69e4bd),
	.w3(32'hbd0a2a5e),
	.w4(32'hbbe26c20),
	.w5(32'h3c4e24fb),
	.w6(32'hbcef766b),
	.w7(32'hbafcb688),
	.w8(32'hbb14efb7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddaf18),
	.w1(32'hb9c58017),
	.w2(32'hbabe36fa),
	.w3(32'h3be663ea),
	.w4(32'hbb12473a),
	.w5(32'hbc6a57ca),
	.w6(32'h3ada8e78),
	.w7(32'hbc007cf6),
	.w8(32'hbbd6dd97),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc412e31),
	.w1(32'h3bea489a),
	.w2(32'hbb128ffc),
	.w3(32'hbc118196),
	.w4(32'h3bd406f8),
	.w5(32'hbab45252),
	.w6(32'hba2a3ce1),
	.w7(32'h3a914e06),
	.w8(32'hbbf2e921),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1128f),
	.w1(32'h3bbad856),
	.w2(32'h3bc2c2fa),
	.w3(32'h3987c566),
	.w4(32'hbbc0dcf0),
	.w5(32'hbc106719),
	.w6(32'hbbd44eb7),
	.w7(32'hbb90a581),
	.w8(32'hbbd15614),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25750b),
	.w1(32'hbb8a567f),
	.w2(32'h3bdccfe0),
	.w3(32'hba1f0cc8),
	.w4(32'hbbb724f5),
	.w5(32'h3c179000),
	.w6(32'hbbe85188),
	.w7(32'hbc0e2e20),
	.w8(32'h3bb72c28),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99ba72),
	.w1(32'hbc08d732),
	.w2(32'hbd0126e7),
	.w3(32'h3b76e075),
	.w4(32'hbc991831),
	.w5(32'hbd1d46bc),
	.w6(32'h3b84f07c),
	.w7(32'hbc62d11e),
	.w8(32'hbd062f87),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcde2303),
	.w1(32'hbc88e6df),
	.w2(32'hbc278446),
	.w3(32'hbd0a4af0),
	.w4(32'hbc8dfcab),
	.w5(32'hbc64de5c),
	.w6(32'hbcb1c9a8),
	.w7(32'hbc2209b2),
	.w8(32'hbc65379b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902e32d),
	.w1(32'h3ba53288),
	.w2(32'h3b240873),
	.w3(32'hbc49b7e0),
	.w4(32'h3bb9bc80),
	.w5(32'h3c15d271),
	.w6(32'hbc54872b),
	.w7(32'h3a9d6997),
	.w8(32'h3c08fc62),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3e8c0),
	.w1(32'hbc457932),
	.w2(32'hbc2dff61),
	.w3(32'hbbd6cfe4),
	.w4(32'hbc679a02),
	.w5(32'h3b85d27f),
	.w6(32'hbaf8de0b),
	.w7(32'hbbe93d34),
	.w8(32'hb9df0a02),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fef54),
	.w1(32'h3c041e9f),
	.w2(32'h3c62db47),
	.w3(32'hbb269d14),
	.w4(32'hbb9b307c),
	.w5(32'h3b43b704),
	.w6(32'hbaea93ec),
	.w7(32'hbc4617e3),
	.w8(32'hbae2369d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76bcb6),
	.w1(32'h3c0a3e5b),
	.w2(32'h3b2159a6),
	.w3(32'h3b115669),
	.w4(32'h3c3c633b),
	.w5(32'h3b7a080f),
	.w6(32'hbb805964),
	.w7(32'h3c6e32b8),
	.w8(32'h3c7afb6f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e34e8),
	.w1(32'hba8831a9),
	.w2(32'h3c2cffbf),
	.w3(32'hbc068786),
	.w4(32'h3b19612d),
	.w5(32'h3c836c1b),
	.w6(32'h394213dc),
	.w7(32'h3ba243ce),
	.w8(32'h3c633cb9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d7042),
	.w1(32'hbbe4f57f),
	.w2(32'hbb9386de),
	.w3(32'h3c39ba1b),
	.w4(32'hbc0363c6),
	.w5(32'hbc1c1484),
	.w6(32'h3c688320),
	.w7(32'hb94fa4a1),
	.w8(32'h3aaf0b23),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1e0e1),
	.w1(32'h3b0c8501),
	.w2(32'h3c249178),
	.w3(32'hbbd988eb),
	.w4(32'h3c2debec),
	.w5(32'h3cee7fe3),
	.w6(32'hbc1d1d7b),
	.w7(32'h3a93f5d3),
	.w8(32'h3bf4412c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d8ad9),
	.w1(32'hbb3f8702),
	.w2(32'hb9a35f85),
	.w3(32'h3bb79d6d),
	.w4(32'h3a6cde01),
	.w5(32'h3bff01f0),
	.w6(32'hbb75526a),
	.w7(32'h39fa46b8),
	.w8(32'h3ab57c48),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc228a1),
	.w1(32'hbc4a430e),
	.w2(32'hbc06d129),
	.w3(32'hbc451efd),
	.w4(32'h3b14c02a),
	.w5(32'h3b5a0ea5),
	.w6(32'hbc0a747b),
	.w7(32'hbc331588),
	.w8(32'h3ac46775),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe29895),
	.w1(32'hb9f2c5fa),
	.w2(32'hbb47defe),
	.w3(32'hb978c9ab),
	.w4(32'h3bc930e3),
	.w5(32'hba5f4cf3),
	.w6(32'h39ccc05c),
	.w7(32'hba37ac67),
	.w8(32'hb8979e02),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc122736),
	.w1(32'hbb8cffde),
	.w2(32'hbbb9c864),
	.w3(32'h3a025af1),
	.w4(32'hbc4acf83),
	.w5(32'hbc393da7),
	.w6(32'hbc134ddf),
	.w7(32'hbc1fc5c7),
	.w8(32'hbbda3415),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cc037),
	.w1(32'hbb1a1f06),
	.w2(32'h3b3b4d4d),
	.w3(32'hbb99e09a),
	.w4(32'h3bd56ec2),
	.w5(32'h3bff6671),
	.w6(32'hbc0f3b98),
	.w7(32'h3ac61f39),
	.w8(32'h3c2201d4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd06e0e),
	.w1(32'hbc1b78cf),
	.w2(32'hbb3bc127),
	.w3(32'h3ae07dc6),
	.w4(32'hb944ff49),
	.w5(32'h3c333ce9),
	.w6(32'hbbcea633),
	.w7(32'h3a403c3d),
	.w8(32'h3b50c4ae),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc50fee),
	.w1(32'h3be70a36),
	.w2(32'h3aa224d2),
	.w3(32'h3a468bbe),
	.w4(32'h3b9e9fd6),
	.w5(32'hbc258301),
	.w6(32'h3c159a7d),
	.w7(32'h3c5f4c8d),
	.w8(32'h3b8b9f88),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386d740b),
	.w1(32'h3b91e8ba),
	.w2(32'h3b4a0e4c),
	.w3(32'hbbc6302e),
	.w4(32'hbb23c003),
	.w5(32'hbab74732),
	.w6(32'hbb578b4b),
	.w7(32'hbbc64ee5),
	.w8(32'hbb29c75c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80544b),
	.w1(32'h3a929403),
	.w2(32'hbbb48891),
	.w3(32'hbbf79b9d),
	.w4(32'hbb9d4a53),
	.w5(32'hbc216ab1),
	.w6(32'h3b8475b9),
	.w7(32'h3abf141f),
	.w8(32'hbbce529d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b849827),
	.w1(32'hbbbfcdb7),
	.w2(32'hb99bc6ce),
	.w3(32'hba7b2a07),
	.w4(32'hbbfe8d34),
	.w5(32'hbaa1cc0c),
	.w6(32'h3b9662b9),
	.w7(32'hbc07d1e7),
	.w8(32'hbc0be890),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77207d),
	.w1(32'hbc2c9e20),
	.w2(32'hbc31ffcd),
	.w3(32'hbb522778),
	.w4(32'hbc18bc70),
	.w5(32'hbc857661),
	.w6(32'hbc02ea8d),
	.w7(32'h38c1659e),
	.w8(32'hbc13a2aa),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40247a),
	.w1(32'h3c2a3552),
	.w2(32'h3c5aeda2),
	.w3(32'hbac779cd),
	.w4(32'h3c0145f7),
	.w5(32'h3bba40e1),
	.w6(32'hba09eda5),
	.w7(32'h3b2466f2),
	.w8(32'h3c18ed9f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9fe22),
	.w1(32'h3b687948),
	.w2(32'h3b7cd9c0),
	.w3(32'h3b5e7672),
	.w4(32'hbb23eb6b),
	.w5(32'hbc528b06),
	.w6(32'h3ba0afa3),
	.w7(32'hbc143d6e),
	.w8(32'hbc34c57b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41b351),
	.w1(32'hbbd09353),
	.w2(32'hbbb54c04),
	.w3(32'hbc3bef63),
	.w4(32'hbb05cd4b),
	.w5(32'h3c28ed54),
	.w6(32'hbc17ffb2),
	.w7(32'hbc2223ab),
	.w8(32'h3a81201b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5e41e),
	.w1(32'hbbdea4a2),
	.w2(32'h3b9dc416),
	.w3(32'hbb1fc314),
	.w4(32'hbb4cf253),
	.w5(32'h3c89ca65),
	.w6(32'h3b3b3246),
	.w7(32'hbb667747),
	.w8(32'h3bf8372e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc271556),
	.w1(32'hbc11f54a),
	.w2(32'h3a6d8d3e),
	.w3(32'hbc42c48f),
	.w4(32'hbc2d63e5),
	.w5(32'hbc9318a1),
	.w6(32'hbbb10fed),
	.w7(32'hb9e4b46e),
	.w8(32'hbbf73f25),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25f74f),
	.w1(32'hbc39764b),
	.w2(32'hbc87d1aa),
	.w3(32'hbb577120),
	.w4(32'hbc49dfb8),
	.w5(32'hbcbd8a00),
	.w6(32'hb957896d),
	.w7(32'hbbe657e2),
	.w8(32'hbccc4f74),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0521b9),
	.w1(32'hbc419479),
	.w2(32'hbcdff4bd),
	.w3(32'hbbcf913b),
	.w4(32'hbc0f2bf4),
	.w5(32'hbceb6d17),
	.w6(32'hbb9e7719),
	.w7(32'hbb2b98ad),
	.w8(32'hbcc51f90),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc641626),
	.w1(32'h3b80b7a3),
	.w2(32'h3c0efb22),
	.w3(32'hbc89a3b1),
	.w4(32'h3a8b9d47),
	.w5(32'h3ba96dff),
	.w6(32'hbca4945e),
	.w7(32'h3ad6bcec),
	.w8(32'h3bfaa3f5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d0591),
	.w1(32'h3b7c1bda),
	.w2(32'h3b6911b8),
	.w3(32'h3b1f11fc),
	.w4(32'h3bcedb3a),
	.w5(32'h3c00478a),
	.w6(32'h3b82cb00),
	.w7(32'hbb206f41),
	.w8(32'hb991e71b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5abb1),
	.w1(32'h3b88647f),
	.w2(32'h3b7af1d8),
	.w3(32'hbba6c9e7),
	.w4(32'h3b49c615),
	.w5(32'h3ba27f33),
	.w6(32'hbb09306a),
	.w7(32'h3bf025ae),
	.w8(32'h3be66d3e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5a8e4),
	.w1(32'h3b273b95),
	.w2(32'h3bd3d7d6),
	.w3(32'h3aa5f0bb),
	.w4(32'hbae17605),
	.w5(32'h3b5dd257),
	.w6(32'h380f9e07),
	.w7(32'h3bb9828a),
	.w8(32'h3be78f01),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95fb4d),
	.w1(32'hbc17686a),
	.w2(32'hbc30f40d),
	.w3(32'hbbde4157),
	.w4(32'h3a9258c6),
	.w5(32'hbaf9778d),
	.w6(32'h3c2625d9),
	.w7(32'h3c3732fd),
	.w8(32'h3b6b0676),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3114dd),
	.w1(32'h3c5e4d61),
	.w2(32'h3bfac6bb),
	.w3(32'hbbbfa536),
	.w4(32'h3c6a74aa),
	.w5(32'h3ba0f6d6),
	.w6(32'hbb1294b0),
	.w7(32'h3c5759a5),
	.w8(32'h3c087c14),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c37cb),
	.w1(32'hbc27f3bf),
	.w2(32'hbc496ba4),
	.w3(32'h3bcebc65),
	.w4(32'hbc32aef5),
	.w5(32'hbbd700af),
	.w6(32'h3b927532),
	.w7(32'hbbd29d7d),
	.w8(32'hbc096fcf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb117bd3),
	.w1(32'hbb91a9e8),
	.w2(32'hbc5a25f4),
	.w3(32'hbbabb99d),
	.w4(32'hbc6281e8),
	.w5(32'hbcb21b56),
	.w6(32'hba2e97e6),
	.w7(32'hbc17dd3d),
	.w8(32'hbc2b7fc0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8797e4),
	.w1(32'h3b6acfcc),
	.w2(32'hbc262741),
	.w3(32'hbcc6e920),
	.w4(32'h3c5b9897),
	.w5(32'hbba1f55d),
	.w6(32'hbc9d66bc),
	.w7(32'h3c239490),
	.w8(32'hbbb3e0c8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66d7c9),
	.w1(32'hbb0e33e4),
	.w2(32'hbbcfe78c),
	.w3(32'hbc8ebeac),
	.w4(32'h3bbdf221),
	.w5(32'h3c258dae),
	.w6(32'hbc8a3591),
	.w7(32'hbbec114f),
	.w8(32'hba494ef6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd56d8a),
	.w1(32'hbb13dc8f),
	.w2(32'hbb86e989),
	.w3(32'h3bc990a8),
	.w4(32'h3bfedeb3),
	.w5(32'h3c64bc7f),
	.w6(32'hbb9183ba),
	.w7(32'h3affddab),
	.w8(32'h3b16f7c7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c0aa9),
	.w1(32'h3a37bfa6),
	.w2(32'h3ba0d9c1),
	.w3(32'h3ba185e2),
	.w4(32'h3b82b553),
	.w5(32'h3c3375a6),
	.w6(32'hbb1618fb),
	.w7(32'hbb802027),
	.w8(32'h3b4be460),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15fbdb),
	.w1(32'hbc39cc15),
	.w2(32'hbc6134fd),
	.w3(32'hbb612b17),
	.w4(32'hba125b5b),
	.w5(32'hbbfdd30b),
	.w6(32'hbb0609d6),
	.w7(32'hbab1db02),
	.w8(32'hbc369a8c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942adb),
	.w1(32'hbb2e783f),
	.w2(32'hbb0bed46),
	.w3(32'hba94ef51),
	.w4(32'hbb6dc3cf),
	.w5(32'h3b827c13),
	.w6(32'h3ab66720),
	.w7(32'hbba8e1ff),
	.w8(32'h3997a47b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc460c67),
	.w1(32'hbae0fa34),
	.w2(32'hbb28d34b),
	.w3(32'hbbe6830e),
	.w4(32'h3c35c90d),
	.w5(32'h3c9cd958),
	.w6(32'hbaacccc7),
	.w7(32'h3b0bf351),
	.w8(32'h3b039b0a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ebc66),
	.w1(32'hbad6f461),
	.w2(32'hbba115c2),
	.w3(32'h3ac3c512),
	.w4(32'h3b2f72ba),
	.w5(32'hbb8533b6),
	.w6(32'hb9d279d4),
	.w7(32'h3c16f59d),
	.w8(32'h3b50d374),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb920320),
	.w1(32'h3ae97d9f),
	.w2(32'h3a6a6430),
	.w3(32'hbb623a17),
	.w4(32'hbb8b076a),
	.w5(32'hbbe54968),
	.w6(32'hbb96810d),
	.w7(32'h3bb8d250),
	.w8(32'hba3991a1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96e36a),
	.w1(32'h3b113c8b),
	.w2(32'h3b228a7b),
	.w3(32'hbb981090),
	.w4(32'hbbb347c0),
	.w5(32'hbaa3b141),
	.w6(32'hba2268fc),
	.w7(32'hbb712535),
	.w8(32'hbb2544f2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcf876),
	.w1(32'h3c267481),
	.w2(32'hbb892e04),
	.w3(32'hbc37cbcb),
	.w4(32'h3c538ace),
	.w5(32'hb96a49ec),
	.w6(32'hbb703771),
	.w7(32'h3c1a2a96),
	.w8(32'h3b9e49e0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd110cd),
	.w1(32'h3b051e6f),
	.w2(32'h3b3bf297),
	.w3(32'hba5c84a9),
	.w4(32'hbb9d2e4d),
	.w5(32'hbb74cc6d),
	.w6(32'hbbbecff5),
	.w7(32'h3b37f343),
	.w8(32'h3aa0c8ed),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dae9d),
	.w1(32'hbc19438b),
	.w2(32'hba25c256),
	.w3(32'hbb21755d),
	.w4(32'hbb832e04),
	.w5(32'hb914e768),
	.w6(32'h3c0d3505),
	.w7(32'hbaa92584),
	.w8(32'h3b46953c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2583fb),
	.w1(32'hb9a93b39),
	.w2(32'h3b6e4e82),
	.w3(32'hbb439844),
	.w4(32'h3bc4d3a7),
	.w5(32'h3c179722),
	.w6(32'hbbde6a1b),
	.w7(32'h3b01331e),
	.w8(32'h3b89a4f9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc136066),
	.w1(32'h3ab34007),
	.w2(32'h3aecf4cf),
	.w3(32'hbc1f1ff4),
	.w4(32'h3b650e12),
	.w5(32'hbc03108e),
	.w6(32'hbbae7440),
	.w7(32'h3bb598e2),
	.w8(32'h3b007097),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f71f7),
	.w1(32'h3c521851),
	.w2(32'h3c7d9ded),
	.w3(32'h3b0f4efe),
	.w4(32'h3c05bd93),
	.w5(32'h3c2eea66),
	.w6(32'hbb49fb8b),
	.w7(32'h3c510971),
	.w8(32'h3c8af120),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92bfd0),
	.w1(32'hbc0b160e),
	.w2(32'h38a9c2e2),
	.w3(32'h3c51bb40),
	.w4(32'hbb9e69b6),
	.w5(32'h3c15e7e9),
	.w6(32'h3c9743c6),
	.w7(32'hbbbf66a7),
	.w8(32'h3b9424e4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fed59),
	.w1(32'hbbb7f493),
	.w2(32'hbb6eb8f6),
	.w3(32'h3c175fde),
	.w4(32'h3a774a83),
	.w5(32'h3c020ad4),
	.w6(32'h3bf51363),
	.w7(32'hbb3fbba0),
	.w8(32'hb994faa6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc431245),
	.w1(32'hbbfcaeb2),
	.w2(32'hbb74d5a7),
	.w3(32'hbb04fbe1),
	.w4(32'hbc226481),
	.w5(32'hbbd09182),
	.w6(32'hbbc5005d),
	.w7(32'hbb9f4a09),
	.w8(32'hbb8f561d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20d328),
	.w1(32'h3be7ac54),
	.w2(32'hbad36e4f),
	.w3(32'hbc8e1b9e),
	.w4(32'h3996ac53),
	.w5(32'h398d7540),
	.w6(32'hbb9adbcd),
	.w7(32'h3b81c57d),
	.w8(32'h3b07152f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc779cf),
	.w1(32'hbaad98a4),
	.w2(32'hbbab8cdf),
	.w3(32'h3ad39dab),
	.w4(32'hbbcb4df8),
	.w5(32'hbc36acf4),
	.w6(32'hbc2b0237),
	.w7(32'hbc37265f),
	.w8(32'hb94f83d0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba261a9),
	.w1(32'hbc2b416e),
	.w2(32'hbad99db5),
	.w3(32'hbbac016a),
	.w4(32'hb950d734),
	.w5(32'hbbc9a014),
	.w6(32'hb94c04aa),
	.w7(32'h3a2d9b46),
	.w8(32'hbb08ab4a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8da0b),
	.w1(32'hbb57041f),
	.w2(32'hbc246cd0),
	.w3(32'h3ba36a1f),
	.w4(32'hb9a56a97),
	.w5(32'hbbfee3f8),
	.w6(32'h3af4841f),
	.w7(32'hb98176e9),
	.w8(32'hbb80390f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafab9b9),
	.w1(32'hbba6ffbc),
	.w2(32'hbb04a2f2),
	.w3(32'hbb9da20f),
	.w4(32'hbc5c6bc0),
	.w5(32'hbc5e45dc),
	.w6(32'hbbc1843e),
	.w7(32'hbc6a18e1),
	.w8(32'hbb17eb0d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb14411),
	.w1(32'h3c96db52),
	.w2(32'h3c6e2684),
	.w3(32'hbbe00ed8),
	.w4(32'h3cadcf30),
	.w5(32'h3c79ca38),
	.w6(32'hbb786213),
	.w7(32'h3ca6e42e),
	.w8(32'h3b03a6ff),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf869e),
	.w1(32'hb98fb486),
	.w2(32'hbaa6ef65),
	.w3(32'h3c4a03a7),
	.w4(32'hbab3eb83),
	.w5(32'h3a205484),
	.w6(32'h3b4e9368),
	.w7(32'hbbbc53ef),
	.w8(32'hbc1fbd5c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb3f4),
	.w1(32'h3a80caeb),
	.w2(32'h3c137ea1),
	.w3(32'h3ac40c67),
	.w4(32'hba838694),
	.w5(32'h3aad4de8),
	.w6(32'hb9fac000),
	.w7(32'h3b0b80f4),
	.w8(32'hba69341d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c024dfc),
	.w1(32'hbbf6dc7c),
	.w2(32'hba6ec403),
	.w3(32'hb92038e4),
	.w4(32'h3c291e7e),
	.w5(32'h3c9a3b77),
	.w6(32'hbbb5c87b),
	.w7(32'h3a5093e5),
	.w8(32'h3b7e0c7e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84a184),
	.w1(32'hbbe5c7f5),
	.w2(32'hbbfe32d6),
	.w3(32'h3c0d399c),
	.w4(32'hba7a8d82),
	.w5(32'h3c9553db),
	.w6(32'h3c12d811),
	.w7(32'h3b490615),
	.w8(32'h3bbb0077),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc632d4e),
	.w1(32'hbb103261),
	.w2(32'h3bb4f899),
	.w3(32'hbc00c56d),
	.w4(32'h3a55687c),
	.w5(32'h3b77b544),
	.w6(32'hbb5c30ac),
	.w7(32'h3bc91faf),
	.w8(32'hbae2be1c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8755ed),
	.w1(32'hbc86f3a1),
	.w2(32'hbcb6d0b4),
	.w3(32'h3b130e72),
	.w4(32'h3ab1de82),
	.w5(32'h3bd294cf),
	.w6(32'hbb1a473c),
	.w7(32'hbc23b9b2),
	.w8(32'hbcb5221b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e77e5),
	.w1(32'h3ba68863),
	.w2(32'hba81cd31),
	.w3(32'hbc1395cc),
	.w4(32'h3af7e5e9),
	.w5(32'h3bf188cd),
	.w6(32'hba286697),
	.w7(32'h3c23203c),
	.w8(32'h3b000341),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58e24d),
	.w1(32'hbbedebc2),
	.w2(32'hbbea4869),
	.w3(32'hbb59c7c5),
	.w4(32'hbc22878a),
	.w5(32'hbc62b40b),
	.w6(32'h39eedb31),
	.w7(32'h37fccc35),
	.w8(32'hbb6fe72d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc356d7f),
	.w1(32'hbc24f389),
	.w2(32'hbc457a6a),
	.w3(32'hbc074349),
	.w4(32'hbc537c7f),
	.w5(32'hbbc45c1f),
	.w6(32'hbbd3edcd),
	.w7(32'hbbd7b614),
	.w8(32'hbc008775),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06ad4b),
	.w1(32'hba2f27ee),
	.w2(32'hbb0f875a),
	.w3(32'hbb882b95),
	.w4(32'hba3b2d21),
	.w5(32'hba51646b),
	.w6(32'hb9896116),
	.w7(32'h3bbf4000),
	.w8(32'h3b4f2e00),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18cefa),
	.w1(32'h3acaa90b),
	.w2(32'hba62082e),
	.w3(32'h3b250328),
	.w4(32'h3c1938c1),
	.w5(32'h3ba9693a),
	.w6(32'h3b7e31a3),
	.w7(32'h388cdce2),
	.w8(32'h3afbfe2d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba82bf0),
	.w1(32'hbb917ed6),
	.w2(32'h3c18712e),
	.w3(32'h3b9e335f),
	.w4(32'h3ae7584f),
	.w5(32'hbc091b55),
	.w6(32'h3b73313f),
	.w7(32'h3a5c2b0c),
	.w8(32'hbbbfd768),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00170f),
	.w1(32'h3c3c8074),
	.w2(32'h3c91e8f6),
	.w3(32'hba890101),
	.w4(32'h3bca7e5c),
	.w5(32'h3c9bec7a),
	.w6(32'hb75e64c7),
	.w7(32'hbbc21ed4),
	.w8(32'h3adcc051),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3683dc),
	.w1(32'h3a2eff6c),
	.w2(32'hba720214),
	.w3(32'h3c7ec939),
	.w4(32'h3a0d907d),
	.w5(32'hbb586df9),
	.w6(32'h3c28ac03),
	.w7(32'hbb8543d9),
	.w8(32'hbc1d5ad1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d6f5b),
	.w1(32'h3c00de24),
	.w2(32'h3b16c298),
	.w3(32'hbb1e8c6e),
	.w4(32'hba62ec30),
	.w5(32'hbcca0a3e),
	.w6(32'hbb88bf5b),
	.w7(32'h3c77f4f5),
	.w8(32'h3c609252),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04614c),
	.w1(32'h3c50ccba),
	.w2(32'h3c66833d),
	.w3(32'hbc0df2ab),
	.w4(32'hbbc38a07),
	.w5(32'hbcca48f6),
	.w6(32'hb9fe8c84),
	.w7(32'h3c9442d0),
	.w8(32'h3cc92a99),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1218fe),
	.w1(32'hbbb0849d),
	.w2(32'h3b62ae46),
	.w3(32'hbbb6be5f),
	.w4(32'h3bbf05b0),
	.w5(32'hbbe85125),
	.w6(32'h3c4a61dc),
	.w7(32'hbae7ab85),
	.w8(32'hbc3b99a5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc8cbc),
	.w1(32'h3bea4570),
	.w2(32'h3b19814c),
	.w3(32'hbb05a2aa),
	.w4(32'h3c0c8131),
	.w5(32'h3b9cc9bc),
	.w6(32'hba333d72),
	.w7(32'h3c171423),
	.w8(32'h3b186a50),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddb97d),
	.w1(32'h3afc9ad8),
	.w2(32'h3a7ecfe4),
	.w3(32'h3b9a1d99),
	.w4(32'h3a82bcfe),
	.w5(32'hbc13c63a),
	.w6(32'h3ae18039),
	.w7(32'hbb23501b),
	.w8(32'hbb00f25c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89cb12),
	.w1(32'h3bc00e8e),
	.w2(32'h3c2f626c),
	.w3(32'hbac85285),
	.w4(32'hbc151e8d),
	.w5(32'hbba7fc78),
	.w6(32'h3c1d39c0),
	.w7(32'h3b999d38),
	.w8(32'h3c1e5dcf),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fdf88),
	.w1(32'h3b91792b),
	.w2(32'hbbb37df5),
	.w3(32'h3a77d6ff),
	.w4(32'h3bc86fb7),
	.w5(32'h3bfaa463),
	.w6(32'hbaa80fea),
	.w7(32'h3b4c23c6),
	.w8(32'hbbd59c77),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb915d64),
	.w1(32'hbc332063),
	.w2(32'hbc1e89f9),
	.w3(32'h3bf2230b),
	.w4(32'hbb0013a9),
	.w5(32'h39a4b581),
	.w6(32'h3b482c73),
	.w7(32'hba78cf69),
	.w8(32'h3a943634),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc181943),
	.w1(32'h3be2c4dd),
	.w2(32'h3bc7fa16),
	.w3(32'hbc825756),
	.w4(32'hbb05440b),
	.w5(32'hbb784127),
	.w6(32'hbbfdfd3c),
	.w7(32'hba87217b),
	.w8(32'hbb451e12),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e95ad),
	.w1(32'hbb584234),
	.w2(32'hbc27d6ee),
	.w3(32'hbb899296),
	.w4(32'hbbecdb87),
	.w5(32'hbc9cda59),
	.w6(32'hbba6abc1),
	.w7(32'hbc416540),
	.w8(32'hbc971c93),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7262a),
	.w1(32'h3bca7ad3),
	.w2(32'h3bc78a57),
	.w3(32'hbc3fc039),
	.w4(32'hbbfdd559),
	.w5(32'h3a89509c),
	.w6(32'hbc210a8d),
	.w7(32'h3bafc1d0),
	.w8(32'h3ca15a97),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc518be),
	.w1(32'h3aef94bd),
	.w2(32'hbb5633ae),
	.w3(32'h3b07b1e1),
	.w4(32'hb900660e),
	.w5(32'hbab10a5d),
	.w6(32'h3c4d14cc),
	.w7(32'h3af8bba2),
	.w8(32'hbb314157),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3c734),
	.w1(32'h3baac09e),
	.w2(32'hba59847e),
	.w3(32'hbb3af4e7),
	.w4(32'h3bd1b126),
	.w5(32'h3abb7a48),
	.w6(32'h3c0bd8e1),
	.w7(32'h3c1e5b99),
	.w8(32'h3c455a99),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c421f),
	.w1(32'hbbd165a9),
	.w2(32'h3bd6ad6a),
	.w3(32'hbc0920cc),
	.w4(32'h3bd63959),
	.w5(32'h3cb4fb32),
	.w6(32'hbb744f95),
	.w7(32'hbbc762a8),
	.w8(32'h3c2ea9f1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec531f),
	.w1(32'h3b941275),
	.w2(32'h3c125d64),
	.w3(32'h3b82bb57),
	.w4(32'hbc16a9cd),
	.w5(32'hbbc99e4c),
	.w6(32'h396bf6bf),
	.w7(32'hb9d08813),
	.w8(32'h3c03f9f3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1f2a0),
	.w1(32'h3cb9e4c0),
	.w2(32'h3a32a1bf),
	.w3(32'hbbfda6d6),
	.w4(32'h3c87e4bf),
	.w5(32'h3b64db33),
	.w6(32'h392ed313),
	.w7(32'h3c3d3093),
	.w8(32'h3c0bbd5e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf00ab4),
	.w1(32'hbc7a7493),
	.w2(32'h3b3a7dcd),
	.w3(32'h3ac270c8),
	.w4(32'hbb777a49),
	.w5(32'h3c23d7a2),
	.w6(32'h3c82d8eb),
	.w7(32'hbaaefe34),
	.w8(32'hba4e1248),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e5c3),
	.w1(32'h39614cfa),
	.w2(32'h3b26d00b),
	.w3(32'hbb703f33),
	.w4(32'hbc017498),
	.w5(32'h3bbdaf10),
	.w6(32'hbc3a5e29),
	.w7(32'hbc7713ba),
	.w8(32'hbc4b3ae3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab088d),
	.w1(32'hbc58151c),
	.w2(32'hbb8bf6a1),
	.w3(32'hbc25e436),
	.w4(32'h3be468cb),
	.w5(32'h3c0b35a8),
	.w6(32'hbb3669cc),
	.w7(32'h3bbfd17c),
	.w8(32'h3bbc1749),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb927edc),
	.w1(32'hbbd764df),
	.w2(32'hbbd95b04),
	.w3(32'h3b826b60),
	.w4(32'h3a908979),
	.w5(32'hba672098),
	.w6(32'hba423238),
	.w7(32'h3b6c0c3c),
	.w8(32'hb9aad1e4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7ca90),
	.w1(32'hbb0c634f),
	.w2(32'hbba6ecc7),
	.w3(32'h3b522f28),
	.w4(32'hbb4b86c4),
	.w5(32'hbb8b3e36),
	.w6(32'h3be40ad1),
	.w7(32'hbc6e71f7),
	.w8(32'hbc167f34),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc196fc7),
	.w1(32'hba3ea5bc),
	.w2(32'h3b376e4a),
	.w3(32'hbb899744),
	.w4(32'h389c3360),
	.w5(32'h3c270fb2),
	.w6(32'hbc01c4c8),
	.w7(32'hbc0c229c),
	.w8(32'h3b559b73),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e163b),
	.w1(32'h3b7ffafa),
	.w2(32'hbba07e93),
	.w3(32'h3c068793),
	.w4(32'h3cae68ee),
	.w5(32'h3c32a1cc),
	.w6(32'h3c067153),
	.w7(32'h3c9cf890),
	.w8(32'h3cc3d357),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b993593),
	.w1(32'h3b9197f1),
	.w2(32'hbb89e720),
	.w3(32'h3c25b9cb),
	.w4(32'h3c2993c2),
	.w5(32'h39f021e1),
	.w6(32'h3c539b4a),
	.w7(32'hbc2359cd),
	.w8(32'hbb995748),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf11e3f),
	.w1(32'h3c3baf68),
	.w2(32'hb9bd735e),
	.w3(32'h3bc57156),
	.w4(32'hb96067b3),
	.w5(32'h3b8ca4f7),
	.w6(32'h3b83ee3d),
	.w7(32'h3bcd2112),
	.w8(32'hbb8b96c7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab60c6),
	.w1(32'hbb248c28),
	.w2(32'hbbbd5c22),
	.w3(32'h3b53007d),
	.w4(32'h3a04650a),
	.w5(32'hbb8f3593),
	.w6(32'hbc1b0309),
	.w7(32'h3bfe6d60),
	.w8(32'h3be0bef2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb128db2),
	.w1(32'h3b54b1ae),
	.w2(32'h3c932220),
	.w3(32'hb9e69d10),
	.w4(32'h3bbf11ac),
	.w5(32'h3c8bd14a),
	.w6(32'h3b3c093f),
	.w7(32'hbb9dff79),
	.w8(32'hbb694762),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f8e645),
	.w1(32'h3b1f079b),
	.w2(32'h3c0ac088),
	.w3(32'h3b94cc95),
	.w4(32'h3c1c98f0),
	.w5(32'h3c5acae2),
	.w6(32'h3a5d7354),
	.w7(32'h3b4527de),
	.w8(32'h3af8fdae),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84492e),
	.w1(32'hbadc1f13),
	.w2(32'hbadf2da4),
	.w3(32'h3aab669b),
	.w4(32'h3b17bf91),
	.w5(32'hbaf0c0ad),
	.w6(32'hbbd054ee),
	.w7(32'h3be2663f),
	.w8(32'hbb827495),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1d441),
	.w1(32'h395aaaf9),
	.w2(32'hbbae36c8),
	.w3(32'hbab1a7bc),
	.w4(32'hbbc396bd),
	.w5(32'hbb4d5619),
	.w6(32'h3a571f2f),
	.w7(32'hbbe1cca6),
	.w8(32'hbbd9c872),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023fd1),
	.w1(32'h3bec5940),
	.w2(32'h3c4e5169),
	.w3(32'hbb1abea8),
	.w4(32'h39f9b84e),
	.w5(32'hbb36578e),
	.w6(32'hba65520f),
	.w7(32'hbb382c50),
	.w8(32'hbb8da1a2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a7094),
	.w1(32'hbbb3eeab),
	.w2(32'hbc8a4fe0),
	.w3(32'h3bd98142),
	.w4(32'h3bd30b98),
	.w5(32'h3b9b487c),
	.w6(32'h3b405b00),
	.w7(32'hbb907dc7),
	.w8(32'hbbe812d0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe34ec),
	.w1(32'h3ae3265a),
	.w2(32'h3c1cd598),
	.w3(32'h3b4f0ff8),
	.w4(32'hbc064c07),
	.w5(32'hbc96e0a4),
	.w6(32'h3c029cb8),
	.w7(32'h3c180f53),
	.w8(32'h3b8f49ec),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a169878),
	.w1(32'hbc2eecc5),
	.w2(32'hbc6167d8),
	.w3(32'hbbcd28d0),
	.w4(32'hbbe6737f),
	.w5(32'hbbcb94aa),
	.w6(32'h3b4fca0d),
	.w7(32'hbc646bd7),
	.w8(32'hbc8f87bf),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c9292),
	.w1(32'h3c010bc5),
	.w2(32'h3bb69809),
	.w3(32'hbbe5bce0),
	.w4(32'h3af526b3),
	.w5(32'hbc311ba9),
	.w6(32'hbc6288b4),
	.w7(32'hbb68356f),
	.w8(32'hbc3c553d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911fd1c),
	.w1(32'hbc2d24eb),
	.w2(32'hbbcff12b),
	.w3(32'hbacfa679),
	.w4(32'hb9e74229),
	.w5(32'h3b8d3e40),
	.w6(32'hbb2c2551),
	.w7(32'hbb03024e),
	.w8(32'h3c0bce9f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c9ce4),
	.w1(32'h3c07abbd),
	.w2(32'h3c02a052),
	.w3(32'h3b9f7b3d),
	.w4(32'hbb12fbcd),
	.w5(32'hbc7cd03b),
	.w6(32'h3bf9f633),
	.w7(32'h3ae6a4aa),
	.w8(32'h3b64fc2c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96ce9b),
	.w1(32'h3c42cc7b),
	.w2(32'h3bf49eaa),
	.w3(32'h3904fecf),
	.w4(32'h3c3a48d0),
	.w5(32'h3b56b74f),
	.w6(32'h3b79e17c),
	.w7(32'h3bb4088f),
	.w8(32'h3bd817ef),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89d4b2),
	.w1(32'h3cea5a71),
	.w2(32'h3c7b4ebe),
	.w3(32'h3b5a2d21),
	.w4(32'h3cc4f910),
	.w5(32'h3c796fb2),
	.w6(32'h3c1a524b),
	.w7(32'h3cca1014),
	.w8(32'h3c803772),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca9d746),
	.w1(32'h3be64e41),
	.w2(32'h3c0e0a86),
	.w3(32'h3caa0872),
	.w4(32'h3c2093d0),
	.w5(32'h3ab6b04a),
	.w6(32'h3ce45bc6),
	.w7(32'h3b937466),
	.w8(32'hba1551c7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7f006),
	.w1(32'hbb3abac3),
	.w2(32'hbbe697be),
	.w3(32'h3c48f283),
	.w4(32'hb7c0b43a),
	.w5(32'hbbb0b28e),
	.w6(32'hbaa01feb),
	.w7(32'h3bf03c9d),
	.w8(32'h3c42618f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc854682),
	.w1(32'hbc5dd7bc),
	.w2(32'hbb88089c),
	.w3(32'hbacb72b0),
	.w4(32'hba7a300f),
	.w5(32'hba9470d4),
	.w6(32'h3b6c0c96),
	.w7(32'hbb9043ea),
	.w8(32'hbc2436d3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc237836),
	.w1(32'hbb92948b),
	.w2(32'hbb47921a),
	.w3(32'hbc3bd717),
	.w4(32'h3b9131d6),
	.w5(32'h3a12238c),
	.w6(32'hbc507488),
	.w7(32'h3bfd5e54),
	.w8(32'h3b2cf3de),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb181271),
	.w1(32'h3b5d8ba8),
	.w2(32'h3bca10fb),
	.w3(32'hba4e9c11),
	.w4(32'h388d0108),
	.w5(32'hba4e2100),
	.w6(32'h3b2356d9),
	.w7(32'h3be88d44),
	.w8(32'hbb3790a9),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1470f),
	.w1(32'h3b84313b),
	.w2(32'h3a606539),
	.w3(32'h3b0ccd42),
	.w4(32'h3c225356),
	.w5(32'h3bea1315),
	.w6(32'hbb88dc69),
	.w7(32'h3a6405cb),
	.w8(32'h3be2c050),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d26f9),
	.w1(32'h3c08238e),
	.w2(32'hbab90fe5),
	.w3(32'hbbffd223),
	.w4(32'h3c5498ae),
	.w5(32'h3c8969c1),
	.w6(32'hbaa6a44f),
	.w7(32'h3cd2bc83),
	.w8(32'h3c81052c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8cb29),
	.w1(32'h3c089474),
	.w2(32'hbbbec360),
	.w3(32'h3bd31373),
	.w4(32'h3c5db258),
	.w5(32'h3c02f341),
	.w6(32'h3c433d6b),
	.w7(32'h3c0adcae),
	.w8(32'h3c8d472b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c8ced),
	.w1(32'hbb940cfa),
	.w2(32'hbaff6fd3),
	.w3(32'hbb50c489),
	.w4(32'hbacbdf57),
	.w5(32'hbbe6e2f1),
	.w6(32'h3c3ba6fc),
	.w7(32'hb9946d9c),
	.w8(32'hbbd8878f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21eba7),
	.w1(32'hbc62e8f7),
	.w2(32'hbc69ad4f),
	.w3(32'hbc49311f),
	.w4(32'hbb084711),
	.w5(32'h3c4b1960),
	.w6(32'h3b792157),
	.w7(32'hbb9cf586),
	.w8(32'hbba791d4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aaa97),
	.w1(32'hbb2c7538),
	.w2(32'hbbc45c10),
	.w3(32'hbc0d6ee8),
	.w4(32'hbbe0e13a),
	.w5(32'hbc56d4a0),
	.w6(32'hbbc46b2d),
	.w7(32'h3abf7085),
	.w8(32'h3bb449f1),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada38c6),
	.w1(32'hbc32bc64),
	.w2(32'hbc30748b),
	.w3(32'hbb8334f2),
	.w4(32'hbbe71006),
	.w5(32'h3aaf84cc),
	.w6(32'h3c00a6a2),
	.w7(32'hbb61f707),
	.w8(32'hbb07e195),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc161318),
	.w1(32'h3b59b628),
	.w2(32'hbb16bf84),
	.w3(32'hbc018ec2),
	.w4(32'h3c02424c),
	.w5(32'h3b21ec5c),
	.w6(32'hbb997f01),
	.w7(32'h3c771eba),
	.w8(32'h3caea690),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee8b91),
	.w1(32'h3987a72a),
	.w2(32'h3a923f06),
	.w3(32'hbaa44602),
	.w4(32'h3c608586),
	.w5(32'h3c6b7027),
	.w6(32'h3c351b10),
	.w7(32'hbadb6c3a),
	.w8(32'h3b9d90e8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed41ad),
	.w1(32'h3bbdc987),
	.w2(32'hbacf6558),
	.w3(32'h39d784e5),
	.w4(32'h3b1f0f41),
	.w5(32'hbb1cb969),
	.w6(32'hbb4d7607),
	.w7(32'h3b6f235c),
	.w8(32'hbb79a68f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbc625),
	.w1(32'hbc2077a5),
	.w2(32'hbc8d90fe),
	.w3(32'h3b158f48),
	.w4(32'hbb5675cf),
	.w5(32'hbc25eaa0),
	.w6(32'hba7c2e21),
	.w7(32'hbae5986f),
	.w8(32'hbc90606e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f4436),
	.w1(32'hb9e88f1d),
	.w2(32'hbb8af738),
	.w3(32'hbbc724fc),
	.w4(32'hba544933),
	.w5(32'h3a198158),
	.w6(32'hbc5cdde4),
	.w7(32'hbc23241d),
	.w8(32'hbb44253e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03b5b0),
	.w1(32'h3c35a415),
	.w2(32'h3c458975),
	.w3(32'h3ac97c31),
	.w4(32'h3c868397),
	.w5(32'h3c750aeb),
	.w6(32'h3bfdc461),
	.w7(32'h3c945413),
	.w8(32'h3c9a6517),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fb496),
	.w1(32'h3b932b97),
	.w2(32'h3ae8cdf1),
	.w3(32'h3c20d407),
	.w4(32'h394f8576),
	.w5(32'h3c065bfb),
	.w6(32'h3be9cbea),
	.w7(32'hbb3c3b38),
	.w8(32'hba7ae3f0),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05cf83),
	.w1(32'h3c188f22),
	.w2(32'h3c2e7b23),
	.w3(32'h3b8154ff),
	.w4(32'h3c143a27),
	.w5(32'h3bb15405),
	.w6(32'hba822ca5),
	.w7(32'hbb8c7933),
	.w8(32'hbc12efa8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa65a06),
	.w1(32'h3b8e8e77),
	.w2(32'hba04f9ad),
	.w3(32'h3bd0b1ab),
	.w4(32'hbbc7f05d),
	.w5(32'hbc0cf6a0),
	.w6(32'hbc0d5d7f),
	.w7(32'h3bd5c808),
	.w8(32'h3a344ec1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64b378),
	.w1(32'h3b95e6e5),
	.w2(32'h3c0adf9a),
	.w3(32'h3a81ce34),
	.w4(32'h3bda085a),
	.w5(32'h3c071df3),
	.w6(32'h3b7bd207),
	.w7(32'hbab24069),
	.w8(32'h3a509814),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae295d),
	.w1(32'hbbb97cdf),
	.w2(32'hbb84b3ad),
	.w3(32'h3bd776d9),
	.w4(32'hbc03f2a7),
	.w5(32'h3bae4171),
	.w6(32'h3bf19d01),
	.w7(32'h3b014f8f),
	.w8(32'hbb9c5560),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922f0d),
	.w1(32'hba881a13),
	.w2(32'h3b3780b5),
	.w3(32'h3b08c266),
	.w4(32'hba395a36),
	.w5(32'hbb89cfbb),
	.w6(32'h3b689d21),
	.w7(32'hbbc07c55),
	.w8(32'hbc038856),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffaf0c),
	.w1(32'hbbb59f46),
	.w2(32'hbbf10759),
	.w3(32'hbb244fee),
	.w4(32'hbbe9f881),
	.w5(32'hbbd7f9c6),
	.w6(32'hbb20f9e0),
	.w7(32'h3b2724ac),
	.w8(32'hbba47cf6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04ad49),
	.w1(32'hbb5f5919),
	.w2(32'hbc501a88),
	.w3(32'hbb83b293),
	.w4(32'hbab8cc4d),
	.w5(32'hbb151d8e),
	.w6(32'hbc0e8fbc),
	.w7(32'h3b3e23c5),
	.w8(32'hbb3724bf),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbba4c),
	.w1(32'hbbd023af),
	.w2(32'hbbc95dce),
	.w3(32'hbc3f75f5),
	.w4(32'h3b689b63),
	.w5(32'h3be10a9d),
	.w6(32'hbb526aab),
	.w7(32'hbb5020d9),
	.w8(32'hbb23eaaf),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5842f3),
	.w1(32'h3b99fc1c),
	.w2(32'hbbb416a8),
	.w3(32'hbbd187cf),
	.w4(32'h3c30966f),
	.w5(32'hbc1f87c0),
	.w6(32'hbc1afe06),
	.w7(32'h3b874536),
	.w8(32'h3b3fd40a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04a36c),
	.w1(32'hba4414f0),
	.w2(32'hb8a38c40),
	.w3(32'hbbcc0337),
	.w4(32'hbbf70515),
	.w5(32'h3b7ace54),
	.w6(32'h3ac8270a),
	.w7(32'hbbfe10d3),
	.w8(32'hbbdbc457),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1d4cf),
	.w1(32'h3a8247f1),
	.w2(32'hbbc86792),
	.w3(32'hbb9a1c95),
	.w4(32'h3af2b76a),
	.w5(32'hbb4315e8),
	.w6(32'hbbf4de6e),
	.w7(32'h3b0bfb53),
	.w8(32'hbb58d2a2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc042ac5),
	.w1(32'hb899f813),
	.w2(32'hba0c1e67),
	.w3(32'hbc1c5f80),
	.w4(32'hb83e7cbd),
	.w5(32'hbbbd5084),
	.w6(32'hbbe9a24f),
	.w7(32'hbb972715),
	.w8(32'hbbd8ec45),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef1865),
	.w1(32'hbbab981e),
	.w2(32'h3bf45bbc),
	.w3(32'h3b52ac2d),
	.w4(32'h3b9e63a9),
	.w5(32'h3bc93c90),
	.w6(32'h3b2be806),
	.w7(32'h3b08f2cb),
	.w8(32'h3a4850a7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baec68c),
	.w1(32'h3be62980),
	.w2(32'h3b53795c),
	.w3(32'hba1bbe6c),
	.w4(32'h3b84c415),
	.w5(32'hbad72c10),
	.w6(32'h38ff9b86),
	.w7(32'h3b27816f),
	.w8(32'hbaf4ada4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55c093),
	.w1(32'h3aeca36c),
	.w2(32'h3aceb4c1),
	.w3(32'h3af20591),
	.w4(32'h3b050852),
	.w5(32'h3bf99817),
	.w6(32'h3c0ccbc4),
	.w7(32'hb9df1874),
	.w8(32'hbb84fb1e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a11ba),
	.w1(32'hbac5e9a1),
	.w2(32'hbb8105a9),
	.w3(32'h3beb7504),
	.w4(32'h3a89cf61),
	.w5(32'h3a9d601d),
	.w6(32'hb95d51e7),
	.w7(32'hba534f07),
	.w8(32'hbb0b85c7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2abe06),
	.w1(32'h3b80c8bc),
	.w2(32'h3a38af10),
	.w3(32'hbb58ee47),
	.w4(32'hbbe94684),
	.w5(32'hbc20b536),
	.w6(32'h3b0c9781),
	.w7(32'h3c0f763a),
	.w8(32'hba041c9a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba89839),
	.w1(32'hbaf1f3d1),
	.w2(32'h39ce566a),
	.w3(32'hbbf2b378),
	.w4(32'hbb3d0be6),
	.w5(32'h3a6d252d),
	.w6(32'h3a298840),
	.w7(32'hbbeb03ff),
	.w8(32'hbc8992f1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3de3e6),
	.w1(32'hbb078089),
	.w2(32'hbc23fbca),
	.w3(32'hbb8c683a),
	.w4(32'h3c0e69e0),
	.w5(32'h39b2ff7b),
	.w6(32'hbc099158),
	.w7(32'h3b0d52c5),
	.w8(32'hbb90eb04),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb707781),
	.w1(32'h3b11de82),
	.w2(32'hbb8d6a8a),
	.w3(32'h3bda9459),
	.w4(32'h3be75f40),
	.w5(32'h3bc4668f),
	.w6(32'h3a4ea57e),
	.w7(32'h3c0ceea1),
	.w8(32'h3b11999f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79a660),
	.w1(32'hbbc776e0),
	.w2(32'hbb604c41),
	.w3(32'h3c2d4f49),
	.w4(32'hbb9b5f9d),
	.w5(32'h3c62f786),
	.w6(32'h3b67fa8a),
	.w7(32'hbcd84159),
	.w8(32'hbbec325d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01c3be),
	.w1(32'hbc12bed3),
	.w2(32'hbbf1971b),
	.w3(32'h3aaf1a64),
	.w4(32'hbb78b798),
	.w5(32'h3abb49e8),
	.w6(32'hbb1db4d4),
	.w7(32'h3a228514),
	.w8(32'hb9a81fd3),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba83d30),
	.w1(32'hbb677d51),
	.w2(32'hba9d3a70),
	.w3(32'hbb9e8d7a),
	.w4(32'h3b4cdcf2),
	.w5(32'h3b5f11e0),
	.w6(32'h3b995f9c),
	.w7(32'hbc022d39),
	.w8(32'hbb0b402a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03c971),
	.w1(32'hbb14326f),
	.w2(32'hbb8d22a5),
	.w3(32'hbb1a2eb8),
	.w4(32'h3b13f58a),
	.w5(32'h3ba64f87),
	.w6(32'h3b25e1c2),
	.w7(32'h3c558f44),
	.w8(32'h3c8487fa),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0223b),
	.w1(32'hbc216791),
	.w2(32'h3c021643),
	.w3(32'h3b1c3f4e),
	.w4(32'hbbd85798),
	.w5(32'h3be9911d),
	.w6(32'h3be9e75e),
	.w7(32'h3ba44c3a),
	.w8(32'hbb9e599d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33d37f),
	.w1(32'h3c465ea9),
	.w2(32'h3c0c323e),
	.w3(32'h3bfdeba6),
	.w4(32'h3b7ec538),
	.w5(32'h3ab52a45),
	.w6(32'h3a0fb6ee),
	.w7(32'h3bebc9b3),
	.w8(32'h3c4553a5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78899d),
	.w1(32'h3bfcbb74),
	.w2(32'h3bd578d1),
	.w3(32'hba274d7f),
	.w4(32'h3c3047f3),
	.w5(32'h3c6e4f02),
	.w6(32'h3a8979e2),
	.w7(32'h3c501de4),
	.w8(32'hbba30b35),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c954921),
	.w1(32'h39e344d5),
	.w2(32'hbbd02817),
	.w3(32'h3bcabfb9),
	.w4(32'h3b00af7f),
	.w5(32'hbb1f89ac),
	.w6(32'hbbae18ca),
	.w7(32'h3b77ac9d),
	.w8(32'h3b1e03bf),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03bb86),
	.w1(32'h3b65fbc6),
	.w2(32'h3c1d2898),
	.w3(32'hbb8e2335),
	.w4(32'hb9196f0a),
	.w5(32'h3b4b9efc),
	.w6(32'hb9c90f5f),
	.w7(32'h3ad35806),
	.w8(32'hbaa10206),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942d99f),
	.w1(32'h3b5736a6),
	.w2(32'hb8a17a64),
	.w3(32'h380c073f),
	.w4(32'hbbe09e41),
	.w5(32'h3bc9f8db),
	.w6(32'h3ae2c90a),
	.w7(32'hbbd934ae),
	.w8(32'h3bb06a91),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba1003),
	.w1(32'hbba299f9),
	.w2(32'hbad79913),
	.w3(32'hbbd5f765),
	.w4(32'h3be35c2c),
	.w5(32'h3b64b20f),
	.w6(32'hbbc54086),
	.w7(32'hbb4d7c8b),
	.w8(32'hba782a72),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafab1b8),
	.w1(32'hbb86a75e),
	.w2(32'hbc112c64),
	.w3(32'hba82fc87),
	.w4(32'h3b5508d6),
	.w5(32'hba9f7802),
	.w6(32'hbb859181),
	.w7(32'hbae37d25),
	.w8(32'h3ad244a4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8946eb),
	.w1(32'h3aeca0a3),
	.w2(32'hbb26499a),
	.w3(32'hbc0a6815),
	.w4(32'h3bd56140),
	.w5(32'h3b575301),
	.w6(32'h393a71fc),
	.w7(32'h3c623a4e),
	.w8(32'h3c3ab165),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be31e88),
	.w1(32'h3c2226f4),
	.w2(32'hbb1b818f),
	.w3(32'h3bd64c40),
	.w4(32'h3bd1e4e2),
	.w5(32'h3ae87a71),
	.w6(32'h3c73c065),
	.w7(32'h3bf1b7ca),
	.w8(32'hba883abd),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51300e),
	.w1(32'hbb0dc1ed),
	.w2(32'hbb3f9d58),
	.w3(32'h3c47921f),
	.w4(32'hbae88f30),
	.w5(32'hbb2a97b3),
	.w6(32'h3bef0a0b),
	.w7(32'h3b29d9a3),
	.w8(32'hbb7929b8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b8f06),
	.w1(32'h3b69c0bc),
	.w2(32'h3b34cefa),
	.w3(32'hbb2d7b90),
	.w4(32'h3ad67214),
	.w5(32'h3bbbec02),
	.w6(32'h32b93100),
	.w7(32'hbbfc59b6),
	.w8(32'hbb242d5c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d314c),
	.w1(32'hbaf567b4),
	.w2(32'h3c00009b),
	.w3(32'hb9c3a759),
	.w4(32'hbbdb0720),
	.w5(32'hbc25985c),
	.w6(32'h38cbf04b),
	.w7(32'h3b6c5e41),
	.w8(32'h3b9db485),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a54c4),
	.w1(32'h3c02f506),
	.w2(32'h3b86d151),
	.w3(32'hbc1aa0b3),
	.w4(32'hba9685e9),
	.w5(32'hbc20d993),
	.w6(32'h3977cb2c),
	.w7(32'h3c32cd8b),
	.w8(32'h3c68e807),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadae30b),
	.w1(32'hbc218f8b),
	.w2(32'hbc2dd4a8),
	.w3(32'hbbfc92b3),
	.w4(32'hbb882690),
	.w5(32'hbbad9849),
	.w6(32'h3c1bc3e4),
	.w7(32'hbb16f96f),
	.w8(32'h3ba3be1a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c59452),
	.w1(32'h3bec20e6),
	.w2(32'h3bd95295),
	.w3(32'hbc066f1b),
	.w4(32'h3bc2922b),
	.w5(32'h3ae2858e),
	.w6(32'hba17aa18),
	.w7(32'h3bc54ddc),
	.w8(32'h3ab05622),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0d425),
	.w1(32'h3bced1aa),
	.w2(32'h3aedd001),
	.w3(32'hbc2c7adc),
	.w4(32'h3b985212),
	.w5(32'h3bdf5d52),
	.w6(32'hbb133934),
	.w7(32'h39d0667f),
	.w8(32'hbb227b48),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a747b),
	.w1(32'hbb35c96f),
	.w2(32'hbae7015e),
	.w3(32'hbbefd568),
	.w4(32'hbb0aef3a),
	.w5(32'h3be39ded),
	.w6(32'h399bcdff),
	.w7(32'hbbb48c4d),
	.w8(32'h3afef5f7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ecc41),
	.w1(32'h3a91b62c),
	.w2(32'h3b8bb839),
	.w3(32'h3ae9d0c9),
	.w4(32'h3bb3b49b),
	.w5(32'h3b9b84da),
	.w6(32'hbb0a39b5),
	.w7(32'h3b278ba0),
	.w8(32'hbb06700f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb403b67),
	.w1(32'hbc12abb0),
	.w2(32'hbc074f50),
	.w3(32'hbbc21b1b),
	.w4(32'h3b6e8f72),
	.w5(32'hbbcc8925),
	.w6(32'hbc86e924),
	.w7(32'hbb40508c),
	.w8(32'h39bea8a1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc50216),
	.w1(32'h3c9fa639),
	.w2(32'h3c3baf2f),
	.w3(32'hbaa4dfc2),
	.w4(32'hba6980f6),
	.w5(32'hbc1281c2),
	.w6(32'hba4ba9b3),
	.w7(32'h3c27ae2b),
	.w8(32'h3bce22fc),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c031ea3),
	.w1(32'h3bcb6a2e),
	.w2(32'h3c222161),
	.w3(32'hbb89ecde),
	.w4(32'h3b941793),
	.w5(32'h3b752918),
	.w6(32'hba339cb2),
	.w7(32'hbb654496),
	.w8(32'hb9af7325),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c299a18),
	.w1(32'h3be5cb5e),
	.w2(32'h3bcc08cc),
	.w3(32'h3c00ec5a),
	.w4(32'h3b895028),
	.w5(32'h3c25808b),
	.w6(32'h399cd60a),
	.w7(32'h3c4d0204),
	.w8(32'h3bcf7a66),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c512bff),
	.w1(32'h3bd71344),
	.w2(32'h3bdd4e2c),
	.w3(32'h3c1a4035),
	.w4(32'h3b24cf56),
	.w5(32'h3795b99a),
	.w6(32'h3b346b09),
	.w7(32'hb930a5bb),
	.w8(32'hbb942322),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72886b),
	.w1(32'hbbe25cc8),
	.w2(32'hbbf61dde),
	.w3(32'h3b9a6ecc),
	.w4(32'hb642934c),
	.w5(32'h39643ac0),
	.w6(32'h3a174466),
	.w7(32'h3bd93030),
	.w8(32'h3bc9657a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfefa7a),
	.w1(32'h3900f99f),
	.w2(32'hbb7ce3c3),
	.w3(32'h3b94260e),
	.w4(32'hbb2a0023),
	.w5(32'h3b232f93),
	.w6(32'h3c3d8923),
	.w7(32'hbb7b0fd5),
	.w8(32'hb8257548),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0df45),
	.w1(32'hbbf7a6b9),
	.w2(32'hba01d644),
	.w3(32'hbb13ea84),
	.w4(32'hbbeea7fb),
	.w5(32'hbb3feb72),
	.w6(32'h3b85de7d),
	.w7(32'h3acc6549),
	.w8(32'h3b23459b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4a01a),
	.w1(32'hbbd86436),
	.w2(32'hbc202201),
	.w3(32'hbb863806),
	.w4(32'h3be33d57),
	.w5(32'hbb6f7cbb),
	.w6(32'h3a207dc9),
	.w7(32'h3bfa9cb4),
	.w8(32'h3c0e7c41),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97782d),
	.w1(32'hbc278e4a),
	.w2(32'hbbf9750e),
	.w3(32'hba106095),
	.w4(32'hbba6e8a7),
	.w5(32'hbc16a077),
	.w6(32'h3c4d35f8),
	.w7(32'hbb542648),
	.w8(32'hbbcb23d3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c0753),
	.w1(32'hbaba01b6),
	.w2(32'hbb5fd929),
	.w3(32'hbbebaa1d),
	.w4(32'h399b0b2e),
	.w5(32'hba1c327f),
	.w6(32'hba107a38),
	.w7(32'h3a8c244d),
	.w8(32'hb9efdec5),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba843bae),
	.w1(32'hba78f615),
	.w2(32'h398c2d8e),
	.w3(32'h38bdd498),
	.w4(32'hb79f6146),
	.w5(32'hb942349d),
	.w6(32'h3a7475d5),
	.w7(32'h3a706fd1),
	.w8(32'hba486195),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965d8e1),
	.w1(32'hb9736565),
	.w2(32'hb90f09a1),
	.w3(32'hb8784a9f),
	.w4(32'h3a01305e),
	.w5(32'hba94bf84),
	.w6(32'h39257682),
	.w7(32'h3a128a85),
	.w8(32'h39737752),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91831b),
	.w1(32'hbb826f72),
	.w2(32'hba4d0efc),
	.w3(32'hbb413b9e),
	.w4(32'h3abadc33),
	.w5(32'h3b8d99c8),
	.w6(32'hbaacdfd3),
	.w7(32'h3b477f1d),
	.w8(32'h3b9ae9b9),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba593a),
	.w1(32'h3950960a),
	.w2(32'hb847598d),
	.w3(32'h398aad45),
	.w4(32'h39384827),
	.w5(32'h371d8dc1),
	.w6(32'h39f7701a),
	.w7(32'h39dfcffb),
	.w8(32'h39bfb212),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcf8bb),
	.w1(32'hba61572b),
	.w2(32'hbaca4f43),
	.w3(32'hba4121e0),
	.w4(32'h39b879f1),
	.w5(32'h3a25e399),
	.w6(32'h3aa934a5),
	.w7(32'h3a96bc7e),
	.w8(32'h39a1af2e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b2576),
	.w1(32'hb6933390),
	.w2(32'hbb4ba846),
	.w3(32'h3a8ceb49),
	.w4(32'h3aa49761),
	.w5(32'hbb50a87d),
	.w6(32'h3a3e24d4),
	.w7(32'h3a6740aa),
	.w8(32'hbb8fd678),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a2e6f),
	.w1(32'hb9f96b4e),
	.w2(32'hbaec4061),
	.w3(32'hba02f201),
	.w4(32'h3a1ef234),
	.w5(32'hb9b5bb4c),
	.w6(32'h3a61903c),
	.w7(32'h3afba623),
	.w8(32'hb98b6511),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4556e),
	.w1(32'h3a9a5281),
	.w2(32'h3a7fe616),
	.w3(32'h3a2d2141),
	.w4(32'h3a42a33e),
	.w5(32'hb944fedf),
	.w6(32'h3a45c306),
	.w7(32'h39597154),
	.w8(32'h39d9b0c8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8c662),
	.w1(32'h3a27240d),
	.w2(32'hbb86d776),
	.w3(32'hbac41f66),
	.w4(32'h3a6ebcb4),
	.w5(32'hbabd33b6),
	.w6(32'h3aa365dd),
	.w7(32'h3a23bad7),
	.w8(32'hbb5a92ed),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56e622),
	.w1(32'hbad19406),
	.w2(32'hbb49eebf),
	.w3(32'hbb723da0),
	.w4(32'h397e7395),
	.w5(32'hba59f266),
	.w6(32'hba71fa08),
	.w7(32'h3b136146),
	.w8(32'h3aef21b6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf178fe),
	.w1(32'hbb375dd3),
	.w2(32'hbb8e17a8),
	.w3(32'h3a07e785),
	.w4(32'hba50a139),
	.w5(32'hbb2db8a1),
	.w6(32'h3a1c1452),
	.w7(32'h38b9948d),
	.w8(32'hba829a0d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3791b3ed),
	.w1(32'hb9bf2366),
	.w2(32'hb90a4242),
	.w3(32'hb9ae04a2),
	.w4(32'hba1f8551),
	.w5(32'hb91ec648),
	.w6(32'h3893b7a2),
	.w7(32'hb986b831),
	.w8(32'hb994ab59),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb868af58),
	.w1(32'h39445ffa),
	.w2(32'h398a1bc4),
	.w3(32'h39d8bbd0),
	.w4(32'h39a6e547),
	.w5(32'hb941ec62),
	.w6(32'h39227773),
	.w7(32'hb78c7f08),
	.w8(32'hb9d4dcb4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e1d41),
	.w1(32'hbb6623a0),
	.w2(32'hba941d5b),
	.w3(32'h3b88c6f2),
	.w4(32'h3b81dae0),
	.w5(32'h3b0110b2),
	.w6(32'h39c1b096),
	.w7(32'h3a9239e1),
	.w8(32'h3a6bfb95),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7724b),
	.w1(32'hbade550d),
	.w2(32'hba073be9),
	.w3(32'hb9c5569b),
	.w4(32'h3b20849e),
	.w5(32'h3a86a9df),
	.w6(32'hbb144eb6),
	.w7(32'h3afb25e9),
	.w8(32'h3b0bdcde),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb288784),
	.w1(32'hbacfa2bb),
	.w2(32'hbb68ca8a),
	.w3(32'hb8270819),
	.w4(32'h39965299),
	.w5(32'hbac2dce3),
	.w6(32'hb781db49),
	.w7(32'h3878d204),
	.w8(32'hbaf15e94),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cde0e7),
	.w1(32'hb90f3ccb),
	.w2(32'h3a604c93),
	.w3(32'hbbb3c340),
	.w4(32'hbbb8186d),
	.w5(32'hbae46354),
	.w6(32'h3ba5f36c),
	.w7(32'hba98ac21),
	.w8(32'h3ac3d339),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6116c0),
	.w1(32'hb9a5ab03),
	.w2(32'hb84e1edc),
	.w3(32'hba386703),
	.w4(32'hb9ba13f6),
	.w5(32'h3abb6a73),
	.w6(32'hba659aaa),
	.w7(32'hba7ae133),
	.w8(32'h3a56c325),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac84ed7),
	.w1(32'hbaef0a25),
	.w2(32'h370dfc74),
	.w3(32'hbaa0eb22),
	.w4(32'h39962143),
	.w5(32'h3b09cd5a),
	.w6(32'hba1b7ea3),
	.w7(32'h3a94f9d6),
	.w8(32'h3aa30f30),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f68c4),
	.w1(32'hbbada9fc),
	.w2(32'h3a114601),
	.w3(32'h3a61d582),
	.w4(32'hbb830b90),
	.w5(32'hbb3422f4),
	.w6(32'hba72a98d),
	.w7(32'hb995da8c),
	.w8(32'h3b283a1e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecf41c),
	.w1(32'hbb23120b),
	.w2(32'hba83fca7),
	.w3(32'hbb0d060e),
	.w4(32'h3a0bf33e),
	.w5(32'h3ad6d721),
	.w6(32'hbb4affa9),
	.w7(32'h3affe2d8),
	.w8(32'h3a9283c9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8ced1),
	.w1(32'hbb4483fe),
	.w2(32'h3b5dad0e),
	.w3(32'hbb634c54),
	.w4(32'hba4a02a9),
	.w5(32'h3ba3569c),
	.w6(32'hbb1318aa),
	.w7(32'h3b148e9d),
	.w8(32'h3bf08dc4),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878d2e),
	.w1(32'h3a0bdf21),
	.w2(32'hba928cb3),
	.w3(32'h3abc26c9),
	.w4(32'hba31ab3e),
	.w5(32'hbb13cf14),
	.w6(32'h3aa92805),
	.w7(32'hbac8a4a3),
	.w8(32'hbb7c00b8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0b1c8),
	.w1(32'hba34585f),
	.w2(32'hbbb3eeb0),
	.w3(32'hbaf092a5),
	.w4(32'h379daf36),
	.w5(32'hbb2e7d39),
	.w6(32'hb9663542),
	.w7(32'h3a24fa44),
	.w8(32'hbb8caeda),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f93c73),
	.w1(32'h37ae8ff2),
	.w2(32'hb9b3aebc),
	.w3(32'hb8659fb6),
	.w4(32'hb9ad9dfd),
	.w5(32'hb97640ae),
	.w6(32'h39aaa1b6),
	.w7(32'hba22b86d),
	.w8(32'hba8fc273),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38db7084),
	.w1(32'h398f998f),
	.w2(32'h39b81675),
	.w3(32'h39f2a97c),
	.w4(32'hb89612ba),
	.w5(32'hb714eee6),
	.w6(32'hb98ba1f7),
	.w7(32'hb5d62b14),
	.w8(32'hb9b94c71),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa18809),
	.w1(32'h3a790f07),
	.w2(32'h39dad7ba),
	.w3(32'h3b1e547b),
	.w4(32'h3b1f8f96),
	.w5(32'h3a956e0e),
	.w6(32'h3aa998b8),
	.w7(32'hb8ce244b),
	.w8(32'hba1e6d28),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946d780),
	.w1(32'hba075dbb),
	.w2(32'hb8c6175d),
	.w3(32'hb9d7f51b),
	.w4(32'hba3adc7e),
	.w5(32'hb95917a0),
	.w6(32'hb9ee0454),
	.w7(32'hba8a645d),
	.w8(32'h38f765ad),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4c56),
	.w1(32'hbb650dd4),
	.w2(32'hbb21c7e7),
	.w3(32'hbb05df07),
	.w4(32'hbb722474),
	.w5(32'hbb05ff73),
	.w6(32'hbac39053),
	.w7(32'hb91527a3),
	.w8(32'hbacbd0f4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd210f1),
	.w1(32'hbb856919),
	.w2(32'hbaa15b30),
	.w3(32'hbac2d171),
	.w4(32'h3b03207d),
	.w5(32'h3b0397a9),
	.w6(32'hbb234627),
	.w7(32'hba1b03a9),
	.w8(32'h3b7b0829),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e2a8a),
	.w1(32'hba352469),
	.w2(32'hbafa30c8),
	.w3(32'hb9652ea7),
	.w4(32'h3a76036e),
	.w5(32'h3a790d05),
	.w6(32'hb9d8f955),
	.w7(32'h3a48a6f7),
	.w8(32'hb5a16709),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956c18a),
	.w1(32'hb98bd14b),
	.w2(32'hb917ca0a),
	.w3(32'hb8237a72),
	.w4(32'hb99f4049),
	.w5(32'h3a01c404),
	.w6(32'hb99ac757),
	.w7(32'hb975c5f2),
	.w8(32'hb6e7bdf7),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c1743),
	.w1(32'hbbda1225),
	.w2(32'hbb14db74),
	.w3(32'hbb9f8755),
	.w4(32'h3a977f3c),
	.w5(32'h3c08ec29),
	.w6(32'hbb97a16c),
	.w7(32'h3a81ad8a),
	.w8(32'h3c1dab1e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb106df3),
	.w1(32'hbabb50d3),
	.w2(32'hba09016c),
	.w3(32'hb9488e79),
	.w4(32'h399bbbaa),
	.w5(32'h396a2f57),
	.w6(32'h393c9844),
	.w7(32'h3a70e3c3),
	.w8(32'h3aa8e792),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86b2f4),
	.w1(32'h3a065368),
	.w2(32'h3a2fc8cd),
	.w3(32'h39e3981e),
	.w4(32'h3a4b42e8),
	.w5(32'h3a84c29a),
	.w6(32'h399062c1),
	.w7(32'h3a815131),
	.w8(32'h3a81db75),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafba6d9),
	.w1(32'hbb05aa02),
	.w2(32'hbb0af93f),
	.w3(32'hbb0d89f9),
	.w4(32'hbaab2835),
	.w5(32'hb9a2c7b2),
	.w6(32'h3958651c),
	.w7(32'h38f50bf8),
	.w8(32'h3a87ca30),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bf37b),
	.w1(32'hb9114e82),
	.w2(32'h3959b7a0),
	.w3(32'h384dc66a),
	.w4(32'hb7a329e8),
	.w5(32'h39873015),
	.w6(32'h3974714c),
	.w7(32'hb9b37c6c),
	.w8(32'hba668726),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b2cbc3),
	.w1(32'h39ca3d09),
	.w2(32'h39285e00),
	.w3(32'hb9db960f),
	.w4(32'h399cd31a),
	.w5(32'h3a02934d),
	.w6(32'hbac1b82d),
	.w7(32'h39d57acc),
	.w8(32'h38cf5016),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3955ce30),
	.w1(32'hb8a79934),
	.w2(32'h38b68fe8),
	.w3(32'h3abdc866),
	.w4(32'h3a0e95e6),
	.w5(32'h39c3ce18),
	.w6(32'h3aaa3fae),
	.w7(32'h3a534a22),
	.w8(32'h39e245b0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365f55bf),
	.w1(32'hb994cba4),
	.w2(32'h3982d87f),
	.w3(32'h3930aca1),
	.w4(32'hba1a92ad),
	.w5(32'hb8e7c056),
	.w6(32'hb88e30ff),
	.w7(32'h387b66e9),
	.w8(32'hb7bf6ba3),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35cdde),
	.w1(32'h39fdb211),
	.w2(32'h3a2a98e6),
	.w3(32'h3a844dc4),
	.w4(32'h393cae56),
	.w5(32'h3a78907e),
	.w6(32'h3aa69999),
	.w7(32'h37b1ec7c),
	.w8(32'h39b49a54),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7a618),
	.w1(32'hba4da904),
	.w2(32'hbbb9cc1b),
	.w3(32'hbc01e6bb),
	.w4(32'h3a9f98de),
	.w5(32'hba3976bb),
	.w6(32'h3b26d603),
	.w7(32'h3c01c26c),
	.w8(32'h3b42d205),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9249cf),
	.w1(32'hbb40cc59),
	.w2(32'hbb86d355),
	.w3(32'hbb1a9c0d),
	.w4(32'h3a030067),
	.w5(32'h391c8d9b),
	.w6(32'h395876fc),
	.w7(32'h3b0d7d38),
	.w8(32'h3af4698e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fd33a),
	.w1(32'hbaf8a3f2),
	.w2(32'hbb801e75),
	.w3(32'hbb6cd6d5),
	.w4(32'h3ab7112b),
	.w5(32'hba3ee161),
	.w6(32'h3ad32307),
	.w7(32'h3b77945d),
	.w8(32'h3b04ce21),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b3a1fd),
	.w1(32'hba29d340),
	.w2(32'hb9c6df69),
	.w3(32'hb9810124),
	.w4(32'hb933f7a9),
	.w5(32'hb9a01024),
	.w6(32'h395cd707),
	.w7(32'hba427cc3),
	.w8(32'h39c10228),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba325d06),
	.w1(32'hb709699c),
	.w2(32'hb868149a),
	.w3(32'h39821f24),
	.w4(32'h3a0b237f),
	.w5(32'h39f78673),
	.w6(32'hb88b8530),
	.w7(32'h39c62468),
	.w8(32'h3a30dcd0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81fc213),
	.w1(32'hb9f0d81e),
	.w2(32'hb9e8d3e5),
	.w3(32'h39b28f8b),
	.w4(32'hb9b159b7),
	.w5(32'hb97bae1f),
	.w6(32'h3a71df23),
	.w7(32'hb9eac5fc),
	.w8(32'hb980d194),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f057dd),
	.w1(32'hb9904ad8),
	.w2(32'hb9f26bc2),
	.w3(32'hba0f97c1),
	.w4(32'h3940a8bf),
	.w5(32'hb9babe37),
	.w6(32'hba09c006),
	.w7(32'h381e9d6f),
	.w8(32'hb98d0d29),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefbfb5),
	.w1(32'hba5f634a),
	.w2(32'hb972769b),
	.w3(32'hbb75f1ca),
	.w4(32'h3b350c71),
	.w5(32'h3bb849bd),
	.w6(32'h382adc84),
	.w7(32'h3ba4325c),
	.w8(32'h3baeb858),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6cedb),
	.w1(32'h395233d9),
	.w2(32'hba0c21d2),
	.w3(32'hba0ec254),
	.w4(32'h3959091b),
	.w5(32'hb9da57d9),
	.w6(32'h3833423e),
	.w7(32'h38c9f656),
	.w8(32'h3a24bebb),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967850e),
	.w1(32'h3a46011d),
	.w2(32'h3aa53fb0),
	.w3(32'h3989f9ed),
	.w4(32'h3a9ec77b),
	.w5(32'h3a85d154),
	.w6(32'h3a50a351),
	.w7(32'h3aa7216c),
	.w8(32'h3aa9383c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19e3a6),
	.w1(32'hba860368),
	.w2(32'hba556ee6),
	.w3(32'hbb172335),
	.w4(32'hba917c89),
	.w5(32'h3a27e2e7),
	.w6(32'hba94e508),
	.w7(32'h3a9ead50),
	.w8(32'h3adb22f1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39093b62),
	.w1(32'h3a07d7c6),
	.w2(32'h39cd3d32),
	.w3(32'h39b7d1d1),
	.w4(32'h398fbcd2),
	.w5(32'h39359dd9),
	.w6(32'h39e5de93),
	.w7(32'hb9bd4a7e),
	.w8(32'hb9c06843),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5482f7),
	.w1(32'h39d1ba02),
	.w2(32'h3a135ffa),
	.w3(32'hba223f1d),
	.w4(32'h39ff6262),
	.w5(32'h3774dc64),
	.w6(32'h398af0dd),
	.w7(32'hb7866337),
	.w8(32'h38c01d49),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba418fea),
	.w1(32'hb934d0d7),
	.w2(32'hb97200bb),
	.w3(32'hb997623d),
	.w4(32'h3a59fcfe),
	.w5(32'hba02a0ea),
	.w6(32'hb9153b41),
	.w7(32'h3a718b03),
	.w8(32'hba025497),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd86db),
	.w1(32'hba95be7f),
	.w2(32'hbbaf34d2),
	.w3(32'hbc2127dc),
	.w4(32'h3b932c86),
	.w5(32'h3bcdd9d3),
	.w6(32'h3802cfa6),
	.w7(32'h3c35ac83),
	.w8(32'h3c2abc9d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a65bd),
	.w1(32'hbab96541),
	.w2(32'h380dd40c),
	.w3(32'h3a0445c0),
	.w4(32'hba991d7c),
	.w5(32'hb9f41155),
	.w6(32'h39c0e6ac),
	.w7(32'hbab7db57),
	.w8(32'hbac8c95c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb842c2),
	.w1(32'hbb5e2261),
	.w2(32'hba58a13a),
	.w3(32'h3a63df07),
	.w4(32'h3af1d9dc),
	.w5(32'hba2e13f9),
	.w6(32'h3a5ea68f),
	.w7(32'hbb534182),
	.w8(32'hbb4cb5be),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule