module layer_8_featuremap_32(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb301611),
	.w1(32'hbb602b80),
	.w2(32'hbb439481),
	.w3(32'hbb177622),
	.w4(32'hbb18e368),
	.w5(32'hbb15c857),
	.w6(32'hbbb99e79),
	.w7(32'hbb9cd34b),
	.w8(32'hbb81d798),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a08f29),
	.w1(32'hba062678),
	.w2(32'hba3dbb6f),
	.w3(32'hba28f068),
	.w4(32'hba96c6c7),
	.w5(32'hba7e89ef),
	.w6(32'hbb061a87),
	.w7(32'hbad82a76),
	.w8(32'hba90a0e8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d73d2),
	.w1(32'h3a5db9e0),
	.w2(32'hba1b048c),
	.w3(32'h3aacb1a4),
	.w4(32'h3a0e8754),
	.w5(32'hb9dd6f1d),
	.w6(32'h3b0a4e04),
	.w7(32'h3ab2a2da),
	.w8(32'h39fb7d69),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7e67d),
	.w1(32'hba99e480),
	.w2(32'hba98ae07),
	.w3(32'h398f39b7),
	.w4(32'hbb16c575),
	.w5(32'hbad07a19),
	.w6(32'h3af23134),
	.w7(32'h3b18a929),
	.w8(32'hbb01e6fc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3f15c),
	.w1(32'h3a33ecb8),
	.w2(32'hb83a3e2f),
	.w3(32'h3ab150aa),
	.w4(32'h3accea64),
	.w5(32'h3a85ff34),
	.w6(32'hb9f3ed04),
	.w7(32'hb9f51f1f),
	.w8(32'hbbb63a9f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b4e69),
	.w1(32'hbbf4bec5),
	.w2(32'hbba2c181),
	.w3(32'hbbe2753d),
	.w4(32'hbc04d59b),
	.w5(32'hbb9af1ed),
	.w6(32'hbb09c97c),
	.w7(32'hbb5075ad),
	.w8(32'h3b2254a8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5645fd),
	.w1(32'hbb6b798f),
	.w2(32'hbb4f11ab),
	.w3(32'hbb4d6a82),
	.w4(32'hbb51508e),
	.w5(32'hbb48e9b5),
	.w6(32'hbb6ed8a1),
	.w7(32'hbb371b4d),
	.w8(32'hbb1ccd2d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac905cc),
	.w1(32'h3af2f59a),
	.w2(32'h3988cc82),
	.w3(32'h3b0ecbc8),
	.w4(32'h3b3d089b),
	.w5(32'h3a715ac1),
	.w6(32'h3ac49b50),
	.w7(32'h3ae7c025),
	.w8(32'hbb011970),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade98e2),
	.w1(32'hb950ea25),
	.w2(32'h397fce28),
	.w3(32'h3a9cdff8),
	.w4(32'h3a357591),
	.w5(32'h36cf0b29),
	.w6(32'hb9898786),
	.w7(32'hba64a836),
	.w8(32'h3bf5754c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d1b26),
	.w1(32'hb9470b30),
	.w2(32'hbace6fd6),
	.w3(32'hbb6aab6d),
	.w4(32'hbb6b7f1e),
	.w5(32'hba77c919),
	.w6(32'h3984582f),
	.w7(32'hb9572e1c),
	.w8(32'hbb822645),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18b80c),
	.w1(32'hba97b308),
	.w2(32'hbb0edaf2),
	.w3(32'hba6e262e),
	.w4(32'h3a99a5c0),
	.w5(32'hba658a29),
	.w6(32'hbb1989a1),
	.w7(32'hba245798),
	.w8(32'hbaefa990),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c370e),
	.w1(32'hbabc470b),
	.w2(32'hbad58bd3),
	.w3(32'h393c729e),
	.w4(32'hba1d8978),
	.w5(32'hba14f00f),
	.w6(32'hbb198411),
	.w7(32'hbb61dc0d),
	.w8(32'hbb7ff56e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c2e41),
	.w1(32'hb905dab2),
	.w2(32'hba250077),
	.w3(32'h39d98c96),
	.w4(32'hba8f8c4a),
	.w5(32'hbac171f8),
	.w6(32'hb9980dd6),
	.w7(32'hbab31a7f),
	.w8(32'hbbde59f4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be05b),
	.w1(32'hbbc81720),
	.w2(32'hbbd10823),
	.w3(32'hbc105cf9),
	.w4(32'hbbd651b4),
	.w5(32'hbbcdeaad),
	.w6(32'hbbb2e0c5),
	.w7(32'hbba17b5e),
	.w8(32'hbb3c64db),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936922),
	.w1(32'hbb629d0e),
	.w2(32'hbb909f59),
	.w3(32'hbbbee334),
	.w4(32'hbb9be108),
	.w5(32'hbbab6d9e),
	.w6(32'hbb8c5227),
	.w7(32'hbba0e90b),
	.w8(32'hba41f7ea),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84d840),
	.w1(32'h39e91c01),
	.w2(32'h39b7c3e6),
	.w3(32'h3a94dbb0),
	.w4(32'h3a0778c8),
	.w5(32'h39f0f901),
	.w6(32'h3a6d25b2),
	.w7(32'h3a30b5cf),
	.w8(32'h3b1f1a72),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f8263),
	.w1(32'hbba76a96),
	.w2(32'hbb53de5c),
	.w3(32'hbbae6431),
	.w4(32'hbb30c349),
	.w5(32'h3a9e3695),
	.w6(32'h3aa3556b),
	.w7(32'h3bef0d5a),
	.w8(32'hba80aa2c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37b7fc),
	.w1(32'h3acfa108),
	.w2(32'hba8b7554),
	.w3(32'h3a152682),
	.w4(32'h3a819bb2),
	.w5(32'h3a352b5e),
	.w6(32'h3ac38fca),
	.w7(32'hb9d00f31),
	.w8(32'hb974c54e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb353078),
	.w1(32'h3b0a3036),
	.w2(32'hbb722e7b),
	.w3(32'h3b27bf0f),
	.w4(32'h3c09c8e9),
	.w5(32'h3b7d5bb3),
	.w6(32'hbc14aba8),
	.w7(32'hbb9f41d2),
	.w8(32'hbb7417ee),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba537b8),
	.w1(32'h3baede76),
	.w2(32'h3c6c6ffa),
	.w3(32'h3b970fa1),
	.w4(32'h3b8ab43e),
	.w5(32'h3c15018b),
	.w6(32'h3c056ad5),
	.w7(32'h3c5328ae),
	.w8(32'h3b556577),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04f318),
	.w1(32'h39915ca9),
	.w2(32'h3b3b3695),
	.w3(32'hbb111c5f),
	.w4(32'hbb9192e5),
	.w5(32'h3af77186),
	.w6(32'hbb9f717e),
	.w7(32'hbbbe6b84),
	.w8(32'hbb4f0aae),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b085d81),
	.w1(32'hbb040495),
	.w2(32'h39c5bd39),
	.w3(32'hbb050533),
	.w4(32'hbb8d4d34),
	.w5(32'hba1aa292),
	.w6(32'hbb460447),
	.w7(32'hbb8a86f2),
	.w8(32'h3c84cd19),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53c3ab),
	.w1(32'h3c574900),
	.w2(32'h3c08ea76),
	.w3(32'h3c9a91b6),
	.w4(32'h3cbfd4a6),
	.w5(32'h3c8bb2e0),
	.w6(32'h3c1de916),
	.w7(32'h3c323223),
	.w8(32'hba6e95f2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ead191),
	.w1(32'h3b05bda0),
	.w2(32'h3a9d671f),
	.w3(32'hb94d0b4b),
	.w4(32'h3ac02077),
	.w5(32'h3ac1751b),
	.w6(32'hba18c9cf),
	.w7(32'h39b75796),
	.w8(32'h3b3a16b2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b303b2c),
	.w1(32'h3b1f5e7c),
	.w2(32'h3b370c95),
	.w3(32'h3b762910),
	.w4(32'h3b16a71a),
	.w5(32'h3b1ae751),
	.w6(32'h3afe1980),
	.w7(32'h3ba9bc90),
	.w8(32'h3c861fd1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10f36f),
	.w1(32'h3be6c9e5),
	.w2(32'h3bcf2862),
	.w3(32'h3c5ab200),
	.w4(32'h3c660240),
	.w5(32'h3c5a7190),
	.w6(32'h3bf2163c),
	.w7(32'h3c10c0ce),
	.w8(32'h3c2cd919),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba21035),
	.w1(32'h3b6dec3f),
	.w2(32'h3b48dc8e),
	.w3(32'h3c04856a),
	.w4(32'h3bea24db),
	.w5(32'h3bc1eb88),
	.w6(32'h3bd2d8c5),
	.w7(32'h3baea3e8),
	.w8(32'hbb990537),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcae266),
	.w1(32'h3bb53426),
	.w2(32'h3c21c894),
	.w3(32'h3b5e6a79),
	.w4(32'h3cd402e0),
	.w5(32'h3cb824a1),
	.w6(32'hbca205c5),
	.w7(32'hbc87a187),
	.w8(32'h3c69c37e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d4ff5),
	.w1(32'hba264c3a),
	.w2(32'h3a8bf6c0),
	.w3(32'h3b58bf7b),
	.w4(32'h3a196d12),
	.w5(32'h3ab26304),
	.w6(32'hba8d0a70),
	.w7(32'hba9a4e0c),
	.w8(32'hba51b233),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea396c),
	.w1(32'h3aa3d6fd),
	.w2(32'h3accec72),
	.w3(32'h3a860eb2),
	.w4(32'h39cec12c),
	.w5(32'h3ac47ace),
	.w6(32'h3afcb178),
	.w7(32'h3ac5aefa),
	.w8(32'hba264025),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0aec6f),
	.w1(32'hbc21eb60),
	.w2(32'hbb828e20),
	.w3(32'hbbd0779f),
	.w4(32'hbc491fc0),
	.w5(32'hbc466f69),
	.w6(32'hbbba7c36),
	.w7(32'hbbc815cc),
	.w8(32'h39146a2f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11afd4),
	.w1(32'h3c2845a9),
	.w2(32'h3b8869bb),
	.w3(32'h3bb6c9ec),
	.w4(32'h3bff9db9),
	.w5(32'h3bfff2fe),
	.w6(32'h3b788c38),
	.w7(32'hbaae18d8),
	.w8(32'hbac95018),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02c63b),
	.w1(32'h3a901ab8),
	.w2(32'h3aca0a46),
	.w3(32'hbacbcc3c),
	.w4(32'hbaf011f2),
	.w5(32'h36f3d077),
	.w6(32'hba9de1f4),
	.w7(32'h3a5ba911),
	.w8(32'hbb482881),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad117c5),
	.w1(32'hbbb9e2a9),
	.w2(32'hbb62244b),
	.w3(32'h3a4b99ed),
	.w4(32'h3b5322a2),
	.w5(32'h3b529d85),
	.w6(32'hbb669846),
	.w7(32'hbba9c82a),
	.w8(32'hbbe5ec67),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0e45a),
	.w1(32'hbbb11f9e),
	.w2(32'hbba7a4a2),
	.w3(32'hbc158311),
	.w4(32'hbc00216c),
	.w5(32'hbbd23f61),
	.w6(32'hbb977ab8),
	.w7(32'hbb9d050c),
	.w8(32'hba8b2c7f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bd78c),
	.w1(32'hbad58c8e),
	.w2(32'hbb17ab51),
	.w3(32'hbb3182ae),
	.w4(32'hba4de20b),
	.w5(32'hbab06749),
	.w6(32'hbbc8d863),
	.w7(32'hbba3e099),
	.w8(32'h3b127d74),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9a805),
	.w1(32'hbafaca07),
	.w2(32'hbb9200d2),
	.w3(32'h3c0dd6df),
	.w4(32'h3b4e7c5d),
	.w5(32'hb9107a59),
	.w6(32'h3af1852f),
	.w7(32'hba00987f),
	.w8(32'hbac045ef),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4f99e),
	.w1(32'h3a85bffc),
	.w2(32'h3a86d81c),
	.w3(32'hb8371605),
	.w4(32'hba2183af),
	.w5(32'hb8ca41ab),
	.w6(32'hba762b6e),
	.w7(32'hbad7dfcd),
	.w8(32'hbc0d8299),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0de4b7),
	.w1(32'hbbe3846f),
	.w2(32'hbc12d45b),
	.w3(32'hbc3bf889),
	.w4(32'hbc1eedd6),
	.w5(32'hbc1fbf13),
	.w6(32'hbc146456),
	.w7(32'hbc309c45),
	.w8(32'hbb1a6fc1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d858f),
	.w1(32'hbc3450f6),
	.w2(32'hbc417343),
	.w3(32'hbb0c7d0f),
	.w4(32'hbbdd638f),
	.w5(32'hbbf4ff44),
	.w6(32'hbc0bafbc),
	.w7(32'hbc291637),
	.w8(32'h3b6fccdc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73ca45),
	.w1(32'h3b44aa7d),
	.w2(32'h3baa0eb3),
	.w3(32'h3c0fcb25),
	.w4(32'h3c09a8f2),
	.w5(32'h3c22421f),
	.w6(32'h3bd0f774),
	.w7(32'h3b975de6),
	.w8(32'h3b846460),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12b27b),
	.w1(32'h3aa730a1),
	.w2(32'h39975d96),
	.w3(32'h3a12f346),
	.w4(32'h3a5be40a),
	.w5(32'h38ac52e9),
	.w6(32'hbade5d19),
	.w7(32'hb9f1b2cf),
	.w8(32'h3abe97f3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbca7f),
	.w1(32'hbb071b39),
	.w2(32'hbb0c8468),
	.w3(32'h39f7b17c),
	.w4(32'h3935ebdd),
	.w5(32'hbb2f4457),
	.w6(32'h3b1399b9),
	.w7(32'hb9c6c90c),
	.w8(32'hba168823),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a878991),
	.w1(32'h3a1a979a),
	.w2(32'h3a189a03),
	.w3(32'h3b1467fb),
	.w4(32'h3b22e71d),
	.w5(32'h3abdc36b),
	.w6(32'hb976c44f),
	.w7(32'h3a664074),
	.w8(32'h3ae1238b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c763a),
	.w1(32'h3b33cf34),
	.w2(32'h3b0ca24e),
	.w3(32'h3b6dbd5a),
	.w4(32'h3b9bd05d),
	.w5(32'h3b70dbb9),
	.w6(32'hbab32883),
	.w7(32'h3af58c31),
	.w8(32'h3b55f3ce),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91897a8),
	.w1(32'hb9eba357),
	.w2(32'h3a1a196a),
	.w3(32'h38776790),
	.w4(32'h3a6b348a),
	.w5(32'h3a77da50),
	.w6(32'hbb1901fd),
	.w7(32'hbaaaade1),
	.w8(32'hba24a28e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa70c42),
	.w1(32'hbb2e1550),
	.w2(32'hbb814a17),
	.w3(32'hbb46da43),
	.w4(32'hbb7c186d),
	.w5(32'hbb0b635f),
	.w6(32'h3a500bb4),
	.w7(32'hb976f535),
	.w8(32'hba1d5b89),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87c389),
	.w1(32'h3bc17d0e),
	.w2(32'h3ba78316),
	.w3(32'h3bd6ef84),
	.w4(32'h3c08f492),
	.w5(32'h3bca8b8c),
	.w6(32'hba5e356d),
	.w7(32'h3b3ec032),
	.w8(32'h3a3fedb1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965336b),
	.w1(32'h3ab630b2),
	.w2(32'h38a190e9),
	.w3(32'hba83545e),
	.w4(32'hb872e183),
	.w5(32'hba0e5687),
	.w6(32'h3a0988d9),
	.w7(32'hb94e62fb),
	.w8(32'h3a730ef9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94b94c),
	.w1(32'h389257a9),
	.w2(32'h3a43268b),
	.w3(32'h3b92a0a3),
	.w4(32'h3b304451),
	.w5(32'h3ac3d444),
	.w6(32'h3aabed0d),
	.w7(32'h3abacca6),
	.w8(32'h3a0c17ad),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fd3a6),
	.w1(32'hbad46917),
	.w2(32'h3a3cd6b1),
	.w3(32'hba3c93cb),
	.w4(32'hbb134f5e),
	.w5(32'h3a929adc),
	.w6(32'hbb19fb17),
	.w7(32'hbb83ba79),
	.w8(32'hbb1af275),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad42cec),
	.w1(32'h3b705d4b),
	.w2(32'h3ba23391),
	.w3(32'h3c0ad337),
	.w4(32'h3c3d4cd9),
	.w5(32'h3c25c8f2),
	.w6(32'h3b97ee8f),
	.w7(32'h3c2ba312),
	.w8(32'h3c593e0c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989c69),
	.w1(32'h38be8c25),
	.w2(32'hbbcd4bd9),
	.w3(32'hba0d8350),
	.w4(32'h3b3137c7),
	.w5(32'hba17625a),
	.w6(32'h3c0a1797),
	.w7(32'h3acf7218),
	.w8(32'h3b01ea26),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96d31d),
	.w1(32'h3bcbee04),
	.w2(32'h3bbc8f7b),
	.w3(32'h3b417bee),
	.w4(32'h3b2cd0d7),
	.w5(32'h3b50ab7b),
	.w6(32'h3b291949),
	.w7(32'h3abf9d1a),
	.w8(32'h3ad12cb6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b233113),
	.w1(32'hbb8636cd),
	.w2(32'hbb89d328),
	.w3(32'h3a6863e9),
	.w4(32'hbad0f1d5),
	.w5(32'hbb1d14bc),
	.w6(32'h395029ef),
	.w7(32'hbb13291e),
	.w8(32'h39fb86eb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c308219),
	.w1(32'h3c26eac3),
	.w2(32'h3c1b006e),
	.w3(32'h3c200048),
	.w4(32'h3c68c9f8),
	.w5(32'h3c42112b),
	.w6(32'hb9e1b94a),
	.w7(32'hb9dee8a3),
	.w8(32'hbb858027),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c6f4e),
	.w1(32'hbb8eb18d),
	.w2(32'hb88fa7a2),
	.w3(32'hb9a45fbe),
	.w4(32'hbb17c549),
	.w5(32'hba042b56),
	.w6(32'hb9e6359c),
	.w7(32'hba80522c),
	.w8(32'h3a8f7dbe),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaea926),
	.w1(32'hbb94ef12),
	.w2(32'hbb9f70a2),
	.w3(32'h3bb32cb0),
	.w4(32'h3b7512c8),
	.w5(32'hba447592),
	.w6(32'h3b21f638),
	.w7(32'h3b12770d),
	.w8(32'h3a75f3a5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a650bf9),
	.w1(32'h3ae23c08),
	.w2(32'h3af1002e),
	.w3(32'h3aa72d71),
	.w4(32'h3b273861),
	.w5(32'h3b0cbb0e),
	.w6(32'h3a84fb3a),
	.w7(32'h3b225a0a),
	.w8(32'hba7c2325),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b817c),
	.w1(32'hbb644de2),
	.w2(32'hbb690c60),
	.w3(32'hbb30843d),
	.w4(32'hbb3cf456),
	.w5(32'hbb55c329),
	.w6(32'h3abb599d),
	.w7(32'hbabd7105),
	.w8(32'hbb1f420f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a01e1),
	.w1(32'hb9f0fdc4),
	.w2(32'hba01fbbc),
	.w3(32'h3ba4aa12),
	.w4(32'h3b6dd8e1),
	.w5(32'hbad3880d),
	.w6(32'h3ae8770c),
	.w7(32'h3b0382ba),
	.w8(32'h3ada48f6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9136d8),
	.w1(32'h3a863298),
	.w2(32'h3af1fccb),
	.w3(32'h3acf5692),
	.w4(32'h3b078eae),
	.w5(32'h3ae93d2d),
	.w6(32'hb985e765),
	.w7(32'h3a9e881c),
	.w8(32'hb9fcbe92),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952551e),
	.w1(32'hbaa9f617),
	.w2(32'hba385c60),
	.w3(32'h3b8d27ca),
	.w4(32'h3b8671bc),
	.w5(32'h3b6dc3c2),
	.w6(32'hbae3d2a3),
	.w7(32'hba83c6d8),
	.w8(32'hb84876a0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf73337),
	.w1(32'hbb445c0e),
	.w2(32'hbbd022e7),
	.w3(32'hbb3901d7),
	.w4(32'hba9e1421),
	.w5(32'hbb78cd4b),
	.w6(32'hbaa330e1),
	.w7(32'hbaa5173a),
	.w8(32'h3a2ffd62),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc7be7),
	.w1(32'hbaf15b92),
	.w2(32'hbaccd8f9),
	.w3(32'hba39935e),
	.w4(32'hba600a67),
	.w5(32'hba95b9b5),
	.w6(32'hbac598b7),
	.w7(32'hb9d28b83),
	.w8(32'hbaabf103),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff7c1e),
	.w1(32'h3aed7219),
	.w2(32'h3a14b0b0),
	.w3(32'h3b2cbaa5),
	.w4(32'h3b78c701),
	.w5(32'h3b1a9075),
	.w6(32'h3a95efaf),
	.w7(32'h3b14e23f),
	.w8(32'h3a944731),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83acd9),
	.w1(32'h3b271a6b),
	.w2(32'h3b498243),
	.w3(32'h3ba0fd37),
	.w4(32'h3b845953),
	.w5(32'h3b8e2baa),
	.w6(32'h3b7fa594),
	.w7(32'h3b66742b),
	.w8(32'h3ba1bed8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd8151),
	.w1(32'h3b09d0ca),
	.w2(32'h3ac181e7),
	.w3(32'h3677dd0a),
	.w4(32'h3b28e522),
	.w5(32'h3b4d8c0f),
	.w6(32'h3a5d8bf9),
	.w7(32'h3a8cc672),
	.w8(32'h39cdbf9c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e91f3),
	.w1(32'h39e5127f),
	.w2(32'h3a244490),
	.w3(32'h3b014b0e),
	.w4(32'h3a776940),
	.w5(32'hba0a88f7),
	.w6(32'h3a874de5),
	.w7(32'h39ddae84),
	.w8(32'hbb2236fd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33133b),
	.w1(32'hb84722ad),
	.w2(32'h3ab47446),
	.w3(32'h3b928d46),
	.w4(32'h3bcd2ae8),
	.w5(32'h3b99c667),
	.w6(32'h3a6ffa08),
	.w7(32'h3b87f7ad),
	.w8(32'h3b4cb136),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba339ab9),
	.w1(32'hbad4fc7d),
	.w2(32'hbaa48eb5),
	.w3(32'hbad74c83),
	.w4(32'hbb14322f),
	.w5(32'hbaffb129),
	.w6(32'hbaf79cf8),
	.w7(32'hbb05a93f),
	.w8(32'hb8b8a94c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03579f),
	.w1(32'h3a9a25ad),
	.w2(32'h3abc3ba4),
	.w3(32'h3b3532d5),
	.w4(32'h3b7c8e9e),
	.w5(32'h3b5fdb7e),
	.w6(32'h3b127170),
	.w7(32'h3b82ce8b),
	.w8(32'h3b1b89e1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c48c0),
	.w1(32'hba0bee29),
	.w2(32'hba86eaa2),
	.w3(32'h3a40450d),
	.w4(32'hba1efa03),
	.w5(32'hbac02a66),
	.w6(32'h3a6331f7),
	.w7(32'hb87d393d),
	.w8(32'h39a6015d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be76102),
	.w1(32'h3bf36171),
	.w2(32'h3c0757fe),
	.w3(32'h3bc37aaf),
	.w4(32'h3c1c5097),
	.w5(32'h3bf1bf18),
	.w6(32'h3c387b69),
	.w7(32'h3c0fe415),
	.w8(32'h3ae1a324),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb863a203),
	.w1(32'hb835f495),
	.w2(32'h3903504b),
	.w3(32'hb9a7a008),
	.w4(32'hb97a66e6),
	.w5(32'hb9e1faaa),
	.w6(32'hb740dd50),
	.w7(32'h39c28d72),
	.w8(32'hba29a616),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dbc4b),
	.w1(32'h3b3aeb37),
	.w2(32'h3b5963cb),
	.w3(32'h3b6d70b6),
	.w4(32'h3b7def3b),
	.w5(32'h3b71af62),
	.w6(32'h3aefed1d),
	.w7(32'h3b26e9f3),
	.w8(32'h3b4275e3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26e511),
	.w1(32'h3a22e936),
	.w2(32'h39e23711),
	.w3(32'h397a8f2a),
	.w4(32'h38b13ce2),
	.w5(32'hb9d8017d),
	.w6(32'h38dc3fcb),
	.w7(32'h39e9663e),
	.w8(32'h3974d850),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920ffdc),
	.w1(32'hba2f7cfb),
	.w2(32'h3a29c0c4),
	.w3(32'h3b86e017),
	.w4(32'h3bb1b696),
	.w5(32'h3ba38d30),
	.w6(32'hbb0f184e),
	.w7(32'h3a94f4dc),
	.w8(32'h3ab7c9d0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3526a9),
	.w1(32'h3b387c0d),
	.w2(32'h3ad4ff28),
	.w3(32'h3b83e332),
	.w4(32'h3b90e371),
	.w5(32'h3b764180),
	.w6(32'h3a124fea),
	.w7(32'h3a7bdd40),
	.w8(32'hba2f0dbe),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ecb95),
	.w1(32'h3b3fd6da),
	.w2(32'h3b5ab60a),
	.w3(32'h3ad82668),
	.w4(32'h3a039b70),
	.w5(32'h3a8c1c03),
	.w6(32'h3b329a18),
	.w7(32'h3b0a8972),
	.w8(32'hb8945ef8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5920ef),
	.w1(32'hba289864),
	.w2(32'hbb24a0c2),
	.w3(32'hbb308fa2),
	.w4(32'hbb1af9e7),
	.w5(32'hbaf3849e),
	.w6(32'hbb227457),
	.w7(32'hba99f43c),
	.w8(32'hba0297d7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e27c6),
	.w1(32'h3b27822e),
	.w2(32'h3b18c1d7),
	.w3(32'h3af88aed),
	.w4(32'h3a75cf86),
	.w5(32'hb8d7d129),
	.w6(32'h3b508afd),
	.w7(32'h3b94ef6d),
	.w8(32'h3baea30d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82b44e),
	.w1(32'h3b5325e1),
	.w2(32'h3b928732),
	.w3(32'h3bcbac44),
	.w4(32'h3bee6b32),
	.w5(32'h3bdaa052),
	.w6(32'h3b0a190c),
	.w7(32'h3b76477a),
	.w8(32'h3ada2f2e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3c06a),
	.w1(32'hbbcb3ed9),
	.w2(32'h3adefc76),
	.w3(32'h3adb64d5),
	.w4(32'hbbbf7517),
	.w5(32'hba5c42de),
	.w6(32'h3b339cc2),
	.w7(32'h3a2e0b63),
	.w8(32'h3b86773a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b891edb),
	.w1(32'h3b459188),
	.w2(32'h3a994d91),
	.w3(32'h3c21e0f2),
	.w4(32'h3c44a94d),
	.w5(32'h3be849cf),
	.w6(32'h3afc32e1),
	.w7(32'h3afa07a4),
	.w8(32'h391f3b5e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390469f8),
	.w1(32'hb916471e),
	.w2(32'h3a33d32f),
	.w3(32'h3b6c219d),
	.w4(32'h3b7ff868),
	.w5(32'h3a9599a0),
	.w6(32'h3b185101),
	.w7(32'h3bc8cbe5),
	.w8(32'h39a0f4f6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba910ab2),
	.w1(32'h3ad20a79),
	.w2(32'h3916daf9),
	.w3(32'hbb3b9dd2),
	.w4(32'hba52f4e9),
	.w5(32'hbab39e29),
	.w6(32'hba260149),
	.w7(32'hba78cc1d),
	.w8(32'hb9c46246),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05b1fc),
	.w1(32'hbab0d0dc),
	.w2(32'h3a380ff9),
	.w3(32'hb9df3123),
	.w4(32'hba4d9f92),
	.w5(32'h3a3486a4),
	.w6(32'hba4f6b0b),
	.w7(32'h3a54a169),
	.w8(32'hbb391fac),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b3896),
	.w1(32'hbb68ddca),
	.w2(32'hbb802b60),
	.w3(32'hbbad03d2),
	.w4(32'hbbe0af0b),
	.w5(32'hbbb35206),
	.w6(32'hbb57dc7c),
	.w7(32'hbb5a53c4),
	.w8(32'hba55dd03),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39c614),
	.w1(32'h3a1ae1d7),
	.w2(32'hb9a0609b),
	.w3(32'hbb5f8718),
	.w4(32'hba1883ff),
	.w5(32'hbaa2a005),
	.w6(32'hbae2d342),
	.w7(32'hba25ec1c),
	.w8(32'hba8ac044),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42e41a),
	.w1(32'h3b582dcc),
	.w2(32'h3b3b2596),
	.w3(32'hba814ade),
	.w4(32'h3a69c6d5),
	.w5(32'h3a91f9c1),
	.w6(32'h3a302e1e),
	.w7(32'h3a7dd73e),
	.w8(32'h3b6095a3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bd8a5),
	.w1(32'hb91508f5),
	.w2(32'h3a4dea73),
	.w3(32'hbaaac4eb),
	.w4(32'hbb1af73b),
	.w5(32'hbaa68d66),
	.w6(32'hbab4e68d),
	.w7(32'hbb028fcf),
	.w8(32'hba1e80e1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb970f32),
	.w1(32'hbc06f99d),
	.w2(32'hba0efedf),
	.w3(32'hbbb64495),
	.w4(32'hbc117d2e),
	.w5(32'hbbc5020c),
	.w6(32'h3a69a02c),
	.w7(32'hb8824981),
	.w8(32'hba524794),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b587871),
	.w1(32'h3b578990),
	.w2(32'h3b4d85a6),
	.w3(32'h3b670969),
	.w4(32'h3b57dc96),
	.w5(32'h3b62f39d),
	.w6(32'h3b8a8301),
	.w7(32'h3b9bbd92),
	.w8(32'h3ba48ddb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba915577),
	.w1(32'h3a833ba7),
	.w2(32'h38f3efff),
	.w3(32'hbb526df2),
	.w4(32'hbb2632f1),
	.w5(32'hbb01844d),
	.w6(32'h39534d8e),
	.w7(32'h399258d4),
	.w8(32'h3b625658),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12ef61),
	.w1(32'h3a3a9894),
	.w2(32'h3a2e274b),
	.w3(32'hbb0ae7a7),
	.w4(32'hbac1fe65),
	.w5(32'hb95ee81b),
	.w6(32'hbb81302c),
	.w7(32'hbb412f98),
	.w8(32'hba884c85),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4536ee),
	.w1(32'h3ae484dd),
	.w2(32'h3adf8fcd),
	.w3(32'h3bc76e2c),
	.w4(32'h3bd22afb),
	.w5(32'h3badcaea),
	.w6(32'h3a450538),
	.w7(32'h3b186fea),
	.w8(32'h3b4cd521),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c12cb),
	.w1(32'h3bcff41e),
	.w2(32'h3b4c413d),
	.w3(32'hbb1d9578),
	.w4(32'hb9c49845),
	.w5(32'hba1e5ab4),
	.w6(32'hbaa51f8a),
	.w7(32'hba55b854),
	.w8(32'h395091e8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dadf91),
	.w1(32'hba4d3d8c),
	.w2(32'h39d278e5),
	.w3(32'h3a9c04d3),
	.w4(32'h39a3e6b7),
	.w5(32'h3a592eb7),
	.w6(32'hb9f7fc48),
	.w7(32'h3a7fcb42),
	.w8(32'h3a9a4c26),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbfc60),
	.w1(32'h3a9199f2),
	.w2(32'h3adc3cec),
	.w3(32'h3a84ba5b),
	.w4(32'h3a646fcc),
	.w5(32'h3a83efec),
	.w6(32'h3a3222a6),
	.w7(32'h3ae47bdc),
	.w8(32'h39603137),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92ec1f),
	.w1(32'hbb2b935d),
	.w2(32'hbaeb853f),
	.w3(32'hbab7e696),
	.w4(32'hbb3e3705),
	.w5(32'hbb0d9e12),
	.w6(32'hba361552),
	.w7(32'hbaf124b1),
	.w8(32'hba5eea29),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbad207),
	.w1(32'h3b89c447),
	.w2(32'h3b8eea2c),
	.w3(32'h3b508314),
	.w4(32'h3b2b85cd),
	.w5(32'h3b82edd5),
	.w6(32'h3b047259),
	.w7(32'h3a842eea),
	.w8(32'h3badc5ce),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3f58),
	.w1(32'h39e8ae92),
	.w2(32'h3b800891),
	.w3(32'h3b8ac275),
	.w4(32'h3b85570c),
	.w5(32'h3ba26e1a),
	.w6(32'h3a7181d6),
	.w7(32'h3b8d756a),
	.w8(32'h3ae443a2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b5027),
	.w1(32'h3b4811d7),
	.w2(32'h3b33bcee),
	.w3(32'h3ad71bcf),
	.w4(32'h39f9874e),
	.w5(32'h39a87fd6),
	.w6(32'h3b3a0959),
	.w7(32'h3b2404f1),
	.w8(32'h3b1d585a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94eea8a),
	.w1(32'h3a1ace90),
	.w2(32'h397820c1),
	.w3(32'hba8987d1),
	.w4(32'hba396aad),
	.w5(32'hba799aab),
	.w6(32'h39a20017),
	.w7(32'hb94d2b8e),
	.w8(32'hb849610d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b681a),
	.w1(32'h3b3dead4),
	.w2(32'hba68bd20),
	.w3(32'h3c20e492),
	.w4(32'h3c32bf8d),
	.w5(32'h3b4fc9d4),
	.w6(32'h3beb6eb8),
	.w7(32'h3beaba6d),
	.w8(32'h39844aa3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b68ad),
	.w1(32'h3ad1fe50),
	.w2(32'h3b4a7983),
	.w3(32'h3aa55d35),
	.w4(32'h3aece2ba),
	.w5(32'h3b600eca),
	.w6(32'h379bdb33),
	.w7(32'h3a24307f),
	.w8(32'h3b63e424),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19f27c),
	.w1(32'h3b2e9506),
	.w2(32'h3b1dae0e),
	.w3(32'h3af645f8),
	.w4(32'h3aa2147b),
	.w5(32'h3b0dbbeb),
	.w6(32'h3ab58d93),
	.w7(32'h3ac6cddb),
	.w8(32'h3b3d4065),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b4704),
	.w1(32'hbb35cb90),
	.w2(32'hbac87fc9),
	.w3(32'hbb1f5a3a),
	.w4(32'hbb726594),
	.w5(32'hbb47e7d1),
	.w6(32'hba8fc703),
	.w7(32'hbb458985),
	.w8(32'hbb136747),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be318da),
	.w1(32'h3bb84a6f),
	.w2(32'h3bad0842),
	.w3(32'h3ba5d5a2),
	.w4(32'h3ba58288),
	.w5(32'h3ba9a9c1),
	.w6(32'h3b794bf0),
	.w7(32'h3b97d6f6),
	.w8(32'h3b87a431),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49286b),
	.w1(32'h3b2be56e),
	.w2(32'h3b4f5a15),
	.w3(32'h3aa4090c),
	.w4(32'h3a8e8a60),
	.w5(32'h3b0d6429),
	.w6(32'h3a720651),
	.w7(32'h38e37691),
	.w8(32'h3b02e51e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83910f),
	.w1(32'h3b14924a),
	.w2(32'h3b8eadd2),
	.w3(32'h3b0b119b),
	.w4(32'hb80cd49d),
	.w5(32'h3b08b7ae),
	.w6(32'h3b03f6fb),
	.w7(32'h3a677881),
	.w8(32'h3b4f96bb),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba791125),
	.w1(32'hbafb86f9),
	.w2(32'hbaf1029d),
	.w3(32'hbab2b128),
	.w4(32'hbb24fa3b),
	.w5(32'hbb3f8d20),
	.w6(32'h3a321a96),
	.w7(32'hba743721),
	.w8(32'hba6aef4f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b80d0e),
	.w1(32'hb932254e),
	.w2(32'hb9411014),
	.w3(32'h38b04550),
	.w4(32'h396fe37a),
	.w5(32'h38f1a552),
	.w6(32'hb84331c7),
	.w7(32'h39113da7),
	.w8(32'hb8cfb051),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11a590),
	.w1(32'hb7f81c78),
	.w2(32'hb954014c),
	.w3(32'h398d42af),
	.w4(32'h39e35688),
	.w5(32'h3a09ceb8),
	.w6(32'h38ee8e9b),
	.w7(32'h3a2abece),
	.w8(32'h3a3fea51),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c4f43),
	.w1(32'h3b2090ab),
	.w2(32'h3b43871d),
	.w3(32'h3b159f6e),
	.w4(32'h3b1d4ccd),
	.w5(32'h3b347bd1),
	.w6(32'h3b061022),
	.w7(32'h3b0ec2af),
	.w8(32'h3b10b2bd),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2260d),
	.w1(32'h3a74a9b1),
	.w2(32'h3aaed25a),
	.w3(32'hba009841),
	.w4(32'hbab2daa9),
	.w5(32'h395c7a6e),
	.w6(32'h39a42b3f),
	.w7(32'hba4399a1),
	.w8(32'h3a307f24),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42a003),
	.w1(32'h3993498c),
	.w2(32'h3ac34b78),
	.w3(32'h3ab912b0),
	.w4(32'h3aaf03b6),
	.w5(32'h3b0567fa),
	.w6(32'h3ab532bb),
	.w7(32'h39593d8a),
	.w8(32'h3adcaa40),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83995f9),
	.w1(32'hb76abb8c),
	.w2(32'hb7d6acf8),
	.w3(32'hb81a4a21),
	.w4(32'hb745ec5e),
	.w5(32'hb7fdb3fb),
	.w6(32'hb802577c),
	.w7(32'hb6a7a0ef),
	.w8(32'hb7ffdf3d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a6043),
	.w1(32'h38bee582),
	.w2(32'hb905d9a5),
	.w3(32'hb9214dc5),
	.w4(32'hb78741f6),
	.w5(32'hb8474c40),
	.w6(32'hb936c4a9),
	.w7(32'hb96a4f05),
	.w8(32'hb9a10eac),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec624a),
	.w1(32'h3aed7410),
	.w2(32'h3af3cae7),
	.w3(32'h3a15c52c),
	.w4(32'hb8789b41),
	.w5(32'hb9ac95f5),
	.w6(32'h3b23a016),
	.w7(32'h3b01ebfb),
	.w8(32'h3a867d80),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1e43b),
	.w1(32'h3bdef4d6),
	.w2(32'h3bd6f914),
	.w3(32'h3b7c1b55),
	.w4(32'h3bb55f9c),
	.w5(32'h3bae404b),
	.w6(32'h3a834aaf),
	.w7(32'h3b3f7c99),
	.w8(32'h3b97b8c9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef2b3a),
	.w1(32'h39a33b29),
	.w2(32'h3a3a9bbf),
	.w3(32'h3931ca2a),
	.w4(32'hb98bcb9e),
	.w5(32'hb921a497),
	.w6(32'h39349ae4),
	.w7(32'hb94feffc),
	.w8(32'hba281bed),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a554302),
	.w1(32'hb98b55ff),
	.w2(32'h3a6a60bf),
	.w3(32'hba0e4a7e),
	.w4(32'hbabd1def),
	.w5(32'hb942b266),
	.w6(32'h3a4c1680),
	.w7(32'hb8dbe153),
	.w8(32'h3a8022eb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8832e5),
	.w1(32'h3b3d53d2),
	.w2(32'h3b158857),
	.w3(32'h3b566a46),
	.w4(32'h3aabcf32),
	.w5(32'h3ae9f617),
	.w6(32'h3b02a657),
	.w7(32'h398c8932),
	.w8(32'h3ac1f707),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a199a72),
	.w1(32'h389d8d33),
	.w2(32'h3a3931ac),
	.w3(32'h39037a9b),
	.w4(32'hba2bf28f),
	.w5(32'h3a1247d4),
	.w6(32'hb9319b70),
	.w7(32'hba5d9d1c),
	.w8(32'h39abe2d2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81bbcf),
	.w1(32'h3b7bea21),
	.w2(32'h3ba6c67d),
	.w3(32'h3b157fff),
	.w4(32'h3b698703),
	.w5(32'h3ba75b46),
	.w6(32'h3aa33b80),
	.w7(32'h3b417c8d),
	.w8(32'h3b5bdb7a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6d0bc),
	.w1(32'hb82485cf),
	.w2(32'h39f1bcae),
	.w3(32'hbae1fe77),
	.w4(32'hb99c203d),
	.w5(32'h3a045210),
	.w6(32'hbb099e42),
	.w7(32'hb9a62a79),
	.w8(32'h3a06400a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule