module layer_6_featuremap_121(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61c9e5),
	.w1(32'hbace382e),
	.w2(32'h3a02bce2),
	.w3(32'h3a34382d),
	.w4(32'h3b0f0c2c),
	.w5(32'h3b7c9217),
	.w6(32'hba65a362),
	.w7(32'h3b05938f),
	.w8(32'h3b9c270b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba719f1b),
	.w1(32'hbb553700),
	.w2(32'hb9a0e1b0),
	.w3(32'hbc6a48fc),
	.w4(32'hbc363538),
	.w5(32'hbbe0047e),
	.w6(32'hbcb72b10),
	.w7(32'hbcb092fa),
	.w8(32'hbc9bf5a0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6937c),
	.w1(32'h3abacfec),
	.w2(32'h3c2cd3c1),
	.w3(32'h3c0a9cb7),
	.w4(32'h3c7fc07b),
	.w5(32'h3c5c5115),
	.w6(32'hbd01d38e),
	.w7(32'hbc2fee11),
	.w8(32'hbb9e3ebe),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e0c2d),
	.w1(32'h3bb1c3ab),
	.w2(32'hbae384e7),
	.w3(32'h3c09591f),
	.w4(32'h3b96a263),
	.w5(32'hb9b06b60),
	.w6(32'h3a3c00d9),
	.w7(32'hbc0c02d1),
	.w8(32'hbbe0dd56),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60f384),
	.w1(32'hbd114d6d),
	.w2(32'hbd732cb6),
	.w3(32'hbbef89d9),
	.w4(32'hbcc0a5aa),
	.w5(32'hbbe7599d),
	.w6(32'h3c4694d6),
	.w7(32'h3d21b78d),
	.w8(32'h3cbeb3b2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd748d3f),
	.w1(32'hbb78c356),
	.w2(32'hbb89c6c9),
	.w3(32'h3b33e35d),
	.w4(32'h3a820a39),
	.w5(32'h3b83802c),
	.w6(32'h3a8210ec),
	.w7(32'h3b0fd4af),
	.w8(32'h3b5772f3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb58275),
	.w1(32'h3b86ffe7),
	.w2(32'h3bdb17e5),
	.w3(32'h3bc6f799),
	.w4(32'h3c2b16e8),
	.w5(32'h3bbb5d07),
	.w6(32'hbb2a251d),
	.w7(32'hbba39401),
	.w8(32'hbbc47b4c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58f0bd),
	.w1(32'h3cba0ea4),
	.w2(32'h3c5c14f8),
	.w3(32'h3bf1935f),
	.w4(32'hbc23a2c7),
	.w5(32'hbc1c2e6a),
	.w6(32'hbccefbe7),
	.w7(32'h3ad55820),
	.w8(32'h3bbd2cee),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a904e3d),
	.w1(32'hbc26b708),
	.w2(32'hbd25fbad),
	.w3(32'hbd0cc72e),
	.w4(32'hbd600396),
	.w5(32'hbcd2163b),
	.w6(32'h3d8906d7),
	.w7(32'h3dba4c93),
	.w8(32'h3d605205),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfc222e),
	.w1(32'hbc075fe8),
	.w2(32'hbbec2f23),
	.w3(32'h390b9d27),
	.w4(32'h3b184e71),
	.w5(32'h3ae8248f),
	.w6(32'hbbb7be9e),
	.w7(32'hbaebb350),
	.w8(32'hbb6f9862),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb920b12),
	.w1(32'h3a895f45),
	.w2(32'h3b6465f0),
	.w3(32'h3abbcc4c),
	.w4(32'h3b23e384),
	.w5(32'hbaa36062),
	.w6(32'hbc95abb6),
	.w7(32'h3bb04b6f),
	.w8(32'h3c8159bd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85d4e6),
	.w1(32'hbbc1bdd1),
	.w2(32'hba7f02f1),
	.w3(32'hbbdd10d3),
	.w4(32'hbb891926),
	.w5(32'hbc2eb47f),
	.w6(32'h3bebf4b1),
	.w7(32'h3b3b757a),
	.w8(32'hba0c1efa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64814a),
	.w1(32'h3b270a66),
	.w2(32'h3bc4ba16),
	.w3(32'hb83a50b6),
	.w4(32'h3ba32398),
	.w5(32'h3b1ca233),
	.w6(32'hbba1b2a6),
	.w7(32'hbb2517fc),
	.w8(32'hbb5dce04),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaef78c),
	.w1(32'hbc807f68),
	.w2(32'hbc985c82),
	.w3(32'h3d1bda5a),
	.w4(32'h3d183c0e),
	.w5(32'hbba06b74),
	.w6(32'h3c1c3fc4),
	.w7(32'h3d3c9e96),
	.w8(32'h3d322ec6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf56d93),
	.w1(32'hbb76fe5f),
	.w2(32'h3ae82fb3),
	.w3(32'hbc12a0ad),
	.w4(32'hbc133359),
	.w5(32'hbb51d43c),
	.w6(32'hbb5a1c74),
	.w7(32'hbc763716),
	.w8(32'hbc572f83),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc2766),
	.w1(32'h3a360737),
	.w2(32'h39d1ed98),
	.w3(32'hbbfb6b80),
	.w4(32'hbbc83962),
	.w5(32'hbbc22383),
	.w6(32'hbbf0846e),
	.w7(32'hbb841da1),
	.w8(32'hbba51d01),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca047cc),
	.w1(32'hbcda7951),
	.w2(32'hbd0282e0),
	.w3(32'hbd2f9572),
	.w4(32'hbd3df461),
	.w5(32'hbc0c962c),
	.w6(32'hbd320b4c),
	.w7(32'hbd4f6761),
	.w8(32'hbcef6c72),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91a7f1),
	.w1(32'hbb3bbf3f),
	.w2(32'hb9906162),
	.w3(32'hbb6de9d4),
	.w4(32'hba614ad7),
	.w5(32'hb9a91a61),
	.w6(32'hbb9bf666),
	.w7(32'hbbd2d393),
	.w8(32'hbb44850a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e7d8e),
	.w1(32'hbc030be5),
	.w2(32'hbc22edc4),
	.w3(32'hbb8b2bee),
	.w4(32'hbbd2c36c),
	.w5(32'hbbccdab2),
	.w6(32'hbc4c758d),
	.w7(32'hbc5491c5),
	.w8(32'hbc2904f3),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7cba),
	.w1(32'hbbce0e42),
	.w2(32'hbba6e555),
	.w3(32'h3bd2a416),
	.w4(32'h3b622455),
	.w5(32'h3bbc01a3),
	.w6(32'hbcbbaaed),
	.w7(32'hbb87de6f),
	.w8(32'hbb585fcd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a0c69),
	.w1(32'hbadaf9e9),
	.w2(32'hba8d7ec8),
	.w3(32'hbb773c51),
	.w4(32'hbb02c4da),
	.w5(32'hbacfe920),
	.w6(32'hbb0097c8),
	.w7(32'hbbb30651),
	.w8(32'hbb454f73),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06933e),
	.w1(32'hbb7ee301),
	.w2(32'hb8efe398),
	.w3(32'hbb56a8ec),
	.w4(32'hbb2ac4cb),
	.w5(32'hba7ee450),
	.w6(32'hbb5c6925),
	.w7(32'h3a09b102),
	.w8(32'hba11e696),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b864fbf),
	.w1(32'hbc1f0e6d),
	.w2(32'h3b4a1076),
	.w3(32'h3c86fc87),
	.w4(32'h3c235cd7),
	.w5(32'hbc347858),
	.w6(32'hbb007c28),
	.w7(32'h3c1b625f),
	.w8(32'h3c815f90),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4238b7),
	.w1(32'hba2593dc),
	.w2(32'h3cad8e32),
	.w3(32'h3c99dd08),
	.w4(32'h3d00bc7b),
	.w5(32'h3d01e701),
	.w6(32'hbd61701e),
	.w7(32'hbd66f15f),
	.w8(32'hbd4b857c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c940ff9),
	.w1(32'hbb9a77ca),
	.w2(32'h3acb4571),
	.w3(32'h3aa4f999),
	.w4(32'h3ba1b351),
	.w5(32'h3c7c30e6),
	.w6(32'hbce95e6b),
	.w7(32'hbc9adf0b),
	.w8(32'hbcb19a70),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ba44e),
	.w1(32'hbc9950c3),
	.w2(32'hbcc675a4),
	.w3(32'hbc817707),
	.w4(32'hbcd9d9cc),
	.w5(32'hbc9f09b6),
	.w6(32'hbc5f3489),
	.w7(32'hbd16d74d),
	.w8(32'hbceb8ce4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ecb623),
	.w1(32'h3b9167ae),
	.w2(32'h3b6aac0d),
	.w3(32'h3c279e7e),
	.w4(32'h3c5e1fc9),
	.w5(32'h3ab6a373),
	.w6(32'h3bc0b4e6),
	.w7(32'h3b0a9bff),
	.w8(32'h3c4b40f8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc669bf),
	.w1(32'hb9d3bb9b),
	.w2(32'hbad568e6),
	.w3(32'h3b6a55eb),
	.w4(32'h3bc5dedb),
	.w5(32'h3b89b8a9),
	.w6(32'hbba30405),
	.w7(32'hbb7543a6),
	.w8(32'hbacc1c91),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba241c65),
	.w1(32'h3b2251b5),
	.w2(32'h37f8d27f),
	.w3(32'hbae88546),
	.w4(32'hbb7fe8a8),
	.w5(32'hbb72b1c8),
	.w6(32'h3b4594ae),
	.w7(32'h3b27fa3e),
	.w8(32'h3b2ef659),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03b605),
	.w1(32'h3c15f6d8),
	.w2(32'h3c73e1fa),
	.w3(32'hbc3ea94e),
	.w4(32'hbc6f426e),
	.w5(32'hbc0adf82),
	.w6(32'hbd0d22db),
	.w7(32'hbd40625b),
	.w8(32'hbcb1923c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc339f3d),
	.w1(32'h3c1b6871),
	.w2(32'h3c753b2c),
	.w3(32'h3ca96bf0),
	.w4(32'h3c401458),
	.w5(32'h3c75c539),
	.w6(32'hbd146ef2),
	.w7(32'hbd325375),
	.w8(32'hbd495d6d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24d8af),
	.w1(32'hbbafc3a9),
	.w2(32'h3c4e70ce),
	.w3(32'hbcdcb3ca),
	.w4(32'hbcdafef0),
	.w5(32'hbb538d7b),
	.w6(32'hbccf1ccb),
	.w7(32'hbce71bb9),
	.w8(32'hbc638248),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c921079),
	.w1(32'h3c3551d0),
	.w2(32'h3c80e1b9),
	.w3(32'hbc36a1f4),
	.w4(32'hbbdf9e44),
	.w5(32'h3c0a6a60),
	.w6(32'hbcae572d),
	.w7(32'hbce44911),
	.w8(32'hbcd041b5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51aad9),
	.w1(32'hbc1223c3),
	.w2(32'hbc0ff032),
	.w3(32'hbc29dd78),
	.w4(32'h3bc78b72),
	.w5(32'h3c88080d),
	.w6(32'h3c4e3caf),
	.w7(32'hbb0c0e26),
	.w8(32'hbc71f52f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb399a53),
	.w1(32'hbb860fa4),
	.w2(32'hbb5b5c06),
	.w3(32'h3a30af50),
	.w4(32'h3a9b19d7),
	.w5(32'h3bbf0f63),
	.w6(32'h3beb9360),
	.w7(32'h3be3b610),
	.w8(32'h3bf54e5c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec3fe8),
	.w1(32'hbbe6c944),
	.w2(32'hbc454454),
	.w3(32'hbbb8a6b0),
	.w4(32'hbb25f8f9),
	.w5(32'hbbd381bc),
	.w6(32'hbb085f33),
	.w7(32'h38d31722),
	.w8(32'hbb0c64c9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20939a),
	.w1(32'hbc1d10da),
	.w2(32'hbc3f5e2d),
	.w3(32'hbb5cb787),
	.w4(32'hbbecf15f),
	.w5(32'hbb072ed0),
	.w6(32'h3a9d3859),
	.w7(32'hbb709efd),
	.w8(32'hbb425280),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e7f23),
	.w1(32'hbbbbc361),
	.w2(32'hbc1ea8eb),
	.w3(32'hbb90eaac),
	.w4(32'hbb9d2179),
	.w5(32'hbbb119b1),
	.w6(32'hbc179420),
	.w7(32'hbc4d2132),
	.w8(32'hbc1d6eab),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94bc55),
	.w1(32'h3d11d065),
	.w2(32'h3cda36f8),
	.w3(32'hbc788cfc),
	.w4(32'hbc9a0c11),
	.w5(32'h3b1ea683),
	.w6(32'hbcec33e0),
	.w7(32'hbc88a745),
	.w8(32'hbcfd9b42),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc01fc),
	.w1(32'h3a0c4379),
	.w2(32'hbc93c68e),
	.w3(32'hbd233bb1),
	.w4(32'hbc29e750),
	.w5(32'h3c5f4dbb),
	.w6(32'hbbc2690e),
	.w7(32'h3aa664ed),
	.w8(32'hbc980f18),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2cf13),
	.w1(32'hbc236970),
	.w2(32'hbcf47430),
	.w3(32'hbc799791),
	.w4(32'hbc23f094),
	.w5(32'hbb33b870),
	.w6(32'hbcec1f2b),
	.w7(32'hbcd0e09a),
	.w8(32'hbb31923f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1cd641),
	.w1(32'hbb13c4d5),
	.w2(32'hbb82d3b7),
	.w3(32'hbb3cf313),
	.w4(32'hba9c51bd),
	.w5(32'hbb8de080),
	.w6(32'hbbbf1341),
	.w7(32'hbc1e76bd),
	.w8(32'hbc060043),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92b722),
	.w1(32'h3b3e687d),
	.w2(32'hb9d4c1b0),
	.w3(32'h3b890901),
	.w4(32'h3a65aeed),
	.w5(32'h3a05b1ac),
	.w6(32'hbb025deb),
	.w7(32'hbbb935ce),
	.w8(32'hbbf9bd4d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0441c3),
	.w1(32'hb93dfbaf),
	.w2(32'hbc36cb89),
	.w3(32'hbc64f276),
	.w4(32'hbca72a6a),
	.w5(32'hbcb81785),
	.w6(32'hbc1af8b5),
	.w7(32'hbc6b24a4),
	.w8(32'hbc6cbc34),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fa501),
	.w1(32'hbb93b3af),
	.w2(32'hbb812551),
	.w3(32'hbc1992f3),
	.w4(32'hbb899b6b),
	.w5(32'hbb21565c),
	.w6(32'hbb360f51),
	.w7(32'hbaf48e7f),
	.w8(32'hbb17525b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb462),
	.w1(32'hbd0ef2fa),
	.w2(32'hbd1710d9),
	.w3(32'h3a6b85a9),
	.w4(32'hbc87998a),
	.w5(32'hbc30efb3),
	.w6(32'hbc00dff8),
	.w7(32'h3c0e3166),
	.w8(32'hbc034658),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2edaf9),
	.w1(32'h3c40a5c6),
	.w2(32'h3c84011d),
	.w3(32'h3b30253b),
	.w4(32'h3c54780f),
	.w5(32'h3cb4c9b9),
	.w6(32'hbcaa8bc1),
	.w7(32'hbc92c96c),
	.w8(32'hbbdbdd83),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d3a08),
	.w1(32'hbb5a33d8),
	.w2(32'h3b2aa91b),
	.w3(32'hbc13e135),
	.w4(32'h3a25cecf),
	.w5(32'hbc1a546b),
	.w6(32'hba9b34e6),
	.w7(32'hbc601c5d),
	.w8(32'hbbcaf21d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a706a0f),
	.w1(32'h3b7eae1a),
	.w2(32'h3b62ea04),
	.w3(32'hba93b058),
	.w4(32'h377e1720),
	.w5(32'h3aad2f6f),
	.w6(32'h3a03a1c6),
	.w7(32'h3ad70bc9),
	.w8(32'h3aaf3245),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc202133),
	.w1(32'hbc7cddad),
	.w2(32'hb8d7644d),
	.w3(32'h3c8e8dcb),
	.w4(32'h3d0afacf),
	.w5(32'h3cdf8082),
	.w6(32'hbdaf8eae),
	.w7(32'hbe141a6e),
	.w8(32'hbdc4b438),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a6cd3),
	.w1(32'h3b14f985),
	.w2(32'hbac737aa),
	.w3(32'hbb1ee3a7),
	.w4(32'hbaefe7f0),
	.w5(32'hbc1c319d),
	.w6(32'hbbaf9fec),
	.w7(32'hbc469e01),
	.w8(32'hbc519816),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d276),
	.w1(32'hbbc6f593),
	.w2(32'hbae2ba1e),
	.w3(32'hbc120850),
	.w4(32'hbb7ce2f6),
	.w5(32'h3a321cdd),
	.w6(32'hbc8daef1),
	.w7(32'hbc0ca86a),
	.w8(32'hbb773a08),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ee375),
	.w1(32'hbc5f6ac1),
	.w2(32'hbccbad5b),
	.w3(32'hbcd6b7c0),
	.w4(32'hbce1ffeb),
	.w5(32'hbcb6deeb),
	.w6(32'hbd0b6ba4),
	.w7(32'hbd049c20),
	.w8(32'hbced7490),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ad525),
	.w1(32'h3a855cae),
	.w2(32'h3a11f1f9),
	.w3(32'hbc08897d),
	.w4(32'hbbe1eb96),
	.w5(32'hbbb1a0be),
	.w6(32'hbc01e729),
	.w7(32'hbc2550b0),
	.w8(32'hbc299223),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce8526),
	.w1(32'h3be2c104),
	.w2(32'h3c00e69f),
	.w3(32'hbb70095e),
	.w4(32'hbadfdc90),
	.w5(32'hbba05580),
	.w6(32'hbb44b679),
	.w7(32'hbbde001e),
	.w8(32'hbbdef2be),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38be3f),
	.w1(32'h3a6b06a0),
	.w2(32'hbae7aaec),
	.w3(32'hbb946ba4),
	.w4(32'h3b48d8e1),
	.w5(32'hbbe4b1fa),
	.w6(32'hbc83abd2),
	.w7(32'hbcebc23d),
	.w8(32'hbb9cb3ef),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55fb02),
	.w1(32'hbb8aa9ad),
	.w2(32'hbbaff065),
	.w3(32'hbbc7bee7),
	.w4(32'hbab0045a),
	.w5(32'hbbd2847b),
	.w6(32'hbb1da613),
	.w7(32'hba210641),
	.w8(32'hbab1562d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d5946),
	.w1(32'hbc49a9d7),
	.w2(32'hbbae3115),
	.w3(32'hbc4bece2),
	.w4(32'hba6b69e7),
	.w5(32'hbc6a3471),
	.w6(32'h3b5c338e),
	.w7(32'hbcccedb0),
	.w8(32'hbbcbaa4e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2d725),
	.w1(32'h3b100b89),
	.w2(32'hba9d6181),
	.w3(32'hbb248051),
	.w4(32'h3b07d45a),
	.w5(32'h3a39ec4b),
	.w6(32'hba383060),
	.w7(32'h3957ceff),
	.w8(32'hbb01e8ff),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32baee),
	.w1(32'hbb24fcfc),
	.w2(32'hbba3562a),
	.w3(32'hbba60752),
	.w4(32'hbc3e65da),
	.w5(32'hbc0c5c8c),
	.w6(32'hbc5df9e4),
	.w7(32'hbc97d856),
	.w8(32'hbc83887b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3937899b),
	.w1(32'hbc35a9c5),
	.w2(32'hbb3b07e1),
	.w3(32'hbc0f31cb),
	.w4(32'hbb8edd78),
	.w5(32'hbc0184ce),
	.w6(32'hbb8c05ff),
	.w7(32'hbbe2c593),
	.w8(32'hba9d9142),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37f6e5),
	.w1(32'h3c0b5ab0),
	.w2(32'hbcc5a2f1),
	.w3(32'hbcacc37f),
	.w4(32'hbcd223c1),
	.w5(32'hbca41775),
	.w6(32'hbc7a61ea),
	.w7(32'hbd205a2d),
	.w8(32'hbcc5e014),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c049144),
	.w1(32'h3b6be702),
	.w2(32'h3b629274),
	.w3(32'h3c8ed662),
	.w4(32'h3d6099cd),
	.w5(32'h3ccba7dc),
	.w6(32'h3d358735),
	.w7(32'hbd564c9b),
	.w8(32'hbd35ecd3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf4db0),
	.w1(32'hbb4269d5),
	.w2(32'h3b0a067d),
	.w3(32'hbb83d2b5),
	.w4(32'h3a7f9984),
	.w5(32'h3ae80810),
	.w6(32'hbbaa2ff9),
	.w7(32'h3adb8ddc),
	.w8(32'h3a9615c7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule