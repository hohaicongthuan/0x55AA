module layer_10_featuremap_246(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16f0c5),
	.w1(32'hba095afb),
	.w2(32'h38a916a4),
	.w3(32'h3860ad90),
	.w4(32'h3a826585),
	.w5(32'h3a346496),
	.w6(32'hb89fa8db),
	.w7(32'h3a5e692e),
	.w8(32'h3a940f8d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ea7a9),
	.w1(32'h3af150da),
	.w2(32'hba4ae041),
	.w3(32'h3a95740c),
	.w4(32'h3b307502),
	.w5(32'hb9f3eaa3),
	.w6(32'h3aa4b788),
	.w7(32'h3b170439),
	.w8(32'hbb19e266),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a507cfd),
	.w1(32'h39d8acf2),
	.w2(32'h39a28791),
	.w3(32'hba7ed574),
	.w4(32'hb9942dea),
	.w5(32'h397eb11f),
	.w6(32'hb98a717e),
	.w7(32'hb8d2d899),
	.w8(32'h39459f0b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7319c5),
	.w1(32'h3ab2d028),
	.w2(32'h3a02165b),
	.w3(32'h38ece3b2),
	.w4(32'hb990c3e9),
	.w5(32'h39212496),
	.w6(32'h3a69b830),
	.w7(32'h39c0a8e3),
	.w8(32'h39398294),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d96e95),
	.w1(32'hb9c432ae),
	.w2(32'h39c13900),
	.w3(32'hba71d273),
	.w4(32'hba51aa6c),
	.w5(32'hb912d327),
	.w6(32'hba0b0b39),
	.w7(32'h39751f16),
	.w8(32'hb9af150d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967187c),
	.w1(32'hb9fe44ed),
	.w2(32'hb89ecbe9),
	.w3(32'h3809f220),
	.w4(32'h38919b50),
	.w5(32'h3a81ce94),
	.w6(32'h38982357),
	.w7(32'h38d83875),
	.w8(32'h39ff018a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1ee11),
	.w1(32'hba8629d9),
	.w2(32'hbb8640f1),
	.w3(32'h38c9a8e7),
	.w4(32'hbb4b7e01),
	.w5(32'hbb91622f),
	.w6(32'h3a9169a7),
	.w7(32'hbb0f6d2e),
	.w8(32'hbb5e9215),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb415600),
	.w1(32'hba898df4),
	.w2(32'hbb2d4bb8),
	.w3(32'hbc042121),
	.w4(32'hbb44dcd0),
	.w5(32'hbacd0e7d),
	.w6(32'hbbe188e5),
	.w7(32'hbb8ca3a6),
	.w8(32'hbbb8b496),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64157d),
	.w1(32'hb9ca23da),
	.w2(32'hba8fb499),
	.w3(32'hbace6cf6),
	.w4(32'hba404b99),
	.w5(32'hbae34bea),
	.w6(32'hbad39c6e),
	.w7(32'hbaf4872c),
	.w8(32'hbb0c230a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ad253),
	.w1(32'hbbc1b29d),
	.w2(32'hbc514f5d),
	.w3(32'hbbb4d3a3),
	.w4(32'hbaefd0c4),
	.w5(32'hbbf46b8f),
	.w6(32'hbbb17a49),
	.w7(32'hbac18360),
	.w8(32'hbbecc21a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9871e94),
	.w1(32'hb8806251),
	.w2(32'hba473163),
	.w3(32'h39c52898),
	.w4(32'h39afaf67),
	.w5(32'hb9d7a755),
	.w6(32'h3a3cf647),
	.w7(32'h3a086ddb),
	.w8(32'h3a5ea7e3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3f127),
	.w1(32'h3ba7a6c5),
	.w2(32'hbab25ad4),
	.w3(32'hba54e53f),
	.w4(32'h3ab67982),
	.w5(32'hbbacccb0),
	.w6(32'hbad1a448),
	.w7(32'h3af2ba06),
	.w8(32'hbbf14696),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4da4d),
	.w1(32'hbbc09a56),
	.w2(32'hbc26f661),
	.w3(32'hbb8b6339),
	.w4(32'hbab18676),
	.w5(32'hbbc46873),
	.w6(32'hbb9e9011),
	.w7(32'hbafc396d),
	.w8(32'hbbc1387a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7269b),
	.w1(32'h394fef70),
	.w2(32'hba90b1c8),
	.w3(32'h39c73c96),
	.w4(32'h3acc0eb0),
	.w5(32'hb913b2e4),
	.w6(32'h3aa48690),
	.w7(32'h3b11dd73),
	.w8(32'hbaa354e4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8ffe3),
	.w1(32'h3881fc0a),
	.w2(32'hbb7cf886),
	.w3(32'h38fb3003),
	.w4(32'h3b23fef0),
	.w5(32'hbb055302),
	.w6(32'hbadaaa8d),
	.w7(32'h3aa511e6),
	.w8(32'hbb37af3d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe09b67),
	.w1(32'hbba27695),
	.w2(32'hbc0df9fb),
	.w3(32'hbb790ff0),
	.w4(32'h3aa333ce),
	.w5(32'hbb687846),
	.w6(32'hbbc2d6d3),
	.w7(32'hbac3dc4d),
	.w8(32'hbbcffbd3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9930929),
	.w1(32'hb8e75d48),
	.w2(32'h3a115434),
	.w3(32'hba397be2),
	.w4(32'h398c96b1),
	.w5(32'h39ff925e),
	.w6(32'hba891517),
	.w7(32'h3a26c0b8),
	.w8(32'h39d210c2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96d1b6),
	.w1(32'hbb807817),
	.w2(32'hbc12ff21),
	.w3(32'hbbaff9c8),
	.w4(32'hbb24f54f),
	.w5(32'hbbb29ea7),
	.w6(32'hbbb15910),
	.w7(32'hbb4458f1),
	.w8(32'hbbc58b0b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbbb8b),
	.w1(32'hbad48be8),
	.w2(32'hbb9d1032),
	.w3(32'hbaedf3d1),
	.w4(32'hba89dbf8),
	.w5(32'hbb85bc3b),
	.w6(32'hbaf29301),
	.w7(32'hba81b03c),
	.w8(32'hbba91be6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba123b21),
	.w1(32'hba28c8de),
	.w2(32'h3a3abf77),
	.w3(32'h3a636723),
	.w4(32'h39b7102b),
	.w5(32'hba6b4688),
	.w6(32'hba36d40c),
	.w7(32'h3a0471bc),
	.w8(32'hb9a97203),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9946b45),
	.w1(32'hb9afb3fd),
	.w2(32'h3779aed7),
	.w3(32'hba13693b),
	.w4(32'hb9f3544c),
	.w5(32'h3a8c8322),
	.w6(32'h3906c461),
	.w7(32'h3a4f0eea),
	.w8(32'h3a6dae83),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d85fe),
	.w1(32'h3b28dcb9),
	.w2(32'hba00c858),
	.w3(32'h3b020583),
	.w4(32'h3b29de1f),
	.w5(32'h395beaf5),
	.w6(32'h3a39f0d7),
	.w7(32'h3acfbcfb),
	.w8(32'hb984418d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf1970),
	.w1(32'hbb065595),
	.w2(32'hbc13b0a7),
	.w3(32'hbb79c07e),
	.w4(32'h3acb3517),
	.w5(32'hbc274b4d),
	.w6(32'hbc2037cc),
	.w7(32'hbbc379e9),
	.w8(32'hbca367df),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7ecaa),
	.w1(32'hbb51e5c2),
	.w2(32'hbc4c18ed),
	.w3(32'hbb0748b3),
	.w4(32'h3aaf94ae),
	.w5(32'hbbbd16f5),
	.w6(32'hbb1b0e3c),
	.w7(32'hb9886fbd),
	.w8(32'hbbe4d3a4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b1dd2),
	.w1(32'h3ab3b620),
	.w2(32'hbbeaf9ea),
	.w3(32'hbad06957),
	.w4(32'h3b9ff265),
	.w5(32'hbbb0dc87),
	.w6(32'hbc009acb),
	.w7(32'h3a985233),
	.w8(32'hbc0b7a6b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05f319),
	.w1(32'hba80203c),
	.w2(32'h394403b7),
	.w3(32'hba9336f7),
	.w4(32'hba89599d),
	.w5(32'hb9f714f2),
	.w6(32'hba381c29),
	.w7(32'hba004ca9),
	.w8(32'hba571b52),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0952cc),
	.w1(32'h3948a98d),
	.w2(32'h3a528b73),
	.w3(32'hb9aee506),
	.w4(32'h38d8e405),
	.w5(32'hba5faa29),
	.w6(32'h3811c71d),
	.w7(32'h390913f8),
	.w8(32'hba53b61b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2364f4),
	.w1(32'h3a90480d),
	.w2(32'hbaac39cc),
	.w3(32'hbb073188),
	.w4(32'h3b34f963),
	.w5(32'h3a78ea97),
	.w6(32'hbacd81de),
	.w7(32'h3b58ed49),
	.w8(32'h3b23a6b9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a9fb91),
	.w1(32'h3b6c082b),
	.w2(32'h3b0185cc),
	.w3(32'h39a25e44),
	.w4(32'h3b734f6d),
	.w5(32'h38c80fd4),
	.w6(32'hb925b716),
	.w7(32'h3b89680a),
	.w8(32'h3a265cb5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce9550),
	.w1(32'hbad80ea7),
	.w2(32'hbbaa72b4),
	.w3(32'hbbc3b817),
	.w4(32'hb9cc48e6),
	.w5(32'hbb5d8509),
	.w6(32'hbbab95cd),
	.w7(32'h387b972e),
	.w8(32'hbb0b2ba1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff18d9),
	.w1(32'hb907eda9),
	.w2(32'h3a73aa00),
	.w3(32'h3a0114d2),
	.w4(32'h39db81e4),
	.w5(32'h3a15b7cc),
	.w6(32'hba1227f3),
	.w7(32'hb9ab5a89),
	.w8(32'hb8d9eec7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f61ed),
	.w1(32'h3a3350d2),
	.w2(32'h3a6a0641),
	.w3(32'hba7bcf4e),
	.w4(32'hba64d684),
	.w5(32'h3b0feb5a),
	.w6(32'hbabdefa6),
	.w7(32'h39a029ba),
	.w8(32'h3ab2f19c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb098a4a),
	.w1(32'hbab41dd0),
	.w2(32'hbb92bfbf),
	.w3(32'h398ed8d9),
	.w4(32'h3a047aeb),
	.w5(32'hbb810849),
	.w6(32'hbaba9670),
	.w7(32'hba6087b1),
	.w8(32'hbb495358),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86fa9f),
	.w1(32'hba931f56),
	.w2(32'hbb4b8d46),
	.w3(32'hbb19fb73),
	.w4(32'hba676a2a),
	.w5(32'hbada4db0),
	.w6(32'hbb6641e9),
	.w7(32'hbb0cdb71),
	.w8(32'hbb03714d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0a1bc),
	.w1(32'h3a14f8e3),
	.w2(32'h3a805149),
	.w3(32'hbb0d38ca),
	.w4(32'hba9230f4),
	.w5(32'hb9e8107e),
	.w6(32'hbad2dd06),
	.w7(32'hb98fe98e),
	.w8(32'hb9b176ad),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba395c60),
	.w1(32'hb9fe18d9),
	.w2(32'hbb2a1b00),
	.w3(32'hba6961fc),
	.w4(32'hbab5ff34),
	.w5(32'hba698eba),
	.w6(32'hb9a45d12),
	.w7(32'hba825881),
	.w8(32'hbad01d5d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9478a2),
	.w1(32'hbb532d63),
	.w2(32'hbc131651),
	.w3(32'h3a1e6286),
	.w4(32'h3a94baa3),
	.w5(32'hbba5747b),
	.w6(32'hbab9c4eb),
	.w7(32'h3b08fb08),
	.w8(32'hbc0e0bec),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46d595),
	.w1(32'h3c047402),
	.w2(32'h3a283ce2),
	.w3(32'h3944901d),
	.w4(32'h3c41d2c5),
	.w5(32'h3b228087),
	.w6(32'hbb740ca3),
	.w7(32'h3bafdee5),
	.w8(32'hbba2e3e7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba313bcc),
	.w1(32'h3c4f55e5),
	.w2(32'h3a8f42d5),
	.w3(32'hbb5f1082),
	.w4(32'h3c09c108),
	.w5(32'hbb74c33f),
	.w6(32'hbbf913e3),
	.w7(32'h3b1cf574),
	.w8(32'hbc1c5a77),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b5046),
	.w1(32'h3aabaeb1),
	.w2(32'hbb11c220),
	.w3(32'h3adb09b9),
	.w4(32'h3b118e40),
	.w5(32'h3a2365b0),
	.w6(32'h3a497091),
	.w7(32'h3a407004),
	.w8(32'hba6141a5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38217d25),
	.w1(32'h3903c40c),
	.w2(32'h38cfece8),
	.w3(32'hb9b8d5bb),
	.w4(32'h3a0dccc3),
	.w5(32'hba692790),
	.w6(32'hb7d83622),
	.w7(32'h39b32ce8),
	.w8(32'hba8b10d1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6ca8d),
	.w1(32'h3900f305),
	.w2(32'h389edb94),
	.w3(32'hb97d4747),
	.w4(32'hba063cf6),
	.w5(32'h3985b62e),
	.w6(32'h399e0d33),
	.w7(32'hba11b788),
	.w8(32'h39aa69db),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e5f49),
	.w1(32'hb913daa3),
	.w2(32'h3a5df6b3),
	.w3(32'hbb8ebaee),
	.w4(32'hba0c393a),
	.w5(32'hb9958d88),
	.w6(32'hbadeefa0),
	.w7(32'hb8d02bb8),
	.w8(32'hb9d8c498),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07ff56),
	.w1(32'hbb9ebeb1),
	.w2(32'hbc188958),
	.w3(32'hbc0ae0e1),
	.w4(32'hba9c7e7e),
	.w5(32'hbbe7f63c),
	.w6(32'hbc1b9873),
	.w7(32'hbb50c8c1),
	.w8(32'hbc1ea3b4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e03ee),
	.w1(32'hbb6648da),
	.w2(32'hbc2ef5c2),
	.w3(32'hbb9a8535),
	.w4(32'h3a90ea7c),
	.w5(32'hbbe2a933),
	.w6(32'hbbdb6a8a),
	.w7(32'hba6ec502),
	.w8(32'hbc038843),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13eb7e),
	.w1(32'hbb8ad138),
	.w2(32'hbc547c69),
	.w3(32'hbb943192),
	.w4(32'h3a63295c),
	.w5(32'hbbf746ad),
	.w6(32'hbc0a66d7),
	.w7(32'hbb12fe4d),
	.w8(32'hbc1471da),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe6f33),
	.w1(32'hbafedb0f),
	.w2(32'hbbd1416a),
	.w3(32'hbbd5d2ce),
	.w4(32'hba28ac74),
	.w5(32'hbb9ba6c2),
	.w6(32'hbbd9c480),
	.w7(32'hbb34c7a9),
	.w8(32'hbbfe74d1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f11679),
	.w1(32'hbb7841fb),
	.w2(32'hbbfaf6a1),
	.w3(32'hbb8d3cea),
	.w4(32'hbb928dd9),
	.w5(32'hbc08dae3),
	.w6(32'hbbb3c8c4),
	.w7(32'hbbb0a0eb),
	.w8(32'hbc1d3911),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb4bb6),
	.w1(32'hb985ec85),
	.w2(32'hbab27784),
	.w3(32'h399ce38e),
	.w4(32'hb9a066cb),
	.w5(32'h39e8f2d8),
	.w6(32'h3a0c0b9d),
	.w7(32'hba4937ce),
	.w8(32'hb912f0a9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae2842),
	.w1(32'h3ab507f9),
	.w2(32'h39bbbdda),
	.w3(32'h3a24428e),
	.w4(32'hb951b3be),
	.w5(32'hba12b4ca),
	.w6(32'hb8e0db2b),
	.w7(32'hbae33a5c),
	.w8(32'hbb11e0e0),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a681f06),
	.w1(32'hb8e3395a),
	.w2(32'hb801cfe6),
	.w3(32'h3afbdc5c),
	.w4(32'h3a941baf),
	.w5(32'hba47a052),
	.w6(32'h3ab55267),
	.w7(32'h3a25b5fc),
	.w8(32'hba18a467),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926567),
	.w1(32'hbb33ed44),
	.w2(32'hbb8ed460),
	.w3(32'hbaaf4255),
	.w4(32'h3a638d70),
	.w5(32'hbb09cdb2),
	.w6(32'hba90f1cc),
	.w7(32'hb886ad22),
	.w8(32'hbaf20707),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43b0ea),
	.w1(32'h3acb09bc),
	.w2(32'hba65154a),
	.w3(32'h3a37064b),
	.w4(32'h3a9867e5),
	.w5(32'hbb05890a),
	.w6(32'h3a603ad5),
	.w7(32'h39f88bae),
	.w8(32'hbafd357b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b8907),
	.w1(32'hbb56469b),
	.w2(32'hbc3de9b7),
	.w3(32'hbb4bad19),
	.w4(32'hbb4cac38),
	.w5(32'hbbf575ee),
	.w6(32'hbb6c2921),
	.w7(32'hbad4459c),
	.w8(32'hbbcbc575),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa57187),
	.w1(32'h3a8572fa),
	.w2(32'h387024a3),
	.w3(32'h39fbcb5c),
	.w4(32'h38c4141a),
	.w5(32'hb97d9a73),
	.w6(32'hba22cc1c),
	.w7(32'hb9c2cb6e),
	.w8(32'hbab4992f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39799ef3),
	.w1(32'h3910f369),
	.w2(32'h39b288be),
	.w3(32'h39f6e934),
	.w4(32'h3985914d),
	.w5(32'hba1ee61a),
	.w6(32'hba17d046),
	.w7(32'h39aa0edf),
	.w8(32'hba0eea0b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8d365),
	.w1(32'hb9e0a43d),
	.w2(32'hb980fa54),
	.w3(32'hba198af6),
	.w4(32'hb85cf1b8),
	.w5(32'hb9c0daf0),
	.w6(32'hba566c3d),
	.w7(32'hb8b35299),
	.w8(32'hb9eb9725),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a27de),
	.w1(32'hba4c11cb),
	.w2(32'hba1a79d1),
	.w3(32'hb7935225),
	.w4(32'h38628199),
	.w5(32'h3a5bc1f7),
	.w6(32'hb8412df2),
	.w7(32'hb9bce92b),
	.w8(32'h39a6ce7e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a063f4c),
	.w1(32'h3af5be45),
	.w2(32'h3a260cf5),
	.w3(32'h39c57a72),
	.w4(32'h3a8d7054),
	.w5(32'h3aa5a251),
	.w6(32'hb98cc86b),
	.w7(32'hb975c5ba),
	.w8(32'hbad799f4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94778d),
	.w1(32'hbb18032c),
	.w2(32'hbaf2396f),
	.w3(32'hba97ba69),
	.w4(32'hbadc54ba),
	.w5(32'hba9e2d29),
	.w6(32'hbb4499e9),
	.w7(32'hbb4994e5),
	.w8(32'hba80f075),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb758ef4),
	.w1(32'hbac0c9ca),
	.w2(32'hbb85121f),
	.w3(32'hbb865a95),
	.w4(32'hba1dfa85),
	.w5(32'hbb862d5d),
	.w6(32'hbb8d6d5a),
	.w7(32'h39d74a91),
	.w8(32'hbb8924bb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749330),
	.w1(32'hbb8a5f33),
	.w2(32'hbb4330c7),
	.w3(32'hbb8faea8),
	.w4(32'hbb269a33),
	.w5(32'hbb27b98b),
	.w6(32'hbb818ca1),
	.w7(32'hbb5b8cc4),
	.w8(32'hbb2f76d2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc388f),
	.w1(32'h3a42b10a),
	.w2(32'h3a53d52f),
	.w3(32'hba2cad60),
	.w4(32'hb9e727a5),
	.w5(32'hb782e5b1),
	.w6(32'hba71ce9c),
	.w7(32'hb9c1312d),
	.w8(32'h3a1ee22e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39230946),
	.w1(32'h390fa8d0),
	.w2(32'h3a3af262),
	.w3(32'hb8f097a0),
	.w4(32'h39b3ccf0),
	.w5(32'hb9be4426),
	.w6(32'hb61d4097),
	.w7(32'h3a40e293),
	.w8(32'hba0673c7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b8a7a),
	.w1(32'hb9822c68),
	.w2(32'h39957a4f),
	.w3(32'hba128bde),
	.w4(32'hba74d297),
	.w5(32'h3a3fd515),
	.w6(32'hba5570f4),
	.w7(32'hba221774),
	.w8(32'h3a4de731),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f2f45),
	.w1(32'h3aa73621),
	.w2(32'h3a9e3566),
	.w3(32'h3a0408cd),
	.w4(32'h3a030898),
	.w5(32'h38fc3ff9),
	.w6(32'h394219ee),
	.w7(32'h3a286c1b),
	.w8(32'hb9666a2c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b83a3),
	.w1(32'hbb17be15),
	.w2(32'hbbcc4fbe),
	.w3(32'hbb722e09),
	.w4(32'hbb526790),
	.w5(32'hbb1a88da),
	.w6(32'hbb7d0400),
	.w7(32'hbb8710bd),
	.w8(32'hbb81fb28),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ee508),
	.w1(32'hba86cb80),
	.w2(32'hbc2866b2),
	.w3(32'hbb017b69),
	.w4(32'hbad79256),
	.w5(32'hbc20670c),
	.w6(32'hbb6ac4f3),
	.w7(32'hbb062ce5),
	.w8(32'hbc374c0f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a89ae),
	.w1(32'h3b3f0199),
	.w2(32'hbb9adbf4),
	.w3(32'h39aa111b),
	.w4(32'h3b96545d),
	.w5(32'hbb97680d),
	.w6(32'hbb6c87ab),
	.w7(32'h3627596c),
	.w8(32'hbbf8850a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf94c2),
	.w1(32'h3adf766b),
	.w2(32'hbc7b18f9),
	.w3(32'hbaa1739d),
	.w4(32'h3c09d7fa),
	.w5(32'hbbaa5e99),
	.w6(32'hbbeb31bb),
	.w7(32'h3b7515d5),
	.w8(32'hbc2c2772),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39819153),
	.w1(32'hba27e091),
	.w2(32'h3955929a),
	.w3(32'hb9e6afab),
	.w4(32'hb84bfe2d),
	.w5(32'h38841527),
	.w6(32'hb9f55786),
	.w7(32'hb8d6d939),
	.w8(32'hb981918b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2395b7),
	.w1(32'h3aa9636d),
	.w2(32'h39e94f35),
	.w3(32'h3a3d7216),
	.w4(32'h3959a46c),
	.w5(32'h3a6a8ae6),
	.w6(32'h3ab3e315),
	.w7(32'h3a8db810),
	.w8(32'h3a95da21),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f34133),
	.w1(32'h3a627928),
	.w2(32'h3a0dc905),
	.w3(32'hb82578fd),
	.w4(32'h395562c2),
	.w5(32'hba4bb588),
	.w6(32'h3a47f2a5),
	.w7(32'h39b45745),
	.w8(32'hb96e453f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7dcb1),
	.w1(32'hba2a5039),
	.w2(32'hba8397ba),
	.w3(32'hba0c3884),
	.w4(32'hb9608df0),
	.w5(32'hba7f57ee),
	.w6(32'hbb0c25ec),
	.w7(32'h39a2849e),
	.w8(32'hbabe7ff0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22e835),
	.w1(32'h3a005dff),
	.w2(32'h38f10ad4),
	.w3(32'h3916754b),
	.w4(32'hb84a1bd9),
	.w5(32'hba8d1385),
	.w6(32'h3a37720b),
	.w7(32'h39b3a3de),
	.w8(32'hba6084ea),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f0579),
	.w1(32'hbabb157e),
	.w2(32'hbb425443),
	.w3(32'hbb151477),
	.w4(32'hbaddb11d),
	.w5(32'hbad30120),
	.w6(32'hbb204765),
	.w7(32'hba9a9d08),
	.w8(32'hba8393b1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc066faa),
	.w1(32'hbaa2609d),
	.w2(32'hbb7aa7d3),
	.w3(32'hbbb5a21b),
	.w4(32'h3a5359e2),
	.w5(32'hbb0c32ff),
	.w6(32'hbbc5bac6),
	.w7(32'hba3c8698),
	.w8(32'hbbce2347),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0a420),
	.w1(32'hbba5b2a0),
	.w2(32'hbbfbd5bc),
	.w3(32'hbbb09566),
	.w4(32'hba9bd879),
	.w5(32'hbb883555),
	.w6(32'hbbb80457),
	.w7(32'hbb130f30),
	.w8(32'hbb918ad4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2583a4),
	.w1(32'hba915274),
	.w2(32'hbbd23df1),
	.w3(32'hba93269f),
	.w4(32'h3a7d1fd8),
	.w5(32'hbb7b7443),
	.w6(32'hbaf4bf36),
	.w7(32'hba96115e),
	.w8(32'hbba7b679),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75e6c8),
	.w1(32'hbb15b021),
	.w2(32'hbb863597),
	.w3(32'hbb2a5c97),
	.w4(32'hbb0e1e00),
	.w5(32'hbb882fce),
	.w6(32'hbac347ad),
	.w7(32'hba6ef5bd),
	.w8(32'hbb5a7999),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc08c1),
	.w1(32'hbb1bf452),
	.w2(32'hbba64e1a),
	.w3(32'hbb590a8b),
	.w4(32'hbaa73e7c),
	.w5(32'hbb22f38a),
	.w6(32'hbaeccac8),
	.w7(32'hba3dd66c),
	.w8(32'hbae44f68),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fe1fa),
	.w1(32'hbb1b0758),
	.w2(32'hbb807ec3),
	.w3(32'hbb132b5f),
	.w4(32'hbb070497),
	.w5(32'hbb3338dc),
	.w6(32'hbb3d4d48),
	.w7(32'hbb04be3d),
	.w8(32'hbb24f9ff),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978f3b0),
	.w1(32'hb9c2215d),
	.w2(32'h3912b9a8),
	.w3(32'hb7a9fe1f),
	.w4(32'hb9dee06e),
	.w5(32'h3a680520),
	.w6(32'hb905d92d),
	.w7(32'hb9af30a8),
	.w8(32'h3a3d687c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3a778),
	.w1(32'h3ab006be),
	.w2(32'h3b034ac2),
	.w3(32'h3a6f46eb),
	.w4(32'h3998e1a1),
	.w5(32'h392e2b00),
	.w6(32'h3afad9f8),
	.w7(32'h3a34da52),
	.w8(32'h38efb4bb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h320b59e4),
	.w1(32'hb927b89e),
	.w2(32'h38be24f0),
	.w3(32'hb91f8e2c),
	.w4(32'hb9854a35),
	.w5(32'hba8ebd30),
	.w6(32'hb9e140b2),
	.w7(32'hb98ce4de),
	.w8(32'hbaf979f8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b4f44),
	.w1(32'hba1537cc),
	.w2(32'h39c37c40),
	.w3(32'hbadf2a92),
	.w4(32'hb8248877),
	.w5(32'hb9e65e75),
	.w6(32'hbadc5cb7),
	.w7(32'h3a0cd0d2),
	.w8(32'h37b7fd9e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3193df),
	.w1(32'h393cbb39),
	.w2(32'hbb8321d6),
	.w3(32'hbb268d9c),
	.w4(32'h3b09b6e0),
	.w5(32'hbae9110f),
	.w6(32'hba839de1),
	.w7(32'h3adf3da0),
	.w8(32'hbb133c84),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f4d84e),
	.w1(32'h3a5b4778),
	.w2(32'h399f579b),
	.w3(32'hb852a5fc),
	.w4(32'h3a9a40ae),
	.w5(32'h39a46f2b),
	.w6(32'hbaf018ae),
	.w7(32'h39f929f9),
	.w8(32'hba063ccf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a54cc),
	.w1(32'hbad04d2e),
	.w2(32'hbba6257f),
	.w3(32'hba976e9d),
	.w4(32'h3a06aee9),
	.w5(32'hbb406a1d),
	.w6(32'hba81f290),
	.w7(32'h3a9c6e3f),
	.w8(32'hbb0a3f5e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb760d2d),
	.w1(32'hb970fdfc),
	.w2(32'hbb27fb04),
	.w3(32'hbb83fbd7),
	.w4(32'hb9e13c72),
	.w5(32'hbb6059b6),
	.w6(32'hbbddb28a),
	.w7(32'hbb76d0fd),
	.w8(32'hbbbfb0eb),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389a3654),
	.w1(32'h3b5b28c0),
	.w2(32'hba750e3b),
	.w3(32'hb9db668b),
	.w4(32'h3b57194b),
	.w5(32'hba811899),
	.w6(32'h38ee639d),
	.w7(32'h3afeff94),
	.w8(32'hbaf81a83),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3adb6f),
	.w1(32'hbaaa439f),
	.w2(32'hbba28348),
	.w3(32'hbb4122db),
	.w4(32'h3a6ea797),
	.w5(32'hbbba870c),
	.w6(32'hbb2020bd),
	.w7(32'hbb2aa5ae),
	.w8(32'hbc2f48b5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e7672),
	.w1(32'h3b58b195),
	.w2(32'hbb0715e7),
	.w3(32'h3b1d0d05),
	.w4(32'h3b7e2731),
	.w5(32'hba10f122),
	.w6(32'h3a74ce81),
	.w7(32'h3ba9f526),
	.w8(32'h3a80ff45),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf60239),
	.w1(32'hba9ec59e),
	.w2(32'hbbf24750),
	.w3(32'hba467889),
	.w4(32'h3b7c8971),
	.w5(32'hbb760201),
	.w6(32'hbb362341),
	.w7(32'hb95a1290),
	.w8(32'hbc01bf35),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42850c),
	.w1(32'h3ac55a7a),
	.w2(32'hbb73a74f),
	.w3(32'h3b094f8c),
	.w4(32'h3b8d454c),
	.w5(32'hb8d40ba4),
	.w6(32'h3b47b198),
	.w7(32'h3b66bfea),
	.w8(32'hba6b55be),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8273c9),
	.w1(32'h3b43d177),
	.w2(32'hbaecbac5),
	.w3(32'hba33647e),
	.w4(32'h3b92a610),
	.w5(32'hbb8a1e91),
	.w6(32'hbb42b8a6),
	.w7(32'h3b46e92e),
	.w8(32'hbb89b38e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37580eb3),
	.w1(32'hb9e00264),
	.w2(32'hbaf55f4d),
	.w3(32'h3938f9cf),
	.w4(32'hb878a074),
	.w5(32'h38dcd34f),
	.w6(32'hba261c7f),
	.w7(32'hbad96dd1),
	.w8(32'hba2096b0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7dcab),
	.w1(32'hba341188),
	.w2(32'hbbfa12e7),
	.w3(32'hb98c0df4),
	.w4(32'h3ad9d4dc),
	.w5(32'hbbc7d202),
	.w6(32'hbb43e2b9),
	.w7(32'hbb1eed7d),
	.w8(32'hbc1ffc1d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf8fc8),
	.w1(32'h3b1fb25c),
	.w2(32'hbb46d421),
	.w3(32'h3b0ead2a),
	.w4(32'h3b168da3),
	.w5(32'hbb870b1c),
	.w6(32'hb93174b4),
	.w7(32'hbafc247a),
	.w8(32'hbc14b3cb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4780a2),
	.w1(32'hba0682b3),
	.w2(32'hbc24de4b),
	.w3(32'hbb269122),
	.w4(32'hbb1c3147),
	.w5(32'hbc1eda13),
	.w6(32'hbbc5e176),
	.w7(32'hbb03cb57),
	.w8(32'hbc4ef95f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b045dac),
	.w1(32'h3c468348),
	.w2(32'h3b4a4b3d),
	.w3(32'h3b9925d5),
	.w4(32'h3c67bf4d),
	.w5(32'hbb7db5ec),
	.w6(32'h3a1b1db4),
	.w7(32'h3b813fc5),
	.w8(32'hbc0c2f57),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadac953),
	.w1(32'hb91978e4),
	.w2(32'hbbd78b56),
	.w3(32'hbba692a4),
	.w4(32'hbb0ed882),
	.w5(32'hbbba538b),
	.w6(32'hbad64d45),
	.w7(32'h3abbfd92),
	.w8(32'hbba4dd76),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba368103),
	.w1(32'h389048ac),
	.w2(32'hbb8a865f),
	.w3(32'h3a9ddb09),
	.w4(32'h3b3dbc0c),
	.w5(32'hbb6217c4),
	.w6(32'h3b07b36f),
	.w7(32'h3abee43f),
	.w8(32'hbb858315),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392dd0e2),
	.w1(32'hb9c25892),
	.w2(32'hba344bcb),
	.w3(32'h3a582cd9),
	.w4(32'hb96f24c9),
	.w5(32'h39d11d29),
	.w6(32'h3b0ec379),
	.w7(32'h3a8b2243),
	.w8(32'h3a01c230),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038c50),
	.w1(32'hbb3eb455),
	.w2(32'hbc2c1a36),
	.w3(32'hbabeac5c),
	.w4(32'hba6f97dc),
	.w5(32'hbc155cab),
	.w6(32'hbb4effb9),
	.w7(32'h392eec48),
	.w8(32'hbbd752be),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48a989),
	.w1(32'hbb122f8c),
	.w2(32'hbbb9442e),
	.w3(32'hb9b45a4f),
	.w4(32'hbba9aa1f),
	.w5(32'hbba96a66),
	.w6(32'h3a3a93ac),
	.w7(32'hb95aa17d),
	.w8(32'hbb96363e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba784e24),
	.w1(32'hb9ac368e),
	.w2(32'hbac41495),
	.w3(32'hbb62e5ba),
	.w4(32'hbb42369a),
	.w5(32'h39d1eef3),
	.w6(32'hbaa643b9),
	.w7(32'hba320ffe),
	.w8(32'h3aca4115),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc302b),
	.w1(32'hb99e705c),
	.w2(32'hba300d79),
	.w3(32'h39aa0694),
	.w4(32'h3aa48a17),
	.w5(32'hbb0deecb),
	.w6(32'h3aa301b1),
	.w7(32'h3a015e40),
	.w8(32'hbb38e4f6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb540580),
	.w1(32'hbb885d4c),
	.w2(32'hbbcb9269),
	.w3(32'hbba0cd17),
	.w4(32'hbb8545cf),
	.w5(32'hbb6a79c1),
	.w6(32'hbbfa56d7),
	.w7(32'hbbbbf6a9),
	.w8(32'hbbc79f3b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3abbf),
	.w1(32'hbaaee8c3),
	.w2(32'hbbe4be09),
	.w3(32'h3a08ea8f),
	.w4(32'h3b144ff6),
	.w5(32'hbb99119a),
	.w6(32'hba129438),
	.w7(32'h3b20544f),
	.w8(32'hbb5a17f8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba575308),
	.w1(32'h3adeac77),
	.w2(32'hbb99e590),
	.w3(32'hbaaecc2e),
	.w4(32'h3b141801),
	.w5(32'h39bccf7e),
	.w6(32'hbb3416f8),
	.w7(32'hbb135ddd),
	.w8(32'hbbcf3797),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57b8be),
	.w1(32'hba21e116),
	.w2(32'hbaf41a03),
	.w3(32'hbaaee7a5),
	.w4(32'h3a2a47ce),
	.w5(32'h39545591),
	.w6(32'hbb9ab8f8),
	.w7(32'hbb23079a),
	.w8(32'hbb3ad7aa),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10d096),
	.w1(32'h3acbfe36),
	.w2(32'hbb3bb286),
	.w3(32'hbae747a5),
	.w4(32'h3ad388f4),
	.w5(32'hbb0a1450),
	.w6(32'hbb8c72a6),
	.w7(32'hba04e6c2),
	.w8(32'hbb1d03cd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa692e6),
	.w1(32'h3b0b745b),
	.w2(32'hbb079480),
	.w3(32'hbb3c184c),
	.w4(32'hba3be3f6),
	.w5(32'hbb156a62),
	.w6(32'h39aa452a),
	.w7(32'hbb1b3386),
	.w8(32'hbb37d2f4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02b307),
	.w1(32'hba6ee36c),
	.w2(32'hbb526c2f),
	.w3(32'hbac39489),
	.w4(32'h38a03ac6),
	.w5(32'hbab31ceb),
	.w6(32'hbb05fda6),
	.w7(32'hbaea0326),
	.w8(32'hbb8de148),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb0949),
	.w1(32'hba19e3ad),
	.w2(32'hb97b51db),
	.w3(32'hb9599d8c),
	.w4(32'hbaabf1fb),
	.w5(32'h3a8950a6),
	.w6(32'hbaf4dd78),
	.w7(32'hba3b24d2),
	.w8(32'h3a310bd8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba869a68),
	.w1(32'hbb0d5426),
	.w2(32'hba0df23f),
	.w3(32'hb91dd0c1),
	.w4(32'hb8bdb3b7),
	.w5(32'h3a322623),
	.w6(32'hbacf6f6a),
	.w7(32'hb7431a41),
	.w8(32'hb948fc55),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac70648),
	.w1(32'h3b2d487b),
	.w2(32'h3b02eb2f),
	.w3(32'hb887ebca),
	.w4(32'hbb36e1de),
	.w5(32'h3a2b4e27),
	.w6(32'h3b5bab1e),
	.w7(32'h3a94b5c8),
	.w8(32'h39e1545f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8aab7),
	.w1(32'h39ee2a97),
	.w2(32'h39d179a7),
	.w3(32'h394c24a5),
	.w4(32'h3acab6b8),
	.w5(32'hbbaddee6),
	.w6(32'hb90a0a0c),
	.w7(32'h3aa5c380),
	.w8(32'hbb6cba95),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d6186),
	.w1(32'hbbd737a2),
	.w2(32'hbc2ac1c1),
	.w3(32'hbbcd110e),
	.w4(32'hbaebc1f5),
	.w5(32'h3be1109b),
	.w6(32'hbbc44d3e),
	.w7(32'hbacd751b),
	.w8(32'hbab4bd29),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13f27e),
	.w1(32'hbb25eacd),
	.w2(32'hbb743385),
	.w3(32'h3bd84b05),
	.w4(32'h3b9fb62e),
	.w5(32'hbb67d010),
	.w6(32'hba2f6719),
	.w7(32'h3a2fcdf8),
	.w8(32'hbb292086),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba931bee),
	.w1(32'hbb646c1e),
	.w2(32'hbb3400e5),
	.w3(32'hbb6fcc2d),
	.w4(32'hbb0b8c67),
	.w5(32'hbb979348),
	.w6(32'hbb5d90ff),
	.w7(32'hbac0ec25),
	.w8(32'hbba4b733),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d4a08),
	.w1(32'h3b45bd42),
	.w2(32'h3a952b47),
	.w3(32'hbb6d3a9f),
	.w4(32'hbaae8702),
	.w5(32'hbab7f31f),
	.w6(32'hbb9d0420),
	.w7(32'hbb1d86a0),
	.w8(32'hbbf4ebb1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4c146),
	.w1(32'hbac0505c),
	.w2(32'hb9221175),
	.w3(32'h3ac98144),
	.w4(32'h3b4a692d),
	.w5(32'h3ab5c0b7),
	.w6(32'h3b2e2003),
	.w7(32'h3b687f3f),
	.w8(32'hbb520e9a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8de874),
	.w1(32'h3b75fb3a),
	.w2(32'h3a485f89),
	.w3(32'h3b202393),
	.w4(32'h3a84a3f9),
	.w5(32'hbb24591c),
	.w6(32'hbb5a3cc8),
	.w7(32'hbb22a33f),
	.w8(32'h3b861ffc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c051b58),
	.w1(32'h3bb59024),
	.w2(32'h3b61c7cd),
	.w3(32'hba5445c9),
	.w4(32'hba8e7409),
	.w5(32'hba956c06),
	.w6(32'h3bb18322),
	.w7(32'h3b0d1951),
	.w8(32'hba1be4c8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba909a),
	.w1(32'hba68ff08),
	.w2(32'hba56786b),
	.w3(32'hbab6a028),
	.w4(32'hbb0ad8f7),
	.w5(32'h3a0d229f),
	.w6(32'h394e1756),
	.w7(32'hba22c4b2),
	.w8(32'hba33a8bb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b02e0),
	.w1(32'hbb82852f),
	.w2(32'hbb0e0da0),
	.w3(32'hba492cf6),
	.w4(32'hbb875a80),
	.w5(32'hbbc927fe),
	.w6(32'hbaa1fa08),
	.w7(32'hbaf81912),
	.w8(32'hbb67c9ec),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6575c4),
	.w1(32'hbb64c75a),
	.w2(32'hbc26734d),
	.w3(32'hbb5907f2),
	.w4(32'hbaef9f15),
	.w5(32'hbb14838d),
	.w6(32'hbb074e90),
	.w7(32'hbb0be96c),
	.w8(32'hbbdf973b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dbe72),
	.w1(32'h3ae175a5),
	.w2(32'h3b795b3e),
	.w3(32'h3b415d82),
	.w4(32'h3b01ad18),
	.w5(32'h3b048d12),
	.w6(32'h3aada0c2),
	.w7(32'h3a95d92d),
	.w8(32'hbb077e4c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cacb1),
	.w1(32'h3a711338),
	.w2(32'h3a958a32),
	.w3(32'hba5941d4),
	.w4(32'hba4c44d4),
	.w5(32'hbb57b8b2),
	.w6(32'hbb81eeab),
	.w7(32'hba9fcaf0),
	.w8(32'hbb967e9a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95192e),
	.w1(32'hbac405c8),
	.w2(32'hbb584d44),
	.w3(32'hbb527f0b),
	.w4(32'hbad838df),
	.w5(32'hbb8001fd),
	.w6(32'hbb860a68),
	.w7(32'hbad68cba),
	.w8(32'hbbc0e3b7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31879d),
	.w1(32'hbbddaecc),
	.w2(32'hbb4f4782),
	.w3(32'hbb82972f),
	.w4(32'hba4411f8),
	.w5(32'hbaa1e2ae),
	.w6(32'hbba0d7bd),
	.w7(32'h39e7ab9d),
	.w8(32'hbb49225e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bfd4c),
	.w1(32'hbb16bb08),
	.w2(32'hbbc86e32),
	.w3(32'hbaa920f2),
	.w4(32'h3a81e0f7),
	.w5(32'hbac78adc),
	.w6(32'hbb1b268a),
	.w7(32'hb96e22d7),
	.w8(32'hbb289670),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74b021),
	.w1(32'hbb6a9023),
	.w2(32'hbbfd15fa),
	.w3(32'hbb57b9d0),
	.w4(32'hbb4a88cf),
	.w5(32'hbc0666cf),
	.w6(32'hbb8710fb),
	.w7(32'hbb45cbc6),
	.w8(32'hbc061271),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec8df0),
	.w1(32'hbb84af71),
	.w2(32'hbbbfbea5),
	.w3(32'hbb81beab),
	.w4(32'hbb8d2512),
	.w5(32'hb953a0fc),
	.w6(32'hbb9920c6),
	.w7(32'hbb884af4),
	.w8(32'hbb212c2d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf30f86),
	.w1(32'hbb77432e),
	.w2(32'hbbb0089f),
	.w3(32'h3ad4416f),
	.w4(32'h3b02a3d2),
	.w5(32'hbb1d136c),
	.w6(32'h3a03f854),
	.w7(32'h3a6df496),
	.w8(32'hbb81a6c3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f560b),
	.w1(32'hbb1c1103),
	.w2(32'hbbb55478),
	.w3(32'hbae7433f),
	.w4(32'hb9b32bed),
	.w5(32'hbbadb942),
	.w6(32'hbb6318fc),
	.w7(32'hba2919b4),
	.w8(32'hbbe55d7f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba55211),
	.w1(32'hbb12915b),
	.w2(32'hbb7e4e03),
	.w3(32'hbb29e193),
	.w4(32'h3af6238f),
	.w5(32'hba02008c),
	.w6(32'hbbafa9e8),
	.w7(32'hba8e3097),
	.w8(32'hbb8edca2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51776d),
	.w1(32'hba613093),
	.w2(32'hbba85450),
	.w3(32'hbb396f32),
	.w4(32'hbadff3a7),
	.w5(32'hbba7b8fe),
	.w6(32'hbad7e0ac),
	.w7(32'hbade8464),
	.w8(32'hbba5ff20),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed2a44),
	.w1(32'hbaf22b0c),
	.w2(32'hbb50b7d4),
	.w3(32'hbb7b8942),
	.w4(32'hbab92aa3),
	.w5(32'hba8885eb),
	.w6(32'h3781b84b),
	.w7(32'hb9c23e84),
	.w8(32'h3aa1843b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb014e0c),
	.w1(32'h3b33dc81),
	.w2(32'h3ac6c7eb),
	.w3(32'hbbb53ca9),
	.w4(32'h3b301595),
	.w5(32'hbb065848),
	.w6(32'hbb23f546),
	.w7(32'h3aa3fe4b),
	.w8(32'hbb988509),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b072324),
	.w1(32'h3b64da74),
	.w2(32'hb9e954dc),
	.w3(32'h3af19e43),
	.w4(32'h3b89425c),
	.w5(32'h3a893a72),
	.w6(32'hba90b22b),
	.w7(32'hb82f763f),
	.w8(32'hba8045f6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10f0b8),
	.w1(32'h39545644),
	.w2(32'hb971c13c),
	.w3(32'hbabbbd9c),
	.w4(32'hba6590af),
	.w5(32'hba6ee3fd),
	.w6(32'h39fd1a83),
	.w7(32'hbb1229a2),
	.w8(32'hba390cd6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39509a78),
	.w1(32'h3a8d170f),
	.w2(32'hb9cb9316),
	.w3(32'hba454be9),
	.w4(32'hba463286),
	.w5(32'hbac0c146),
	.w6(32'h38fcddda),
	.w7(32'hba67b984),
	.w8(32'hbabeb53b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4de2b1),
	.w1(32'hbb92b7d0),
	.w2(32'hbb6a4c56),
	.w3(32'hbb2ebe93),
	.w4(32'hbadde371),
	.w5(32'hbb4e5913),
	.w6(32'hbad2f652),
	.w7(32'hba6f6bb5),
	.w8(32'hbab77728),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48328f),
	.w1(32'h3a16bb21),
	.w2(32'hbb874387),
	.w3(32'h38c165bf),
	.w4(32'h3b7d5c8d),
	.w5(32'hbb3f27c6),
	.w6(32'h3a7813d7),
	.w7(32'h3b418f10),
	.w8(32'hbab927e7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49d9bb),
	.w1(32'h3ae04d38),
	.w2(32'hbb351b0c),
	.w3(32'hbb90cb02),
	.w4(32'h3b4df111),
	.w5(32'hba1e38a3),
	.w6(32'hbb778f5c),
	.w7(32'h3a130711),
	.w8(32'hbb97b72b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b6d15),
	.w1(32'h397cb63f),
	.w2(32'h3a46067b),
	.w3(32'h3673e192),
	.w4(32'hbad17f87),
	.w5(32'h399205c0),
	.w6(32'hba5a9968),
	.w7(32'hbafe8a14),
	.w8(32'h3746d8f4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9f394),
	.w1(32'hbbad8c4b),
	.w2(32'hbc11b897),
	.w3(32'hbb7bed01),
	.w4(32'hbaccc3d3),
	.w5(32'hbbad4a16),
	.w6(32'hbbd4d1f5),
	.w7(32'hbb1405bb),
	.w8(32'hbba93be5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49c903),
	.w1(32'h39a0124b),
	.w2(32'hbb3a0e38),
	.w3(32'hba150bd9),
	.w4(32'hba05e63f),
	.w5(32'hbb547580),
	.w6(32'hbad96566),
	.w7(32'hba8a0a0f),
	.w8(32'hbaa5cca8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb4cf9),
	.w1(32'hbbd62897),
	.w2(32'hbc0bddc6),
	.w3(32'hbbd60e5a),
	.w4(32'hbb57ac0e),
	.w5(32'hbbcacc7e),
	.w6(32'hbb75b56b),
	.w7(32'hbbc3aacc),
	.w8(32'hbbae3e3f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac23d07),
	.w1(32'h3b880afa),
	.w2(32'hbb574d62),
	.w3(32'h39fac315),
	.w4(32'h3b251208),
	.w5(32'hbbcc957a),
	.w6(32'h3b804d17),
	.w7(32'h3bdf7d57),
	.w8(32'hbae3c67f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e576b),
	.w1(32'h3b9cfc8e),
	.w2(32'hba52217a),
	.w3(32'h3a8a67a1),
	.w4(32'h3b36621e),
	.w5(32'hbab89a14),
	.w6(32'h3b0a098f),
	.w7(32'h39aaeb31),
	.w8(32'hbb47ecb3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe7401),
	.w1(32'hba91d76f),
	.w2(32'hba9dc17c),
	.w3(32'h3b0fb8fd),
	.w4(32'h3a131523),
	.w5(32'hb91e2110),
	.w6(32'h3a32b593),
	.w7(32'hbac222a4),
	.w8(32'hbaa0313c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf22b39),
	.w1(32'hbadcd63c),
	.w2(32'hbb8f28e3),
	.w3(32'hbb7bedf6),
	.w4(32'h3a4c855e),
	.w5(32'hbb44180d),
	.w6(32'hbb96b5ee),
	.w7(32'h38c3090c),
	.w8(32'hbad62d3b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12fa52),
	.w1(32'h3bcf36a1),
	.w2(32'h3b954518),
	.w3(32'h3b5dccc7),
	.w4(32'h3c0f108f),
	.w5(32'hbb2734e1),
	.w6(32'h3c049b9f),
	.w7(32'h3c18fc69),
	.w8(32'hbbd9675d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb257c64),
	.w1(32'h3ac413c8),
	.w2(32'h3ad2737e),
	.w3(32'hbb243528),
	.w4(32'h3b8dfe0e),
	.w5(32'h3b05022a),
	.w6(32'hbb5a5496),
	.w7(32'h3b838c46),
	.w8(32'h3a0311e5),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a859909),
	.w1(32'hba52b5f0),
	.w2(32'hbb10c4c6),
	.w3(32'h38f8d681),
	.w4(32'hbb3c39a7),
	.w5(32'h3a963004),
	.w6(32'h3b53dfd9),
	.w7(32'hbacf2dc8),
	.w8(32'hbb217fc4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a91ef),
	.w1(32'hba3a2fb4),
	.w2(32'hbacd0a3e),
	.w3(32'h3b5a2c62),
	.w4(32'h3b83711b),
	.w5(32'hbad60b9f),
	.w6(32'h3b05067a),
	.w7(32'hbabe1486),
	.w8(32'hb984bfce),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fef3c),
	.w1(32'hbb628828),
	.w2(32'hbbaae8b2),
	.w3(32'hb92810b9),
	.w4(32'hba5951dd),
	.w5(32'hbbbb6f48),
	.w6(32'hbab02e4d),
	.w7(32'hbb9520ea),
	.w8(32'hbbddd99d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94326b8),
	.w1(32'hbb543d3a),
	.w2(32'hbb55933d),
	.w3(32'hba75b9f0),
	.w4(32'hbb133b16),
	.w5(32'hb9dd7f1a),
	.w6(32'hb993d314),
	.w7(32'hbb081ea5),
	.w8(32'hb930aabc),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad76539),
	.w1(32'hbacfb629),
	.w2(32'hbb406a24),
	.w3(32'hba5f0742),
	.w4(32'h3b8c63a9),
	.w5(32'hba8eeed1),
	.w6(32'hbae07d1b),
	.w7(32'h3aafbf43),
	.w8(32'h3a30adca),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22e08e),
	.w1(32'hbac8e513),
	.w2(32'hb9abbe44),
	.w3(32'h39d28abd),
	.w4(32'hba88851e),
	.w5(32'h3a74077b),
	.w6(32'h3ad9cecc),
	.w7(32'h3acc3197),
	.w8(32'hb993ca93),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caa435),
	.w1(32'h3b859ceb),
	.w2(32'hbb1bccab),
	.w3(32'h3a386de4),
	.w4(32'h3b39efad),
	.w5(32'hbae7df82),
	.w6(32'h39d4291a),
	.w7(32'h3b333937),
	.w8(32'hbb26e039),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6b98f),
	.w1(32'hbaad840e),
	.w2(32'h38abf193),
	.w3(32'hb9a53a3e),
	.w4(32'hb7a9c755),
	.w5(32'h3b4ee6fd),
	.w6(32'hbb16cdd2),
	.w7(32'hba85f27c),
	.w8(32'hb98ed2cc),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a201a),
	.w1(32'h3a025a29),
	.w2(32'hb8156de0),
	.w3(32'h3bc79298),
	.w4(32'h3b94e1d6),
	.w5(32'h39ec9c15),
	.w6(32'h3b16037f),
	.w7(32'h3b2972c4),
	.w8(32'h3ae7cce8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb474c2a),
	.w1(32'hba79e56a),
	.w2(32'hbb27753e),
	.w3(32'h3a63c0f5),
	.w4(32'h3b4158a7),
	.w5(32'hba5297b3),
	.w6(32'h3ad63323),
	.w7(32'h3aea50ee),
	.w8(32'hbb1c1fb5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0081ca),
	.w1(32'hbb8c9254),
	.w2(32'hbc2c2aad),
	.w3(32'hbbb308aa),
	.w4(32'hbb81ff09),
	.w5(32'hbc64b3ae),
	.w6(32'hbbeaa2cb),
	.w7(32'hbb40c53a),
	.w8(32'hbc238be6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1224a7),
	.w1(32'h3b626644),
	.w2(32'h3a077af9),
	.w3(32'hbae2b30b),
	.w4(32'h3a03ef61),
	.w5(32'h3a1cb022),
	.w6(32'hba8442a3),
	.w7(32'h3b19bb0d),
	.w8(32'hb92b0bc1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde0c68),
	.w1(32'hbbbfd2bd),
	.w2(32'hbc05344f),
	.w3(32'hbb759dea),
	.w4(32'h3ae02201),
	.w5(32'hbac7e63a),
	.w6(32'hbb9a56de),
	.w7(32'h396dd022),
	.w8(32'hbbdb3f4c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa337f),
	.w1(32'hbac9bd52),
	.w2(32'hba48318c),
	.w3(32'h3a3a60b4),
	.w4(32'h3aab68c3),
	.w5(32'hbb87ab9e),
	.w6(32'h3a5bdc7c),
	.w7(32'hb98a0b50),
	.w8(32'hbb015231),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec366b),
	.w1(32'hbb82e383),
	.w2(32'hbc7ee247),
	.w3(32'hbb9bc94e),
	.w4(32'hba86ebca),
	.w5(32'hbc26f7f2),
	.w6(32'hbbedad38),
	.w7(32'hbb028a8f),
	.w8(32'hbc43c88e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd05b58),
	.w1(32'h38a3cea5),
	.w2(32'hbbff65a6),
	.w3(32'hbb85ca64),
	.w4(32'hba797ec8),
	.w5(32'hbbbfc152),
	.w6(32'hbb6732a1),
	.w7(32'hbb1cd13b),
	.w8(32'hbc1971db),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfd33d),
	.w1(32'hbb95b252),
	.w2(32'hbc31896e),
	.w3(32'hbbb68769),
	.w4(32'hbb7d02f6),
	.w5(32'hbbb67eec),
	.w6(32'hbbd16ef6),
	.w7(32'hbbb9a4cb),
	.w8(32'hbbb9f868),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f49cd9),
	.w1(32'h3a8b4bf9),
	.w2(32'h3aad0dff),
	.w3(32'h3aafd783),
	.w4(32'h3b6fcd06),
	.w5(32'hb9fe7b44),
	.w6(32'hbafdbbcc),
	.w7(32'h3b13cf3b),
	.w8(32'hb99fad1f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0c072),
	.w1(32'hbb17fdf9),
	.w2(32'hbbb83357),
	.w3(32'hba903d80),
	.w4(32'hb9be6647),
	.w5(32'hbb06c8d9),
	.w6(32'hba02994f),
	.w7(32'hb993cfb1),
	.w8(32'hbadf76d4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96dba6),
	.w1(32'hbaac983f),
	.w2(32'h38494989),
	.w3(32'h38cbc57f),
	.w4(32'hb955acf3),
	.w5(32'hb454be0a),
	.w6(32'hbabb2b60),
	.w7(32'hba6eae06),
	.w8(32'hbaa22934),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30f5cf),
	.w1(32'hbb3259be),
	.w2(32'hbb64c2e0),
	.w3(32'hba3aadb4),
	.w4(32'hbb05c4d3),
	.w5(32'hba39304d),
	.w6(32'hbb5854e4),
	.w7(32'hba9de42e),
	.w8(32'hbb25a54b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d8c29),
	.w1(32'h3b421ac1),
	.w2(32'h3a8e1a03),
	.w3(32'hb9018b80),
	.w4(32'hb9802ff7),
	.w5(32'h3ad5bfc9),
	.w6(32'h382d8305),
	.w7(32'h3b1dfef5),
	.w8(32'hbb00bfdc),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a019a),
	.w1(32'hbb75332a),
	.w2(32'hbbfed2ca),
	.w3(32'hbada3c74),
	.w4(32'h3b0116d5),
	.w5(32'hbbb92331),
	.w6(32'hbbcfe821),
	.w7(32'hbb8338fe),
	.w8(32'hbbd4658f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c90cb),
	.w1(32'h3ac91a1c),
	.w2(32'hba3f25ff),
	.w3(32'hba71a0ee),
	.w4(32'h39a05b48),
	.w5(32'hba212314),
	.w6(32'h394d4901),
	.w7(32'h3a478df6),
	.w8(32'h3a0b91a9),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadc033),
	.w1(32'h3b11989c),
	.w2(32'h3a2aa3a9),
	.w3(32'h39e36494),
	.w4(32'h3ae4d5df),
	.w5(32'h3986c8bc),
	.w6(32'h3ac6cfb1),
	.w7(32'hba7717ad),
	.w8(32'h3a13815f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e2a8d),
	.w1(32'hba8a1354),
	.w2(32'h3a156e4d),
	.w3(32'hbb41a8cc),
	.w4(32'h390d9c07),
	.w5(32'h3a266d46),
	.w6(32'hb8fe173b),
	.w7(32'h3a5e709f),
	.w8(32'h3ab79d2c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986a187),
	.w1(32'hbb155de9),
	.w2(32'hbb4d027b),
	.w3(32'h3a2c52d4),
	.w4(32'h39a666f3),
	.w5(32'hb9417686),
	.w6(32'hbb0b4439),
	.w7(32'hbb2bc8d2),
	.w8(32'hbb62113a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43cec3),
	.w1(32'h3a54c680),
	.w2(32'hba7a4d9f),
	.w3(32'hba281dd3),
	.w4(32'h3a3e3c20),
	.w5(32'hba84ed27),
	.w6(32'h38bb7426),
	.w7(32'h3af54fa4),
	.w8(32'hbaa9a663),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8127c8),
	.w1(32'hba8fcf04),
	.w2(32'hba520c83),
	.w3(32'hba1de921),
	.w4(32'h39b05758),
	.w5(32'h3aaf4025),
	.w6(32'hbae13789),
	.w7(32'h3994650e),
	.w8(32'hbaf275a7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7216d0),
	.w1(32'hbc041363),
	.w2(32'hbc8f2adb),
	.w3(32'hbbadb60d),
	.w4(32'h3ab35b5a),
	.w5(32'hbc2665f2),
	.w6(32'hbb40a0d6),
	.w7(32'h3b454834),
	.w8(32'hbb920b98),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01928),
	.w1(32'h3b10717b),
	.w2(32'hbb8d09d9),
	.w3(32'h39b5e9b9),
	.w4(32'h3c127e1b),
	.w5(32'hbb994252),
	.w6(32'h3b164fa9),
	.w7(32'h3bd196a3),
	.w8(32'hbb83ba06),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3d695),
	.w1(32'h3b16c0b8),
	.w2(32'hb9e00ef9),
	.w3(32'hbb21b13d),
	.w4(32'hbb686d00),
	.w5(32'h3ae1ff29),
	.w6(32'h3b628f4c),
	.w7(32'hba383994),
	.w8(32'hbb214cd7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6d0ce),
	.w1(32'hba50db17),
	.w2(32'hb9a9e5a6),
	.w3(32'h3b9bbe07),
	.w4(32'h3be5f821),
	.w5(32'hb9685d35),
	.w6(32'h3a2228ad),
	.w7(32'hb9537467),
	.w8(32'h3a10ef88),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d845a),
	.w1(32'h39ce2068),
	.w2(32'h3a9df0e4),
	.w3(32'h3a8113ee),
	.w4(32'h3b576192),
	.w5(32'hba8c234d),
	.w6(32'h39193365),
	.w7(32'h3a8d3ecd),
	.w8(32'hbac1db97),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894686e),
	.w1(32'hba8a5c84),
	.w2(32'hba9f7dfb),
	.w3(32'h3aa03df7),
	.w4(32'h3bf4ae0c),
	.w5(32'hb9611f9b),
	.w6(32'h36f34155),
	.w7(32'hba461141),
	.w8(32'hbac0e4e7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e8c3e),
	.w1(32'h37aedf0a),
	.w2(32'hbae590a6),
	.w3(32'h3b0a885a),
	.w4(32'h3a4fea98),
	.w5(32'hbb4ae7af),
	.w6(32'h3af6e13f),
	.w7(32'hbb2a77f9),
	.w8(32'hbb524409),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34433f),
	.w1(32'h3aa51515),
	.w2(32'hbb8fca5f),
	.w3(32'hbb1d50f3),
	.w4(32'hb9dd7d9a),
	.w5(32'hbb0760bc),
	.w6(32'hba3021fb),
	.w7(32'h3784d690),
	.w8(32'hbb5da080),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe4308),
	.w1(32'hbb12ea8f),
	.w2(32'hbbec9f65),
	.w3(32'hbb97c262),
	.w4(32'h3b2fea75),
	.w5(32'hbb8a0251),
	.w6(32'hbbfff98a),
	.w7(32'h38d433da),
	.w8(32'hbb901fec),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0517da),
	.w1(32'hbaa219f4),
	.w2(32'hba5feff5),
	.w3(32'hbae844fd),
	.w4(32'hba1bec79),
	.w5(32'hbb1443ad),
	.w6(32'hbb5d9d73),
	.w7(32'hbb5feb54),
	.w8(32'hbb673a56),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c4af5),
	.w1(32'hbbfe7ac2),
	.w2(32'hbc517f8f),
	.w3(32'hbb657207),
	.w4(32'hbbc06115),
	.w5(32'hbbcc6b2e),
	.w6(32'hbbe51dd3),
	.w7(32'hbbaa5faa),
	.w8(32'hbbb56382),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcbf0f),
	.w1(32'hbb1c100c),
	.w2(32'hbb3732f5),
	.w3(32'hb81d93e1),
	.w4(32'hb8f674b1),
	.w5(32'hbb0f8a08),
	.w6(32'hba9997a6),
	.w7(32'hba452ade),
	.w8(32'hbac9629a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d5032),
	.w1(32'h3ad46254),
	.w2(32'h3a5f7ce2),
	.w3(32'h39eb1409),
	.w4(32'hbac206e6),
	.w5(32'h3a231489),
	.w6(32'h3ad3eb1b),
	.w7(32'h38a904fe),
	.w8(32'h3b5fed2c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06e208),
	.w1(32'hba182969),
	.w2(32'hb8b90dfb),
	.w3(32'h39f244a1),
	.w4(32'h3aea4118),
	.w5(32'hb90f2d92),
	.w6(32'h3bac1aa3),
	.w7(32'h3ba509d2),
	.w8(32'hba809a4d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3d3c9),
	.w1(32'hba5d7ad2),
	.w2(32'hba88fe6d),
	.w3(32'h3b80fa30),
	.w4(32'h3b47336c),
	.w5(32'h39e58d76),
	.w6(32'h3b1d7348),
	.w7(32'h3b730bb6),
	.w8(32'hb6fb3e2b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b46ff),
	.w1(32'h3ac92be4),
	.w2(32'hbacec5f9),
	.w3(32'h3a81c70f),
	.w4(32'h3afe8e57),
	.w5(32'hb9fea2b0),
	.w6(32'hbb16cf6f),
	.w7(32'hb9b15e30),
	.w8(32'hbb06d93e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacd6b3),
	.w1(32'h3b8c3fe0),
	.w2(32'hbaf272f6),
	.w3(32'h3adc5e59),
	.w4(32'h3c112fa8),
	.w5(32'hba0abeae),
	.w6(32'h3ac5aaa6),
	.w7(32'h3bdf022a),
	.w8(32'hbb1dcb20),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb961190),
	.w1(32'hbb2829b4),
	.w2(32'hbbb4ad14),
	.w3(32'hba842c58),
	.w4(32'h3b002382),
	.w5(32'hbb838970),
	.w6(32'hbb87baa0),
	.w7(32'hbb22b9d5),
	.w8(32'hbbcf98d5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b098b33),
	.w1(32'h3aa52a10),
	.w2(32'hba72cd4a),
	.w3(32'hbb615672),
	.w4(32'hbb71e495),
	.w5(32'hbab799d2),
	.w6(32'hbb1f0b83),
	.w7(32'hbb6a395f),
	.w8(32'hbaf16f24),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1f54c),
	.w1(32'hbac239ab),
	.w2(32'hbbbd43b5),
	.w3(32'hbacb99f5),
	.w4(32'h3a6fb576),
	.w5(32'hbb702435),
	.w6(32'hbae4c985),
	.w7(32'hbaaab8ae),
	.w8(32'hbbb88e85),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27bf86),
	.w1(32'hb9f0d9ae),
	.w2(32'hbb8fbf80),
	.w3(32'hbad103b9),
	.w4(32'hba4170e6),
	.w5(32'hbaaf19b9),
	.w6(32'hbb22e0ca),
	.w7(32'hba846db5),
	.w8(32'h3ad134fe),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba065a9),
	.w1(32'hbaf4e43f),
	.w2(32'hbbc7d0cf),
	.w3(32'hbc0d0b32),
	.w4(32'hb9d3a98e),
	.w5(32'hbc028414),
	.w6(32'hbbe93f44),
	.w7(32'h3b003692),
	.w8(32'hbbe92279),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3ec56),
	.w1(32'hbb1bbf72),
	.w2(32'hbb20cbf0),
	.w3(32'hba3f6011),
	.w4(32'hbb1bff9c),
	.w5(32'hb9ec2893),
	.w6(32'h3a1bc388),
	.w7(32'h3a9e2e47),
	.w8(32'hb9e35c32),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3ed90),
	.w1(32'h3ac2f28e),
	.w2(32'h3b61c552),
	.w3(32'hb98d8f13),
	.w4(32'hb9fe7d09),
	.w5(32'h39f6c5b9),
	.w6(32'hb9dba798),
	.w7(32'h39596eef),
	.w8(32'h3a0e9e90),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004916),
	.w1(32'hb771dfa9),
	.w2(32'hbb957d63),
	.w3(32'hbb739df9),
	.w4(32'h39f0750f),
	.w5(32'hbbb9db45),
	.w6(32'hbb878275),
	.w7(32'hb81f7ff9),
	.w8(32'hbc021cdb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24375a),
	.w1(32'h3b8981b2),
	.w2(32'hbb3ab7d4),
	.w3(32'hbb48c47f),
	.w4(32'hbb0fa2d8),
	.w5(32'hbc157648),
	.w6(32'hba816f6a),
	.w7(32'h3a80a4b8),
	.w8(32'hbc0da7ca),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1e67d),
	.w1(32'hb907a817),
	.w2(32'hbc0166ea),
	.w3(32'hbaf8000e),
	.w4(32'hb87157d0),
	.w5(32'hbbdda1a0),
	.w6(32'hb94344e2),
	.w7(32'hb8e7947e),
	.w8(32'hbbef8aec),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae853a6),
	.w1(32'h398dbc21),
	.w2(32'hba83dcfc),
	.w3(32'hbb9e8bf4),
	.w4(32'hbbc01473),
	.w5(32'hba810a80),
	.w6(32'hba86ef4e),
	.w7(32'hbb574083),
	.w8(32'hb9a91c3b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b076a67),
	.w1(32'h3a9fd162),
	.w2(32'h3a970539),
	.w3(32'h3a7859bd),
	.w4(32'hba1f0ee4),
	.w5(32'hb9eaaebc),
	.w6(32'h3b6dab58),
	.w7(32'h3adf4653),
	.w8(32'hb9edb941),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab11094),
	.w1(32'hbb0c741c),
	.w2(32'hbae529a1),
	.w3(32'hbae136e1),
	.w4(32'hbadaede9),
	.w5(32'hbb3ff760),
	.w6(32'hbb1883f8),
	.w7(32'hbb3d63a0),
	.w8(32'hbb1290bf),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2d420),
	.w1(32'hbaff81b4),
	.w2(32'hbba11a8b),
	.w3(32'hbb47a49d),
	.w4(32'hbb9d4c8b),
	.w5(32'hbc1481ae),
	.w6(32'hbae9d7f6),
	.w7(32'hb9b314a0),
	.w8(32'hbb8ed35d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6cb46),
	.w1(32'hbb2f7baf),
	.w2(32'hbc0f2d15),
	.w3(32'hbc16587a),
	.w4(32'hbaec04cf),
	.w5(32'hbc1e539c),
	.w6(32'hbc2b4e2d),
	.w7(32'hbb0b2e16),
	.w8(32'hbc08a390),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359794),
	.w1(32'hbaabc5c3),
	.w2(32'hba5a59ae),
	.w3(32'hbab39ed6),
	.w4(32'h3a0338ea),
	.w5(32'hbbb1681a),
	.w6(32'hb8a72117),
	.w7(32'h3abf4282),
	.w8(32'hbb91ba39),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e2f5),
	.w1(32'h3b8106d4),
	.w2(32'h3a78049c),
	.w3(32'hbad69b07),
	.w4(32'h3b81b694),
	.w5(32'h3a023f42),
	.w6(32'hbb4159c0),
	.w7(32'h38088839),
	.w8(32'hbb0e5f10),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeeac9),
	.w1(32'h396f4a13),
	.w2(32'hbb03fbaf),
	.w3(32'hbaece298),
	.w4(32'h3b9e3384),
	.w5(32'hbb3e25d6),
	.w6(32'hbb10f441),
	.w7(32'h3b51fbc7),
	.w8(32'hbb83bb6a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39863609),
	.w1(32'h3a0a9918),
	.w2(32'h3a791519),
	.w3(32'hb86bf087),
	.w4(32'h3911ba76),
	.w5(32'h3a810f38),
	.w6(32'hba80a08c),
	.w7(32'hb9817e1a),
	.w8(32'hbaa9b675),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73970e),
	.w1(32'h39e6c20b),
	.w2(32'hba08242b),
	.w3(32'hb99fcb97),
	.w4(32'h3a7f956d),
	.w5(32'h3b3df338),
	.w6(32'hba9dcc91),
	.w7(32'h3a221928),
	.w8(32'h3b3509b6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7e004),
	.w1(32'h3b1ad006),
	.w2(32'h3b800b28),
	.w3(32'h3b3a149e),
	.w4(32'h3a9f9fb4),
	.w5(32'hba6b297e),
	.w6(32'h3ba00f51),
	.w7(32'h3b6acd4e),
	.w8(32'h3b6ee2dc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f1e85),
	.w1(32'hbb2c9787),
	.w2(32'hbaaae0d8),
	.w3(32'h3affa307),
	.w4(32'h3b4a8329),
	.w5(32'h39f89aa7),
	.w6(32'h3988d788),
	.w7(32'hbb125bd8),
	.w8(32'h384911ed),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b283d4),
	.w1(32'hbadbd2d1),
	.w2(32'hbac52dec),
	.w3(32'hb9ccfc38),
	.w4(32'hbb1beb68),
	.w5(32'hb9c0b738),
	.w6(32'hbaff2f1e),
	.w7(32'hbb1250e9),
	.w8(32'hbaa69859),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb412356),
	.w1(32'hbb5abb24),
	.w2(32'hbb9d93f8),
	.w3(32'hb9e598c0),
	.w4(32'hba819e4a),
	.w5(32'hbbda56eb),
	.w6(32'hbb0186b2),
	.w7(32'hbb184dd2),
	.w8(32'hbbb854ae),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e6612),
	.w1(32'hbaeec8f0),
	.w2(32'hbb5325bd),
	.w3(32'hbb2d358e),
	.w4(32'hbae7b554),
	.w5(32'h38d78d65),
	.w6(32'hbb53ce0d),
	.w7(32'hbab959c6),
	.w8(32'hba234640),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b473750),
	.w1(32'h3ad36fc4),
	.w2(32'h3ae88128),
	.w3(32'h3b4ca230),
	.w4(32'h3b70ada1),
	.w5(32'h3a1aa399),
	.w6(32'h3b584650),
	.w7(32'h39e95b47),
	.w8(32'h394e3e6a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0af485),
	.w1(32'hbab3babc),
	.w2(32'hbbd9b0ec),
	.w3(32'hbb37cb8b),
	.w4(32'hbb55f46c),
	.w5(32'hbbcf88b4),
	.w6(32'hbaa1d021),
	.w7(32'hbb46fb54),
	.w8(32'hbbd2bd37),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ffac91),
	.w1(32'h39259c9b),
	.w2(32'hbb3153ac),
	.w3(32'h39ee4ec0),
	.w4(32'h39963bcd),
	.w5(32'h38686d28),
	.w6(32'hbac17e6d),
	.w7(32'h39e17810),
	.w8(32'h3730f877),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9baf2e),
	.w1(32'h3abf74cb),
	.w2(32'h3a203ee0),
	.w3(32'hbab67159),
	.w4(32'hbb0b8dc7),
	.w5(32'hba15df00),
	.w6(32'hbaa9d4f6),
	.w7(32'h3871d2e4),
	.w8(32'hba841582),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82b863),
	.w1(32'hbb0a1941),
	.w2(32'hbafe5976),
	.w3(32'hbb0bbeda),
	.w4(32'hb9fcba21),
	.w5(32'hb9a69efa),
	.w6(32'hbad11c3b),
	.w7(32'hbab27d50),
	.w8(32'hbb4cd219),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90a610),
	.w1(32'h3a104c1c),
	.w2(32'h3b6d21a5),
	.w3(32'h3b1aee7c),
	.w4(32'h3b557559),
	.w5(32'h3af70272),
	.w6(32'h3b08ad23),
	.w7(32'h3b1468d7),
	.w8(32'h3b0ad21e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db4b4a),
	.w1(32'hba8252b0),
	.w2(32'h398b4b69),
	.w3(32'h3a226301),
	.w4(32'h3973cbdc),
	.w5(32'h3a1f2def),
	.w6(32'hba0b6cd9),
	.w7(32'h39120446),
	.w8(32'hb9b7b7c6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b223c0),
	.w1(32'hb9c9d8a7),
	.w2(32'hbab77d9f),
	.w3(32'h3981882e),
	.w4(32'hba4efdce),
	.w5(32'hb9847a47),
	.w6(32'hbacbfbe1),
	.w7(32'hba6e7a1f),
	.w8(32'h39ec9dec),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d012d),
	.w1(32'hb98efa79),
	.w2(32'hb83fca0d),
	.w3(32'hb986d175),
	.w4(32'h36fb4507),
	.w5(32'h395bf982),
	.w6(32'hb7488f7f),
	.w7(32'h38844bf4),
	.w8(32'h3912099b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73f92c),
	.w1(32'h3b4a7a34),
	.w2(32'h3b074ab3),
	.w3(32'h3a470804),
	.w4(32'h3b36c37c),
	.w5(32'hba32582b),
	.w6(32'hbab537a0),
	.w7(32'h3af068d0),
	.w8(32'hb9da51f4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1d55d),
	.w1(32'hbbbeec1d),
	.w2(32'hbc280418),
	.w3(32'hbbb72b52),
	.w4(32'hbb16be3f),
	.w5(32'hbc007f35),
	.w6(32'hbb70df08),
	.w7(32'hbb1dc338),
	.w8(32'hbbf0bb16),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2e86c),
	.w1(32'hbb563199),
	.w2(32'hbbb77eac),
	.w3(32'hbb9dbfb7),
	.w4(32'hbb0ba9fd),
	.w5(32'hbb371ad6),
	.w6(32'hbb56b05f),
	.w7(32'hba856f3c),
	.w8(32'hbb6a221a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb878708),
	.w1(32'hbb84c410),
	.w2(32'hbbd53447),
	.w3(32'hbb866a98),
	.w4(32'hbb42b6d1),
	.w5(32'hbbac5975),
	.w6(32'hbb5e1377),
	.w7(32'hbabbeab7),
	.w8(32'hbb9fe912),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace3155),
	.w1(32'hbaaa173c),
	.w2(32'h3a932b8a),
	.w3(32'hb92c555c),
	.w4(32'h3a352cce),
	.w5(32'h391efaac),
	.w6(32'hbaa303a4),
	.w7(32'hba019fd9),
	.w8(32'h3b012439),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39506f96),
	.w1(32'h38e3bdcb),
	.w2(32'h3b182159),
	.w3(32'h3a81cee1),
	.w4(32'h3a8daf88),
	.w5(32'hba3b27bc),
	.w6(32'h3b0f95e6),
	.w7(32'h396e0d42),
	.w8(32'hb987d861),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f999f4),
	.w1(32'h3a0a9fa5),
	.w2(32'h3936c9cd),
	.w3(32'hba12ec10),
	.w4(32'hba14de58),
	.w5(32'h3a845606),
	.w6(32'hba106b57),
	.w7(32'hb80f988b),
	.w8(32'h3a8ee21d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a738cb5),
	.w1(32'h3a873926),
	.w2(32'h39794c89),
	.w3(32'h3af7c174),
	.w4(32'h3a95afe9),
	.w5(32'hb92956ad),
	.w6(32'h3a2d5635),
	.w7(32'h39eb5aaa),
	.w8(32'hba05a19b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb961761),
	.w1(32'hbb6adba0),
	.w2(32'hbc03838f),
	.w3(32'hba3b84a1),
	.w4(32'hba3ef4fa),
	.w5(32'hbaca8e70),
	.w6(32'hbb4769ea),
	.w7(32'hbb24fcde),
	.w8(32'hbb769b4d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a06b4),
	.w1(32'h37b29289),
	.w2(32'hb9ae608e),
	.w3(32'h3ad28c52),
	.w4(32'h39d7528f),
	.w5(32'hb9aa53c6),
	.w6(32'h3a03af8f),
	.w7(32'hba870208),
	.w8(32'h38c28061),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ac630),
	.w1(32'h3ae5d8f6),
	.w2(32'hbace7edd),
	.w3(32'hba92114e),
	.w4(32'h3aeb412b),
	.w5(32'h3a356a91),
	.w6(32'h3ae543c1),
	.w7(32'h3a9291dd),
	.w8(32'hba7a02a9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafabb66),
	.w1(32'hba98a003),
	.w2(32'h39d483d3),
	.w3(32'hbaa4fc46),
	.w4(32'hb94ce978),
	.w5(32'hbaa16548),
	.w6(32'hba90e661),
	.w7(32'h3a8acb6c),
	.w8(32'hba447faa),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a902c19),
	.w1(32'h3abff4d4),
	.w2(32'h3adad4a2),
	.w3(32'hbade0fdb),
	.w4(32'hb98c725a),
	.w5(32'h3980fac4),
	.w6(32'h3b103ea5),
	.w7(32'h3b3ac61f),
	.w8(32'h39a65ec6),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e4975),
	.w1(32'hb9df33a0),
	.w2(32'hba9b073c),
	.w3(32'hba66ecb2),
	.w4(32'h3aceb8fe),
	.w5(32'hbaa8d178),
	.w6(32'hb9aac3bf),
	.w7(32'hbac2a078),
	.w8(32'hbae4dfdd),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d0b7a),
	.w1(32'h3ae2e595),
	.w2(32'h3b1c7bce),
	.w3(32'hba9a588a),
	.w4(32'hba96c63a),
	.w5(32'h3a8a6576),
	.w6(32'h3a8e0d26),
	.w7(32'h3a2f4b5e),
	.w8(32'h3adacb06),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f2741),
	.w1(32'hbb3138c1),
	.w2(32'hbbd86199),
	.w3(32'hbad7a734),
	.w4(32'hba92ee17),
	.w5(32'hba5099c4),
	.w6(32'hba83a957),
	.w7(32'hba975fae),
	.w8(32'hbb2e70c6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b2cdb),
	.w1(32'h3a243d4c),
	.w2(32'h3ac48518),
	.w3(32'h38d1e9ae),
	.w4(32'hb9d38cad),
	.w5(32'h3a82b17b),
	.w6(32'hb9815370),
	.w7(32'h39a79216),
	.w8(32'h3a4043e9),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e4357),
	.w1(32'h3bd67717),
	.w2(32'h3b71a595),
	.w3(32'h3b57fd51),
	.w4(32'h3bd9bc8f),
	.w5(32'h3b288309),
	.w6(32'hbb73ab65),
	.w7(32'h3b2d066d),
	.w8(32'hba9d3a32),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule