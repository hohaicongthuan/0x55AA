module layer_8_featuremap_118(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf167c),
	.w1(32'h3b3dc014),
	.w2(32'h3bb7ac5a),
	.w3(32'h3a4e217f),
	.w4(32'h3c644ddb),
	.w5(32'hbacd12ee),
	.w6(32'h3a5c580d),
	.w7(32'h3c066bb6),
	.w8(32'hbb92bd6e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf34292),
	.w1(32'h3c5584f7),
	.w2(32'h3c3fa9b3),
	.w3(32'hbbfb6ea8),
	.w4(32'hb8f8bfa8),
	.w5(32'h3c3166f5),
	.w6(32'hb9bd2b50),
	.w7(32'hb794a98e),
	.w8(32'h3a2d7e7a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12bf72),
	.w1(32'h3b9f3326),
	.w2(32'hbb3f6424),
	.w3(32'h3b927512),
	.w4(32'h3b4f3834),
	.w5(32'hbac74284),
	.w6(32'h3bc379a6),
	.w7(32'h3c98e2e2),
	.w8(32'hbc894c20),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c386e63),
	.w1(32'hbb6f3f6d),
	.w2(32'h3c00da65),
	.w3(32'h3b2512b0),
	.w4(32'hba0d0db4),
	.w5(32'hbc00f9b4),
	.w6(32'hbae8f846),
	.w7(32'hbacd54dc),
	.w8(32'h3c0e3d42),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35b358),
	.w1(32'hbbce6622),
	.w2(32'h3ce11a92),
	.w3(32'hba5c95a2),
	.w4(32'h3b7ce642),
	.w5(32'hbd0e6b26),
	.w6(32'h3c9b8258),
	.w7(32'h3b90f365),
	.w8(32'hbc933f1b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcefeb9e),
	.w1(32'hbce19e0b),
	.w2(32'hbc461576),
	.w3(32'h3b9466dc),
	.w4(32'h3b9c16aa),
	.w5(32'hba979f89),
	.w6(32'hbc717994),
	.w7(32'h3c25ea01),
	.w8(32'hbcb82dc4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1b340),
	.w1(32'hbca94837),
	.w2(32'hbc96803f),
	.w3(32'hbc11a7c3),
	.w4(32'h3bb60d6b),
	.w5(32'hbc85b8ea),
	.w6(32'h3c44388d),
	.w7(32'hbd35a51d),
	.w8(32'h3c6dc086),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb991500),
	.w1(32'hbc0a3b0b),
	.w2(32'h3bcf1ff4),
	.w3(32'hbcd6c255),
	.w4(32'h3bfa10f5),
	.w5(32'hbc32c061),
	.w6(32'hbc7daa6c),
	.w7(32'hbcbc9c34),
	.w8(32'hbc143ee9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51f987),
	.w1(32'hbbe4c65b),
	.w2(32'h3bbc1e73),
	.w3(32'hbc8a319c),
	.w4(32'hbbae6e75),
	.w5(32'h3bc0332c),
	.w6(32'h3bbaa408),
	.w7(32'hbc6a5c0d),
	.w8(32'h3ca056f1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb305b77),
	.w1(32'h3b7ac752),
	.w2(32'hbb7fc731),
	.w3(32'hbc0f4586),
	.w4(32'hbb7e7339),
	.w5(32'hbcacb500),
	.w6(32'hbc1cfaa1),
	.w7(32'hb9ea2f94),
	.w8(32'h3d6adaa4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca50e32),
	.w1(32'hbb9eadcd),
	.w2(32'hbc6f023a),
	.w3(32'h39bbad98),
	.w4(32'hbbd7dd4f),
	.w5(32'h3aad12c1),
	.w6(32'hbc1610ff),
	.w7(32'h3b3482df),
	.w8(32'hbc346272),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12ae24),
	.w1(32'h3b456f76),
	.w2(32'hbba0644c),
	.w3(32'hbc7bd543),
	.w4(32'hbbfdc57d),
	.w5(32'hbbc0de46),
	.w6(32'h3bc891d9),
	.w7(32'hbb8fd7db),
	.w8(32'hbc8ef0c2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2c5c2),
	.w1(32'hbb39f118),
	.w2(32'h396f95e1),
	.w3(32'hbbcbe495),
	.w4(32'hbac7d9a7),
	.w5(32'h3af1b72b),
	.w6(32'h3b9834d9),
	.w7(32'h3ba737ee),
	.w8(32'h3c86b703),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fe6a4),
	.w1(32'h3b4e5b0c),
	.w2(32'hbb573262),
	.w3(32'h3c0a8eec),
	.w4(32'hba9dbe53),
	.w5(32'hbb5b6e39),
	.w6(32'hbade77c0),
	.w7(32'hbadd1449),
	.w8(32'h3a73a2cd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f92a3a),
	.w1(32'h3b0ecc2a),
	.w2(32'hbadf8d35),
	.w3(32'h3ac7de35),
	.w4(32'h3a0f7c00),
	.w5(32'h3a222b06),
	.w6(32'hbb85f07c),
	.w7(32'h3ac54584),
	.w8(32'h3a86443e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90f1966),
	.w1(32'hbac51086),
	.w2(32'h3b950913),
	.w3(32'h3b9e6161),
	.w4(32'h3b140d4e),
	.w5(32'h3a49b220),
	.w6(32'h3abcaa78),
	.w7(32'hbcadf006),
	.w8(32'hbc302fa2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07b303),
	.w1(32'hbac5a53a),
	.w2(32'hbbc21d5b),
	.w3(32'hbc76c6be),
	.w4(32'h3b70cf55),
	.w5(32'h3c848816),
	.w6(32'hba6c2227),
	.w7(32'h3c82b22f),
	.w8(32'hbbeb09a8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c766786),
	.w1(32'h3c112968),
	.w2(32'hbc5aedfd),
	.w3(32'h3bf0c4f1),
	.w4(32'hbc878490),
	.w5(32'hbbe12247),
	.w6(32'hba6ed0cd),
	.w7(32'h3bcc3c9e),
	.w8(32'hbc33883d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f3dbd),
	.w1(32'hbb16b75d),
	.w2(32'h3b0a7005),
	.w3(32'hbbafb050),
	.w4(32'h3c14c899),
	.w5(32'hbab77377),
	.w6(32'h3bd7b476),
	.w7(32'hbb29defa),
	.w8(32'hbbabe110),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b5751),
	.w1(32'hbb279021),
	.w2(32'hbca4efd7),
	.w3(32'h3b086a4b),
	.w4(32'hbb195bf8),
	.w5(32'hbcdf6288),
	.w6(32'hbc020232),
	.w7(32'h3cb0350c),
	.w8(32'h3d245a58),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1719a9),
	.w1(32'h3bbc5c1c),
	.w2(32'h3b87e958),
	.w3(32'hbc008e22),
	.w4(32'hbbbe3858),
	.w5(32'h3c80d4d1),
	.w6(32'hbcd5aa33),
	.w7(32'hbc8ae8fd),
	.w8(32'hbc1434b4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddd62f),
	.w1(32'h3be3f50a),
	.w2(32'h3c9ddc22),
	.w3(32'hbb459ed1),
	.w4(32'hbbec1d2b),
	.w5(32'h3b4d8e68),
	.w6(32'hbc96d0c8),
	.w7(32'hbb5b9594),
	.w8(32'hbbd78114),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c211a30),
	.w1(32'hbb07b245),
	.w2(32'hbc7e40c4),
	.w3(32'hbb59bc2e),
	.w4(32'h3b843ad1),
	.w5(32'hb991e1af),
	.w6(32'hbb350081),
	.w7(32'h3b4b69a2),
	.w8(32'hb8b274cc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dbaa6),
	.w1(32'h3c12eb3e),
	.w2(32'hbb1b964e),
	.w3(32'hbc1c652c),
	.w4(32'h3b559378),
	.w5(32'h3b8c7508),
	.w6(32'h3c0909f6),
	.w7(32'h3c05332d),
	.w8(32'h3b248e33),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed67a2),
	.w1(32'hbc0fbd9f),
	.w2(32'hbbd3b179),
	.w3(32'h3928a439),
	.w4(32'hbbd9bbdc),
	.w5(32'h3b856ba7),
	.w6(32'hbab8b243),
	.w7(32'h3b8127a2),
	.w8(32'hbbd5e7a3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d260a),
	.w1(32'hbaa8df51),
	.w2(32'h3c868bbd),
	.w3(32'hbc100193),
	.w4(32'h3bc100cc),
	.w5(32'h3cae212c),
	.w6(32'hbb505a54),
	.w7(32'hbcd4d284),
	.w8(32'hbd8ea277),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d57851f),
	.w1(32'h3c612f59),
	.w2(32'hbbcef3b6),
	.w3(32'hbb415c0d),
	.w4(32'hbc36b71c),
	.w5(32'hbbfafa4a),
	.w6(32'h3cd54333),
	.w7(32'hb9a1f883),
	.w8(32'h3b1bd3db),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca19198),
	.w1(32'hbcb804a6),
	.w2(32'hbc2ece50),
	.w3(32'h3b393753),
	.w4(32'hba61b7cf),
	.w5(32'hbbc53125),
	.w6(32'h39c3c4eb),
	.w7(32'hbcad5460),
	.w8(32'hbcd0b937),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc7c5a3),
	.w1(32'h3c0ae4c3),
	.w2(32'hbbc24b64),
	.w3(32'hbc974e79),
	.w4(32'h3b3815ee),
	.w5(32'hbb928b51),
	.w6(32'h3b4628c7),
	.w7(32'h3c7401a7),
	.w8(32'hbcbb3789),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc143145),
	.w1(32'h3cab25bd),
	.w2(32'hbcd4a13a),
	.w3(32'hba30dc96),
	.w4(32'h3b7cd06d),
	.w5(32'h3c6eab9f),
	.w6(32'h3c1e6918),
	.w7(32'h3d56a17a),
	.w8(32'hbd034f0c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf93ef2),
	.w1(32'h3ca77a40),
	.w2(32'h3bb22e84),
	.w3(32'h3c6dddfb),
	.w4(32'h3bc5997a),
	.w5(32'h3b88dc14),
	.w6(32'hbd57213b),
	.w7(32'h3b6dd97b),
	.w8(32'h3b75ada5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93adf8a),
	.w1(32'h3b725f22),
	.w2(32'hbc948189),
	.w3(32'h3c091131),
	.w4(32'hbb8c5749),
	.w5(32'hbca3b483),
	.w6(32'h3b2145b9),
	.w7(32'hbc9b73e1),
	.w8(32'h3d714391),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd6780),
	.w1(32'h3bf12963),
	.w2(32'hbcc33522),
	.w3(32'hbcac2e54),
	.w4(32'hbc8c8c3f),
	.w5(32'h3d04cd1a),
	.w6(32'hbc378242),
	.w7(32'h3d665424),
	.w8(32'h3b3f0f92),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0fa4f9),
	.w1(32'h3c2fdd63),
	.w2(32'h3c005de8),
	.w3(32'h3c93d182),
	.w4(32'hbc533f73),
	.w5(32'h3c0f274d),
	.w6(32'hbd153a35),
	.w7(32'h3a31a858),
	.w8(32'hbc785064),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd23f28),
	.w1(32'h3b26d46d),
	.w2(32'h3b77f8aa),
	.w3(32'h3b8a23e1),
	.w4(32'h3b8addfd),
	.w5(32'h3a1bf55c),
	.w6(32'h3cdd5d73),
	.w7(32'h3a609691),
	.w8(32'hbad61d6c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9af3a),
	.w1(32'h3bb2b1ae),
	.w2(32'hbcb89b7d),
	.w3(32'h3c1c0b80),
	.w4(32'hbc1b8cc7),
	.w5(32'h3b8d512b),
	.w6(32'h3b54c55e),
	.w7(32'h3cbced0b),
	.w8(32'h3c1e988d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1332c),
	.w1(32'hbcc5079a),
	.w2(32'hbab144e1),
	.w3(32'h3a4994df),
	.w4(32'hbc6bd2fd),
	.w5(32'hbad4e5eb),
	.w6(32'h3d01423f),
	.w7(32'hbca479aa),
	.w8(32'h3b983215),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc275490),
	.w1(32'hbc400e7e),
	.w2(32'h3c820416),
	.w3(32'h3bdff440),
	.w4(32'hbbc031a1),
	.w5(32'hbbeeda2e),
	.w6(32'hbb3abbb5),
	.w7(32'hbc145797),
	.w8(32'hbc477145),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cf261),
	.w1(32'h3bf25381),
	.w2(32'hbbf9205c),
	.w3(32'hbb8663d1),
	.w4(32'hbaeb8d73),
	.w5(32'hbc4fcb50),
	.w6(32'h3add84a3),
	.w7(32'hbb977c9c),
	.w8(32'hbb34d65e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea519d),
	.w1(32'h3c60f4e2),
	.w2(32'h3b6d59d8),
	.w3(32'hbc32361c),
	.w4(32'h3bb3c846),
	.w5(32'hbb1d9aeb),
	.w6(32'hbb15e9a4),
	.w7(32'hbb3ea209),
	.w8(32'hbb7fbfc0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baed063),
	.w1(32'hbb92b7a7),
	.w2(32'h3c138683),
	.w3(32'hbb5e0a67),
	.w4(32'h3c86d4bd),
	.w5(32'hbcd91f25),
	.w6(32'hbc191b4c),
	.w7(32'hbc9b35c3),
	.w8(32'h3d27d420),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1efd23),
	.w1(32'h3b5d1ff0),
	.w2(32'hbbdb784f),
	.w3(32'hbc5237fd),
	.w4(32'h39a5b66b),
	.w5(32'h3bc43f71),
	.w6(32'h3c2d4ce4),
	.w7(32'hbbcf9499),
	.w8(32'hbb6d6465),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc109047),
	.w1(32'hbc4ec579),
	.w2(32'hbcb61faf),
	.w3(32'hbc242839),
	.w4(32'hbc246e40),
	.w5(32'hbad1f4c1),
	.w6(32'h3c21d4a5),
	.w7(32'h3cf0cd17),
	.w8(32'h3d750079),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9b1b21),
	.w1(32'hbb9f081b),
	.w2(32'hba5ceef1),
	.w3(32'h3c8187fd),
	.w4(32'hba7f2342),
	.w5(32'h3b289261),
	.w6(32'hbcb3f597),
	.w7(32'h3b3921a6),
	.w8(32'h3c22e51c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb442ebb),
	.w1(32'h3b6006f0),
	.w2(32'hbc510f2f),
	.w3(32'h3c04ae61),
	.w4(32'hbaa511fc),
	.w5(32'hbc0098a6),
	.w6(32'hbbedeb43),
	.w7(32'h3c5c53e7),
	.w8(32'hbbccf8e4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19f3bf),
	.w1(32'h3c447714),
	.w2(32'hbca2813b),
	.w3(32'hbb57e819),
	.w4(32'h3bafedad),
	.w5(32'hbb0aad90),
	.w6(32'h3b13a7c2),
	.w7(32'h3cc5878b),
	.w8(32'h3d30d7d9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabae84),
	.w1(32'hbc879455),
	.w2(32'h3bc9120b),
	.w3(32'h3bdf463e),
	.w4(32'h3b71bf76),
	.w5(32'h3b7dd291),
	.w6(32'h3c0e89ea),
	.w7(32'hbc034726),
	.w8(32'hbc761c07),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb263c2),
	.w1(32'h3c74f6e7),
	.w2(32'hbb8e1c52),
	.w3(32'hba1ea53a),
	.w4(32'hba5f6776),
	.w5(32'h3ca3b644),
	.w6(32'h3a5b5afe),
	.w7(32'h3c91badc),
	.w8(32'hbc568b04),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a858843),
	.w1(32'h3c580e6b),
	.w2(32'h3c63b580),
	.w3(32'hbb116d1d),
	.w4(32'hbc81fc9b),
	.w5(32'hba8896d6),
	.w6(32'hbcc08a73),
	.w7(32'h3ba98e4e),
	.w8(32'hbd2cbb30),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c54a5),
	.w1(32'hbd373cee),
	.w2(32'hbc80dc32),
	.w3(32'hbc00b7bf),
	.w4(32'hbd0028aa),
	.w5(32'hbcff863b),
	.w6(32'hbbc1efb1),
	.w7(32'hbcf248dd),
	.w8(32'hbbf83692),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53d678),
	.w1(32'hbcbcac80),
	.w2(32'h3c014f8d),
	.w3(32'hbcefc417),
	.w4(32'hbb8e65cd),
	.w5(32'h3bf79084),
	.w6(32'hbcb32254),
	.w7(32'hbb07c0ca),
	.w8(32'hbd101364),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfd57bc),
	.w1(32'h3c1ba116),
	.w2(32'h3be20396),
	.w3(32'hbb3f52d6),
	.w4(32'h3ac86b0b),
	.w5(32'h3a791659),
	.w6(32'hbba551bc),
	.w7(32'hbd065f8c),
	.w8(32'hbc94bf59),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb760a19),
	.w1(32'h3cb73057),
	.w2(32'hbc2a91c6),
	.w3(32'hbc58b45d),
	.w4(32'h3c782084),
	.w5(32'hbcd820c8),
	.w6(32'hbc908a75),
	.w7(32'hbcbf3895),
	.w8(32'h3ce0f226),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd2379),
	.w1(32'h3c7c827d),
	.w2(32'hbb382eb5),
	.w3(32'hbbee75b9),
	.w4(32'h38e5b802),
	.w5(32'h3b31a63a),
	.w6(32'hbbb7c72d),
	.w7(32'h3b2f0ee5),
	.w8(32'h3bf12266),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6434ed),
	.w1(32'h3b19354f),
	.w2(32'hbc430748),
	.w3(32'h3c0a52c4),
	.w4(32'h3c501e2f),
	.w5(32'h3c5d50c5),
	.w6(32'hbb7177b1),
	.w7(32'h3a818507),
	.w8(32'hbd01166b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359f74),
	.w1(32'hbc18f87d),
	.w2(32'h3c29f6cb),
	.w3(32'h3ba4a8e9),
	.w4(32'h3b56ddd6),
	.w5(32'hbc8bc97e),
	.w6(32'hbbbaba81),
	.w7(32'h38e9ff02),
	.w8(32'h3b071772),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b38e6),
	.w1(32'hbb05228e),
	.w2(32'hbac0ba97),
	.w3(32'hbb0856ef),
	.w4(32'h3a3516c0),
	.w5(32'h3b021ce2),
	.w6(32'hbaa7d70e),
	.w7(32'hbaad0719),
	.w8(32'hba89527b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8f20c),
	.w1(32'hb91587eb),
	.w2(32'hbc51c3bd),
	.w3(32'hb67aec7b),
	.w4(32'h3c9fe901),
	.w5(32'h3c6a8dea),
	.w6(32'hbaec35b2),
	.w7(32'h3b42b788),
	.w8(32'hbd0142f9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb282ed),
	.w1(32'h3ce43e6f),
	.w2(32'hbb09a2fc),
	.w3(32'hbbb41a36),
	.w4(32'h3988ca51),
	.w5(32'h3b1fe7d3),
	.w6(32'hbc556c53),
	.w7(32'h3b560887),
	.w8(32'h3bebaf5d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c35b9),
	.w1(32'h3ac4e159),
	.w2(32'h3c921116),
	.w3(32'h3bfc86c6),
	.w4(32'h3b471cd3),
	.w5(32'hbc9fe402),
	.w6(32'hbbd90721),
	.w7(32'hbd5d5625),
	.w8(32'h3d10dfae),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47936a),
	.w1(32'hbc221421),
	.w2(32'hbc6a2ebf),
	.w3(32'hbc92cd46),
	.w4(32'hbbf3a3b8),
	.w5(32'hbd2c9913),
	.w6(32'h3d3c62a0),
	.w7(32'hbc656674),
	.w8(32'h3d2bf362),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b34b8),
	.w1(32'h3c402e71),
	.w2(32'hbb92ceef),
	.w3(32'hbbe0d28b),
	.w4(32'hbba7919f),
	.w5(32'hbbee5266),
	.w6(32'h3caacece),
	.w7(32'hbbb6c1cc),
	.w8(32'hbbfd6975),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafae8b9),
	.w1(32'h3ab11f92),
	.w2(32'h3c3ebd4d),
	.w3(32'hbbb47d15),
	.w4(32'hbae4d7da),
	.w5(32'h3bc5b02d),
	.w6(32'hbb0e6c66),
	.w7(32'hbb136c90),
	.w8(32'hbb8819e7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba82c70),
	.w1(32'hbb6d9d8a),
	.w2(32'h3b1966f7),
	.w3(32'h3b907c13),
	.w4(32'h3b663ee0),
	.w5(32'hbc153f56),
	.w6(32'hbc532707),
	.w7(32'h3c8d45bc),
	.w8(32'h3cc13594),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bc890),
	.w1(32'h3c6c3583),
	.w2(32'h3b731d86),
	.w3(32'hbaedac72),
	.w4(32'h3bf8a79c),
	.w5(32'h3c66f2fb),
	.w6(32'hbb0eb10b),
	.w7(32'h3952c730),
	.w8(32'hbc2935c3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cd997),
	.w1(32'h3c1d9010),
	.w2(32'hbb7c0c91),
	.w3(32'h3ba219d0),
	.w4(32'hbc0de417),
	.w5(32'h3c5e0a70),
	.w6(32'hbc26b370),
	.w7(32'h3c21c84e),
	.w8(32'hbb39445b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dadd3),
	.w1(32'h3a40d054),
	.w2(32'hbb323ae9),
	.w3(32'h3c2e2b73),
	.w4(32'hbba05f04),
	.w5(32'h3ad4fae6),
	.w6(32'h3b8e8da1),
	.w7(32'hbc5911dd),
	.w8(32'hbb986386),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5b7c5),
	.w1(32'h3c5c3ea3),
	.w2(32'h3bb4d3bd),
	.w3(32'hbbde36c6),
	.w4(32'hbc951963),
	.w5(32'hb90b6f02),
	.w6(32'h3c43f2a4),
	.w7(32'hbbb7885b),
	.w8(32'h3d97c1a7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13ae19),
	.w1(32'hbc83fd75),
	.w2(32'hbc60ec93),
	.w3(32'h3a937337),
	.w4(32'h3c2e67bb),
	.w5(32'h3c89988e),
	.w6(32'hbba1b04d),
	.w7(32'hbcb2f2b3),
	.w8(32'h3b4925bd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48497c),
	.w1(32'h3c15b9c6),
	.w2(32'h3b19f4d9),
	.w3(32'hbbbd8293),
	.w4(32'h3b74104c),
	.w5(32'h3bbfb65f),
	.w6(32'hbb1c6d93),
	.w7(32'h3b837522),
	.w8(32'h3b82956a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4fdc4),
	.w1(32'h3c444a98),
	.w2(32'hbc8d8ca5),
	.w3(32'h3c1a7197),
	.w4(32'hbc7e8960),
	.w5(32'hbcc7353c),
	.w6(32'hbcc0c08b),
	.w7(32'hbc975b77),
	.w8(32'h3ced0ad4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b0693),
	.w1(32'hbbed2804),
	.w2(32'h3b73dc46),
	.w3(32'hbbd853ef),
	.w4(32'hbb8f6888),
	.w5(32'hbbca486b),
	.w6(32'hbcc45add),
	.w7(32'h3baf2044),
	.w8(32'hbbdeeed4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b685414),
	.w1(32'hbc3a7393),
	.w2(32'hb995125b),
	.w3(32'h3b3eb71d),
	.w4(32'h3b332052),
	.w5(32'h3c4ce280),
	.w6(32'h3c6aa9fb),
	.w7(32'h3abeb070),
	.w8(32'h3d401688),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f1fb8),
	.w1(32'hbba726c2),
	.w2(32'hbc0a91c2),
	.w3(32'h3c3d0e0d),
	.w4(32'h3b9d6706),
	.w5(32'hbbb3a67d),
	.w6(32'hba01a694),
	.w7(32'h3c08c4ff),
	.w8(32'h3d02736c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed6baa),
	.w1(32'hbc139290),
	.w2(32'h3c086e32),
	.w3(32'h3c3d90c7),
	.w4(32'hbc7fbd3e),
	.w5(32'hbb234f12),
	.w6(32'hbb904c0a),
	.w7(32'hbbaa7910),
	.w8(32'hbc63b2c7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c830703),
	.w1(32'h3bff07d8),
	.w2(32'hbae46f3b),
	.w3(32'hbb04afd4),
	.w4(32'h3b795eb9),
	.w5(32'hbb9516bc),
	.w6(32'h3b3e4c9d),
	.w7(32'hb9006401),
	.w8(32'h3c848b1d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7722b8),
	.w1(32'hbb76e9e9),
	.w2(32'h3ad1fbc9),
	.w3(32'h3c9c8f5a),
	.w4(32'h3b2ff52a),
	.w5(32'h3a197a02),
	.w6(32'hbc51d5c7),
	.w7(32'h3c370a70),
	.w8(32'h3bc56da7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b756c28),
	.w1(32'h3a4f0ca5),
	.w2(32'hb91b3828),
	.w3(32'h3a4a9cc7),
	.w4(32'h39adb758),
	.w5(32'h3c12707e),
	.w6(32'h3a728940),
	.w7(32'h3b4f2641),
	.w8(32'h3bb21697),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47d970),
	.w1(32'h3af3fbde),
	.w2(32'h3b003ff5),
	.w3(32'h3b8e7abf),
	.w4(32'h38bece94),
	.w5(32'h3a017698),
	.w6(32'h3b703169),
	.w7(32'h3b3f9816),
	.w8(32'h3afdf6ec),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b396651),
	.w1(32'h3a8db362),
	.w2(32'h3c43278b),
	.w3(32'h3af08835),
	.w4(32'h3c280521),
	.w5(32'h3b6e59d3),
	.w6(32'hbaa14ead),
	.w7(32'h3c71ff3a),
	.w8(32'h3b963486),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc542e5c),
	.w1(32'hbbbff323),
	.w2(32'h3ac22c7f),
	.w3(32'h3b6c83ef),
	.w4(32'h3c6ec157),
	.w5(32'hbc5b688d),
	.w6(32'h3b096a69),
	.w7(32'h3cc3204e),
	.w8(32'h3d1b9d9d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97d433),
	.w1(32'hb8ad7af5),
	.w2(32'h3c089ac5),
	.w3(32'hbc87d65a),
	.w4(32'h3a8d4753),
	.w5(32'hbc695679),
	.w6(32'hbbcac43a),
	.w7(32'hba963f7a),
	.w8(32'hbc92c1db),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadba47a),
	.w1(32'hbbe61ee1),
	.w2(32'hbcab84c0),
	.w3(32'hbb9dcc4b),
	.w4(32'h3c76fbf1),
	.w5(32'h3ab6d91f),
	.w6(32'hbc3c2238),
	.w7(32'h3bdc474e),
	.w8(32'h3c231a5e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d16d32f),
	.w1(32'h3ab9a260),
	.w2(32'hbc4689ba),
	.w3(32'h3b2ea706),
	.w4(32'hbaf11201),
	.w5(32'hbc14af49),
	.w6(32'h3bdd0e37),
	.w7(32'h3a1b202d),
	.w8(32'hbc6b771f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b773ffc),
	.w1(32'h3b2b2dfe),
	.w2(32'hbc452197),
	.w3(32'h3ae223d5),
	.w4(32'h3bf33ca3),
	.w5(32'h3cc7245c),
	.w6(32'hbca49eae),
	.w7(32'hbccf57a2),
	.w8(32'h3d95dd99),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafa186),
	.w1(32'h3bfeb151),
	.w2(32'hbaef27fc),
	.w3(32'hbafe5c22),
	.w4(32'hbc0007a8),
	.w5(32'h3c40aab0),
	.w6(32'h3c3dd141),
	.w7(32'hbc02203d),
	.w8(32'h3c987f4a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc935b7c),
	.w1(32'hbb49b3f5),
	.w2(32'h3ad54275),
	.w3(32'hbc0b2cc9),
	.w4(32'hbb4e14d3),
	.w5(32'hbc3a41b3),
	.w6(32'h3ad3a24e),
	.w7(32'hbb9ac8aa),
	.w8(32'hba0a9e68),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fd382),
	.w1(32'hbbeae4d1),
	.w2(32'h3c7ae6bf),
	.w3(32'hb9f61668),
	.w4(32'h3b81ba72),
	.w5(32'h3b82a7d4),
	.w6(32'hbc8a2471),
	.w7(32'h3c1cf33b),
	.w8(32'h3b8ea8a1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b6c5e),
	.w1(32'hbacb1baa),
	.w2(32'hbad425e6),
	.w3(32'hbc1325d5),
	.w4(32'h3c1d0933),
	.w5(32'h3b305625),
	.w6(32'hb9b24022),
	.w7(32'h3b68f8ea),
	.w8(32'h3aeee8fa),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6f12d),
	.w1(32'h3b2a5d1b),
	.w2(32'hbcaa514a),
	.w3(32'h39a798b6),
	.w4(32'hbad63d2a),
	.w5(32'h3b547f45),
	.w6(32'h39a01767),
	.w7(32'h3bd48ccb),
	.w8(32'h3c828aa4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc686cc1),
	.w1(32'hbbfec4a2),
	.w2(32'hbadb00b6),
	.w3(32'h3baa0c5e),
	.w4(32'h3bd6f1be),
	.w5(32'hbc25a29c),
	.w6(32'h3c37d9f1),
	.w7(32'h3cfbdcc6),
	.w8(32'hbcc83364),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99136f),
	.w1(32'h3c8ed93d),
	.w2(32'h3c0cc3cb),
	.w3(32'h3bec1070),
	.w4(32'h3bb42e15),
	.w5(32'hbc83a821),
	.w6(32'h3c319e84),
	.w7(32'hbb227671),
	.w8(32'hbca67753),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce6590f),
	.w1(32'h3b6c85f6),
	.w2(32'hbb406f7b),
	.w3(32'hbc0bd461),
	.w4(32'hbb259343),
	.w5(32'hbc98da3e),
	.w6(32'hbba6cd29),
	.w7(32'h3c019215),
	.w8(32'hbcc35a6a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b279893),
	.w1(32'hbba0d2d2),
	.w2(32'h3b4f02a0),
	.w3(32'hbb2fe387),
	.w4(32'hbbbe7839),
	.w5(32'h3b9853b0),
	.w6(32'hbb810ab4),
	.w7(32'hbbb57282),
	.w8(32'hbb987907),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd17c8da),
	.w1(32'hbbd8ccc3),
	.w2(32'hba42ff3b),
	.w3(32'h3be8873f),
	.w4(32'h39f96d12),
	.w5(32'hbacaa0c8),
	.w6(32'h3c9e7eee),
	.w7(32'h3a0236a5),
	.w8(32'hbafade5f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940d52d),
	.w1(32'hb8aa4c95),
	.w2(32'h3cda8ff5),
	.w3(32'hba0fb6ec),
	.w4(32'h3b430ef2),
	.w5(32'h3ac3023c),
	.w6(32'hbb1db3d0),
	.w7(32'h3ac09d56),
	.w8(32'hbb48d04b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf45b60),
	.w1(32'hbaacfa4a),
	.w2(32'h3b058587),
	.w3(32'hbabdb7a1),
	.w4(32'hbd05367b),
	.w5(32'h3bffdeb5),
	.w6(32'h3c9596b2),
	.w7(32'hbc66d0b7),
	.w8(32'h3c9ee91e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d080ae2),
	.w1(32'hbc47d802),
	.w2(32'hba210212),
	.w3(32'hbb9a113a),
	.w4(32'hbb3dc359),
	.w5(32'hb840a9db),
	.w6(32'hbc5eecf5),
	.w7(32'hbbb4d7b8),
	.w8(32'h3ccab9e4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addae49),
	.w1(32'hbac08bfe),
	.w2(32'hbc3b736e),
	.w3(32'hbc3b6a7a),
	.w4(32'hbb273fc3),
	.w5(32'h3a353c0e),
	.w6(32'hbab75a43),
	.w7(32'hbc20ab95),
	.w8(32'h3b3a7d89),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb445d03),
	.w1(32'h3c0545ec),
	.w2(32'h3c506c5c),
	.w3(32'h3b644a03),
	.w4(32'h3a97e451),
	.w5(32'hbbc0fc08),
	.w6(32'h3b67bfb2),
	.w7(32'h3b9cd214),
	.w8(32'hbc1f3482),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d59f7),
	.w1(32'hbba8f41a),
	.w2(32'hbb877238),
	.w3(32'h3c02512e),
	.w4(32'hbbbfe6ac),
	.w5(32'h3a1c4d7c),
	.w6(32'hbcb0fd55),
	.w7(32'h3c160ca3),
	.w8(32'h3c235420),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277ff0),
	.w1(32'hb9c2070e),
	.w2(32'h3b6bd565),
	.w3(32'hb9e4e580),
	.w4(32'h3b186311),
	.w5(32'hbc9ee43f),
	.w6(32'hbb83fd8d),
	.w7(32'h3c66cf1a),
	.w8(32'hbc498315),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1c28b),
	.w1(32'hbb63d78e),
	.w2(32'hbab45e7e),
	.w3(32'hbc0bd074),
	.w4(32'h3a392134),
	.w5(32'hbc00f553),
	.w6(32'h3aa8d2b0),
	.w7(32'hbb1d8777),
	.w8(32'h3c9ddb8f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee08aa),
	.w1(32'hbaf2a3fe),
	.w2(32'hbbfd35ec),
	.w3(32'hbc31fd0e),
	.w4(32'hbaf2391b),
	.w5(32'hbb1c5b5a),
	.w6(32'hbb5601bf),
	.w7(32'hbb89dc67),
	.w8(32'hbc0ccbc5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07c378),
	.w1(32'h3af5cec2),
	.w2(32'h3b74b2e1),
	.w3(32'h3c4525a7),
	.w4(32'h3a004d6d),
	.w5(32'hbad60b93),
	.w6(32'hba5aa081),
	.w7(32'h3bc6915c),
	.w8(32'hbca49940),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37d8d5),
	.w1(32'h3bb5a3e6),
	.w2(32'hbc32662b),
	.w3(32'h3c31df99),
	.w4(32'hbc7b0188),
	.w5(32'hba8ecf18),
	.w6(32'h3b7daab7),
	.w7(32'hbc9e5442),
	.w8(32'hbce762d2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37549e),
	.w1(32'h3b9f63ff),
	.w2(32'hbbcffdf7),
	.w3(32'h3c1c91ae),
	.w4(32'hbb979735),
	.w5(32'hbb470786),
	.w6(32'h3bceb11c),
	.w7(32'hbc216796),
	.w8(32'h3cdad916),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80b145),
	.w1(32'hbb25ece2),
	.w2(32'hb98e8de2),
	.w3(32'hbbb586dd),
	.w4(32'h39ef4f20),
	.w5(32'hbb3ba624),
	.w6(32'hbbff7903),
	.w7(32'h3c37fb4b),
	.w8(32'h3b347fc2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9acaf5),
	.w1(32'h3a7727df),
	.w2(32'h3c54d358),
	.w3(32'h3a6c9f23),
	.w4(32'hb9e91c1c),
	.w5(32'h3b9e4d68),
	.w6(32'hba356205),
	.w7(32'h3bd6db30),
	.w8(32'h3c44ea4c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88081a),
	.w1(32'h3b7d90be),
	.w2(32'hbb5aee37),
	.w3(32'h3bc9b09e),
	.w4(32'hbc982291),
	.w5(32'hbbbdf1a0),
	.w6(32'h3c2dcb31),
	.w7(32'hbc24601c),
	.w8(32'hbd0b8a7c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc958284),
	.w1(32'hbc1986e2),
	.w2(32'hbb2fcc08),
	.w3(32'h3bf49516),
	.w4(32'hbc8c1b3d),
	.w5(32'hba9544ef),
	.w6(32'hbc4fcc13),
	.w7(32'h3bd435a3),
	.w8(32'hbb91bf94),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b968e30),
	.w1(32'hbc2b3475),
	.w2(32'hbbfabd37),
	.w3(32'h3a548efc),
	.w4(32'hbc5e6405),
	.w5(32'h3c07fe60),
	.w6(32'h3abf2458),
	.w7(32'hbba2b785),
	.w8(32'h3b8856d6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d5ae),
	.w1(32'hbba79949),
	.w2(32'h3c3f8d8c),
	.w3(32'hbc8151b4),
	.w4(32'hbafa605c),
	.w5(32'h3b5b290d),
	.w6(32'hbc05c766),
	.w7(32'h3c14795c),
	.w8(32'hbbbfc583),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d2e10),
	.w1(32'hbbbfcc46),
	.w2(32'h3cd58549),
	.w3(32'hba52799f),
	.w4(32'hbb459775),
	.w5(32'hbca427d4),
	.w6(32'h3b21930b),
	.w7(32'h3ce280d9),
	.w8(32'hbcb2f92d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfffce),
	.w1(32'hbc98a21e),
	.w2(32'hbb571ad3),
	.w3(32'hbc4f799c),
	.w4(32'h3ad4111e),
	.w5(32'hbc0093eb),
	.w6(32'hbb92265d),
	.w7(32'hbc0f2eb6),
	.w8(32'hbc1ed8c5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc091867),
	.w1(32'hba8b8955),
	.w2(32'hbc74bb1f),
	.w3(32'h3b781bae),
	.w4(32'hbbb23014),
	.w5(32'h3c4842f8),
	.w6(32'hbbe62f15),
	.w7(32'hbbf92c69),
	.w8(32'h3d0dbbce),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf80e6),
	.w1(32'h393f8ff2),
	.w2(32'h3cd3d3b6),
	.w3(32'hbca146c5),
	.w4(32'h3c2090a2),
	.w5(32'h3a8cebfc),
	.w6(32'h3c89a3cd),
	.w7(32'h3c93daae),
	.w8(32'hbc711e78),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ca807),
	.w1(32'hbbacafd5),
	.w2(32'h3af2bdc0),
	.w3(32'hbb27c1c8),
	.w4(32'h3b04ba68),
	.w5(32'h3a1f114c),
	.w6(32'h3b78ede5),
	.w7(32'h3bcfc1ab),
	.w8(32'hba333afe),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949da83),
	.w1(32'h3ac19dfd),
	.w2(32'hbb71bab4),
	.w3(32'h3b08dedb),
	.w4(32'h3bbee80b),
	.w5(32'hbb38c846),
	.w6(32'h3b200199),
	.w7(32'h3c923dcf),
	.w8(32'hbc89c6c8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0abb7),
	.w1(32'hbaff6d96),
	.w2(32'h3c45db88),
	.w3(32'h3bc19416),
	.w4(32'h38f5699a),
	.w5(32'hbc9618ba),
	.w6(32'h3bbd9d3a),
	.w7(32'h3c633032),
	.w8(32'hbcf874e3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a860cb),
	.w1(32'hbbcc220f),
	.w2(32'h3bfebb84),
	.w3(32'h3b17b27d),
	.w4(32'hbbb7fbf1),
	.w5(32'hba09d708),
	.w6(32'hbbb786b8),
	.w7(32'hbb6e5502),
	.w8(32'hbb83cc3d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68d18a),
	.w1(32'h3a76e3ef),
	.w2(32'hbc7f5fe6),
	.w3(32'h3b8ce2a9),
	.w4(32'h3c56d315),
	.w5(32'hbc2c803f),
	.w6(32'hbb922e1a),
	.w7(32'h3c39a369),
	.w8(32'h3cb0b158),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54097f),
	.w1(32'h3af73389),
	.w2(32'h3aeb2212),
	.w3(32'hbc3880f4),
	.w4(32'h3ac61e44),
	.w5(32'hbaace6a7),
	.w6(32'hbc758928),
	.w7(32'h3c1af84d),
	.w8(32'h399815b1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2013e2),
	.w1(32'h3a9fe0f8),
	.w2(32'hbae6254e),
	.w3(32'h3a56075e),
	.w4(32'hbb1dee16),
	.w5(32'hbbd6e4f8),
	.w6(32'h396ce588),
	.w7(32'hbc5f3d2f),
	.w8(32'h3c076037),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfaf368),
	.w1(32'hbbb6d7c8),
	.w2(32'hbb1d856f),
	.w3(32'h3b99bc67),
	.w4(32'hbc0ad661),
	.w5(32'h3aa38637),
	.w6(32'hbb6bca5a),
	.w7(32'hbc4d0f26),
	.w8(32'hbd10c549),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a4a41),
	.w1(32'h3c1dba5f),
	.w2(32'h3c131aa0),
	.w3(32'h3ccd5ad2),
	.w4(32'h3c25c140),
	.w5(32'h3b90ef7c),
	.w6(32'h3c0c8a21),
	.w7(32'h3c1f7063),
	.w8(32'h3ca9bb99),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d1db3),
	.w1(32'h3beb1b5c),
	.w2(32'h3ad7a294),
	.w3(32'hbb28e0a7),
	.w4(32'h3b730442),
	.w5(32'h3ba066aa),
	.w6(32'h3b1af6b9),
	.w7(32'h3cb561af),
	.w8(32'hbc7d6909),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4e5a4),
	.w1(32'h3bfb0974),
	.w2(32'h39c97ce8),
	.w3(32'hbc09bf64),
	.w4(32'h3aee0ee6),
	.w5(32'h3b81dc5b),
	.w6(32'h3b401978),
	.w7(32'hb9b8c7ff),
	.w8(32'hbc294cc9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule