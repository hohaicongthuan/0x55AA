module layer_8_featuremap_203(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c500905),
	.w1(32'hbb140718),
	.w2(32'hbc3b6b15),
	.w3(32'h3cb31b7e),
	.w4(32'hba28c711),
	.w5(32'hbc2d53a7),
	.w6(32'hbb7b381d),
	.w7(32'h3c05c115),
	.w8(32'h3bd500b1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a046110),
	.w1(32'hbb832d35),
	.w2(32'hbbd261ce),
	.w3(32'hbc00a5ab),
	.w4(32'h3b067ed9),
	.w5(32'h3b2beccb),
	.w6(32'hbb3605b2),
	.w7(32'hbb5eb89b),
	.w8(32'h3ab4d145),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd61805),
	.w1(32'h3b9ee24b),
	.w2(32'hbb8daf3b),
	.w3(32'hb9b2fdd6),
	.w4(32'h3c3f58fd),
	.w5(32'h3beaf023),
	.w6(32'h3ba745db),
	.w7(32'hbb8d09ba),
	.w8(32'h3a7e5f34),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2d111),
	.w1(32'h3c53140d),
	.w2(32'h3bf95532),
	.w3(32'h3c4819c5),
	.w4(32'h3b9c3195),
	.w5(32'h3c0b0e23),
	.w6(32'h3c401665),
	.w7(32'h3c98eb25),
	.w8(32'h3c596eaa),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4a22d),
	.w1(32'h3b1d984d),
	.w2(32'h3c02f44c),
	.w3(32'h3b6ff148),
	.w4(32'hba712ba9),
	.w5(32'h3b85914e),
	.w6(32'h3ad88a02),
	.w7(32'h3c245d71),
	.w8(32'h3c3fa8d2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f050d),
	.w1(32'hb92c6ddb),
	.w2(32'h3bd60ed5),
	.w3(32'hbc39ceaa),
	.w4(32'hbb8e24a0),
	.w5(32'h3a53582b),
	.w6(32'hbbbd408a),
	.w7(32'hbaea5610),
	.w8(32'h3c5b49d6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8bfc),
	.w1(32'h3bace0c5),
	.w2(32'h3c78be36),
	.w3(32'hbb110b0f),
	.w4(32'hbbb59ef9),
	.w5(32'h39cb859f),
	.w6(32'h3bdc3015),
	.w7(32'h3c9a5791),
	.w8(32'h3c610432),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94ad7b),
	.w1(32'h3a8aeb43),
	.w2(32'hbbb87ccd),
	.w3(32'h3c21f9b0),
	.w4(32'h3c8a0cbb),
	.w5(32'h3b9df89a),
	.w6(32'h3a902c0e),
	.w7(32'hbb3f9854),
	.w8(32'h3bee48d4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53110b),
	.w1(32'hbabc4de8),
	.w2(32'hbc35e7a7),
	.w3(32'h3bcefedc),
	.w4(32'h3baf62d1),
	.w5(32'hbb10a390),
	.w6(32'hb9db044a),
	.w7(32'hbb967bbc),
	.w8(32'hbb7d8aa9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10bcff),
	.w1(32'hbc177006),
	.w2(32'hbc2baa18),
	.w3(32'h3acdfeee),
	.w4(32'hbb8418e2),
	.w5(32'hbc0980b3),
	.w6(32'h3bc7c602),
	.w7(32'hbb643992),
	.w8(32'h3bfd11fa),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4689ce),
	.w1(32'h3c059b57),
	.w2(32'h3be9d613),
	.w3(32'h3b40dc2c),
	.w4(32'h3c172e11),
	.w5(32'h3c09034f),
	.w6(32'h3c8ced52),
	.w7(32'h3c985e71),
	.w8(32'h3b2d50f6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86935b),
	.w1(32'h3c2f8e00),
	.w2(32'h3ca6ecfd),
	.w3(32'h39f5e8f6),
	.w4(32'h3b0d7624),
	.w5(32'h3b6e4fc1),
	.w6(32'h3c210248),
	.w7(32'h3cdcbd30),
	.w8(32'h3c7dae73),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb38608),
	.w1(32'h3bbf7463),
	.w2(32'h3b687b26),
	.w3(32'hbc1a95d1),
	.w4(32'hbbe0266a),
	.w5(32'hbc098272),
	.w6(32'h3c323b92),
	.w7(32'h3bee6a9f),
	.w8(32'h3af5e689),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb831c11),
	.w1(32'h3b9b168f),
	.w2(32'hbc19e8ad),
	.w3(32'hbc0e245d),
	.w4(32'h3bac6d55),
	.w5(32'h3c1c7ddd),
	.w6(32'hbb0a3300),
	.w7(32'hbc0e2c40),
	.w8(32'h3c00d31e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd863e),
	.w1(32'h3ac73b93),
	.w2(32'h3b19deca),
	.w3(32'h3b9e7e4d),
	.w4(32'hbb10b60c),
	.w5(32'hbb612b98),
	.w6(32'h3a6c70f9),
	.w7(32'h3a4a7c37),
	.w8(32'hbb56402e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71d3db),
	.w1(32'h3bc8ff93),
	.w2(32'hbbd0a726),
	.w3(32'hbbaf7aaf),
	.w4(32'h3b89e5e6),
	.w5(32'hbb044683),
	.w6(32'h3bb12b80),
	.w7(32'hbb03faa4),
	.w8(32'h3bf4f00b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8683de),
	.w1(32'hbbd98308),
	.w2(32'hbb1ed0c0),
	.w3(32'h3c5db3f3),
	.w4(32'hbc5053c6),
	.w5(32'hbc53a20a),
	.w6(32'h3c81f0e3),
	.w7(32'h3c4d1ed0),
	.w8(32'h39879485),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b983f53),
	.w1(32'h3c2194e5),
	.w2(32'hbc18e49a),
	.w3(32'hb92df01e),
	.w4(32'h3bda82fb),
	.w5(32'h3c827950),
	.w6(32'h3ba759bd),
	.w7(32'hbbf8c977),
	.w8(32'h3b8c18f4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca75556),
	.w1(32'hbba7b014),
	.w2(32'hbc78f227),
	.w3(32'h3cdbd80b),
	.w4(32'h3b7069ee),
	.w5(32'hbb7d14f0),
	.w6(32'hbb051ba4),
	.w7(32'hbc8bbc41),
	.w8(32'hbc294dfb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68ec93),
	.w1(32'hbb1ba1f3),
	.w2(32'hbb8b01da),
	.w3(32'h3c33d67d),
	.w4(32'hbaa78e45),
	.w5(32'hbb6d4983),
	.w6(32'hbc144df8),
	.w7(32'hbc2c46eb),
	.w8(32'hbba05d6e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6bf5d),
	.w1(32'hbb036d1d),
	.w2(32'h3c3b3985),
	.w3(32'hbc1e663b),
	.w4(32'hbbabca17),
	.w5(32'hbbd2f268),
	.w6(32'hbb80686a),
	.w7(32'h3a5b8732),
	.w8(32'hbb60b3ba),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdbc1e),
	.w1(32'hbc0c86a1),
	.w2(32'hbbc87efd),
	.w3(32'hbc820c05),
	.w4(32'hbb88fcf4),
	.w5(32'hbc0d6b41),
	.w6(32'hbbd02ce7),
	.w7(32'hbab0f87b),
	.w8(32'hbbd80787),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8be06f),
	.w1(32'h3c6173a7),
	.w2(32'hbc1eef4b),
	.w3(32'h3cacdbab),
	.w4(32'h3c973db4),
	.w5(32'h3bee3728),
	.w6(32'h3bcb7616),
	.w7(32'h3b550dff),
	.w8(32'hbc548ded),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91038b),
	.w1(32'hbb71cbe6),
	.w2(32'hbb86d90f),
	.w3(32'h3ba06861),
	.w4(32'h3b96ce7d),
	.w5(32'hbb9ebec9),
	.w6(32'h3b210467),
	.w7(32'h3c640971),
	.w8(32'hbb0d3c20),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a868cc3),
	.w1(32'hbb667283),
	.w2(32'hbbd9fa3d),
	.w3(32'h3a665dba),
	.w4(32'hbb1c8155),
	.w5(32'hbbf07417),
	.w6(32'hba0b08ac),
	.w7(32'h3b70b280),
	.w8(32'h3aa79e17),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb279e3e),
	.w1(32'hbbea5b78),
	.w2(32'hbcd164ad),
	.w3(32'h3bd45287),
	.w4(32'h3b79c73a),
	.w5(32'hbc6dba70),
	.w6(32'h3acc6fbb),
	.w7(32'h3bbd66d0),
	.w8(32'hbb6afd0e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d5657),
	.w1(32'hb9b89075),
	.w2(32'hba755234),
	.w3(32'hbc019bbe),
	.w4(32'hbc12e42f),
	.w5(32'hbc3137a9),
	.w6(32'h3c81791d),
	.w7(32'h3caec3ad),
	.w8(32'h3cbccaf7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c79af),
	.w1(32'h3b9e8385),
	.w2(32'hbbda985c),
	.w3(32'h3d0f5755),
	.w4(32'h3d8559fc),
	.w5(32'h3d691aee),
	.w6(32'hbbff8450),
	.w7(32'h3c43a394),
	.w8(32'hbcadb9e4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fc1ee4),
	.w1(32'hbb825719),
	.w2(32'h3ab55086),
	.w3(32'h3b853f77),
	.w4(32'h3b8c7408),
	.w5(32'h3b574868),
	.w6(32'hbb25be05),
	.w7(32'h3c497173),
	.w8(32'h3acf8c55),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5e3da),
	.w1(32'h3bbc0ce5),
	.w2(32'h3c0ce2d6),
	.w3(32'hbb6b0338),
	.w4(32'hbc3ee1f0),
	.w5(32'hbc4786ba),
	.w6(32'h3b872db2),
	.w7(32'h3c066708),
	.w8(32'h3c925f83),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68d3dd),
	.w1(32'h3b880376),
	.w2(32'h3bc0854d),
	.w3(32'hbba7856f),
	.w4(32'h3be436ae),
	.w5(32'h3bcd6f45),
	.w6(32'h3bf185ec),
	.w7(32'h3c3bc7ba),
	.w8(32'h3c423c27),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abef39c),
	.w1(32'hbc49f89e),
	.w2(32'hbc67ae78),
	.w3(32'h3b95e592),
	.w4(32'hbbd87e96),
	.w5(32'hbbbecd6b),
	.w6(32'hbc7d5c27),
	.w7(32'hbc923b4a),
	.w8(32'hbbdb47d5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a00d),
	.w1(32'h37e0753b),
	.w2(32'hbc5193b3),
	.w3(32'hbbb3a7c2),
	.w4(32'h3c2304a8),
	.w5(32'h3c61d24f),
	.w6(32'hba3fd92f),
	.w7(32'hbc946ec7),
	.w8(32'hbc372334),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeeb17d),
	.w1(32'hbc165d1e),
	.w2(32'h3ba2ae5d),
	.w3(32'h3b8d3d65),
	.w4(32'hbc01f873),
	.w5(32'hbacf7cb5),
	.w6(32'hba8e1e51),
	.w7(32'h3bd894e1),
	.w8(32'h3c4a8ce3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc28af4),
	.w1(32'hbb8bdd26),
	.w2(32'hbc0645a1),
	.w3(32'hbbea6857),
	.w4(32'hbaab1021),
	.w5(32'hbb24e339),
	.w6(32'hbbc86a5b),
	.w7(32'hbc4c47a2),
	.w8(32'hbc3a21e9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83fb64),
	.w1(32'hba8be860),
	.w2(32'h3b3500b4),
	.w3(32'h3bea618b),
	.w4(32'h3c003656),
	.w5(32'h3c309b0f),
	.w6(32'h3baf3fe7),
	.w7(32'h3bba7ca4),
	.w8(32'hbb71886c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6e23e),
	.w1(32'hbb47721e),
	.w2(32'hb83b203d),
	.w3(32'h3b1fb9a6),
	.w4(32'hbb5fdb34),
	.w5(32'hbb753853),
	.w6(32'hba11901b),
	.w7(32'h3aab5c0c),
	.w8(32'h3b2bde69),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19475d),
	.w1(32'hb973d961),
	.w2(32'hbb9ff80a),
	.w3(32'hba96d4bd),
	.w4(32'h3bc97c84),
	.w5(32'h3beeb73c),
	.w6(32'hbc2e56b9),
	.w7(32'hbc9b0bc2),
	.w8(32'hbc8047ee),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf40bd4),
	.w1(32'h3ac8b5f6),
	.w2(32'h3af868a3),
	.w3(32'h39e0a3c3),
	.w4(32'h3bd4b6ef),
	.w5(32'hbb2049d0),
	.w6(32'h3a00c8fa),
	.w7(32'h3be35a7b),
	.w8(32'h3acef683),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916afd3),
	.w1(32'h3b3a67ec),
	.w2(32'h3c468351),
	.w3(32'hbb852f7f),
	.w4(32'hb9d4cfd0),
	.w5(32'hbb13cab5),
	.w6(32'h3af5ec30),
	.w7(32'h3c39d89a),
	.w8(32'h3c367eb6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c854ec6),
	.w1(32'h3c1eb403),
	.w2(32'h3b96634f),
	.w3(32'h3c5d1356),
	.w4(32'h3cbd17c9),
	.w5(32'h3cc7a041),
	.w6(32'h3bdfad58),
	.w7(32'h3a143121),
	.w8(32'h3c930155),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2f0f0),
	.w1(32'hbabb11d6),
	.w2(32'hbbf55f51),
	.w3(32'h3b22aca2),
	.w4(32'h3b823a63),
	.w5(32'hbba19a9e),
	.w6(32'h38d4c92e),
	.w7(32'hba987410),
	.w8(32'h3c08337e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd5acd),
	.w1(32'hbc177c6d),
	.w2(32'hbb34d504),
	.w3(32'hba8712b4),
	.w4(32'hb9edcaca),
	.w5(32'h38c6046f),
	.w6(32'hbc36d370),
	.w7(32'hbaa9c32c),
	.w8(32'hbb43c8ed),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc134f),
	.w1(32'h3c1bfb11),
	.w2(32'h3ba2abcd),
	.w3(32'h3c2c543b),
	.w4(32'h3b76f1db),
	.w5(32'h3b2e31af),
	.w6(32'h3b0790ca),
	.w7(32'h38b93d44),
	.w8(32'h3baf3024),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed7758),
	.w1(32'hba51198e),
	.w2(32'hbc25910b),
	.w3(32'h3c0e12d5),
	.w4(32'hbaf7085a),
	.w5(32'hbbed143e),
	.w6(32'h3bda8a2f),
	.w7(32'hbb94302d),
	.w8(32'hbc919473),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44f890),
	.w1(32'hbb2efc2c),
	.w2(32'hbb722549),
	.w3(32'hbb925382),
	.w4(32'hbbd6bc46),
	.w5(32'hbbf775ff),
	.w6(32'h3b999273),
	.w7(32'h3b00c3dc),
	.w8(32'h3a8cae15),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e6152),
	.w1(32'h3aa1b281),
	.w2(32'h3cdd6224),
	.w3(32'hbaa3f9df),
	.w4(32'hbc99cabe),
	.w5(32'hbc5286f9),
	.w6(32'h3c98514d),
	.w7(32'h3d52cf9d),
	.w8(32'h3d37e720),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d035691),
	.w1(32'h3bc27649),
	.w2(32'h3b77bbf9),
	.w3(32'hbadd65f1),
	.w4(32'h3c0726c6),
	.w5(32'hbb95042c),
	.w6(32'h3b0c1bec),
	.w7(32'hba7110b0),
	.w8(32'hbc18cdc9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c186e05),
	.w1(32'h3c08dd1f),
	.w2(32'hbac3ea42),
	.w3(32'h3bef0144),
	.w4(32'h3c14454a),
	.w5(32'h3bbfdf5c),
	.w6(32'h3aa1c0f4),
	.w7(32'h3a3a070a),
	.w8(32'hbc37d4d3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0453c8),
	.w1(32'hbb16e3be),
	.w2(32'hbb008673),
	.w3(32'h3c2a1ebc),
	.w4(32'h3c1c6039),
	.w5(32'h3bed6a1b),
	.w6(32'h388ec83d),
	.w7(32'hb95ba911),
	.w8(32'hbaa971bd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90dd23),
	.w1(32'hbbf76b1f),
	.w2(32'h3b3a9237),
	.w3(32'hbb56d5e4),
	.w4(32'hbbb5a4c1),
	.w5(32'h3b3326bc),
	.w6(32'hbc59ac60),
	.w7(32'hbb98a85f),
	.w8(32'hbb8d705c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc907b23),
	.w1(32'hbc55b022),
	.w2(32'hbc954992),
	.w3(32'h3c946fee),
	.w4(32'h3c6cef93),
	.w5(32'h3ac98b75),
	.w6(32'hbbe4e911),
	.w7(32'hbbfb7de4),
	.w8(32'hbc0a7a3e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84f6cc),
	.w1(32'h3afa93a0),
	.w2(32'h3ae918ee),
	.w3(32'h3b8c5f78),
	.w4(32'h3c0edbc3),
	.w5(32'h3c0e4394),
	.w6(32'hba97f901),
	.w7(32'h3ac0f150),
	.w8(32'hbb0a1e33),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59bd3a),
	.w1(32'h3c632f07),
	.w2(32'h3c52cb99),
	.w3(32'h3c213835),
	.w4(32'h3c6320e3),
	.w5(32'h3adb7903),
	.w6(32'h3b941d4f),
	.w7(32'hbb3eda78),
	.w8(32'hba366bc3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c008d86),
	.w1(32'h3a01633b),
	.w2(32'hbc64ff57),
	.w3(32'h3b8b61a0),
	.w4(32'h3bc95abe),
	.w5(32'h3b214cdf),
	.w6(32'hbba07bea),
	.w7(32'hbc4e6f15),
	.w8(32'hbbd9f3f9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0c1a8),
	.w1(32'h3b90cc87),
	.w2(32'hbaa89753),
	.w3(32'h3b899b9e),
	.w4(32'h3b4d38a5),
	.w5(32'hba2163ce),
	.w6(32'h3b541ffb),
	.w7(32'h3ac3c6e9),
	.w8(32'hbae7bbdf),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04fd92),
	.w1(32'h3bb0b147),
	.w2(32'hbba1607c),
	.w3(32'h3b9042fd),
	.w4(32'hb982634a),
	.w5(32'hba12e82c),
	.w6(32'h3be9e689),
	.w7(32'h3c46ee4d),
	.w8(32'hbc45c31a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c8ee6),
	.w1(32'hbc158871),
	.w2(32'hbc1b1bbc),
	.w3(32'h3c4dad33),
	.w4(32'h3b26ddfc),
	.w5(32'hbaedb56c),
	.w6(32'hba95f018),
	.w7(32'hbbaa9bd6),
	.w8(32'hbb507e57),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c6363),
	.w1(32'h3b479af0),
	.w2(32'h3b835ac8),
	.w3(32'h3b918cad),
	.w4(32'h3afed2e4),
	.w5(32'h3b5af4fb),
	.w6(32'h3ba635fb),
	.w7(32'h3bbfe693),
	.w8(32'h3acbc711),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb9397),
	.w1(32'h3b735e8f),
	.w2(32'h3c00ebda),
	.w3(32'h3ae092ee),
	.w4(32'h3c1632e2),
	.w5(32'h3c1de3f7),
	.w6(32'h3bc3281a),
	.w7(32'h3c234d6a),
	.w8(32'h3aac6ad9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1eb849),
	.w1(32'hba2205b1),
	.w2(32'hbbd9e6b9),
	.w3(32'h3c0735a9),
	.w4(32'h3b0186c0),
	.w5(32'hbc260d0d),
	.w6(32'h3b20f428),
	.w7(32'h3a8173d7),
	.w8(32'h3b1f62cc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc50012),
	.w1(32'h3b2878cd),
	.w2(32'h3bcf64fd),
	.w3(32'hba2edf36),
	.w4(32'hba952a1e),
	.w5(32'hbafeb88a),
	.w6(32'h3b280142),
	.w7(32'h3c284ca6),
	.w8(32'h3be83e7d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6aa92a),
	.w1(32'hbb631061),
	.w2(32'hbad6a20e),
	.w3(32'h3c5424dc),
	.w4(32'h3c3206be),
	.w5(32'h3c9cbde7),
	.w6(32'hbc56a270),
	.w7(32'hbc93cff7),
	.w8(32'hbb028381),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b752b37),
	.w1(32'h3bd0374d),
	.w2(32'h3a60002c),
	.w3(32'h3c348480),
	.w4(32'h3b8c2d4f),
	.w5(32'h3aa870eb),
	.w6(32'h3c564a6c),
	.w7(32'h3c09a8a1),
	.w8(32'h3bc9427a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc1e08),
	.w1(32'h3ad2746c),
	.w2(32'h3ac0b77d),
	.w3(32'hb70d4405),
	.w4(32'h3b0c6122),
	.w5(32'h3b7a7c70),
	.w6(32'h39d71d9d),
	.w7(32'hbae4b9c7),
	.w8(32'h398d7df4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ae55f),
	.w1(32'hb99fd890),
	.w2(32'h3b83b387),
	.w3(32'h3b893c2a),
	.w4(32'hbb14c526),
	.w5(32'hbafc35f1),
	.w6(32'h3bf0f9c5),
	.w7(32'h3c3c1d70),
	.w8(32'h3b78aec5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa7a54),
	.w1(32'h3a41f81e),
	.w2(32'h3c246ec9),
	.w3(32'hbbba846f),
	.w4(32'hbba014d1),
	.w5(32'hb984ea98),
	.w6(32'h3c463d94),
	.w7(32'h3c8e81b5),
	.w8(32'h3c5909c2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ebc76),
	.w1(32'hbb70e230),
	.w2(32'h3c3b48c0),
	.w3(32'hbc43ecf9),
	.w4(32'hbc8f4889),
	.w5(32'hbc9aa5a8),
	.w6(32'h3c4aaa21),
	.w7(32'h3c984d75),
	.w8(32'h3c6cc10d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c1755),
	.w1(32'h3b92f66c),
	.w2(32'hbbba77b9),
	.w3(32'hbc3c2b40),
	.w4(32'h3c040b9d),
	.w5(32'hba91bde8),
	.w6(32'h3bbb8a5e),
	.w7(32'hbb0eead0),
	.w8(32'h3bc0070d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc81185),
	.w1(32'h3c8364d0),
	.w2(32'hbbafdd4c),
	.w3(32'h3cd3f0fe),
	.w4(32'h3d09e3d9),
	.w5(32'h3d063e65),
	.w6(32'h3ba13614),
	.w7(32'hbc46c42b),
	.w8(32'hbcc9d46e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab228d8),
	.w1(32'hbac1ffdf),
	.w2(32'hbb8a9226),
	.w3(32'h3c8d3d7a),
	.w4(32'hbb1bb07d),
	.w5(32'hbbae7a0f),
	.w6(32'hbb8d1322),
	.w7(32'hbab36643),
	.w8(32'hbb19d66f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152478),
	.w1(32'h3c156264),
	.w2(32'h3c7ee2cc),
	.w3(32'h3abe00e8),
	.w4(32'h3c376185),
	.w5(32'h3c812d8c),
	.w6(32'h3c40d542),
	.w7(32'h3c1888fa),
	.w8(32'h3c7643ea),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3eb26a),
	.w1(32'h3bc091c2),
	.w2(32'h3b8c790c),
	.w3(32'h3ae8a3ce),
	.w4(32'h3b4dabbc),
	.w5(32'h39224cad),
	.w6(32'h3b066396),
	.w7(32'h39406d0f),
	.w8(32'h3b341e9f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ce102),
	.w1(32'hbb869c63),
	.w2(32'hbb7af775),
	.w3(32'h3c13c3e4),
	.w4(32'hba2f403e),
	.w5(32'hb8cc60fe),
	.w6(32'hbb454815),
	.w7(32'hbb145413),
	.w8(32'hbbc7f4c6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e9706),
	.w1(32'h3b61a9a2),
	.w2(32'h3728ffec),
	.w3(32'hba111b46),
	.w4(32'h3b06c9c6),
	.w5(32'hbc0105cf),
	.w6(32'hbb45d216),
	.w7(32'h3bd7aea0),
	.w8(32'h3b0e1a6a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bda19),
	.w1(32'h3bbea24c),
	.w2(32'h3bf4aa66),
	.w3(32'hbc497ca6),
	.w4(32'h3c5aa6e8),
	.w5(32'h3c862d8c),
	.w6(32'hbc406238),
	.w7(32'hbc03ba05),
	.w8(32'hbc0d7940),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb02ee),
	.w1(32'h3aa38a76),
	.w2(32'hbad00aa8),
	.w3(32'h3bb17c2d),
	.w4(32'hbac0a34a),
	.w5(32'hbb0d878e),
	.w6(32'hbbcc79be),
	.w7(32'hbb0aef11),
	.w8(32'hbbbc05f7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19a9c2),
	.w1(32'h3ba4f876),
	.w2(32'h3be4d3d0),
	.w3(32'h3c3f29af),
	.w4(32'h3c38d1dd),
	.w5(32'h3c022e2e),
	.w6(32'hbb63ac85),
	.w7(32'h3bef0558),
	.w8(32'h39f2b88d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1599d3),
	.w1(32'hbc031a24),
	.w2(32'hbc455d98),
	.w3(32'h3c2549eb),
	.w4(32'h39e294f3),
	.w5(32'hbb4742c3),
	.w6(32'hbadb5f32),
	.w7(32'hbc28ee6f),
	.w8(32'hbbcf2a68),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04f05b),
	.w1(32'h3b9c1955),
	.w2(32'h3acc965e),
	.w3(32'h3b79920d),
	.w4(32'h3c2c2f61),
	.w5(32'h3b543eca),
	.w6(32'h3a29537f),
	.w7(32'h3a850f41),
	.w8(32'h3bf98158),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b6338),
	.w1(32'h3b3c45b8),
	.w2(32'hbc2d689f),
	.w3(32'h3b9ae660),
	.w4(32'h3c5cf258),
	.w5(32'h3c2ba9dd),
	.w6(32'h3aff2398),
	.w7(32'hbc08a1e9),
	.w8(32'hba218bc0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b1355),
	.w1(32'h3ab208a8),
	.w2(32'hbb357ac7),
	.w3(32'h3c55e82f),
	.w4(32'h3ba84723),
	.w5(32'h3c014643),
	.w6(32'h3a5a89f8),
	.w7(32'h3bca438d),
	.w8(32'h3bd1a5b4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a69195),
	.w1(32'h3bda642a),
	.w2(32'h3b0e3dda),
	.w3(32'h3bcdfe30),
	.w4(32'h3cb13539),
	.w5(32'h3c950f3a),
	.w6(32'h3b9e8dde),
	.w7(32'hbc4f4155),
	.w8(32'hbc2b2932),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87bc37),
	.w1(32'h3c94826c),
	.w2(32'h3cc1ba33),
	.w3(32'h3cc754d2),
	.w4(32'h3c91e47a),
	.w5(32'h3cb59d51),
	.w6(32'h3c8e0032),
	.w7(32'h3cce6533),
	.w8(32'h3d06765c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c267df5),
	.w1(32'h3c5376e7),
	.w2(32'hbc311a7c),
	.w3(32'h3ccda273),
	.w4(32'h3d26f9f7),
	.w5(32'h3cf911d1),
	.w6(32'h3c064510),
	.w7(32'hbbe6202e),
	.w8(32'h3bb0b8a1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc094a99),
	.w1(32'h3b9a96da),
	.w2(32'h3a05c029),
	.w3(32'h3ca6a114),
	.w4(32'h3c1133aa),
	.w5(32'h3b5e35ca),
	.w6(32'h3bd490c5),
	.w7(32'h3c5c1f24),
	.w8(32'h3c485d38),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7a4f1),
	.w1(32'hbbff1207),
	.w2(32'hbc350de9),
	.w3(32'h39df22ba),
	.w4(32'hbb4b029d),
	.w5(32'hbb7be3b3),
	.w6(32'hbbb10705),
	.w7(32'hbbef3b5c),
	.w8(32'hbb570bb1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd420e9),
	.w1(32'hbc10be42),
	.w2(32'hbbbcfaae),
	.w3(32'hbb9ed3ea),
	.w4(32'hbc06a5fd),
	.w5(32'hbc161892),
	.w6(32'hbbdb2ec7),
	.w7(32'hbc261f89),
	.w8(32'hbc08b07a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17e6b7),
	.w1(32'hb9376722),
	.w2(32'hbb8fbc8e),
	.w3(32'hbc023e17),
	.w4(32'hba1ebe75),
	.w5(32'hbbd103f8),
	.w6(32'h3b8837a3),
	.w7(32'h3b92795e),
	.w8(32'h3b8bb753),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50e6f8),
	.w1(32'h3c03ba0f),
	.w2(32'h3bac2e1e),
	.w3(32'hbb07f726),
	.w4(32'h3c7b8f28),
	.w5(32'h3caccd5e),
	.w6(32'h3c374895),
	.w7(32'h3b2f4052),
	.w8(32'h3bd3a471),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cd31d),
	.w1(32'h3b1e797c),
	.w2(32'h3bb1bbc0),
	.w3(32'h3cb02342),
	.w4(32'hbb6df07e),
	.w5(32'hbae2bcd9),
	.w6(32'hbb703045),
	.w7(32'h3c0bf022),
	.w8(32'h3bce1a4b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c7733),
	.w1(32'hba21ff66),
	.w2(32'h3bf52a2e),
	.w3(32'h3b2ff2b7),
	.w4(32'hbc267767),
	.w5(32'hbb1745fb),
	.w6(32'h3adf6ade),
	.w7(32'h3cb34913),
	.w8(32'h3c16f0c6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2e999),
	.w1(32'hbb24daab),
	.w2(32'h3a5ad2dd),
	.w3(32'h3a85730f),
	.w4(32'h3ae70598),
	.w5(32'h3be47e78),
	.w6(32'h3a231406),
	.w7(32'h3b225aaf),
	.w8(32'h3bda4327),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231ac5),
	.w1(32'hba3826af),
	.w2(32'h3aa2b07b),
	.w3(32'h3b989035),
	.w4(32'hba9e8d7b),
	.w5(32'hb81e8ab6),
	.w6(32'h3b10cbe3),
	.w7(32'h3c239eda),
	.w8(32'h3c341415),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2410b8),
	.w1(32'hbc0b45c5),
	.w2(32'h397e17c4),
	.w3(32'hbb4579c3),
	.w4(32'hbbdf84c0),
	.w5(32'hbc0f276e),
	.w6(32'hbbc72d1d),
	.w7(32'hbb6377dc),
	.w8(32'h3bd09aa0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee6cc5),
	.w1(32'hbbfa2e9f),
	.w2(32'hbc3aa5c3),
	.w3(32'hbb6a8aae),
	.w4(32'hbb804aba),
	.w5(32'hbc2ee219),
	.w6(32'hbc01a51f),
	.w7(32'hbbe9ecf4),
	.w8(32'hbc24a3af),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73cbd4),
	.w1(32'h3bcb6d07),
	.w2(32'h3bdbed3f),
	.w3(32'h39e08557),
	.w4(32'h3ca69458),
	.w5(32'h3c9a556a),
	.w6(32'hbbc7c80e),
	.w7(32'hbc7fbc78),
	.w8(32'hbb34718a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8f50e),
	.w1(32'h3c19f64c),
	.w2(32'h3c59391f),
	.w3(32'h3c7d1981),
	.w4(32'h3c2fbf66),
	.w5(32'h3c3e12a4),
	.w6(32'h3ba3171a),
	.w7(32'h3c3aa722),
	.w8(32'hbb6b0d34),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95bfdc),
	.w1(32'h3b7a43cf),
	.w2(32'h3bce491c),
	.w3(32'h3be2fe06),
	.w4(32'hbb644305),
	.w5(32'hbba141d0),
	.w6(32'hb9c6d754),
	.w7(32'h3c38b80e),
	.w8(32'h3b652abd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb40d2),
	.w1(32'hbad1e760),
	.w2(32'hba276f1c),
	.w3(32'hbb0fe4f7),
	.w4(32'h3b2e11d7),
	.w5(32'h3ba756b7),
	.w6(32'h3bffba40),
	.w7(32'h3c12fd75),
	.w8(32'h3c27dfb4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad35c26),
	.w1(32'h3b221efd),
	.w2(32'h3c82e1eb),
	.w3(32'h3a5b7412),
	.w4(32'hbb241021),
	.w5(32'h3bdc8681),
	.w6(32'h3b979a79),
	.w7(32'h3c3a8185),
	.w8(32'h3bc9a91c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91171c),
	.w1(32'hbb30824e),
	.w2(32'hbb64c94b),
	.w3(32'hbb4deb8e),
	.w4(32'hbb06f27f),
	.w5(32'hbb94205d),
	.w6(32'h3bbba88b),
	.w7(32'hb9d3ecf5),
	.w8(32'h3bb8a206),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8b264),
	.w1(32'hbbd31324),
	.w2(32'h3b80ca8e),
	.w3(32'hbb759f04),
	.w4(32'hbac27796),
	.w5(32'hbb14390d),
	.w6(32'hbb7536d3),
	.w7(32'h3bd14e54),
	.w8(32'h3b91a366),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b98c84),
	.w1(32'hbbe1b26a),
	.w2(32'hbc850f49),
	.w3(32'h3acbd512),
	.w4(32'hbb148b87),
	.w5(32'hbb08ed61),
	.w6(32'h3aff23d8),
	.w7(32'hbbbb2e8b),
	.w8(32'hbc268a20),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32da93),
	.w1(32'h3b833588),
	.w2(32'h3bd9b3a2),
	.w3(32'hbc09ce65),
	.w4(32'hbaa6a19e),
	.w5(32'h39bfdf1d),
	.w6(32'h3c434903),
	.w7(32'h3c43ea45),
	.w8(32'h3ba29c22),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba05fbd),
	.w1(32'h3b004005),
	.w2(32'h39b74756),
	.w3(32'h3c6aeb8f),
	.w4(32'h3bd523a5),
	.w5(32'h3ba147f1),
	.w6(32'h3bcc9e61),
	.w7(32'h3b65172d),
	.w8(32'hbba900f6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde6778),
	.w1(32'hba60198a),
	.w2(32'hbbf260f1),
	.w3(32'h3af19855),
	.w4(32'h3ae7aca6),
	.w5(32'hbb3089ab),
	.w6(32'hbb34daff),
	.w7(32'hbb114364),
	.w8(32'h38aa96b1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ef411),
	.w1(32'hbb8de505),
	.w2(32'hbb4de4f8),
	.w3(32'hbb1d7048),
	.w4(32'h3bb815ae),
	.w5(32'h3a305ee8),
	.w6(32'hbbad1afd),
	.w7(32'hbad61187),
	.w8(32'h3b656adf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd97a94),
	.w1(32'h3bf017cf),
	.w2(32'h3d0ef743),
	.w3(32'hb9dc08ce),
	.w4(32'h3b1aba3e),
	.w5(32'h3c84a839),
	.w6(32'h3bed4dd5),
	.w7(32'h3d03548f),
	.w8(32'h3cfaa88d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d04474c),
	.w1(32'h3b782729),
	.w2(32'h3b8c6387),
	.w3(32'h3c6b533a),
	.w4(32'h3bf41604),
	.w5(32'h3c32a284),
	.w6(32'hba858766),
	.w7(32'h37e95d8d),
	.w8(32'h3b08980f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d8712),
	.w1(32'hbc0bdebe),
	.w2(32'h3b464fea),
	.w3(32'h3919a960),
	.w4(32'hbc1646a0),
	.w5(32'hbc39ea14),
	.w6(32'hbc4c51dc),
	.w7(32'hbc1d1867),
	.w8(32'h3bff3707),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30185a),
	.w1(32'hbbce2e32),
	.w2(32'hbb14a499),
	.w3(32'hbc13c391),
	.w4(32'hbbf609c3),
	.w5(32'hba3a0caa),
	.w6(32'hbb49e2fe),
	.w7(32'h3a8ba0b2),
	.w8(32'h3bcecfdd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d2e26),
	.w1(32'h3c174937),
	.w2(32'h3c008f0a),
	.w3(32'hbba2e9a0),
	.w4(32'h3c3944de),
	.w5(32'h3b597996),
	.w6(32'h3c208fa6),
	.w7(32'h3c2fb577),
	.w8(32'h3c89aa5c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c097041),
	.w1(32'h3b5aa96d),
	.w2(32'hb9bea0c2),
	.w3(32'h3bd3c07f),
	.w4(32'hbb27e67e),
	.w5(32'hbb7f1ae0),
	.w6(32'h3c5986fc),
	.w7(32'h3c177a9f),
	.w8(32'h3c0ae67c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95d877),
	.w1(32'hbae8ccad),
	.w2(32'hbbfc3622),
	.w3(32'h3ace12ca),
	.w4(32'h3b2f6408),
	.w5(32'hbaf0990c),
	.w6(32'hba095118),
	.w7(32'hba4bcc3a),
	.w8(32'h3b99bfea),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac00c20),
	.w1(32'h3b481327),
	.w2(32'h3a8f499d),
	.w3(32'h3abb5e8f),
	.w4(32'h3bb25f80),
	.w5(32'h3bdd062d),
	.w6(32'hba636149),
	.w7(32'hbb5b0fa6),
	.w8(32'hbb0180c8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb514435),
	.w1(32'hbbc8d839),
	.w2(32'hbc09fccc),
	.w3(32'h3b3a2a4c),
	.w4(32'h3981e2d6),
	.w5(32'h3b0ebd76),
	.w6(32'hbbebcc81),
	.w7(32'hbc36a03a),
	.w8(32'hbc102358),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b54ed),
	.w1(32'h3b7c27b5),
	.w2(32'h3b5beb20),
	.w3(32'h3bab2c5b),
	.w4(32'hb97c82ce),
	.w5(32'h3c0cf807),
	.w6(32'h3ba3e74c),
	.w7(32'h3a799197),
	.w8(32'h3b653797),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce02b0),
	.w1(32'hba82bc6f),
	.w2(32'h3ba8e631),
	.w3(32'h3c151a62),
	.w4(32'h3b887772),
	.w5(32'h3ad31a85),
	.w6(32'h3c126f0e),
	.w7(32'h3acdcc64),
	.w8(32'h3c0e4d21),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23944e),
	.w1(32'hbb0da95c),
	.w2(32'hbba1f460),
	.w3(32'h3c15dbc4),
	.w4(32'h39a6f287),
	.w5(32'hbb90a137),
	.w6(32'hbae14c07),
	.w7(32'hb9e43a9f),
	.w8(32'h392c2406),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf83ec),
	.w1(32'hb9d19f56),
	.w2(32'hbc3b4c38),
	.w3(32'h3aeb1430),
	.w4(32'hb9425f01),
	.w5(32'h3b371dd5),
	.w6(32'hbb2e9ec6),
	.w7(32'h3b72d801),
	.w8(32'h3c01beab),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa65ac),
	.w1(32'hbbd651ae),
	.w2(32'hbc42f893),
	.w3(32'hba5fc29d),
	.w4(32'hbbcb7d8a),
	.w5(32'hbb134474),
	.w6(32'hbc1edff5),
	.w7(32'hbc751e2b),
	.w8(32'hbc15a301),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40a29e),
	.w1(32'hbb842188),
	.w2(32'h3888e5bc),
	.w3(32'hbbb8c804),
	.w4(32'hbbd7f877),
	.w5(32'hbb3ebd1d),
	.w6(32'h3b256159),
	.w7(32'h3c0bd525),
	.w8(32'h3c256c39),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e01e93),
	.w1(32'h3c09cf21),
	.w2(32'h3bdc942d),
	.w3(32'hbb157e2e),
	.w4(32'h3b370829),
	.w5(32'h3c375b0d),
	.w6(32'h3c566ef7),
	.w7(32'h3bcc91f5),
	.w8(32'h3b8f7382),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7964e),
	.w1(32'hbae7e50a),
	.w2(32'h3a8fffa1),
	.w3(32'h3b95717d),
	.w4(32'hbacb938f),
	.w5(32'h3c1cdace),
	.w6(32'hbbc6f7ed),
	.w7(32'hbc4197d6),
	.w8(32'h3b269e75),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb48c37),
	.w1(32'hbb980de5),
	.w2(32'h3c14efd2),
	.w3(32'h3bbec2fb),
	.w4(32'h3b23a3e1),
	.w5(32'hb8d757dc),
	.w6(32'h3bcdf308),
	.w7(32'h3b38f059),
	.w8(32'hbbf30fb9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e79ad),
	.w1(32'hbbcfa3ec),
	.w2(32'hbc03d617),
	.w3(32'h3b95c1d0),
	.w4(32'hba4b0bd9),
	.w5(32'hbb866ca2),
	.w6(32'hba3649f3),
	.w7(32'hbb6c55f1),
	.w8(32'h39f5fd1d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9e417),
	.w1(32'hbd42b7db),
	.w2(32'hbd87d2b3),
	.w3(32'h3b39d2b0),
	.w4(32'hbd3245b5),
	.w5(32'hbd5ac33c),
	.w6(32'hbcc0520b),
	.w7(32'hbd26201c),
	.w8(32'hbcf58e68),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule