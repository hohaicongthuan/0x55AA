module layer_10_featuremap_162(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8025aa),
	.w1(32'h3b6a238f),
	.w2(32'h3b065eb9),
	.w3(32'h3a823f3e),
	.w4(32'h3bdfc846),
	.w5(32'h3bd8d2ec),
	.w6(32'h3a372f79),
	.w7(32'hbad91772),
	.w8(32'hbbed5c79),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c813f),
	.w1(32'h3c00d29b),
	.w2(32'h3c19a249),
	.w3(32'hba846472),
	.w4(32'h3bbc44f4),
	.w5(32'h3c0e7573),
	.w6(32'hb9ffa541),
	.w7(32'h3ba2eece),
	.w8(32'h3ad5e5cd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfecfcf),
	.w1(32'h3a74f4cd),
	.w2(32'h3adb9771),
	.w3(32'h3ba2066d),
	.w4(32'hbb012325),
	.w5(32'hb7ace10c),
	.w6(32'hbb36c343),
	.w7(32'hbae33017),
	.w8(32'hbadc1f00),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace6cc9),
	.w1(32'hbb29fefc),
	.w2(32'hbb961388),
	.w3(32'hba5d2ed8),
	.w4(32'hb934263e),
	.w5(32'hbb6617be),
	.w6(32'h3b988c55),
	.w7(32'h3baab8d6),
	.w8(32'h3b8afd13),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa3fb2),
	.w1(32'h3add47df),
	.w2(32'h3be781fd),
	.w3(32'hbb013fb0),
	.w4(32'h39d47392),
	.w5(32'h3be89d90),
	.w6(32'h3b1cbbf3),
	.w7(32'h3bca8c91),
	.w8(32'h3c19a86c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ca226),
	.w1(32'hb7bf493b),
	.w2(32'h3aa3f27b),
	.w3(32'h3c50fae7),
	.w4(32'h3aafe296),
	.w5(32'h3b092e09),
	.w6(32'h3ad543a0),
	.w7(32'h3afbf83a),
	.w8(32'h3b536318),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba066aa),
	.w1(32'h3bc95dcb),
	.w2(32'h3bd58d71),
	.w3(32'h3bc4bf90),
	.w4(32'h3b86a887),
	.w5(32'h3be7bb84),
	.w6(32'hbaef9f35),
	.w7(32'h3aca82bc),
	.w8(32'h3afe295e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff6f92),
	.w1(32'hbc5ad159),
	.w2(32'hbc7f2d1c),
	.w3(32'h3b856f70),
	.w4(32'hbc38a290),
	.w5(32'hbc4bc776),
	.w6(32'hbc1ab818),
	.w7(32'hbc4eafb3),
	.w8(32'hbc0f8b7c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8b179),
	.w1(32'h3a87e189),
	.w2(32'h3a54cf16),
	.w3(32'hbbb1c3eb),
	.w4(32'h3af3f1f7),
	.w5(32'h3aa1b19d),
	.w6(32'h3a9ef485),
	.w7(32'h3a1c5760),
	.w8(32'h3a900daf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba498d9),
	.w1(32'h3b67f802),
	.w2(32'hba1c375c),
	.w3(32'hbb08486b),
	.w4(32'h3ae0adb6),
	.w5(32'hbaf09820),
	.w6(32'hbc0bd8e8),
	.w7(32'h392cf55d),
	.w8(32'hbbdef75c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c191c5d),
	.w1(32'h394c073d),
	.w2(32'hbad73ee8),
	.w3(32'h3c05d757),
	.w4(32'h3b13ef57),
	.w5(32'h3a5829e9),
	.w6(32'h3af3cb59),
	.w7(32'hb7aaf738),
	.w8(32'h39532136),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7917ac),
	.w1(32'h3a7a369b),
	.w2(32'hba256afa),
	.w3(32'hbb13136c),
	.w4(32'h3902c3e1),
	.w5(32'hbb2dee21),
	.w6(32'hbc14eb8c),
	.w7(32'hb9d3c151),
	.w8(32'hbb8fb97f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc467025),
	.w1(32'hbc0604e8),
	.w2(32'hbc69a959),
	.w3(32'hbc3ef5a7),
	.w4(32'hbbb2008a),
	.w5(32'hbc4742f4),
	.w6(32'hbc0e7857),
	.w7(32'hbbd920d3),
	.w8(32'hbbfbebb6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ca2e4),
	.w1(32'hbceb566a),
	.w2(32'hbcf9d95b),
	.w3(32'h3ad69531),
	.w4(32'hbcd63ff5),
	.w5(32'hbcf1e988),
	.w6(32'hbcbd3d3c),
	.w7(32'hbccf0714),
	.w8(32'hbccdbc83),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcecab62),
	.w1(32'h3a8ba31c),
	.w2(32'hba9c55e1),
	.w3(32'hbce05eb7),
	.w4(32'hbb2e7886),
	.w5(32'hbb177441),
	.w6(32'hbb342d16),
	.w7(32'h3b0723fc),
	.w8(32'h3a0830d6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f195b),
	.w1(32'hbb135c8d),
	.w2(32'hbbe72762),
	.w3(32'hbb2ce952),
	.w4(32'hba1e77a8),
	.w5(32'hbbb83054),
	.w6(32'hbb81a6be),
	.w7(32'hbb0f8751),
	.w8(32'hbba2f393),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6db5b1),
	.w1(32'hbb3d7535),
	.w2(32'hbb37d2d6),
	.w3(32'h3aad08af),
	.w4(32'hbb1436f7),
	.w5(32'hbb2f4e09),
	.w6(32'hbb3c3b10),
	.w7(32'hbb4dee28),
	.w8(32'hbb79324e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cd913),
	.w1(32'h3b588678),
	.w2(32'h3a40c9c8),
	.w3(32'hbc064b7d),
	.w4(32'h395890da),
	.w5(32'h39bdb717),
	.w6(32'hbbb0e836),
	.w7(32'hb9b70035),
	.w8(32'hbbd37341),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbec90b),
	.w1(32'hbbd7067d),
	.w2(32'hbc243429),
	.w3(32'h3b9bf6fa),
	.w4(32'hbbd8a2d8),
	.w5(32'hbc137363),
	.w6(32'hbc0c5545),
	.w7(32'hbbe71812),
	.w8(32'hbc3b0ff4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10a14b),
	.w1(32'h3a8397d8),
	.w2(32'h3a606cbe),
	.w3(32'hba6a79de),
	.w4(32'h3acfb024),
	.w5(32'h3a99f1f1),
	.w6(32'h3ad0b774),
	.w7(32'h3a92caf3),
	.w8(32'h3af57491),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc5dc3),
	.w1(32'hbb87aba9),
	.w2(32'hbb8d3784),
	.w3(32'h3afcb77f),
	.w4(32'hbb74d3ef),
	.w5(32'hbb94badf),
	.w6(32'hbb07aa9d),
	.w7(32'hbb69ae94),
	.w8(32'hbb89e486),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc03ef),
	.w1(32'h3a0c4c18),
	.w2(32'h3a6961dd),
	.w3(32'hbbb9f3cf),
	.w4(32'h3b7b9024),
	.w5(32'h3c0f4585),
	.w6(32'hbb92dee9),
	.w7(32'hbaa58cd2),
	.w8(32'hbb5fc787),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1084fe),
	.w1(32'h3c17dd82),
	.w2(32'h39cc9069),
	.w3(32'h3b71ab1a),
	.w4(32'h3b12987e),
	.w5(32'hbc0ef498),
	.w6(32'hbbe9c38f),
	.w7(32'h392612df),
	.w8(32'hbc3e8670),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38be30),
	.w1(32'hbbf12352),
	.w2(32'hbc8ffdca),
	.w3(32'hbb2bcdee),
	.w4(32'hbb91dfeb),
	.w5(32'hbc7340a4),
	.w6(32'hbc0ea86a),
	.w7(32'hbbce1e77),
	.w8(32'hbc3a66f0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d8e92),
	.w1(32'h3bc9585d),
	.w2(32'h3b3d70a1),
	.w3(32'hbc1ee62b),
	.w4(32'h3b51eea2),
	.w5(32'hba71513f),
	.w6(32'hbbaab121),
	.w7(32'h3bda65e9),
	.w8(32'hbb20eee8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afd446),
	.w1(32'h3ad038d9),
	.w2(32'hba97f53f),
	.w3(32'hbb92c610),
	.w4(32'h3b4e9d3a),
	.w5(32'h3907e2f9),
	.w6(32'hba0eced4),
	.w7(32'hba9d7eca),
	.w8(32'hbb0f3695),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0915ae),
	.w1(32'hba014659),
	.w2(32'hba16eb48),
	.w3(32'hba18c4d1),
	.w4(32'hb90d7a48),
	.w5(32'hb9e4e568),
	.w6(32'h39a2c4a4),
	.w7(32'hb85b7789),
	.w8(32'h385e461f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd0852),
	.w1(32'hbbbb7efd),
	.w2(32'hbc11680f),
	.w3(32'hbb36b924),
	.w4(32'hbb816110),
	.w5(32'hbbc5b4ec),
	.w6(32'hbbee6456),
	.w7(32'hbba67592),
	.w8(32'hbb8982c0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50bcbf),
	.w1(32'h3b0ee55d),
	.w2(32'h3b20b39c),
	.w3(32'hbc45412d),
	.w4(32'hb875beac),
	.w5(32'h3a2f2427),
	.w6(32'hbb914255),
	.w7(32'h384960e2),
	.w8(32'hbb426a54),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828a48),
	.w1(32'hbb47078b),
	.w2(32'hbbbde301),
	.w3(32'hbb8c5bd8),
	.w4(32'hbb3af1a3),
	.w5(32'hbbaf42a3),
	.w6(32'hbbe975ea),
	.w7(32'hbb14bda7),
	.w8(32'hbbcdfff0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0296f),
	.w1(32'hbb5beeb3),
	.w2(32'hbb6f2534),
	.w3(32'hbb246c1f),
	.w4(32'hbb43cf64),
	.w5(32'hbb643d2a),
	.w6(32'hbb148eaa),
	.w7(32'hbb4b1632),
	.w8(32'hbb5eb808),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e7c34),
	.w1(32'h38e03d73),
	.w2(32'hba0c50fe),
	.w3(32'hbb627391),
	.w4(32'h3a2e56cf),
	.w5(32'h37e2948a),
	.w6(32'h3acdcd41),
	.w7(32'h39f259b0),
	.w8(32'h39f7185d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a4514c),
	.w1(32'hbaa9bcfe),
	.w2(32'hbc071b6b),
	.w3(32'h3a5237ec),
	.w4(32'hba703d0d),
	.w5(32'hbbe51c6b),
	.w6(32'hbb1456fa),
	.w7(32'hbb116add),
	.w8(32'hbbc146e0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2f2f4),
	.w1(32'hb973778f),
	.w2(32'hbb45b83d),
	.w3(32'hbbd9997b),
	.w4(32'h3b99efb0),
	.w5(32'h3a907f18),
	.w6(32'hbb891d6f),
	.w7(32'hbaa91178),
	.w8(32'h3ad79fc9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba885b5a),
	.w1(32'h3c01c41e),
	.w2(32'h3c32cb46),
	.w3(32'h398594dd),
	.w4(32'h3b9db327),
	.w5(32'h3c18146c),
	.w6(32'hbaf3485e),
	.w7(32'h3b2bb490),
	.w8(32'hb8041709),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9909b),
	.w1(32'hba705ec7),
	.w2(32'hbb2bbce1),
	.w3(32'h3bd58611),
	.w4(32'h3a87e4cf),
	.w5(32'hba6eb596),
	.w6(32'h3acc190a),
	.w7(32'h3a937aa0),
	.w8(32'h39630bbe),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0912ae),
	.w1(32'h3bdd0743),
	.w2(32'h3ae85f82),
	.w3(32'h3b4c0fc8),
	.w4(32'h3b988d03),
	.w5(32'h3b1a6953),
	.w6(32'h3a195ea8),
	.w7(32'h3ba7d37c),
	.w8(32'hbb4fe490),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae76786),
	.w1(32'h3c3d9809),
	.w2(32'h3c70c97e),
	.w3(32'hbad1b27e),
	.w4(32'h3c5255fd),
	.w5(32'h3c80486c),
	.w6(32'hbc5c39bd),
	.w7(32'h3ba784ff),
	.w8(32'h3b807346),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ca3a4),
	.w1(32'h3b822b82),
	.w2(32'h3b809ced),
	.w3(32'hbba54861),
	.w4(32'h3bb713cc),
	.w5(32'h3b5f83e3),
	.w6(32'hbc70a642),
	.w7(32'hba8cb9f8),
	.w8(32'hba92ff2c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2938b),
	.w1(32'h3acf50a7),
	.w2(32'h3ab3ac7f),
	.w3(32'h3aca4dd1),
	.w4(32'h3abf9e4f),
	.w5(32'h3b2c00a6),
	.w6(32'hbbbbdfd5),
	.w7(32'hbb0a0c48),
	.w8(32'hbb0fa2fa),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4538b3),
	.w1(32'hb9c10a58),
	.w2(32'h3a9cebb1),
	.w3(32'h3b6516c1),
	.w4(32'hbaeca11f),
	.w5(32'hb9733a01),
	.w6(32'hba726ee4),
	.w7(32'h3a28a5c8),
	.w8(32'hb9b19fbd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a64153),
	.w1(32'hb893e0d8),
	.w2(32'h3a76f02f),
	.w3(32'hbae7fcaf),
	.w4(32'hbad78a68),
	.w5(32'hbaaabf13),
	.w6(32'hbbc5ad20),
	.w7(32'hbb4577f5),
	.w8(32'hbb8379c0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5700ae),
	.w1(32'h38063025),
	.w2(32'hbab7d0fb),
	.w3(32'hbbbad9bf),
	.w4(32'h39c572be),
	.w5(32'hba9926eb),
	.w6(32'hbb1bb108),
	.w7(32'hb9dd6e1c),
	.w8(32'hbae79054),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe34cb),
	.w1(32'h3adf6cc9),
	.w2(32'h3b9936d0),
	.w3(32'hbbecb148),
	.w4(32'hba8aa57d),
	.w5(32'h3ae6ca7f),
	.w6(32'hbc88e728),
	.w7(32'hbb9f5a39),
	.w8(32'hbc005bcd),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b611e),
	.w1(32'hbbc98477),
	.w2(32'hbc69b5c7),
	.w3(32'h3c0152c9),
	.w4(32'hbb83fa6d),
	.w5(32'hbc3fa4c8),
	.w6(32'hbc371b78),
	.w7(32'hbbf0ed74),
	.w8(32'hbc703424),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc642ebb),
	.w1(32'hbb92a6b8),
	.w2(32'hbc6546c8),
	.w3(32'hbc316944),
	.w4(32'hba70e9f1),
	.w5(32'hbc041724),
	.w6(32'hbc5777b4),
	.w7(32'hbbdfabe2),
	.w8(32'hbc45b87b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad191dd),
	.w1(32'h3b42a20e),
	.w2(32'h3ae59346),
	.w3(32'h3a59fa0b),
	.w4(32'h3a864435),
	.w5(32'hbab2fa32),
	.w6(32'hbc07be4f),
	.w7(32'h3b8385bc),
	.w8(32'hbb0f87f0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c66b15),
	.w1(32'hbbd67607),
	.w2(32'hbc01d7f7),
	.w3(32'hbba55692),
	.w4(32'hbc2100fc),
	.w5(32'hbc4e7566),
	.w6(32'hbc19f50c),
	.w7(32'hbc38dde6),
	.w8(32'hbc56d7e0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f9649),
	.w1(32'hb89b56ea),
	.w2(32'h397b8a2a),
	.w3(32'hb984957d),
	.w4(32'h39ae9a69),
	.w5(32'h3a3969c9),
	.w6(32'h3a6b4437),
	.w7(32'h39c24cd5),
	.w8(32'h3a4f1004),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd6deb),
	.w1(32'hbc2113d6),
	.w2(32'hbc1e8580),
	.w3(32'h39ffb1e6),
	.w4(32'hbc11da11),
	.w5(32'hbc1c6870),
	.w6(32'hbc11959a),
	.w7(32'hbc1d37d9),
	.w8(32'hbc062523),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc260215),
	.w1(32'hbb8807ea),
	.w2(32'hbb987dda),
	.w3(32'hbc13c765),
	.w4(32'hbbbb5a25),
	.w5(32'hbba13c00),
	.w6(32'hbbe3dd91),
	.w7(32'hbbf33b93),
	.w8(32'hbc03bdc7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28a37a),
	.w1(32'h3bef6c4b),
	.w2(32'h397fec9d),
	.w3(32'hbc0c73ff),
	.w4(32'h3b8668a3),
	.w5(32'hbb9916ab),
	.w6(32'hba941b51),
	.w7(32'h3b867a5d),
	.w8(32'hbb213289),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fd3e5),
	.w1(32'h3b803180),
	.w2(32'h3b44c271),
	.w3(32'hbc350d8a),
	.w4(32'h3b273ce1),
	.w5(32'h3aaed81f),
	.w6(32'h3b4dae43),
	.w7(32'h3b975e86),
	.w8(32'h38846e70),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79d5a3),
	.w1(32'hbc1bc08f),
	.w2(32'hbbf06824),
	.w3(32'hbb9828c5),
	.w4(32'hbc108ee5),
	.w5(32'hbc0aa9ae),
	.w6(32'hbc0e1794),
	.w7(32'hbacd411d),
	.w8(32'hbb82e01e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c207a45),
	.w1(32'h3a47bdea),
	.w2(32'h3b85ca5b),
	.w3(32'h3c04ee6f),
	.w4(32'hba043559),
	.w5(32'h3b407bbf),
	.w6(32'hbb3416ac),
	.w7(32'h3a7cf648),
	.w8(32'h370076e7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb194f),
	.w1(32'h3b0bd4b1),
	.w2(32'h3b23f0bd),
	.w3(32'h3a88e9c4),
	.w4(32'h3a9e6172),
	.w5(32'h3b1a6343),
	.w6(32'h3aa19b2f),
	.w7(32'h3adfab08),
	.w8(32'h381490a8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a449fe7),
	.w1(32'hbb3ec066),
	.w2(32'hba89f213),
	.w3(32'hb8f8870a),
	.w4(32'hbbacb65e),
	.w5(32'hbb7bd418),
	.w6(32'hbb8a7327),
	.w7(32'hbb5dd893),
	.w8(32'hbbc4ab46),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994c4c),
	.w1(32'hbb7cb73c),
	.w2(32'hbb4e4ac7),
	.w3(32'hbbddbe76),
	.w4(32'hbb93915c),
	.w5(32'hbafd8ae9),
	.w6(32'hbb9e4642),
	.w7(32'hbb5adc1d),
	.w8(32'hbaf5e6db),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45a1ff),
	.w1(32'h3bcf5aa0),
	.w2(32'h3be14526),
	.w3(32'h39c2518a),
	.w4(32'h3b681e69),
	.w5(32'h3bc45005),
	.w6(32'hbb68144b),
	.w7(32'h39da11a3),
	.w8(32'hba8f0fb0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a6ab6),
	.w1(32'hbb6d0484),
	.w2(32'hbbaafe9a),
	.w3(32'h3ad11163),
	.w4(32'hbadf4322),
	.w5(32'hbb5e2ae2),
	.w6(32'hba0fc988),
	.w7(32'hbb2f4160),
	.w8(32'hbad98fd3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc043abd),
	.w1(32'hbbf036f5),
	.w2(32'hbbbbfe77),
	.w3(32'hbbc7e347),
	.w4(32'hbbfcbb15),
	.w5(32'hbba64109),
	.w6(32'hbc88b98d),
	.w7(32'hbc1a52b9),
	.w8(32'hbc2750ae),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb35f70),
	.w1(32'hbc1323c4),
	.w2(32'hbc2d732b),
	.w3(32'hbb5c15fc),
	.w4(32'hbc0503cd),
	.w5(32'hbc1ce7c9),
	.w6(32'hbc097e02),
	.w7(32'hbc1c5680),
	.w8(32'hbc24dbcc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ac447),
	.w1(32'hbb8ee917),
	.w2(32'hba934e44),
	.w3(32'hbbd84412),
	.w4(32'hbbdddcbc),
	.w5(32'hbaaa9af4),
	.w6(32'hbb6c8683),
	.w7(32'hbb09d226),
	.w8(32'h3a2cf67c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397aed5d),
	.w1(32'h3bbeba87),
	.w2(32'h3c1f9b5c),
	.w3(32'hb94629df),
	.w4(32'h3b7f0808),
	.w5(32'h3c0c9629),
	.w6(32'hbb1418de),
	.w7(32'h3b443318),
	.w8(32'h3b2a700a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14364d),
	.w1(32'hba633007),
	.w2(32'hbb1cab7a),
	.w3(32'h3bf2efca),
	.w4(32'hbb4a1a15),
	.w5(32'hbac5ade6),
	.w6(32'hbac734ab),
	.w7(32'hbb2f56de),
	.w8(32'hba9ab7b0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e9235),
	.w1(32'h3998b2af),
	.w2(32'hbb20f2ac),
	.w3(32'hba18962e),
	.w4(32'hba35540b),
	.w5(32'hbaca7587),
	.w6(32'hb86e6b45),
	.w7(32'hba241650),
	.w8(32'hba80236c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9bd3f),
	.w1(32'hbc2eec52),
	.w2(32'hbc58cae4),
	.w3(32'hbb0890fa),
	.w4(32'hbc2fabce),
	.w5(32'hbc508c8d),
	.w6(32'hbc1b98db),
	.w7(32'hbc1a8c6e),
	.w8(32'hbc3d1f28),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48da6a),
	.w1(32'h3ad6c78e),
	.w2(32'hbbbfc3cd),
	.w3(32'hbc439f87),
	.w4(32'hbb4077b7),
	.w5(32'hbc1d151c),
	.w6(32'hbb51c885),
	.w7(32'h3b10628b),
	.w8(32'hbbfe5fc7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c2a89),
	.w1(32'h3b1f5adf),
	.w2(32'hbaa188d5),
	.w3(32'hbb8a8a21),
	.w4(32'h3ba5d081),
	.w5(32'h3a96c47d),
	.w6(32'hbb39e326),
	.w7(32'h3b9ac1ce),
	.w8(32'h3aaac7f6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ea4ae),
	.w1(32'hbc4c99c8),
	.w2(32'hbcd05520),
	.w3(32'h3b0cbed6),
	.w4(32'hbc25e961),
	.w5(32'hbc9b5c6b),
	.w6(32'hbcab12c4),
	.w7(32'hbc33f390),
	.w8(32'hbc898c05),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46518f),
	.w1(32'h3bce9958),
	.w2(32'h3c0a3c31),
	.w3(32'hbc488951),
	.w4(32'h3b5d517b),
	.w5(32'h3bed4986),
	.w6(32'hba01ffc9),
	.w7(32'h3b08c35a),
	.w8(32'h3a9db3a0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf64840),
	.w1(32'hba6cca05),
	.w2(32'hbb17aa60),
	.w3(32'h3b9ad0a2),
	.w4(32'h399fe707),
	.w5(32'hba807df9),
	.w6(32'h39d4e7e5),
	.w7(32'hba9069e2),
	.w8(32'h3732b986),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925fe6c),
	.w1(32'hbae747a4),
	.w2(32'hbb36897a),
	.w3(32'h3a4b6839),
	.w4(32'hb9800463),
	.w5(32'hba9d5df8),
	.w6(32'h3a2dd1d0),
	.w7(32'hba96026a),
	.w8(32'h38c1b255),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb344c25),
	.w1(32'hb8cb2d60),
	.w2(32'hba6ad0f8),
	.w3(32'hbac75b19),
	.w4(32'h39f9003a),
	.w5(32'hba9f9468),
	.w6(32'hb91274b4),
	.w7(32'h39ed8f6a),
	.w8(32'hb923f1b0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9beb320),
	.w1(32'h3b2efce6),
	.w2(32'h3b9c3aef),
	.w3(32'h39cf20f2),
	.w4(32'hbaaca3f2),
	.w5(32'h3aef5e73),
	.w6(32'hbaf3fc03),
	.w7(32'h3b022634),
	.w8(32'hbafa2ff1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1d250),
	.w1(32'hba33c1f1),
	.w2(32'h3b944b3e),
	.w3(32'hbb5e9c3b),
	.w4(32'h3ab3267f),
	.w5(32'h3b0a8a1d),
	.w6(32'hbc322685),
	.w7(32'hbaa99740),
	.w8(32'hbbcc8930),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97245e),
	.w1(32'hbc1c7ece),
	.w2(32'hbc55fd2b),
	.w3(32'hbc189fd5),
	.w4(32'hbbd6b477),
	.w5(32'hbc28d014),
	.w6(32'hbbbb72b5),
	.w7(32'hbba45f18),
	.w8(32'hbbf1f365),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ae4d9),
	.w1(32'hbb9a8cf2),
	.w2(32'hbb9ea4fe),
	.w3(32'hbc0870b4),
	.w4(32'hbb414fdd),
	.w5(32'hbb47a2c1),
	.w6(32'hbc508615),
	.w7(32'hbbf2976f),
	.w8(32'hbc1f9c20),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08f9e8),
	.w1(32'h3b9200a9),
	.w2(32'h3a8f465b),
	.w3(32'hba405a0e),
	.w4(32'h3bdc888a),
	.w5(32'h3b3321dc),
	.w6(32'h3b64701a),
	.w7(32'h3bb1d3ce),
	.w8(32'h3ac21181),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2e7fc),
	.w1(32'hbb74b705),
	.w2(32'hbc10b46b),
	.w3(32'h3b86ee9d),
	.w4(32'hbba3f730),
	.w5(32'hbc21f1b5),
	.w6(32'hbb36c8f3),
	.w7(32'hbb85b2d7),
	.w8(32'hbbeb5401),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc44f78),
	.w1(32'hb9f75685),
	.w2(32'hba37c7e2),
	.w3(32'hbbb1f23f),
	.w4(32'hbb0ee345),
	.w5(32'hbb21ac76),
	.w6(32'hbb80bce3),
	.w7(32'hb8a843da),
	.w8(32'hbb448eb8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c4a9d),
	.w1(32'hbb429b4f),
	.w2(32'hbab94bae),
	.w3(32'hbb8f55b9),
	.w4(32'hbbfd0784),
	.w5(32'hbbda9c31),
	.w6(32'hbc19649b),
	.w7(32'hbb924b0c),
	.w8(32'hbbdb01d4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acaccb4),
	.w1(32'h3bb89269),
	.w2(32'h3c049e6b),
	.w3(32'hbb03182c),
	.w4(32'h3b35ef96),
	.w5(32'h3b9a48ff),
	.w6(32'h3b8650cf),
	.w7(32'h3be7766a),
	.w8(32'h3b6b549f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dd68d),
	.w1(32'hb9209997),
	.w2(32'h3b2dbf51),
	.w3(32'h38ad4bf4),
	.w4(32'h3a1a4309),
	.w5(32'h3b5520cf),
	.w6(32'hbbd83df5),
	.w7(32'hbb80b3ec),
	.w8(32'hbbd1dd1f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacea0ac),
	.w1(32'h3b306d4b),
	.w2(32'h3ae9a173),
	.w3(32'hba453d29),
	.w4(32'h3b20f87c),
	.w5(32'h3abda9c2),
	.w6(32'h3b9a2841),
	.w7(32'h3b3a8537),
	.w8(32'h3b83fc04),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b275046),
	.w1(32'hb9819633),
	.w2(32'h3aed8634),
	.w3(32'h3b6b70ec),
	.w4(32'hbae992d9),
	.w5(32'hb8d07092),
	.w6(32'hbb22d848),
	.w7(32'hba17b02b),
	.w8(32'hbb0c2344),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09aa03),
	.w1(32'h3b2ce8de),
	.w2(32'hb915e87f),
	.w3(32'hbb0ef097),
	.w4(32'h3b91ffa0),
	.w5(32'hb9c7bb2c),
	.w6(32'hbbe09e8a),
	.w7(32'hbaf69326),
	.w8(32'hbbbb0de4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb41b42),
	.w1(32'hbb11c060),
	.w2(32'hbb4e258e),
	.w3(32'hbbc59ad8),
	.w4(32'hbb1a1ccf),
	.w5(32'hbb3fc274),
	.w6(32'hbb1c7dec),
	.w7(32'hbb059309),
	.w8(32'hbb3be0da),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad39a4d),
	.w1(32'h3a8c2907),
	.w2(32'hba40b7fb),
	.w3(32'hba3b40c1),
	.w4(32'hba8a53db),
	.w5(32'hbb6357b3),
	.w6(32'hba74697f),
	.w7(32'h3b12c80f),
	.w8(32'hbb9fc0fc),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e96ce),
	.w1(32'hbbe6f64c),
	.w2(32'hbbdb13ae),
	.w3(32'hbc3c608b),
	.w4(32'hbbdc0ec8),
	.w5(32'hbbf4f957),
	.w6(32'hbc3fc445),
	.w7(32'hbbf26f59),
	.w8(32'hbc02d5da),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfabdcc),
	.w1(32'hba03cdb7),
	.w2(32'hbae1172b),
	.w3(32'hbbb0c951),
	.w4(32'h3ac78962),
	.w5(32'hba15e545),
	.w6(32'hbb9e802c),
	.w7(32'hb9ca2f80),
	.w8(32'hbb0b8e8a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a872b),
	.w1(32'h3b43383c),
	.w2(32'h3bc46568),
	.w3(32'hbb821a90),
	.w4(32'hba8a53bf),
	.w5(32'h3a862740),
	.w6(32'hbbb9c2f6),
	.w7(32'hba955a1f),
	.w8(32'hbb943182),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb3466),
	.w1(32'h3c10aaf7),
	.w2(32'h3c1f28b5),
	.w3(32'h3bd4c20f),
	.w4(32'h3b9a34f9),
	.w5(32'h3bd51f61),
	.w6(32'h3b1934e3),
	.w7(32'h3c014609),
	.w8(32'h3b3cc4d9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be11835),
	.w1(32'h3b277db0),
	.w2(32'hbb6dad39),
	.w3(32'h3b8dc1a3),
	.w4(32'h3afec8de),
	.w5(32'hbb69b88f),
	.w6(32'hb9b1c1da),
	.w7(32'h3b93e183),
	.w8(32'hbb92e099),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d3162),
	.w1(32'h3b902752),
	.w2(32'h3abf8dad),
	.w3(32'h3b026e2e),
	.w4(32'h3b8b8b15),
	.w5(32'h3a8eccd8),
	.w6(32'hbb0d6691),
	.w7(32'h3a94954f),
	.w8(32'hbb48bbfb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c37c97),
	.w1(32'hba5de42c),
	.w2(32'hbb406c0a),
	.w3(32'h3a08b87a),
	.w4(32'h3bbe3217),
	.w5(32'h3b3f8485),
	.w6(32'hbbf3fcc7),
	.w7(32'hbb302822),
	.w8(32'hbb8d6bd0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b328cec),
	.w1(32'h3b0cf2aa),
	.w2(32'hb88a148e),
	.w3(32'h3c1e5183),
	.w4(32'h3b2e4fce),
	.w5(32'h3a4b740c),
	.w6(32'h3b21cc1b),
	.w7(32'hb9803674),
	.w8(32'h3ab3347e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2df94),
	.w1(32'hba642073),
	.w2(32'hbc453886),
	.w3(32'hba4b49e5),
	.w4(32'hbab4a7dc),
	.w5(32'hbc1984f2),
	.w6(32'hbbc82c0b),
	.w7(32'hbb6755e2),
	.w8(32'hbc2345c3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9abaa0),
	.w1(32'h3a461ca4),
	.w2(32'h3a4f1383),
	.w3(32'hbb4a3d2d),
	.w4(32'hb9da87ad),
	.w5(32'h3a7e5c21),
	.w6(32'hbc03b92d),
	.w7(32'hbabdbef3),
	.w8(32'hbb70a7cb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1cb10),
	.w1(32'h3c1173c6),
	.w2(32'h3bd93d6b),
	.w3(32'hbb206c79),
	.w4(32'h3abeb350),
	.w5(32'hba747535),
	.w6(32'h3acfbaeb),
	.w7(32'h3c0fe91a),
	.w8(32'hbb8871c7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4fcbf),
	.w1(32'h3c6e66a4),
	.w2(32'h3c31d56b),
	.w3(32'h3ac16044),
	.w4(32'h3c812d32),
	.w5(32'h3c430bc2),
	.w6(32'hbb9bf8c2),
	.w7(32'h3bed6def),
	.w8(32'h3b332bd3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84e4e2),
	.w1(32'hbbf4def9),
	.w2(32'hbc25cdfa),
	.w3(32'h3b24e435),
	.w4(32'hbb907c37),
	.w5(32'hbc05d575),
	.w6(32'hbc59771a),
	.w7(32'hbbe1b10b),
	.w8(32'hbc06f73d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb05d7),
	.w1(32'hbb730281),
	.w2(32'hbc3d6673),
	.w3(32'h3bcf82ea),
	.w4(32'hba7cf69a),
	.w5(32'hbc0b3808),
	.w6(32'h3b8b30eb),
	.w7(32'h3af01cb7),
	.w8(32'hbb3c49bb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8c6c1),
	.w1(32'h3a383a80),
	.w2(32'hba8a6b7c),
	.w3(32'hbac052c3),
	.w4(32'h3adb229b),
	.w5(32'h398c5629),
	.w6(32'h3b040d4a),
	.w7(32'h3a10b267),
	.w8(32'h3ab3aa89),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68d323),
	.w1(32'hbbe8d828),
	.w2(32'hbc380901),
	.w3(32'hb9ee3a90),
	.w4(32'hbb780d2c),
	.w5(32'hbc42118b),
	.w6(32'hbab1fb49),
	.w7(32'hbabdb6c8),
	.w8(32'hbb79898b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdb54a),
	.w1(32'hbb3d4e69),
	.w2(32'hbb99ff22),
	.w3(32'hbb82ab29),
	.w4(32'hba9dfb77),
	.w5(32'hbb756423),
	.w6(32'hbae0e8b8),
	.w7(32'hba972a44),
	.w8(32'hbb38a16c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8357b4),
	.w1(32'h3a475a56),
	.w2(32'h3b63ed9d),
	.w3(32'hba859452),
	.w4(32'hbb45826b),
	.w5(32'h3a8c0216),
	.w6(32'hbb18aeac),
	.w7(32'hba7804f0),
	.w8(32'hbabc1d44),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b079d4b),
	.w1(32'hbb952fa7),
	.w2(32'hbbbb1bd5),
	.w3(32'h39a4707c),
	.w4(32'hbb630d5d),
	.w5(32'hbb95771b),
	.w6(32'hbb3dffa9),
	.w7(32'hbb6aadb9),
	.w8(32'hbb98e590),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27dc4e),
	.w1(32'hbc215117),
	.w2(32'hbc43c5e1),
	.w3(32'hbc0e239a),
	.w4(32'hbc019930),
	.w5(32'hbc37bd99),
	.w6(32'hbc18b1bc),
	.w7(32'hbc230b61),
	.w8(32'hbc1f5ace),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba90f9c),
	.w1(32'h391d0922),
	.w2(32'hbb9e1c3c),
	.w3(32'hbb3d837a),
	.w4(32'hbaa14924),
	.w5(32'hbba8f0f2),
	.w6(32'hbbcbc1c9),
	.w7(32'hbb2f9f7b),
	.w8(32'hbbf4daf9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b941f),
	.w1(32'h3accbebb),
	.w2(32'hba8c7f32),
	.w3(32'hbb751ff4),
	.w4(32'h3b6d68f6),
	.w5(32'hba5d7e16),
	.w6(32'hbaffa76b),
	.w7(32'hba5d6eb8),
	.w8(32'hbb80f5bd),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39525eb3),
	.w1(32'h3ba6fa9e),
	.w2(32'h3b1ae4a1),
	.w3(32'h3a892cff),
	.w4(32'h3b4895dd),
	.w5(32'hbaacbbba),
	.w6(32'hba913603),
	.w7(32'h3a004d48),
	.w8(32'hbbaac421),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88d40),
	.w1(32'h3ae215eb),
	.w2(32'hba9887d4),
	.w3(32'hbbf2bc7c),
	.w4(32'h3b4c9e27),
	.w5(32'hb8d101f5),
	.w6(32'h3a6adadc),
	.w7(32'h3b06fcaf),
	.w8(32'h391738cb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9d735),
	.w1(32'hba4a7491),
	.w2(32'hbb9d4667),
	.w3(32'hbb1f27e3),
	.w4(32'hbb7fddab),
	.w5(32'hbbd91360),
	.w6(32'hbb7c4b61),
	.w7(32'hbb6e5c17),
	.w8(32'hbc05f2c4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3478ac),
	.w1(32'hbc49db19),
	.w2(32'hbc633d53),
	.w3(32'hbb7cdc21),
	.w4(32'hbc465f73),
	.w5(32'hbc67452f),
	.w6(32'hbc728bfb),
	.w7(32'hbc4d07ab),
	.w8(32'hbc812da3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc573393),
	.w1(32'hbbb0ad8f),
	.w2(32'hbbd1b055),
	.w3(32'hbc568c83),
	.w4(32'hbb3d28b3),
	.w5(32'hbb9adb2f),
	.w6(32'hb9588b14),
	.w7(32'hbb208867),
	.w8(32'hba92bb51),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d50ac),
	.w1(32'hbba4f9ea),
	.w2(32'hbbcf5b4a),
	.w3(32'hbab1761d),
	.w4(32'hbb621d27),
	.w5(32'hbb97a76d),
	.w6(32'hbb262fd4),
	.w7(32'hbb961c44),
	.w8(32'hbb3f6c7b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ac126),
	.w1(32'hbb07befe),
	.w2(32'hbb68dabc),
	.w3(32'hbb1b1a9b),
	.w4(32'hba0bca76),
	.w5(32'hbaf653c5),
	.w6(32'h3a10ced2),
	.w7(32'hbab3e14f),
	.w8(32'h39a2727a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81d762),
	.w1(32'hbb50337b),
	.w2(32'hbb2b556c),
	.w3(32'h3a2de6fa),
	.w4(32'hbb3cc9c6),
	.w5(32'hbab69efc),
	.w6(32'hbb96343b),
	.w7(32'hbb7a0b1e),
	.w8(32'hbb59d5d1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb149a),
	.w1(32'hba88fe56),
	.w2(32'hbbf616f0),
	.w3(32'hbb3c1253),
	.w4(32'hbac71218),
	.w5(32'hbbafef39),
	.w6(32'hbbbe0eaa),
	.w7(32'hbb88c93f),
	.w8(32'hbc21c103),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ea753),
	.w1(32'h3b10eecb),
	.w2(32'hb90042df),
	.w3(32'hbb556ba9),
	.w4(32'h3b7f0bd0),
	.w5(32'h3ab2cf3b),
	.w6(32'h3b872882),
	.w7(32'h3ae15905),
	.w8(32'h3ab4e937),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bab64),
	.w1(32'hbb82401a),
	.w2(32'hbbaa3aab),
	.w3(32'h3b3b5c63),
	.w4(32'hbb56fd8f),
	.w5(32'hbb8cb6ce),
	.w6(32'hbae2f1f4),
	.w7(32'hbb504772),
	.w8(32'hbb372e69),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbab7e7),
	.w1(32'hbbb77f31),
	.w2(32'hbb88e994),
	.w3(32'hbba08fc8),
	.w4(32'hbb692640),
	.w5(32'hbb907118),
	.w6(32'hbc170050),
	.w7(32'hbbe7d0c6),
	.w8(32'hbbbe9a5e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9df546),
	.w1(32'hbbc3d269),
	.w2(32'hb9af4016),
	.w3(32'hbb4d9b2c),
	.w4(32'hbba37aa8),
	.w5(32'h3a075f9e),
	.w6(32'hbc1a913f),
	.w7(32'hbbeae2b5),
	.w8(32'hbb925797),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3705b5),
	.w1(32'h3b4db754),
	.w2(32'h3be6d53b),
	.w3(32'h3b4d39b8),
	.w4(32'h3b75bed5),
	.w5(32'h3bfad5c2),
	.w6(32'h3ae94be3),
	.w7(32'h3ba4dae3),
	.w8(32'h3b8af306),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee76b9),
	.w1(32'hbb40dd2f),
	.w2(32'hbb3c5755),
	.w3(32'h3c029324),
	.w4(32'hbb13dff5),
	.w5(32'hbb2a1fbd),
	.w6(32'hba9c5116),
	.w7(32'hbb0550e6),
	.w8(32'hbb0b0ca6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66e2be),
	.w1(32'hbb2725f8),
	.w2(32'hb99622d7),
	.w3(32'hbb33ef27),
	.w4(32'hb7b4b595),
	.w5(32'h3b416905),
	.w6(32'hbb3d7c6b),
	.w7(32'h3afb4333),
	.w8(32'hbba66c8f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86feb8),
	.w1(32'h3a79b8b6),
	.w2(32'hbb3f99bf),
	.w3(32'hbb7a8bb8),
	.w4(32'h3a230bf0),
	.w5(32'hbb524393),
	.w6(32'h36552118),
	.w7(32'h39bc7fdb),
	.w8(32'hbbba02b2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c3908),
	.w1(32'hbb24912c),
	.w2(32'hbbe0639e),
	.w3(32'hbb840620),
	.w4(32'hbb7c199b),
	.w5(32'hbc2e419d),
	.w6(32'h386a81ef),
	.w7(32'hbbaaa47d),
	.w8(32'hbc17398a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad22e20),
	.w1(32'hb9adc5bb),
	.w2(32'hba09226b),
	.w3(32'hba0365fd),
	.w4(32'h3a61d6fa),
	.w5(32'h3a0bc926),
	.w6(32'hba51e111),
	.w7(32'hba01e0b5),
	.w8(32'hbaa8bd0c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f08eb),
	.w1(32'hbb05e88e),
	.w2(32'hbb5720ed),
	.w3(32'hbb78bd11),
	.w4(32'hba70c063),
	.w5(32'hbb197c07),
	.w6(32'hbb74daef),
	.w7(32'hbb126ad9),
	.w8(32'hbb86680d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf42664),
	.w1(32'hba2efd44),
	.w2(32'hbb709e3f),
	.w3(32'hbb6b823a),
	.w4(32'hbb7b22bc),
	.w5(32'hb9dacb1d),
	.w6(32'hba9bf4eb),
	.w7(32'h3aec3c39),
	.w8(32'hbb1ed0a7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d6d87),
	.w1(32'hbadaf6ce),
	.w2(32'hbbc81a16),
	.w3(32'hba0ac997),
	.w4(32'h3ab5f364),
	.w5(32'hbb2bd7be),
	.w6(32'hba98e1f6),
	.w7(32'hbb63aff2),
	.w8(32'h3a538f3b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3682c1),
	.w1(32'h3b455669),
	.w2(32'hbb829705),
	.w3(32'h3ba36a6e),
	.w4(32'h3bf8904b),
	.w5(32'h3af682bc),
	.w6(32'h3a68e50c),
	.w7(32'h39f82e97),
	.w8(32'hba9bfad0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21acca),
	.w1(32'hbac1366d),
	.w2(32'hbb9a2eec),
	.w3(32'hbb29c5bb),
	.w4(32'hbb1fdc78),
	.w5(32'hbbc16475),
	.w6(32'hbab7cb27),
	.w7(32'hbaecf5cb),
	.w8(32'hbc19140c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c67db5),
	.w1(32'h3ab47b61),
	.w2(32'hbb02e378),
	.w3(32'hba694226),
	.w4(32'h3b2d02e4),
	.w5(32'hbaa90dbe),
	.w6(32'hbae9de91),
	.w7(32'hb95a69a5),
	.w8(32'hbb90a867),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf551ad),
	.w1(32'h3ab4cce3),
	.w2(32'h39ed60d2),
	.w3(32'hba199e3a),
	.w4(32'h3b46e89f),
	.w5(32'h3a84a8bb),
	.w6(32'h3b32bac0),
	.w7(32'h3ba9f7ab),
	.w8(32'hb9ddf54a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992df73),
	.w1(32'hba6eec96),
	.w2(32'hbc089623),
	.w3(32'hb88b65c6),
	.w4(32'h3af70529),
	.w5(32'hbb8ed830),
	.w6(32'hbac20f8b),
	.w7(32'hbb006755),
	.w8(32'hbba56c7e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf07517),
	.w1(32'h3b4c9d48),
	.w2(32'h3b367ddf),
	.w3(32'h39d5d0b2),
	.w4(32'hbad14b80),
	.w5(32'hbb940bad),
	.w6(32'h3b12ff18),
	.w7(32'h3951eb63),
	.w8(32'hbb24ea03),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38233b),
	.w1(32'h3a030318),
	.w2(32'hbbac986c),
	.w3(32'hbbe78747),
	.w4(32'h3b1536fc),
	.w5(32'hbbbac5b9),
	.w6(32'hbade020e),
	.w7(32'hb9dc3cac),
	.w8(32'hbc08852b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41b5e4),
	.w1(32'hb91536ad),
	.w2(32'hba66ad8e),
	.w3(32'hba91a06f),
	.w4(32'hb9eff47f),
	.w5(32'hba8a2f24),
	.w6(32'hbb266615),
	.w7(32'hb97313a5),
	.w8(32'hbb29f086),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb491b98),
	.w1(32'h3be29c37),
	.w2(32'hbb519480),
	.w3(32'hbb102553),
	.w4(32'h3bd6746c),
	.w5(32'hbb3721c5),
	.w6(32'h3a756849),
	.w7(32'hba80d948),
	.w8(32'hbba93cbd),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1011db),
	.w1(32'h3bac0219),
	.w2(32'h3b56544f),
	.w3(32'hba9b3e7f),
	.w4(32'h3b85a852),
	.w5(32'h3a146091),
	.w6(32'h3b5155cb),
	.w7(32'h3b8b72f3),
	.w8(32'h39ee77b0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae34d6e),
	.w1(32'h3a00c697),
	.w2(32'h3b238f1b),
	.w3(32'h3ac16d5c),
	.w4(32'h3aafcbe4),
	.w5(32'h3b36fe01),
	.w6(32'h3836a95a),
	.w7(32'h3acf747e),
	.w8(32'hbad545a7),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba868f57),
	.w1(32'hb9e1d0be),
	.w2(32'hbb59df6b),
	.w3(32'hbaa6bd27),
	.w4(32'hba89c5c0),
	.w5(32'hbbb01e78),
	.w6(32'h392b9973),
	.w7(32'h3a093259),
	.w8(32'h3c9d5d6c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9853a9),
	.w1(32'hba880432),
	.w2(32'hba07d11f),
	.w3(32'h3c8af142),
	.w4(32'h3ac28450),
	.w5(32'h3b480053),
	.w6(32'hbb203022),
	.w7(32'hb966e904),
	.w8(32'hbaac739e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5db1bd),
	.w1(32'h3ba12bf9),
	.w2(32'h36b25b9e),
	.w3(32'h3b89e9de),
	.w4(32'h3c015572),
	.w5(32'h391ed7d4),
	.w6(32'h3b708dd2),
	.w7(32'h3b9713f2),
	.w8(32'h35897850),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaf399),
	.w1(32'hbb812241),
	.w2(32'hbb53f0b1),
	.w3(32'hbc0611df),
	.w4(32'hbb5c2c98),
	.w5(32'hbb7bb5cc),
	.w6(32'hbc47703b),
	.w7(32'hbb8c8a42),
	.w8(32'hbb93cfd5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dc43f),
	.w1(32'hbb1a9c8c),
	.w2(32'h3ab954eb),
	.w3(32'h3aa5fc2d),
	.w4(32'hba9d0c5e),
	.w5(32'h3b1f0582),
	.w6(32'hbb831b4b),
	.w7(32'h3ab63bed),
	.w8(32'hbb4f2be6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0c21),
	.w1(32'hbb802677),
	.w2(32'hbb9cfc03),
	.w3(32'hbb901c43),
	.w4(32'hbbbd8634),
	.w5(32'hbc1fe7e7),
	.w6(32'hbbb8a4c5),
	.w7(32'hbb6f0663),
	.w8(32'hbbbc3ff7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c603e),
	.w1(32'hbb6c50ed),
	.w2(32'h3c1b6158),
	.w3(32'hbafe55de),
	.w4(32'hbbf8b755),
	.w5(32'h3c7360a7),
	.w6(32'hbbcf8555),
	.w7(32'h3c970d3c),
	.w8(32'hbb97c977),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b69ebf),
	.w1(32'hbb8844e3),
	.w2(32'hbbf28d73),
	.w3(32'hbb1fc2db),
	.w4(32'hbaf5f500),
	.w5(32'hbbea397d),
	.w6(32'hbb1770e6),
	.w7(32'hbb0b095a),
	.w8(32'hbbf269c3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28d948),
	.w1(32'h3a2f025e),
	.w2(32'hbb98557d),
	.w3(32'hbad31342),
	.w4(32'h3ae8432d),
	.w5(32'hbbcd31a9),
	.w6(32'hbb0672f3),
	.w7(32'h3b2aeaf3),
	.w8(32'hba4fc790),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14c475),
	.w1(32'h3bd8cc5e),
	.w2(32'h3b0f2062),
	.w3(32'h39a9409a),
	.w4(32'h3a683b6b),
	.w5(32'hba3ebc40),
	.w6(32'hba8a2c69),
	.w7(32'hbb35cacd),
	.w8(32'hbba466bf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c3c5c),
	.w1(32'h3a2ce707),
	.w2(32'h3ad379d4),
	.w3(32'h3a501d67),
	.w4(32'h3a9ec9d4),
	.w5(32'h3b12f813),
	.w6(32'hba14892b),
	.w7(32'h3ad8a455),
	.w8(32'hbad60eea),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee1f5c),
	.w1(32'h3a921280),
	.w2(32'hbaa92b55),
	.w3(32'hbad1ac43),
	.w4(32'h3ba630f7),
	.w5(32'hbb039a81),
	.w6(32'hbb088290),
	.w7(32'h39e2e46e),
	.w8(32'hbb109ef5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8068ea),
	.w1(32'h3b9d67cf),
	.w2(32'hbb007854),
	.w3(32'h3824b382),
	.w4(32'h3b85b7af),
	.w5(32'hbb0695e8),
	.w6(32'hb9ce2a8b),
	.w7(32'h3b7dfdce),
	.w8(32'h3c346759),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02f179),
	.w1(32'h3a5889e5),
	.w2(32'hbc0f76f7),
	.w3(32'h3b10fb70),
	.w4(32'hb9efb193),
	.w5(32'hbc294bb9),
	.w6(32'hbaedd52f),
	.w7(32'hbbaf673a),
	.w8(32'h3c485d71),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32d3f1),
	.w1(32'hbadfb1a0),
	.w2(32'hb9fa4210),
	.w3(32'h3c018f15),
	.w4(32'hba84cbf3),
	.w5(32'h38480cbc),
	.w6(32'hbb08e6a6),
	.w7(32'h3a4cc84d),
	.w8(32'hbb08a0e6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ef1f7),
	.w1(32'hba763358),
	.w2(32'h368dfa43),
	.w3(32'hba728f57),
	.w4(32'hbaa82532),
	.w5(32'h3a5c4cb4),
	.w6(32'hbb37d9eb),
	.w7(32'hba940122),
	.w8(32'hbb63183d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ceabc),
	.w1(32'h3a0cc53e),
	.w2(32'hbc049079),
	.w3(32'hbb4e69ac),
	.w4(32'hbaa6abca),
	.w5(32'hbbdcf308),
	.w6(32'hba9a866d),
	.w7(32'hbb59c96b),
	.w8(32'h3b09ed75),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd36b54),
	.w1(32'h3b5d0dfd),
	.w2(32'h3bc01204),
	.w3(32'h3bb9fc8a),
	.w4(32'h3a8083be),
	.w5(32'h3b88cac1),
	.w6(32'h3a76bb76),
	.w7(32'h3bb7ab45),
	.w8(32'hbbd831c3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8d44d),
	.w1(32'h3aa69b21),
	.w2(32'hbb50f7b2),
	.w3(32'hbb27ecf4),
	.w4(32'h3b77c06c),
	.w5(32'h37f966f8),
	.w6(32'hba54ca15),
	.w7(32'h39ba1427),
	.w8(32'hbb3c2e86),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba346790),
	.w1(32'hb9531a72),
	.w2(32'h3a20bddf),
	.w3(32'h39a74c64),
	.w4(32'h3a764b8a),
	.w5(32'h3a7cdec2),
	.w6(32'hbb078cca),
	.w7(32'h3a055bc8),
	.w8(32'hbb1e8340),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcce79),
	.w1(32'h3ae6fd34),
	.w2(32'hb957df87),
	.w3(32'hbc2e4146),
	.w4(32'hbab980f6),
	.w5(32'hbb297bbe),
	.w6(32'hbb8d89c2),
	.w7(32'hba5f9af4),
	.w8(32'hbba2f400),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0035bc),
	.w1(32'h3a83293b),
	.w2(32'h3abfbea5),
	.w3(32'hb8f4a75d),
	.w4(32'h3ae64230),
	.w5(32'h3b038d87),
	.w6(32'h3aa1b844),
	.w7(32'h3af8587a),
	.w8(32'h3ad284c3),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2c1ad),
	.w1(32'h3ab9c728),
	.w2(32'h3b15c129),
	.w3(32'h3a5964d8),
	.w4(32'h3b05985f),
	.w5(32'h3b0c2b54),
	.w6(32'h3a7c9c18),
	.w7(32'h3adef47e),
	.w8(32'hbac7be80),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ab823),
	.w1(32'h3b1fa7e1),
	.w2(32'hbaea586b),
	.w3(32'h3b14e7e9),
	.w4(32'h3ba7fa1d),
	.w5(32'h3a3f17aa),
	.w6(32'h3a1cf1de),
	.w7(32'h3a7b56af),
	.w8(32'hbb5480b2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba424c1),
	.w1(32'hbba14546),
	.w2(32'hbc7cc2e5),
	.w3(32'hbb9fc841),
	.w4(32'hbc0f190b),
	.w5(32'hbc8dc1a5),
	.w6(32'hbba3c4e0),
	.w7(32'hbbb87a40),
	.w8(32'hbb8fe06f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0d2a8),
	.w1(32'hbac9d596),
	.w2(32'h3aadf81e),
	.w3(32'hbb77d165),
	.w4(32'hbb0c20d7),
	.w5(32'hbaad96c9),
	.w6(32'hbbe4f19c),
	.w7(32'hb994349c),
	.w8(32'hbb32f81b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6acfe3),
	.w1(32'h39cdb627),
	.w2(32'hbb97f5c0),
	.w3(32'hbb684f4c),
	.w4(32'hba96ddf6),
	.w5(32'hbb623558),
	.w6(32'hbba238b6),
	.w7(32'hbb0cf99e),
	.w8(32'hbbd2f953),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4efcb),
	.w1(32'h3b77a255),
	.w2(32'h397cb7f6),
	.w3(32'hbb0a16d2),
	.w4(32'h3bb3bb96),
	.w5(32'h3aedc195),
	.w6(32'h3b76886b),
	.w7(32'hba43fe15),
	.w8(32'h3a2c4da4),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc086b60),
	.w1(32'hbb36d9f5),
	.w2(32'hbc802d4c),
	.w3(32'hbbb09289),
	.w4(32'h379ff537),
	.w5(32'hbc44b6d3),
	.w6(32'hbb737659),
	.w7(32'hbaa117b9),
	.w8(32'hbb8ab5e5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab573b7),
	.w1(32'hba0024b5),
	.w2(32'hbaed1ac9),
	.w3(32'hbb8587e2),
	.w4(32'h3abeca45),
	.w5(32'hbb227325),
	.w6(32'hbbbb0ef3),
	.w7(32'h39244a9d),
	.w8(32'hbba8dfb5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1cc3a),
	.w1(32'hbb2b8a42),
	.w2(32'hbb931046),
	.w3(32'hbbb1d00d),
	.w4(32'hbbb242d6),
	.w5(32'hbc0866b5),
	.w6(32'h3a3009da),
	.w7(32'h3a90a340),
	.w8(32'hbbc4be1c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44d565),
	.w1(32'h3b8f8bd7),
	.w2(32'hbb88127c),
	.w3(32'h3b2195f6),
	.w4(32'hba9528df),
	.w5(32'hbbb241f3),
	.w6(32'h3b87ac9e),
	.w7(32'hba35e4f6),
	.w8(32'h3c850870),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc01361),
	.w1(32'h3b017885),
	.w2(32'hbb5e532a),
	.w3(32'h3c8ff903),
	.w4(32'h3a8707e5),
	.w5(32'hbb36a465),
	.w6(32'h3b02cafb),
	.w7(32'h3ada9b63),
	.w8(32'hbb793514),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cc7a2),
	.w1(32'h3a1f0992),
	.w2(32'hb91693da),
	.w3(32'hbab92032),
	.w4(32'h3a866a54),
	.w5(32'hba3f7ea7),
	.w6(32'h3a11e9fe),
	.w7(32'hba083005),
	.w8(32'hbb0f26ee),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb346ffd),
	.w1(32'hba989dbb),
	.w2(32'hba106e26),
	.w3(32'hbb5741a6),
	.w4(32'hbb0276cc),
	.w5(32'hbb6ae2c0),
	.w6(32'hbb0009c9),
	.w7(32'hbb1aea31),
	.w8(32'hbbe34557),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d412b),
	.w1(32'hbaddcfd1),
	.w2(32'h3bf400e9),
	.w3(32'hbb9692a9),
	.w4(32'h3b754604),
	.w5(32'h3b0eae50),
	.w6(32'hbac960e2),
	.w7(32'h3b27b759),
	.w8(32'hba2f2e27),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eeae7),
	.w1(32'hbad612ba),
	.w2(32'hbba8a88a),
	.w3(32'hbbaa56d9),
	.w4(32'h3abd5eb1),
	.w5(32'hbb3b1adc),
	.w6(32'hbbc494cb),
	.w7(32'hbb8ebd97),
	.w8(32'hbbdc95d5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5e557),
	.w1(32'h3b9d071c),
	.w2(32'hbbbae54e),
	.w3(32'hbaa9b7e3),
	.w4(32'h3b829abf),
	.w5(32'hbaaa7502),
	.w6(32'h3b7f0ae8),
	.w7(32'hbb7804fa),
	.w8(32'h3aa5a27e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b217cbe),
	.w1(32'h39a806cb),
	.w2(32'hbb7abfcb),
	.w3(32'h3a91593e),
	.w4(32'hbaceb6c5),
	.w5(32'hbb143ded),
	.w6(32'hba00f986),
	.w7(32'hbab1b7ef),
	.w8(32'hba9b24e4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92f0e1),
	.w1(32'hbb9f6adf),
	.w2(32'hbc48490f),
	.w3(32'hbb9e01c7),
	.w4(32'hbb326d08),
	.w5(32'hbc336258),
	.w6(32'hbb1ad222),
	.w7(32'hbc2a4179),
	.w8(32'h3a623e5d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c46cd),
	.w1(32'h3a70db30),
	.w2(32'hbb8acba1),
	.w3(32'hbb800b22),
	.w4(32'h3a11e446),
	.w5(32'hbb12f78b),
	.w6(32'hbac42b11),
	.w7(32'hb851afcd),
	.w8(32'h38130173),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6bd5c),
	.w1(32'h3a04cf92),
	.w2(32'h3ac1bdfa),
	.w3(32'hbb5f9098),
	.w4(32'h3b2ea531),
	.w5(32'hb9895d45),
	.w6(32'h3b19d86b),
	.w7(32'hbacf9775),
	.w8(32'hbb8ae15b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3862fa),
	.w1(32'hba2bc7c5),
	.w2(32'hbac534f5),
	.w3(32'hbb1a1226),
	.w4(32'h3aac9276),
	.w5(32'hb97a0020),
	.w6(32'h395bef01),
	.w7(32'hba2a177a),
	.w8(32'hbad9ef49),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8901db),
	.w1(32'hbc1ac980),
	.w2(32'hbcb4e880),
	.w3(32'hbc80fdab),
	.w4(32'hbb41976e),
	.w5(32'hbc86adab),
	.w6(32'hbbf28074),
	.w7(32'hbb16eff9),
	.w8(32'hbc0f0d8b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18fb11),
	.w1(32'h3b5ae7ec),
	.w2(32'hba573a94),
	.w3(32'hbb105d39),
	.w4(32'h3c158d3d),
	.w5(32'h3b4c2cb1),
	.w6(32'hbb6fa22d),
	.w7(32'h3b9d9847),
	.w8(32'hbb16a06a),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb010524),
	.w1(32'h3aaabfef),
	.w2(32'h3a97387c),
	.w3(32'hbb12bdc6),
	.w4(32'h39d5c967),
	.w5(32'hba0430a6),
	.w6(32'h3b7c970d),
	.w7(32'h3ad80fbf),
	.w8(32'h399aed47),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5236dc),
	.w1(32'h39cab18b),
	.w2(32'hbb4049ed),
	.w3(32'hba8e84fa),
	.w4(32'hba5c31ff),
	.w5(32'h3b5105c8),
	.w6(32'h3ace21ee),
	.w7(32'hbad485db),
	.w8(32'hba6927e1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d4c98),
	.w1(32'h3b261056),
	.w2(32'h39a93e28),
	.w3(32'hba51b597),
	.w4(32'h3b6aef21),
	.w5(32'h3ad2fa57),
	.w6(32'h3b1b42bb),
	.w7(32'hba4239dc),
	.w8(32'h3a31c710),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b4b53),
	.w1(32'hbae19705),
	.w2(32'hba43fff9),
	.w3(32'h3a86dfb2),
	.w4(32'hb9cf10f9),
	.w5(32'hb9d5c1c9),
	.w6(32'hbae54d14),
	.w7(32'hba21d6c2),
	.w8(32'hba4dc05d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fb315),
	.w1(32'h3b94a62e),
	.w2(32'h39653d91),
	.w3(32'h3acf195c),
	.w4(32'h3b9676c9),
	.w5(32'hbb171e5f),
	.w6(32'h3b77050d),
	.w7(32'hbaf3b237),
	.w8(32'hbba0bfaf),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f3b51),
	.w1(32'hb7f67030),
	.w2(32'hbbed3865),
	.w3(32'hb9a76a87),
	.w4(32'h3b53dbda),
	.w5(32'hbbd7db94),
	.w6(32'h3a7b7caf),
	.w7(32'hbab05e8d),
	.w8(32'hb88b3d27),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e1dca),
	.w1(32'hbbc9e785),
	.w2(32'hbc0b1c55),
	.w3(32'hbb93fd92),
	.w4(32'hbc2d0b18),
	.w5(32'hbba8706c),
	.w6(32'hbc2d5e2b),
	.w7(32'h3b1030d0),
	.w8(32'hbbddfdbe),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a957835),
	.w1(32'h3a7259c5),
	.w2(32'h3b759856),
	.w3(32'hbbe5c0eb),
	.w4(32'h3aca1ce5),
	.w5(32'h3b165d6f),
	.w6(32'hbade79a4),
	.w7(32'h3a9140be),
	.w8(32'hbb31c191),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12d840),
	.w1(32'hbc0d0834),
	.w2(32'hbc00b17a),
	.w3(32'hbbf513d0),
	.w4(32'hbbe5801c),
	.w5(32'hbc1219d0),
	.w6(32'hbc21aaef),
	.w7(32'hbbdf2523),
	.w8(32'hbc71f399),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd69b04),
	.w1(32'hba8ddbbb),
	.w2(32'hbaa222b0),
	.w3(32'hbbd35ed4),
	.w4(32'h3a53ffe1),
	.w5(32'h39e55557),
	.w6(32'hba992ae2),
	.w7(32'hb989d66f),
	.w8(32'hb9d9bfb4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8303da),
	.w1(32'h39a44c9c),
	.w2(32'h3b2f8919),
	.w3(32'h39cd86a0),
	.w4(32'h3a46b93d),
	.w5(32'h3b0f9498),
	.w6(32'hb9c67c4e),
	.w7(32'h3af7efe1),
	.w8(32'hbb0e9e61),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4a695),
	.w1(32'h3a766d65),
	.w2(32'h3af76acf),
	.w3(32'hbb2a5cd0),
	.w4(32'h3abf619c),
	.w5(32'h3afe2234),
	.w6(32'h3aa8d592),
	.w7(32'h3afee4b6),
	.w8(32'hba9d62ff),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac3701),
	.w1(32'h38ec8821),
	.w2(32'h3a9d2ec1),
	.w3(32'hba82ff45),
	.w4(32'h39f6b03b),
	.w5(32'h3b019ff6),
	.w6(32'hbb31f083),
	.w7(32'h394cf53f),
	.w8(32'hbb4fa134),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f552c),
	.w1(32'h3a91e2de),
	.w2(32'h39141cd5),
	.w3(32'hbbcc4fb4),
	.w4(32'h3a93a9d6),
	.w5(32'hbb1d589f),
	.w6(32'hbb873533),
	.w7(32'hbb6afe58),
	.w8(32'hbb096107),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc83f24),
	.w1(32'h3c017574),
	.w2(32'h39bb110d),
	.w3(32'hbb5ab171),
	.w4(32'h3c03c048),
	.w5(32'h3b1e4ad0),
	.w6(32'hbb40bdbb),
	.w7(32'h3ba749a8),
	.w8(32'hbb6bc033),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3d5b1),
	.w1(32'h3b2c975a),
	.w2(32'hbb5c040e),
	.w3(32'hbb120168),
	.w4(32'h3b6aad3d),
	.w5(32'hbb1cc93b),
	.w6(32'hba533909),
	.w7(32'hb9d4e9fb),
	.w8(32'hbb880b64),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f55f0),
	.w1(32'h3b365c31),
	.w2(32'h3b175cac),
	.w3(32'hbb666851),
	.w4(32'h3b2d2eef),
	.w5(32'h3b664ad1),
	.w6(32'hba0ba14f),
	.w7(32'h3a23cbc2),
	.w8(32'h3ac758ce),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b376ddf),
	.w1(32'h3b4f5538),
	.w2(32'hbbc5e30f),
	.w3(32'h3ada4245),
	.w4(32'hbb35e933),
	.w5(32'hbb71f119),
	.w6(32'hbbb852ab),
	.w7(32'hbb36622f),
	.w8(32'hbba1758d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10ea7c),
	.w1(32'hbb52ffe1),
	.w2(32'hbb72befd),
	.w3(32'hbad7cdc3),
	.w4(32'hbad8f75b),
	.w5(32'hbb134ca6),
	.w6(32'hbb94d53a),
	.w7(32'h3a922787),
	.w8(32'hbba2b1ea),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e8309),
	.w1(32'hbc35ab97),
	.w2(32'hbc373c83),
	.w3(32'hbc751e7f),
	.w4(32'hbc1c1de7),
	.w5(32'hbba3e9bc),
	.w6(32'hbc5c06e2),
	.w7(32'hba85f04b),
	.w8(32'hbc0c80bd),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf81c6),
	.w1(32'hbb575d2d),
	.w2(32'h3887073e),
	.w3(32'hbb125649),
	.w4(32'hba9d9e13),
	.w5(32'hb83a58d6),
	.w6(32'hbb3e86bd),
	.w7(32'h3822ca49),
	.w8(32'hbaae67df),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fb87c),
	.w1(32'hba602a2e),
	.w2(32'hbad7412c),
	.w3(32'hb9aa8f77),
	.w4(32'hbac87ae8),
	.w5(32'hbb2fa567),
	.w6(32'hbab6d681),
	.w7(32'hbae2ff25),
	.w8(32'h3b6d0bfb),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a768fcc),
	.w1(32'hba7bc479),
	.w2(32'hbb4fdbf1),
	.w3(32'hb99c3030),
	.w4(32'h3b3052e3),
	.w5(32'hbad5401b),
	.w6(32'hbb8a5ec7),
	.w7(32'h398ed8ce),
	.w8(32'hbb87f1e4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1ce7d),
	.w1(32'h3b3cf121),
	.w2(32'hbc035fc2),
	.w3(32'hbaf8cc3a),
	.w4(32'hbb5dc137),
	.w5(32'hbc1b7af7),
	.w6(32'hba65c241),
	.w7(32'h3b9683bc),
	.w8(32'hbc0604c2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb228c07),
	.w1(32'hbb48086b),
	.w2(32'hbb962dba),
	.w3(32'hbbd6874f),
	.w4(32'h3a19575e),
	.w5(32'hbb94f873),
	.w6(32'hbb488a0d),
	.w7(32'h3b1aac14),
	.w8(32'h39c3d239),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98ea0e),
	.w1(32'h3b1f6ade),
	.w2(32'hbb0ff559),
	.w3(32'h3b3a7c8b),
	.w4(32'hba75103a),
	.w5(32'hbb9c574f),
	.w6(32'h3adb7be5),
	.w7(32'hbb2671c0),
	.w8(32'hbb0ed636),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9981831),
	.w1(32'hba979b6f),
	.w2(32'h3a2f42aa),
	.w3(32'h3abfc0f6),
	.w4(32'hb8890ad6),
	.w5(32'h3ae50b90),
	.w6(32'hbb050108),
	.w7(32'h3a810672),
	.w8(32'hba853d55),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb859e18e),
	.w1(32'hbac59093),
	.w2(32'hbb7471db),
	.w3(32'hbab3440a),
	.w4(32'hbac263a6),
	.w5(32'hbb565844),
	.w6(32'hbaa5db62),
	.w7(32'hbb46c092),
	.w8(32'hbae1cf4e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2769c3),
	.w1(32'hbac44478),
	.w2(32'hbac82911),
	.w3(32'hbb82ec32),
	.w4(32'hbb4936ea),
	.w5(32'hba8b2319),
	.w6(32'hbb607fc6),
	.w7(32'h3a612c42),
	.w8(32'hbbb85431),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ab104),
	.w1(32'hbc2a8e31),
	.w2(32'hbc5fae82),
	.w3(32'hbc67c1ea),
	.w4(32'hbc21703e),
	.w5(32'hbc4cb3f0),
	.w6(32'hbc5b2d62),
	.w7(32'hbbd1eebc),
	.w8(32'hbc2ea7b3),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add1d85),
	.w1(32'hba4736fc),
	.w2(32'hbb7d279e),
	.w3(32'h3a8c7a2d),
	.w4(32'h3999f891),
	.w5(32'hbb16a0e1),
	.w6(32'h3aab31c5),
	.w7(32'hb90bf7f4),
	.w8(32'hbac5b480),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae0469),
	.w1(32'h3b7abd32),
	.w2(32'h3a5ca4e9),
	.w3(32'h35678dd6),
	.w4(32'h3bb04dfa),
	.w5(32'h3b045de2),
	.w6(32'hbb823b57),
	.w7(32'h3a948e8f),
	.w8(32'hb99f6495),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde93e7),
	.w1(32'hbbd3d6e6),
	.w2(32'hbbcc5f06),
	.w3(32'hbb84aef7),
	.w4(32'hbb98fcd5),
	.w5(32'hb9845b3e),
	.w6(32'hbbdeebad),
	.w7(32'h3b26f45b),
	.w8(32'h3aa5cb55),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9097ed7),
	.w1(32'hbafe2a30),
	.w2(32'hba4f55e9),
	.w3(32'hbb4d7167),
	.w4(32'hba6b8134),
	.w5(32'hb9c57e55),
	.w6(32'hbb1b885b),
	.w7(32'hbaa418a9),
	.w8(32'hbb19e93c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba951462),
	.w1(32'h3a8a2a4a),
	.w2(32'hba524a76),
	.w3(32'hbacce691),
	.w4(32'hb94b411a),
	.w5(32'hba92d36f),
	.w6(32'hb9a26b6e),
	.w7(32'hbb397099),
	.w8(32'hbb08f594),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88fb36),
	.w1(32'hbaac97dc),
	.w2(32'h3ce747f2),
	.w3(32'hba6d6f24),
	.w4(32'hbc06b7a4),
	.w5(32'h3d0899f8),
	.w6(32'hbb5191b9),
	.w7(32'h3d0643de),
	.w8(32'hbb9daed4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d949e1),
	.w1(32'hba3b9dda),
	.w2(32'hbab28029),
	.w3(32'hbb84a1bc),
	.w4(32'hb997d338),
	.w5(32'hbafbc14d),
	.w6(32'h3a8c6ff1),
	.w7(32'hbb22c270),
	.w8(32'hba101778),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d71d5),
	.w1(32'hbac1e5a5),
	.w2(32'hb9afb39f),
	.w3(32'hbae06167),
	.w4(32'h38afa763),
	.w5(32'h3a5d9e01),
	.w6(32'hbb2c4081),
	.w7(32'hba0e1039),
	.w8(32'hbb177170),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae051ed),
	.w1(32'h3a4c3bee),
	.w2(32'hbc037b4d),
	.w3(32'hbaa23cd7),
	.w4(32'h3b20a983),
	.w5(32'hbbbf9f4b),
	.w6(32'hbaaaf6dc),
	.w7(32'hba929dea),
	.w8(32'hbb491afc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ff306),
	.w1(32'hbb290d2b),
	.w2(32'hbb323268),
	.w3(32'hb8ec2a60),
	.w4(32'hba211a23),
	.w5(32'hbb119ef5),
	.w6(32'hbb908e3e),
	.w7(32'hbbfa143a),
	.w8(32'hbc08f6b7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f6f27),
	.w1(32'hbb0c8dcf),
	.w2(32'h3baa06b8),
	.w3(32'hbb880fe4),
	.w4(32'hb87d0b6d),
	.w5(32'h3b2099b5),
	.w6(32'hbb3eb964),
	.w7(32'h38239a58),
	.w8(32'h3b19e290),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd0789),
	.w1(32'h3a20a8a5),
	.w2(32'hbc07f399),
	.w3(32'hbae4c26e),
	.w4(32'hb93c683b),
	.w5(32'hbc0b1223),
	.w6(32'h3a62243f),
	.w7(32'hbb2ffd7e),
	.w8(32'hbc111bef),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23b723),
	.w1(32'hba20d11a),
	.w2(32'hbac6296c),
	.w3(32'hbb8764b1),
	.w4(32'hba0df69f),
	.w5(32'hbab29277),
	.w6(32'hba826ae5),
	.w7(32'h3a2b2c5e),
	.w8(32'hbb8a0e1a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b1894),
	.w1(32'h3b08cb32),
	.w2(32'hb96cbf5f),
	.w3(32'hbae6f222),
	.w4(32'h3b05f96f),
	.w5(32'hb80fcf68),
	.w6(32'h3b03bcf3),
	.w7(32'h390f0bc3),
	.w8(32'hba5f60c1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb165275),
	.w1(32'hb9aded27),
	.w2(32'hbaa66efe),
	.w3(32'hbb2c6814),
	.w4(32'hb804ceb4),
	.w5(32'hb92b6385),
	.w6(32'hba96af6b),
	.w7(32'h393ce0f6),
	.w8(32'hbb0ec76b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acaa9ce),
	.w1(32'hbac422fa),
	.w2(32'hba7ab7c3),
	.w3(32'h39cf97eb),
	.w4(32'hb9eab383),
	.w5(32'hb9e5308c),
	.w6(32'hbb065ac1),
	.w7(32'hba6ebfe9),
	.w8(32'hbad4ef83),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c2b6f),
	.w1(32'hbaccb72c),
	.w2(32'h3aa50424),
	.w3(32'hbb0bf15c),
	.w4(32'hba816e48),
	.w5(32'h3aeaddb3),
	.w6(32'hbb6a465e),
	.w7(32'h398c659d),
	.w8(32'hbb0cbf49),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1a50f),
	.w1(32'h3ad63ada),
	.w2(32'hb9426aae),
	.w3(32'hba20cd15),
	.w4(32'h3adfd47d),
	.w5(32'hb901275e),
	.w6(32'h3afc4145),
	.w7(32'h38e0e45c),
	.w8(32'hba70bd93),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba589ba4),
	.w1(32'h3b4c9ac7),
	.w2(32'hbb049390),
	.w3(32'hbad1bbd1),
	.w4(32'h3ab9836e),
	.w5(32'hb971e165),
	.w6(32'h3a922785),
	.w7(32'hb9a00477),
	.w8(32'h3a596c36),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b181c9),
	.w1(32'h3ac8f44a),
	.w2(32'h3b3edf5d),
	.w3(32'hbaec3c56),
	.w4(32'h3b75c35f),
	.w5(32'h3b4a3fb0),
	.w6(32'hbaff9fc3),
	.w7(32'h3a4813c6),
	.w8(32'hbad1f785),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2de9f6),
	.w1(32'hb7a39507),
	.w2(32'hbc8cd4c5),
	.w3(32'hbb684f3d),
	.w4(32'hb7b85f78),
	.w5(32'hbc40933d),
	.w6(32'hb9ac4303),
	.w7(32'hbc116337),
	.w8(32'hbbceeeb1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36af43),
	.w1(32'hba4f0ebf),
	.w2(32'hbbb52b79),
	.w3(32'hbab5b154),
	.w4(32'h3a9b0036),
	.w5(32'hbba12574),
	.w6(32'hb8aeb470),
	.w7(32'h3a2af98b),
	.w8(32'hbb9e9933),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc35fc0),
	.w1(32'hbbc2931c),
	.w2(32'hbc01bef2),
	.w3(32'hbbe16572),
	.w4(32'hbb9143e7),
	.w5(32'hbc24d1ed),
	.w6(32'hbbe541df),
	.w7(32'hbbc8cd4a),
	.w8(32'hbc3c92d8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fcfb6),
	.w1(32'h3b6f40a9),
	.w2(32'hbb1ee82d),
	.w3(32'hbb83183b),
	.w4(32'hb976e7e7),
	.w5(32'hbb2576da),
	.w6(32'h3a981a1b),
	.w7(32'hbb3549bc),
	.w8(32'hba2f80c1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f9b93),
	.w1(32'h3b2efec2),
	.w2(32'hb9b3b8c1),
	.w3(32'hba5a5439),
	.w4(32'h3b349da2),
	.w5(32'hb8d89ca8),
	.w6(32'h3b470a0d),
	.w7(32'h395c3662),
	.w8(32'hba95c60e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6000db),
	.w1(32'h3a94f582),
	.w2(32'h3a1fbf31),
	.w3(32'hbb00f419),
	.w4(32'h3ae507a3),
	.w5(32'h3a8c911c),
	.w6(32'h3a0aaa8e),
	.w7(32'h3aa105fb),
	.w8(32'hba3b2a61),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3749a2f6),
	.w1(32'h3b111c10),
	.w2(32'h39d081b0),
	.w3(32'hba86cc9c),
	.w4(32'h3b3983ed),
	.w5(32'h3a68d1c9),
	.w6(32'h3a9b06ee),
	.w7(32'h3a02e0e0),
	.w8(32'hb9e33270),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d8ef7),
	.w1(32'hb8d2407d),
	.w2(32'hbbcffa0a),
	.w3(32'hb80c58a8),
	.w4(32'h3a9b8d15),
	.w5(32'hbbc3f9fa),
	.w6(32'h3ad06a88),
	.w7(32'hbb233d62),
	.w8(32'hbb825115),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86cc00),
	.w1(32'h3a61e760),
	.w2(32'h3b0baa9a),
	.w3(32'hbb38204c),
	.w4(32'h3b320c94),
	.w5(32'h3b08268c),
	.w6(32'h3a9a0c3c),
	.w7(32'h3a9b7ecd),
	.w8(32'h3a087bed),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3895e8f2),
	.w1(32'h3b06746a),
	.w2(32'h39ea2887),
	.w3(32'hb9b9f0b0),
	.w4(32'h3b4ec2a0),
	.w5(32'h3b5198d2),
	.w6(32'hbb711ca1),
	.w7(32'hbb11b35f),
	.w8(32'hbb8df63b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad383c),
	.w1(32'h39817bc7),
	.w2(32'h3b3f1922),
	.w3(32'hbb2d731a),
	.w4(32'h3b32abd6),
	.w5(32'h3b89faea),
	.w6(32'hbb1215eb),
	.w7(32'h3a5be90d),
	.w8(32'hb9f26270),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b038d73),
	.w1(32'h3aaa6e3d),
	.w2(32'h3aa026bb),
	.w3(32'h3aaa5070),
	.w4(32'h3aef32e5),
	.w5(32'h3a9f58a7),
	.w6(32'h3a54c0e3),
	.w7(32'h3a78e5e1),
	.w8(32'hbaec1e44),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b3e5a),
	.w1(32'hbab18f9a),
	.w2(32'h3b392311),
	.w3(32'hbb7cc4e1),
	.w4(32'h3a24061c),
	.w5(32'h38d8ac43),
	.w6(32'hbb2f4fa9),
	.w7(32'hbad18b58),
	.w8(32'hbb47ab1a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94490e),
	.w1(32'h3b811530),
	.w2(32'hbb020544),
	.w3(32'hba7786df),
	.w4(32'h3bc3f968),
	.w5(32'h3a851678),
	.w6(32'h3a52dec6),
	.w7(32'hbae4bf57),
	.w8(32'h3a1c4d5b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa35768),
	.w1(32'hbb4e2e1a),
	.w2(32'hbbc31dcb),
	.w3(32'hba991a19),
	.w4(32'hbac42361),
	.w5(32'hbb29b5a4),
	.w6(32'hbb913d06),
	.w7(32'h3a289edc),
	.w8(32'hbbb28781),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31bf11),
	.w1(32'h3b6a9722),
	.w2(32'hbb81e7ed),
	.w3(32'hba8c2c18),
	.w4(32'h3b6eeff4),
	.w5(32'hbaf0e44a),
	.w6(32'h3b970c19),
	.w7(32'hb9a8f5d0),
	.w8(32'h3a263ff2),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d7af3),
	.w1(32'h3a98d027),
	.w2(32'hba68294c),
	.w3(32'h399989c7),
	.w4(32'h3b817e3f),
	.w5(32'h3b2afe08),
	.w6(32'hbb93ae3e),
	.w7(32'h3b1a62ff),
	.w8(32'h3b7365f9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule