module layer_8_featuremap_95(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a0583),
	.w1(32'h3c042083),
	.w2(32'h3bb3bc1b),
	.w3(32'h3ba112b1),
	.w4(32'h3b9f5b3c),
	.w5(32'h3b30b92d),
	.w6(32'h3a2674c5),
	.w7(32'h3b0dcd9a),
	.w8(32'hb9b0def6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2653b),
	.w1(32'hb973e9d8),
	.w2(32'h3aed980e),
	.w3(32'hbba551c9),
	.w4(32'h3662ca94),
	.w5(32'h3b254f14),
	.w6(32'hbb9e7cbd),
	.w7(32'h395d0d82),
	.w8(32'h3b0e0496),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb88e71),
	.w1(32'h3b5cbbc8),
	.w2(32'h3bc5cd78),
	.w3(32'hbbd1d1ab),
	.w4(32'h3b77e4df),
	.w5(32'h3bd3c186),
	.w6(32'hbbdf87b1),
	.w7(32'h3b2ce274),
	.w8(32'h3bb6c5a0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91d9966),
	.w1(32'h3b3b80cd),
	.w2(32'hbb4bbb97),
	.w3(32'hbb705e11),
	.w4(32'h3aa51649),
	.w5(32'hba8c8121),
	.w6(32'hbb56a84e),
	.w7(32'hbb30b92c),
	.w8(32'hbc0f08a8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fc0b5),
	.w1(32'hbb1b0643),
	.w2(32'hbada19b0),
	.w3(32'hbb6f1381),
	.w4(32'hb9ea76a6),
	.w5(32'hba365cc4),
	.w6(32'hbb99f992),
	.w7(32'hba88d59a),
	.w8(32'hb89bbe36),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc566d24),
	.w1(32'hba113a8b),
	.w2(32'h37e9f4e5),
	.w3(32'hbc395c76),
	.w4(32'h3af0f288),
	.w5(32'h3b2ad460),
	.w6(32'hbc27c150),
	.w7(32'hba05fa3a),
	.w8(32'hbab68488),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3958f441),
	.w1(32'hb660c507),
	.w2(32'h37776139),
	.w3(32'h39570b00),
	.w4(32'h37c4bfee),
	.w5(32'hb7563ed5),
	.w6(32'h3972a3a1),
	.w7(32'h38193e87),
	.w8(32'h36acdc9b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8f0e9),
	.w1(32'h3b390743),
	.w2(32'h3b4170b4),
	.w3(32'hbb4f764e),
	.w4(32'h3b9065f2),
	.w5(32'h3b3bf089),
	.w6(32'hbb3b48bb),
	.w7(32'h3ba5ce96),
	.w8(32'h3b6c2898),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a98e2),
	.w1(32'hba5c55ab),
	.w2(32'h3a8b2548),
	.w3(32'hbb4ff378),
	.w4(32'h3aa61426),
	.w5(32'h3b5c4e58),
	.w6(32'hbb948ab1),
	.w7(32'h39efe8c9),
	.w8(32'h3ab33e74),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ba952),
	.w1(32'h3bed3264),
	.w2(32'h3bf9b1ad),
	.w3(32'h3b0b34da),
	.w4(32'h3c046c62),
	.w5(32'h3c09cbc5),
	.w6(32'hbaa23873),
	.w7(32'h3bc79881),
	.w8(32'h3bc87ddb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce8791),
	.w1(32'h3bb0092a),
	.w2(32'h3b0f6ede),
	.w3(32'h3b696c14),
	.w4(32'h3b93764f),
	.w5(32'h3b1182ab),
	.w6(32'hbabb1c26),
	.w7(32'h39727008),
	.w8(32'hbb712f9f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb05a5a),
	.w1(32'hb9b0f3af),
	.w2(32'hbaf1109b),
	.w3(32'hbbb3b6d8),
	.w4(32'hb8fce0aa),
	.w5(32'hbb2a866b),
	.w6(32'hbbd7c16a),
	.w7(32'hbae68060),
	.w8(32'hbb07ea59),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e22a7),
	.w1(32'h39e1b371),
	.w2(32'hb986043d),
	.w3(32'hbc12ee53),
	.w4(32'hbab763e7),
	.w5(32'hbbed6310),
	.w6(32'hbbedcd28),
	.w7(32'h394d7c70),
	.w8(32'h3c00a2d6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9bf3a),
	.w1(32'h3b25e55c),
	.w2(32'h3b14aada),
	.w3(32'hbb2a4d0a),
	.w4(32'hbb0de1b7),
	.w5(32'h38d4162a),
	.w6(32'h3b28d4db),
	.w7(32'hba6e2ab2),
	.w8(32'h3a7d5f6e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61695f),
	.w1(32'h3b0c1d45),
	.w2(32'h3ba3a281),
	.w3(32'h3b987a49),
	.w4(32'h3b110520),
	.w5(32'hba4df29b),
	.w6(32'h3b621e75),
	.w7(32'h3bc9fea3),
	.w8(32'h3a4bcc0b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a9845),
	.w1(32'h39eb4827),
	.w2(32'hba5cc85b),
	.w3(32'h39091e55),
	.w4(32'h3bdd0b05),
	.w5(32'h3bbf83f8),
	.w6(32'hb7d2da12),
	.w7(32'h3c4b3c8a),
	.w8(32'h3d062de8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb669067),
	.w1(32'hbb9c1dad),
	.w2(32'h3bd88410),
	.w3(32'hbb9649c6),
	.w4(32'h3ab5fcc3),
	.w5(32'h3c1a6fb5),
	.w6(32'h3c792dd9),
	.w7(32'h3b673564),
	.w8(32'hbb1cbaa9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a2633),
	.w1(32'hbc01e0ef),
	.w2(32'h3ab6ccd3),
	.w3(32'hba952b44),
	.w4(32'hb9b68c22),
	.w5(32'hbc354185),
	.w6(32'hbc80f45b),
	.w7(32'h3ca0c8c0),
	.w8(32'hbc1b159c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be28b0a),
	.w1(32'h3c295129),
	.w2(32'h3a81e3d3),
	.w3(32'hbc8d54f3),
	.w4(32'hbc8a24ef),
	.w5(32'hbb80899e),
	.w6(32'hbcb11031),
	.w7(32'hbc39a787),
	.w8(32'hbcc923eb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc201c23),
	.w1(32'hbc000818),
	.w2(32'hbc1cf978),
	.w3(32'hbc6efb8c),
	.w4(32'hbb1355c7),
	.w5(32'hbcc5137e),
	.w6(32'hbcb9f567),
	.w7(32'hbc0b6cfc),
	.w8(32'hbcbcc1f3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c059fc3),
	.w1(32'hbad4b8b3),
	.w2(32'h3b99a7a2),
	.w3(32'hbbe970fc),
	.w4(32'hbcc08797),
	.w5(32'hbae24477),
	.w6(32'hbcbbcfe7),
	.w7(32'hbc3e9755),
	.w8(32'h3c9cc88a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19be47),
	.w1(32'hbc10f390),
	.w2(32'h3c187d5d),
	.w3(32'h3c4bfae7),
	.w4(32'hbbfa674a),
	.w5(32'hbc5d62a5),
	.w6(32'h3cc391a1),
	.w7(32'h3c2a77b7),
	.w8(32'h3c38ce20),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc721d3),
	.w1(32'h3c23d917),
	.w2(32'h3c392b1d),
	.w3(32'h3c570056),
	.w4(32'h3cb2fdbe),
	.w5(32'h3d039c34),
	.w6(32'h3c7f7dc7),
	.w7(32'h3c5b3ffe),
	.w8(32'h3ca3c805),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38fd91),
	.w1(32'hbbe22861),
	.w2(32'h3b3f67e4),
	.w3(32'hbb2d2ad0),
	.w4(32'h3bf5de46),
	.w5(32'h3c00013a),
	.w6(32'hbc3e70ba),
	.w7(32'h3c0e5f0b),
	.w8(32'h3b6d7cd1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b858622),
	.w1(32'hba0d55a7),
	.w2(32'h3b8ee80f),
	.w3(32'hbb5952c1),
	.w4(32'hbaf2ccf9),
	.w5(32'h3b64c502),
	.w6(32'hbb935123),
	.w7(32'hbb8de359),
	.w8(32'h3b28bb06),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c795e1d),
	.w1(32'h3c82260a),
	.w2(32'h3be2acd9),
	.w3(32'h3b879bca),
	.w4(32'h3c9f3bd1),
	.w5(32'h3d0ee71c),
	.w6(32'hbb60e68d),
	.w7(32'hbc94c670),
	.w8(32'hbd8777b7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c4c6e),
	.w1(32'h3c4a68b2),
	.w2(32'h3c672dac),
	.w3(32'h3c42db3b),
	.w4(32'hbc94470c),
	.w5(32'hbc308f06),
	.w6(32'hbd24c85d),
	.w7(32'hb97a9ea0),
	.w8(32'hbba0163c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90ab0c),
	.w1(32'h3ca6cb09),
	.w2(32'hbc652005),
	.w3(32'hbc9e7cf4),
	.w4(32'h3ae9951b),
	.w5(32'h3d0ec151),
	.w6(32'hbd117e6a),
	.w7(32'hbd624767),
	.w8(32'hbc9467f8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc10465),
	.w1(32'hbc521c90),
	.w2(32'h3c4f3516),
	.w3(32'h3c52a6dc),
	.w4(32'h3b04ea57),
	.w5(32'h3b2e512b),
	.w6(32'hbc495588),
	.w7(32'hbb2af31a),
	.w8(32'hbbd8a948),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3483d8),
	.w1(32'hbc1c4223),
	.w2(32'hbce3c767),
	.w3(32'h3c042d8e),
	.w4(32'h3b94bd7c),
	.w5(32'hbba62734),
	.w6(32'hbb802299),
	.w7(32'h3c762660),
	.w8(32'h3cab420b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19981b),
	.w1(32'hbc002031),
	.w2(32'h3b3e5a31),
	.w3(32'h3b62b9cd),
	.w4(32'hbaf339e9),
	.w5(32'hbaa8ffff),
	.w6(32'h3c5e4bea),
	.w7(32'h3b315acf),
	.w8(32'h3ad7020f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54db34),
	.w1(32'h3b16073d),
	.w2(32'hbc879e4b),
	.w3(32'hbb5ba02c),
	.w4(32'hbc36dbc0),
	.w5(32'hbcfa9922),
	.w6(32'hbb6fd6f9),
	.w7(32'h3c04c1f4),
	.w8(32'h3d505b76),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a230b),
	.w1(32'hbc8f5fd4),
	.w2(32'hbbf5782c),
	.w3(32'hbceaf55a),
	.w4(32'hbc80b2c4),
	.w5(32'hbcda9367),
	.w6(32'h3cacde87),
	.w7(32'h3cbfee68),
	.w8(32'h3d063870),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4336e7),
	.w1(32'h3a68d940),
	.w2(32'h3be53c3d),
	.w3(32'hbcb65d33),
	.w4(32'hbbdaa307),
	.w5(32'hbc1a6d6d),
	.w6(32'h3c895a50),
	.w7(32'h3c5015cf),
	.w8(32'hbc3e45ff),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0837dd),
	.w1(32'h3b782dcb),
	.w2(32'hba65030e),
	.w3(32'hbc90df45),
	.w4(32'h3ae85970),
	.w5(32'hbbf8ce02),
	.w6(32'hbc708a3f),
	.w7(32'h3bacd28c),
	.w8(32'hbafe4c03),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad98072),
	.w1(32'h3be551af),
	.w2(32'hbca0550e),
	.w3(32'hbb43b9aa),
	.w4(32'h3c942b07),
	.w5(32'hbc8d89ab),
	.w6(32'h3a14289b),
	.w7(32'h3cfd8893),
	.w8(32'hbb99f4d2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c7533),
	.w1(32'h3cb41089),
	.w2(32'hbccbb850),
	.w3(32'hbcb413c9),
	.w4(32'hbc9fd272),
	.w5(32'hbc31e629),
	.w6(32'hbc198d5e),
	.w7(32'hbb5a0fc7),
	.w8(32'h3d15b06c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc585564),
	.w1(32'hbcc72331),
	.w2(32'h3c42a43e),
	.w3(32'hbcb8da05),
	.w4(32'h3a6e6c1b),
	.w5(32'h3c1e90ad),
	.w6(32'h3cad025b),
	.w7(32'hbbe33e8f),
	.w8(32'h3accbd13),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33510c),
	.w1(32'hbac4fcb0),
	.w2(32'hbb45aed2),
	.w3(32'h3b9fbedb),
	.w4(32'h3b7f73d4),
	.w5(32'h39fbcfb8),
	.w6(32'h3c36ed6d),
	.w7(32'h3c1d6230),
	.w8(32'h3c172380),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f602a),
	.w1(32'hbbddd95f),
	.w2(32'hbb806303),
	.w3(32'h3c28bda3),
	.w4(32'hbc14bd44),
	.w5(32'hbc620e70),
	.w6(32'h3bb1baee),
	.w7(32'hbc5facb5),
	.w8(32'hbc2d484a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf52357),
	.w1(32'hbb7774a1),
	.w2(32'hbbc0fb08),
	.w3(32'hbd3394a2),
	.w4(32'h3ad23da5),
	.w5(32'hbc175494),
	.w6(32'hbd51e73c),
	.w7(32'h3b87341c),
	.w8(32'hbc731e96),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf5f68),
	.w1(32'h3bd33d66),
	.w2(32'hbb42d821),
	.w3(32'hbb3995b6),
	.w4(32'h3a02694e),
	.w5(32'h3ceafd2c),
	.w6(32'hbc4f3484),
	.w7(32'hbbbd21b3),
	.w8(32'h39b5e719),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba99042),
	.w1(32'hb8fd190b),
	.w2(32'h3b918fb9),
	.w3(32'h3c286673),
	.w4(32'hbc9ef2ef),
	.w5(32'hbccae673),
	.w6(32'hbc3f97bd),
	.w7(32'h3c192e75),
	.w8(32'h3d82cf3c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31450f),
	.w1(32'hbbcb69a9),
	.w2(32'hba94d925),
	.w3(32'hbc8a1b3b),
	.w4(32'h3a6c4520),
	.w5(32'hbbd6486f),
	.w6(32'h3cf1b96f),
	.w7(32'hb7b30231),
	.w8(32'h3a7fb7a1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b519906),
	.w1(32'h3be2aefd),
	.w2(32'h39e81b28),
	.w3(32'hbb47db48),
	.w4(32'h3c2e6f2f),
	.w5(32'h3cd09bd9),
	.w6(32'hbbaa39c7),
	.w7(32'hbb77651b),
	.w8(32'hbc4129f8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc851b33),
	.w1(32'hb9973eec),
	.w2(32'hbc05a180),
	.w3(32'h3cb1d2ea),
	.w4(32'h3cc9d227),
	.w5(32'h3c0dc68f),
	.w6(32'hbbbd5f56),
	.w7(32'h3c1fcd9a),
	.w8(32'h3b7bb780),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc342c74),
	.w1(32'h3bb723d6),
	.w2(32'h3b55fefc),
	.w3(32'hbc4e99b8),
	.w4(32'h3bb554c7),
	.w5(32'hbc3fdc76),
	.w6(32'hbc1537cf),
	.w7(32'hbc72a00a),
	.w8(32'hbba5341c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01c73f),
	.w1(32'hbb73c4c2),
	.w2(32'h3c0f2d13),
	.w3(32'hbb92fb08),
	.w4(32'hbb729862),
	.w5(32'h3c8af7d7),
	.w6(32'hbbd309b2),
	.w7(32'h3c009465),
	.w8(32'h3c01adbe),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1de2d),
	.w1(32'hb9be2e1c),
	.w2(32'h3c03f907),
	.w3(32'h3b0bcb3f),
	.w4(32'hba363177),
	.w5(32'h3bf67822),
	.w6(32'h3b85278b),
	.w7(32'hbb323392),
	.w8(32'hbc63335d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72588d),
	.w1(32'h3c48e735),
	.w2(32'hbc8eb251),
	.w3(32'hbb00a600),
	.w4(32'hbbcc8d83),
	.w5(32'h3b4f106d),
	.w6(32'hbcae0729),
	.w7(32'hbcab133f),
	.w8(32'hbc97965a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd362eb),
	.w1(32'hbcc23214),
	.w2(32'h3a9feb89),
	.w3(32'hbcc162e9),
	.w4(32'h3c89a9b8),
	.w5(32'h3d19831e),
	.w6(32'hbcfe79bf),
	.w7(32'hbcab1fa6),
	.w8(32'hbd214c49),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0ac0de),
	.w1(32'hbc3a1789),
	.w2(32'hbbaf1c9e),
	.w3(32'h3c3253c8),
	.w4(32'hbcac23da),
	.w5(32'hbc778a73),
	.w6(32'hbd335d17),
	.w7(32'hbcea4464),
	.w8(32'hbc8fd325),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc21d30),
	.w1(32'hbc861b68),
	.w2(32'hbbe1bdfa),
	.w3(32'h3c415af0),
	.w4(32'hbad3a280),
	.w5(32'hbbd96ae1),
	.w6(32'h3c9213b6),
	.w7(32'hbc2198c1),
	.w8(32'hbc398df1),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03626e),
	.w1(32'h3ba87e08),
	.w2(32'hbb6648ba),
	.w3(32'hbb31ccff),
	.w4(32'hba6e7192),
	.w5(32'hbb806e03),
	.w6(32'hbbd3ab70),
	.w7(32'hbb7c9885),
	.w8(32'hbb5effc5),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1deb10),
	.w1(32'h3a869aa2),
	.w2(32'hbc268691),
	.w3(32'h39d5ae77),
	.w4(32'h3c52ee80),
	.w5(32'h3cb924b8),
	.w6(32'hba3ac20f),
	.w7(32'hbbdfbe9b),
	.w8(32'hbccc4b79),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c91e2),
	.w1(32'h3b25c9a2),
	.w2(32'h3c56c4c1),
	.w3(32'hbc055fa7),
	.w4(32'h3bcd3cdd),
	.w5(32'h3c22d82c),
	.w6(32'hbc9df01e),
	.w7(32'h3bc58333),
	.w8(32'hbc5dbe91),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e4fe6),
	.w1(32'hbb2bb081),
	.w2(32'h3b81d2a5),
	.w3(32'h3b8216f6),
	.w4(32'hbc462f16),
	.w5(32'hbc0d5f4b),
	.w6(32'hbc2a0a03),
	.w7(32'hbb35546a),
	.w8(32'hbb5d9b6b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a497e),
	.w1(32'h3b8a424a),
	.w2(32'hbc6334e2),
	.w3(32'hbc43881d),
	.w4(32'h3cd7dcbb),
	.w5(32'h3d2e0fcf),
	.w6(32'hbc248160),
	.w7(32'hbb66f5d5),
	.w8(32'hba337296),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca026e),
	.w1(32'h3bd683d6),
	.w2(32'h3b888243),
	.w3(32'h3d1ac71b),
	.w4(32'h3b4d1b67),
	.w5(32'h3a2fd2ae),
	.w6(32'hbaa7c369),
	.w7(32'h3b5f78e0),
	.w8(32'h3bdbb5a1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99b4e3),
	.w1(32'hbae2c0a0),
	.w2(32'h3c6294b4),
	.w3(32'hbbe6c8a1),
	.w4(32'hbc0d6f52),
	.w5(32'h3bab7169),
	.w6(32'hbbe0bda3),
	.w7(32'hbc101f84),
	.w8(32'hbce14721),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f7b1e),
	.w1(32'h3c83e4b8),
	.w2(32'hbc049d32),
	.w3(32'h3b253ac6),
	.w4(32'h3c7aac7a),
	.w5(32'h3c2f42b9),
	.w6(32'hbc7478f3),
	.w7(32'h3b6559ff),
	.w8(32'hbcb62dae),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa906ff),
	.w1(32'h3c329824),
	.w2(32'h3b8d5074),
	.w3(32'h3c4026ea),
	.w4(32'hb8054906),
	.w5(32'hbad37ba4),
	.w6(32'hbc91f59f),
	.w7(32'h39b4bf61),
	.w8(32'h3ac84cf0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d9838),
	.w1(32'hbc048c5b),
	.w2(32'h3b22e3a0),
	.w3(32'hbcbce114),
	.w4(32'h3c0aa721),
	.w5(32'hbbda0822),
	.w6(32'hbcb4ef3e),
	.w7(32'hbc48abc6),
	.w8(32'hbccd299e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dc4d9),
	.w1(32'h3ad87097),
	.w2(32'hbbf2852b),
	.w3(32'hbb73cdbb),
	.w4(32'hbb895957),
	.w5(32'hbbe802c0),
	.w6(32'h3bfa8497),
	.w7(32'hbbe8a51f),
	.w8(32'h3baa8878),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66a608),
	.w1(32'hbb0aa75b),
	.w2(32'h389df21a),
	.w3(32'h3bd2520c),
	.w4(32'hbc45a86a),
	.w5(32'hbb7e10c5),
	.w6(32'hbc1069e3),
	.w7(32'hbcac49e2),
	.w8(32'h3a5f1b92),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c1d36),
	.w1(32'h3b1c592c),
	.w2(32'h3bf340bd),
	.w3(32'hbc20f930),
	.w4(32'h3a320ad9),
	.w5(32'hbac67e6c),
	.w6(32'hbc18ac34),
	.w7(32'h3befcf85),
	.w8(32'h3bdf333a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9b652),
	.w1(32'h3c5ade35),
	.w2(32'h3bbf3e89),
	.w3(32'hbc70f8ae),
	.w4(32'h3c48f13a),
	.w5(32'hbb76bf5a),
	.w6(32'hbbac929e),
	.w7(32'hbc209c28),
	.w8(32'hbc807b4d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50b191),
	.w1(32'hbbe86c7f),
	.w2(32'h3c1bcba0),
	.w3(32'hbbb6999f),
	.w4(32'hbcba84f9),
	.w5(32'hbce60850),
	.w6(32'hbc8880c8),
	.w7(32'h3ce07a99),
	.w8(32'h3d06ffcd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0aead),
	.w1(32'h3af35b6a),
	.w2(32'hbc5aaba1),
	.w3(32'hbcd69fc3),
	.w4(32'h3bc9cce0),
	.w5(32'h3c5c84f8),
	.w6(32'h3c42123c),
	.w7(32'hbaec4a25),
	.w8(32'h3a310185),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6a4b),
	.w1(32'hbbd94b95),
	.w2(32'h3c1f3a18),
	.w3(32'h3b365179),
	.w4(32'h3cacb81a),
	.w5(32'h3b788129),
	.w6(32'hbc20cab6),
	.w7(32'h3c1425cc),
	.w8(32'h3ba08ad1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd23e36),
	.w1(32'h3b9a4449),
	.w2(32'h3bc9277a),
	.w3(32'hbbe128c0),
	.w4(32'h3bbcb431),
	.w5(32'hbae7cfa2),
	.w6(32'h3bdc32a7),
	.w7(32'h3bb0d66d),
	.w8(32'h3b89c63b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e8133),
	.w1(32'h3b6a0524),
	.w2(32'hbb8dfe23),
	.w3(32'hbc1b555c),
	.w4(32'h3ba4d025),
	.w5(32'h3a44a225),
	.w6(32'hbc757116),
	.w7(32'h3b6abf09),
	.w8(32'hbc223df8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a4e3e),
	.w1(32'h3c4623fa),
	.w2(32'hbc556384),
	.w3(32'h3bc5b433),
	.w4(32'hbc166151),
	.w5(32'hbc0a5892),
	.w6(32'hbc6b1b45),
	.w7(32'hbbac996d),
	.w8(32'h3ca8aa85),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6810bc),
	.w1(32'hbbcec94d),
	.w2(32'h3c637f92),
	.w3(32'hbca527d3),
	.w4(32'hbbfb63b1),
	.w5(32'hbcac2113),
	.w6(32'hbc6323f3),
	.w7(32'hbb8d5eea),
	.w8(32'hbb736c6e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56c5bd),
	.w1(32'h3bd65874),
	.w2(32'h3bb3d70e),
	.w3(32'hbb26be11),
	.w4(32'h3aa9c12f),
	.w5(32'hbb9976fe),
	.w6(32'h3b6aaa08),
	.w7(32'hbb3e0f83),
	.w8(32'h3b054a39),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cc1b8),
	.w1(32'hbb0cfbc0),
	.w2(32'hbb26f4c9),
	.w3(32'hbcb90e8a),
	.w4(32'hbc1726a5),
	.w5(32'hbbdfdb47),
	.w6(32'hbbc1275d),
	.w7(32'h3b07eb57),
	.w8(32'hbc736a9e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfa4bb),
	.w1(32'hbb266894),
	.w2(32'hbb51483f),
	.w3(32'hbb33da76),
	.w4(32'hbac52029),
	.w5(32'h398e9a17),
	.w6(32'hbc05e1e2),
	.w7(32'hbbfa3078),
	.w8(32'h3b993f9c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b874f8),
	.w1(32'h3c0a567f),
	.w2(32'hbb4ba75e),
	.w3(32'hbae28ad6),
	.w4(32'hbacf4f40),
	.w5(32'h37afbf7e),
	.w6(32'hbbdce689),
	.w7(32'hbb5d50c2),
	.w8(32'hbbe1ccc0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb158b5f),
	.w1(32'h39c4d694),
	.w2(32'h3a7cffbd),
	.w3(32'h3c036ac3),
	.w4(32'h3b8abb0f),
	.w5(32'h3906471c),
	.w6(32'hbb3e58a4),
	.w7(32'h3b21ed28),
	.w8(32'h3b923e25),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba736c05),
	.w1(32'hb9693534),
	.w2(32'hbba13d49),
	.w3(32'hbb5aa1e5),
	.w4(32'h3801e909),
	.w5(32'hbc088b88),
	.w6(32'hbb836908),
	.w7(32'h39e1e158),
	.w8(32'h3a26a0d3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9e31a),
	.w1(32'h3a8d4afe),
	.w2(32'h3bd51564),
	.w3(32'hbc0efde4),
	.w4(32'h3ad22575),
	.w5(32'hbc06de51),
	.w6(32'hbbd22ddf),
	.w7(32'h3c23f56c),
	.w8(32'h3adcc31e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29cb57),
	.w1(32'hba87b194),
	.w2(32'h3ad1406a),
	.w3(32'h3910ea3a),
	.w4(32'h3c861606),
	.w5(32'h3c92bd52),
	.w6(32'hbc015bb5),
	.w7(32'hba9d39cb),
	.w8(32'h3bc008d4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52b69b),
	.w1(32'hbba42b65),
	.w2(32'hbb01d7f8),
	.w3(32'h3af05b29),
	.w4(32'hbc9b3cc6),
	.w5(32'hbc9ce484),
	.w6(32'hbc9d6b28),
	.w7(32'hbbef8628),
	.w8(32'hb90248b3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0db26a),
	.w1(32'hbc892736),
	.w2(32'hbc0ea35c),
	.w3(32'hbd3af75a),
	.w4(32'hbca5dd14),
	.w5(32'hbc262fcd),
	.w6(32'hbd271497),
	.w7(32'hbc1cd87e),
	.w8(32'hbc76cfcf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf84251),
	.w1(32'hbbe66996),
	.w2(32'hbbc9f7d9),
	.w3(32'hbafc25a8),
	.w4(32'hbbb07120),
	.w5(32'h3b6d5100),
	.w6(32'hbd1a64e7),
	.w7(32'hbb77fb79),
	.w8(32'hbc915235),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb2559),
	.w1(32'hbc8021ce),
	.w2(32'hbbcd73f1),
	.w3(32'h3c6f1ebc),
	.w4(32'h3cd1a77c),
	.w5(32'h3d10d9e4),
	.w6(32'hbc0446a8),
	.w7(32'hba8e4047),
	.w8(32'hbd12beb5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c2b1e),
	.w1(32'hbb0b1589),
	.w2(32'hbb3ee8e5),
	.w3(32'h3ab70b5c),
	.w4(32'hbc2a4395),
	.w5(32'hbc24ac52),
	.w6(32'h3cff121c),
	.w7(32'hbb02cb44),
	.w8(32'hbb32fb9a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac53559),
	.w1(32'hbb5488ac),
	.w2(32'hbbe67596),
	.w3(32'hbc0e54ce),
	.w4(32'hbb4e06a3),
	.w5(32'hbb84317f),
	.w6(32'hbc247195),
	.w7(32'hbb53e3a6),
	.w8(32'h3ad2c0a4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a22bf6),
	.w1(32'h3be447b6),
	.w2(32'hbacaf133),
	.w3(32'hbb3b369f),
	.w4(32'h3bc98cc2),
	.w5(32'h3bf27174),
	.w6(32'h3b8d9ae9),
	.w7(32'h3bb3288a),
	.w8(32'h3b91a744),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b0f9c),
	.w1(32'hbbe1197f),
	.w2(32'hbab79830),
	.w3(32'h3af5f75d),
	.w4(32'hbca63815),
	.w5(32'hbc9df62c),
	.w6(32'h3b827f50),
	.w7(32'h3bf3263e),
	.w8(32'h3bf20ba6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d8ed1),
	.w1(32'hbbc65818),
	.w2(32'hbbda5970),
	.w3(32'hbb876246),
	.w4(32'h3be561cf),
	.w5(32'h3c990397),
	.w6(32'h3bc3e5a1),
	.w7(32'hbc47caf2),
	.w8(32'hbafdb2af),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb907af9),
	.w1(32'hbbe90847),
	.w2(32'h3b11e8cf),
	.w3(32'h3c73d361),
	.w4(32'h3bb09d25),
	.w5(32'h3d01e1bc),
	.w6(32'hb9967f7e),
	.w7(32'hbc6fb446),
	.w8(32'hbd3d079d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a640e),
	.w1(32'hbc3fbb84),
	.w2(32'hbaf1a6ae),
	.w3(32'h3b63fe87),
	.w4(32'hbc2c6791),
	.w5(32'hbb62c010),
	.w6(32'hbcd1d440),
	.w7(32'hbc6b11ea),
	.w8(32'hbc909933),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc6dda),
	.w1(32'hbc3c49cf),
	.w2(32'hbc597a74),
	.w3(32'h39b78d5f),
	.w4(32'h3ba547bd),
	.w5(32'h3c27a52a),
	.w6(32'hbc14a2dc),
	.w7(32'hbc15a60a),
	.w8(32'hbcdb4da2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ff687),
	.w1(32'hbb9156f8),
	.w2(32'h3b04cdf2),
	.w3(32'h3c4ec4fb),
	.w4(32'h39fce302),
	.w5(32'hbb729646),
	.w6(32'hbc88d0ca),
	.w7(32'h3b2e9dcd),
	.w8(32'h3a87fd5e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f54d9),
	.w1(32'h3b997ac0),
	.w2(32'hbc5b4f05),
	.w3(32'hbbdee062),
	.w4(32'h3b8fbb4c),
	.w5(32'h3c94968c),
	.w6(32'hbbf047c4),
	.w7(32'hbcf953e8),
	.w8(32'hbd22c173),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf9cc5),
	.w1(32'hbc85368c),
	.w2(32'hbc9033e1),
	.w3(32'h3aa62e5d),
	.w4(32'hbc491ce9),
	.w5(32'hbbe679f2),
	.w6(32'hbd01b987),
	.w7(32'hbb53079a),
	.w8(32'h3d50ae9d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace0f7f),
	.w1(32'h3b498d02),
	.w2(32'hbc0dfc88),
	.w3(32'hbbf8bcfc),
	.w4(32'h3c0a0f62),
	.w5(32'hbc399f8a),
	.w6(32'h3c743958),
	.w7(32'h3bb55c4e),
	.w8(32'h3c8bb84b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61c4b7),
	.w1(32'hba9b5703),
	.w2(32'h3aacca2c),
	.w3(32'hbc82032e),
	.w4(32'hbbfffb6d),
	.w5(32'hbc4e00f0),
	.w6(32'h3c796dd3),
	.w7(32'hbac5d0b4),
	.w8(32'h3b43a515),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b892841),
	.w1(32'h3b6a30cd),
	.w2(32'hbb43c748),
	.w3(32'hbc4ae825),
	.w4(32'h3c61af14),
	.w5(32'hbaa6745a),
	.w6(32'hbaced764),
	.w7(32'hbcae21a3),
	.w8(32'hbc2d66d5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c264a2c),
	.w1(32'h3c560ed7),
	.w2(32'hbc2aa5ba),
	.w3(32'hbc338377),
	.w4(32'h3c2f311e),
	.w5(32'h3ccf5358),
	.w6(32'h3af56e69),
	.w7(32'hbc9b6488),
	.w8(32'h3caf6275),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b11e3),
	.w1(32'hbc963c8b),
	.w2(32'hbb9bc1a0),
	.w3(32'h3c3db03a),
	.w4(32'hbc62d62f),
	.w5(32'hbc85e610),
	.w6(32'h3c24e94a),
	.w7(32'h3b7ffdfa),
	.w8(32'h3c3c3242),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51171e),
	.w1(32'hba9e9300),
	.w2(32'hbad0f640),
	.w3(32'hbb9de70b),
	.w4(32'hbc234d15),
	.w5(32'h3baccd36),
	.w6(32'h3c5068e9),
	.w7(32'hbbf18188),
	.w8(32'hbadf58a1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b39d7),
	.w1(32'hbc454609),
	.w2(32'hbb3529bc),
	.w3(32'hbb7c536b),
	.w4(32'hbc80ada8),
	.w5(32'hbc3331c4),
	.w6(32'hbb75d8d1),
	.w7(32'h3c2ea21b),
	.w8(32'h3c510e42),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb336239),
	.w1(32'hbafd33ce),
	.w2(32'h38644610),
	.w3(32'hbcbcb62f),
	.w4(32'hbb3c84a2),
	.w5(32'hbc2eea8f),
	.w6(32'h3bc8c438),
	.w7(32'hbb855065),
	.w8(32'hbc11b277),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2f29c),
	.w1(32'h3c333c7d),
	.w2(32'h3b5c0421),
	.w3(32'hbae4348b),
	.w4(32'h3b7e93f3),
	.w5(32'h3c4ef268),
	.w6(32'hbc0a1c78),
	.w7(32'h3a95d10f),
	.w8(32'hbc48870d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b840769),
	.w1(32'hbb2312ae),
	.w2(32'hbc84d16f),
	.w3(32'hbbd7472b),
	.w4(32'hbb34834c),
	.w5(32'h3b47d9d0),
	.w6(32'hbca636ef),
	.w7(32'hbbd73edc),
	.w8(32'h3ce693d8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9357bf),
	.w1(32'h3b4c0319),
	.w2(32'hbb9b6277),
	.w3(32'hbb6acd3c),
	.w4(32'h3b2e19b9),
	.w5(32'hbb380ab0),
	.w6(32'h3bc44796),
	.w7(32'hbba1e74d),
	.w8(32'h3ad8b514),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c6e10),
	.w1(32'h3be5ed0a),
	.w2(32'hbb05cba3),
	.w3(32'h3b4674c4),
	.w4(32'h3b39ec32),
	.w5(32'h3c2550ff),
	.w6(32'h3b1a6fd7),
	.w7(32'hba3281d1),
	.w8(32'hbcfeaf97),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd2d1af),
	.w1(32'hbcb81430),
	.w2(32'h3b9f8a6c),
	.w3(32'h3ba186d6),
	.w4(32'h3b21d228),
	.w5(32'h3a814b97),
	.w6(32'hbb6e18cb),
	.w7(32'hbac7f840),
	.w8(32'hbb09eb39),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cc1f7),
	.w1(32'h3b96d7ee),
	.w2(32'hbc262e2f),
	.w3(32'hbc668ed8),
	.w4(32'hba78724a),
	.w5(32'h3c64e242),
	.w6(32'hbca4ea27),
	.w7(32'hbc10951f),
	.w8(32'hbaa3e9c7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38e098),
	.w1(32'h3bd3f86d),
	.w2(32'hba9d9403),
	.w3(32'hbca5dc95),
	.w4(32'hbb8e2a5b),
	.w5(32'hbadeef38),
	.w6(32'hbcf2a789),
	.w7(32'hba312555),
	.w8(32'hbc40af3f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ff93),
	.w1(32'h3c812ced),
	.w2(32'hbbce317e),
	.w3(32'h3ba1385a),
	.w4(32'h3cd9cca3),
	.w5(32'h3d6bfc99),
	.w6(32'h3c6ffb1e),
	.w7(32'hbc26a934),
	.w8(32'hbcbeae34),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb69745),
	.w1(32'hbc2c93c3),
	.w2(32'hbd148334),
	.w3(32'h3d1ceb1e),
	.w4(32'h3b97e167),
	.w5(32'h3cdaee29),
	.w6(32'hbc188a87),
	.w7(32'hbccb0f55),
	.w8(32'hbc3d02a1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa111b),
	.w1(32'hbcc517eb),
	.w2(32'h3c356d7b),
	.w3(32'h3ce9eb04),
	.w4(32'hbc3ac901),
	.w5(32'hbd910cc6),
	.w6(32'hbbc21c10),
	.w7(32'h3ca793b8),
	.w8(32'h3cc0db65),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80cd79),
	.w1(32'h3c51819e),
	.w2(32'h3be8cf5f),
	.w3(32'hbd32ea92),
	.w4(32'hbb3cda20),
	.w5(32'hbc1ae726),
	.w6(32'hbc973acb),
	.w7(32'h3c970c68),
	.w8(32'h3ace3023),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbffb98),
	.w1(32'hbc98f450),
	.w2(32'hbba5a1e8),
	.w3(32'h3c8cab82),
	.w4(32'h3a1c6733),
	.w5(32'hbcb63026),
	.w6(32'hbc5f2bcf),
	.w7(32'hbae942a2),
	.w8(32'hbc5f03d0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63fc6e),
	.w1(32'hbb99ecb5),
	.w2(32'hbb71b05e),
	.w3(32'hbc4c7cdf),
	.w4(32'h3b56ea9b),
	.w5(32'h3b7961c3),
	.w6(32'hbc49f63c),
	.w7(32'hbb5b8020),
	.w8(32'hbae9a235),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16cbb5),
	.w1(32'hbab81df5),
	.w2(32'hbc725873),
	.w3(32'h3be04924),
	.w4(32'hb8da57c3),
	.w5(32'h3b261fa3),
	.w6(32'hb9ea8d32),
	.w7(32'hbc3ab38f),
	.w8(32'hbaea4f3b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03532c),
	.w1(32'hbc64fcad),
	.w2(32'hbc11a090),
	.w3(32'h3c7191d2),
	.w4(32'hbb768c86),
	.w5(32'hbb8c1ac2),
	.w6(32'hb702e2c1),
	.w7(32'h3af3aea1),
	.w8(32'h3af27626),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33c996),
	.w1(32'hbb6007e0),
	.w2(32'hbb64d592),
	.w3(32'h3be49fdd),
	.w4(32'hbbea531c),
	.w5(32'hbbf5386e),
	.w6(32'hbb70a710),
	.w7(32'hba3545d7),
	.w8(32'h3b7af456),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b80b),
	.w1(32'hbabe6e35),
	.w2(32'h3c547192),
	.w3(32'hbc8176fb),
	.w4(32'hbc537496),
	.w5(32'hbd00ce44),
	.w6(32'hbb025c8d),
	.w7(32'hbc2b3de5),
	.w8(32'hbcedb8ad),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a22ca),
	.w1(32'h3bed97ea),
	.w2(32'hbba1be24),
	.w3(32'hbc52727d),
	.w4(32'hb8a1de22),
	.w5(32'hba5fe02f),
	.w6(32'hbc0aae94),
	.w7(32'hbbe4d81b),
	.w8(32'h38719bf4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af64f17),
	.w1(32'h3b9af312),
	.w2(32'hbb254e79),
	.w3(32'h3bdf5e88),
	.w4(32'hbae67df9),
	.w5(32'hbc818097),
	.w6(32'h3b7b77f8),
	.w7(32'h39116d16),
	.w8(32'h3cc64380),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae34d3),
	.w1(32'h3bbf55f4),
	.w2(32'h3befe236),
	.w3(32'hbc291c7d),
	.w4(32'h3b0f3a23),
	.w5(32'hbd076b8b),
	.w6(32'h3bc1e12e),
	.w7(32'h3b905a8c),
	.w8(32'h3b7f6c00),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c343e37),
	.w1(32'h3c3dc556),
	.w2(32'hbb8620fe),
	.w3(32'hbc431449),
	.w4(32'h3b523046),
	.w5(32'h3c12cc72),
	.w6(32'hbafd2cda),
	.w7(32'h3b169cb3),
	.w8(32'h3b6a5170),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde66ca),
	.w1(32'hbb889bf0),
	.w2(32'hbb0abafc),
	.w3(32'hb9925779),
	.w4(32'hb9023b09),
	.w5(32'h3c9d9e25),
	.w6(32'h3b61c3e7),
	.w7(32'h3c707844),
	.w8(32'hbb703250),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d8089),
	.w1(32'h3b8e6584),
	.w2(32'hbb347844),
	.w3(32'h3c2ac581),
	.w4(32'hba146503),
	.w5(32'h3ca22f7c),
	.w6(32'h3b9122a3),
	.w7(32'hbc557336),
	.w8(32'hbac0dba5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule