module layer_10_featuremap_26(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf2c7c),
	.w1(32'h3bb0a11d),
	.w2(32'h3ae8cb0a),
	.w3(32'hbc408771),
	.w4(32'h3bd8031b),
	.w5(32'h3a0a1879),
	.w6(32'hbb9ebad4),
	.w7(32'h3c6aa670),
	.w8(32'hbb05332f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70ab8b),
	.w1(32'hbc1ad6f3),
	.w2(32'hbc175621),
	.w3(32'hb8ac581e),
	.w4(32'hbb2e0dd3),
	.w5(32'hbbbd085f),
	.w6(32'h3bf2a768),
	.w7(32'h3c5a8acb),
	.w8(32'h3b75f792),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d2236),
	.w1(32'h3bccf808),
	.w2(32'h3c0ccfee),
	.w3(32'h3d1121bb),
	.w4(32'h3c78b541),
	.w5(32'h3be77f3e),
	.w6(32'h3c8aecdb),
	.w7(32'h3c2f67e5),
	.w8(32'hbaeb7864),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1abf3f),
	.w1(32'h3b838cc0),
	.w2(32'hbbe6089b),
	.w3(32'hba66487d),
	.w4(32'h3b8123b4),
	.w5(32'hbbefa20f),
	.w6(32'h3c0752fd),
	.w7(32'h3c2292ae),
	.w8(32'h3bfb3415),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb482db),
	.w1(32'h3c8b8844),
	.w2(32'h3b55a147),
	.w3(32'h3c5cd7ce),
	.w4(32'h3cdf09ae),
	.w5(32'h3c2ea407),
	.w6(32'h3cc91ed9),
	.w7(32'h3c12fc4f),
	.w8(32'h3c10ba24),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb171857),
	.w1(32'h3ba16637),
	.w2(32'hbb311f93),
	.w3(32'hbb541f04),
	.w4(32'h3bb4f521),
	.w5(32'hbbaf5efa),
	.w6(32'h3b35242a),
	.w7(32'h3b8dc43d),
	.w8(32'hbb844a21),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9945f8),
	.w1(32'hbb0126ec),
	.w2(32'h3bef2a1c),
	.w3(32'hbba86322),
	.w4(32'hbafb2fa3),
	.w5(32'h3b8f05f1),
	.w6(32'hbb4d9099),
	.w7(32'hbb8a807f),
	.w8(32'h3c1d3061),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d614c),
	.w1(32'h3b8705d1),
	.w2(32'h3be2de9f),
	.w3(32'hbb673a19),
	.w4(32'h3c36f245),
	.w5(32'h3b8854e1),
	.w6(32'hba68d083),
	.w7(32'hbb6e6e56),
	.w8(32'hba6f0005),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d6d29),
	.w1(32'hbb3afe68),
	.w2(32'hbad6e4af),
	.w3(32'hbba9135f),
	.w4(32'h3ae9b417),
	.w5(32'h3bbeb47b),
	.w6(32'h3bf03f1d),
	.w7(32'h3bd0b224),
	.w8(32'h3bf1608c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba01b99),
	.w1(32'h3c3650ac),
	.w2(32'hbaa660d1),
	.w3(32'h3c19699c),
	.w4(32'h3c2ba016),
	.w5(32'h3ac420f8),
	.w6(32'h3c289a5d),
	.w7(32'h3bb756d5),
	.w8(32'h3acc9363),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bb9c0),
	.w1(32'h3b43e32f),
	.w2(32'hba3320f5),
	.w3(32'h3baa8d92),
	.w4(32'h3b599b82),
	.w5(32'h3b6b94a4),
	.w6(32'h3ba2e6aa),
	.w7(32'h3b8ec749),
	.w8(32'h3a8d0fb8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf971a),
	.w1(32'hb90f23ac),
	.w2(32'h3b195ab5),
	.w3(32'h3b17fd8e),
	.w4(32'h3bd80b8f),
	.w5(32'h3909bcb4),
	.w6(32'h3a43ad9d),
	.w7(32'hbaf85355),
	.w8(32'h3ae1eca8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90d1a7),
	.w1(32'h3b3d4eea),
	.w2(32'h3c253821),
	.w3(32'hba567f30),
	.w4(32'h3ba88a1a),
	.w5(32'h3bb42920),
	.w6(32'h3b25c6eb),
	.w7(32'h3bd70cda),
	.w8(32'h3b779a52),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c472ae7),
	.w1(32'h3c0463f5),
	.w2(32'hbc1e8e84),
	.w3(32'h3b868cc3),
	.w4(32'h3c0c8de6),
	.w5(32'hbbd58e73),
	.w6(32'h3c09005f),
	.w7(32'h3ba8aac1),
	.w8(32'hbb72fa84),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc912cf7),
	.w1(32'hbc786644),
	.w2(32'h3ab53930),
	.w3(32'hbc7cdac5),
	.w4(32'hbbf15dcc),
	.w5(32'h3badb9fd),
	.w6(32'hbbe8393f),
	.w7(32'h3b7fec93),
	.w8(32'h3ad5329e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd72870),
	.w1(32'hbb951aee),
	.w2(32'h3aabbe54),
	.w3(32'hb9fc955a),
	.w4(32'hbc053d5f),
	.w5(32'h3ba919d6),
	.w6(32'h3b8b7893),
	.w7(32'hbc0dc577),
	.w8(32'h3badceff),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a0c42),
	.w1(32'h399cfc77),
	.w2(32'h3b0f67ff),
	.w3(32'h3ba689ba),
	.w4(32'h3adc3ffe),
	.w5(32'h3baa153c),
	.w6(32'h3b91c78d),
	.w7(32'h3b04159e),
	.w8(32'h3b7a0825),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbaa5f),
	.w1(32'h3b7caed1),
	.w2(32'h3baecff0),
	.w3(32'h3b5bd88c),
	.w4(32'h3b609de5),
	.w5(32'h3c5022c5),
	.w6(32'h3b1c5171),
	.w7(32'h3ab4faa4),
	.w8(32'h3bfba5d2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6edb9),
	.w1(32'h3af88039),
	.w2(32'hbb022beb),
	.w3(32'h3c3c2be5),
	.w4(32'h3bb68f57),
	.w5(32'hbc02a4ed),
	.w6(32'h3bfb1c63),
	.w7(32'h3be5a93d),
	.w8(32'hbc123dd4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94c1d2),
	.w1(32'h3c29ca85),
	.w2(32'h3bdf7bd7),
	.w3(32'hbc24de31),
	.w4(32'h3b9b5bc0),
	.w5(32'h3be6ea55),
	.w6(32'hbc38bf7c),
	.w7(32'hbbc7e9a7),
	.w8(32'h3bbca446),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfd354),
	.w1(32'h3bc77dc6),
	.w2(32'h3c08bc67),
	.w3(32'h3be4d86d),
	.w4(32'hba806c3f),
	.w5(32'h3ac99fc5),
	.w6(32'h3b97ef59),
	.w7(32'h3a875ab3),
	.w8(32'h3a2c5b3c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bceff),
	.w1(32'h3971ef9a),
	.w2(32'hba46445e),
	.w3(32'hbbda9400),
	.w4(32'h3b29aa73),
	.w5(32'hbc01d264),
	.w6(32'hbac9a32e),
	.w7(32'h3983dab6),
	.w8(32'hba4b2b58),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0cf74),
	.w1(32'h3bba7b11),
	.w2(32'hbbe97175),
	.w3(32'hbc450b30),
	.w4(32'hbb5d65db),
	.w5(32'hbbab41ba),
	.w6(32'hbc0fd1c5),
	.w7(32'hbb064a9e),
	.w8(32'hbb986b57),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0d0d6),
	.w1(32'hba943f4a),
	.w2(32'h3c0487fc),
	.w3(32'hbbbc082b),
	.w4(32'hbb18e0fe),
	.w5(32'h3c286c12),
	.w6(32'hbbb44255),
	.w7(32'h3a18352e),
	.w8(32'h3c0b48f0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b815e94),
	.w1(32'h3b982e5c),
	.w2(32'h3a8f04cf),
	.w3(32'h3b5f80b0),
	.w4(32'h3b08d7da),
	.w5(32'hb8776ed1),
	.w6(32'h3951c56e),
	.w7(32'h3be2b269),
	.w8(32'h3a93950c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b348307),
	.w1(32'h3a32cbc4),
	.w2(32'h3bc85718),
	.w3(32'h3b82e6e3),
	.w4(32'h3c1ae0b8),
	.w5(32'h3c0b51ce),
	.w6(32'hb995efab),
	.w7(32'h3c7097a0),
	.w8(32'hbab9af94),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac6961),
	.w1(32'h3b87dc25),
	.w2(32'hbb88d438),
	.w3(32'h3b2f6775),
	.w4(32'h3bc66136),
	.w5(32'h3b0b44ee),
	.w6(32'hbaa49e1f),
	.w7(32'h3bad8480),
	.w8(32'hbb6728dd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99a161),
	.w1(32'hbb41a2e8),
	.w2(32'h3ac9319e),
	.w3(32'h3cab0034),
	.w4(32'h3ba08f00),
	.w5(32'h3b896a23),
	.w6(32'h3bff8b90),
	.w7(32'hbb3629c2),
	.w8(32'h3b68d2c6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7adc4b),
	.w1(32'hba25afc6),
	.w2(32'h3b24d9b8),
	.w3(32'h3b6bbb98),
	.w4(32'h3b839f34),
	.w5(32'hbb8f0af9),
	.w6(32'h3bdccb2d),
	.w7(32'h3c01393f),
	.w8(32'h3b99df28),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bfdb52),
	.w1(32'hbb52a6de),
	.w2(32'h3c957574),
	.w3(32'hbb3952db),
	.w4(32'hb9fee1da),
	.w5(32'h3b594339),
	.w6(32'hbbcf5636),
	.w7(32'h3a37a1ea),
	.w8(32'h3c5a77df),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07a78d),
	.w1(32'h3c73230f),
	.w2(32'hbaa377c9),
	.w3(32'hbc12b27e),
	.w4(32'h395b37d4),
	.w5(32'h3a1040f9),
	.w6(32'h3ae95398),
	.w7(32'h3c21965d),
	.w8(32'hbb53986b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7837fb),
	.w1(32'hba63ef5d),
	.w2(32'h3abeb2a4),
	.w3(32'h3b2820d0),
	.w4(32'hbb06c885),
	.w5(32'h3a311989),
	.w6(32'h3a9da0c8),
	.w7(32'hbac14ca6),
	.w8(32'h3b1a5cb7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980c582),
	.w1(32'h3b32e088),
	.w2(32'hbb50d57a),
	.w3(32'hba9f2abe),
	.w4(32'hbaf7e8ad),
	.w5(32'hbcf14f87),
	.w6(32'hbaa807e0),
	.w7(32'h3b2eea4c),
	.w8(32'hbc85eb5d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccab0fe),
	.w1(32'hbc3403a0),
	.w2(32'h3b431599),
	.w3(32'hbd7c1c31),
	.w4(32'hbd224896),
	.w5(32'h3b3da7b4),
	.w6(32'hbd3baaf6),
	.w7(32'hbcccfd80),
	.w8(32'hbb084bf8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399299a0),
	.w1(32'hba080db0),
	.w2(32'hbc23f5e9),
	.w3(32'h3a0325f1),
	.w4(32'h3b1aafeb),
	.w5(32'hbb097ebe),
	.w6(32'h39d4e9bc),
	.w7(32'h3b6d2634),
	.w8(32'hbc0764b6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb53987),
	.w1(32'hbc43fc3a),
	.w2(32'h3aba0bb9),
	.w3(32'h3b4e86f8),
	.w4(32'hbb467365),
	.w5(32'h3bb679ad),
	.w6(32'hbb28eba6),
	.w7(32'hbc09c228),
	.w8(32'h39fe9851),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a6c71),
	.w1(32'hba607f6b),
	.w2(32'hbb2851fe),
	.w3(32'h3a048ea2),
	.w4(32'h3b1f2956),
	.w5(32'hbcab7ebd),
	.w6(32'hbaf3185a),
	.w7(32'hbb9c1ec6),
	.w8(32'hbc36867c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5e754),
	.w1(32'hbc495fb5),
	.w2(32'hbb41baea),
	.w3(32'hbd3f95a0),
	.w4(32'hbcf7e447),
	.w5(32'hbaec0a86),
	.w6(32'hbcff0bb2),
	.w7(32'hbc859048),
	.w8(32'hbb93f454),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99abde),
	.w1(32'h3997c6c6),
	.w2(32'hba2f8dfc),
	.w3(32'hbbe8461b),
	.w4(32'hbb8e8984),
	.w5(32'hbba59359),
	.w6(32'h3a08d42b),
	.w7(32'hbb969c49),
	.w8(32'hbb799599),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae97b23),
	.w1(32'h39d2ab39),
	.w2(32'hba552d09),
	.w3(32'h3a41a0fb),
	.w4(32'h3b9c4124),
	.w5(32'hbaa71654),
	.w6(32'h3a7fb803),
	.w7(32'h3b8f0905),
	.w8(32'hbb159fbf),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58cb5a),
	.w1(32'hbbafb3b9),
	.w2(32'hbb7bf3fc),
	.w3(32'hbba3303c),
	.w4(32'hbba0d164),
	.w5(32'h3bbc7ce9),
	.w6(32'hbb3ca2e5),
	.w7(32'hbacc4a03),
	.w8(32'hb991191d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39a826),
	.w1(32'h3b6752b5),
	.w2(32'hba287538),
	.w3(32'h3a203014),
	.w4(32'h3b0f4713),
	.w5(32'hbb3985e4),
	.w6(32'hbadfda5d),
	.w7(32'h3b5ecc96),
	.w8(32'hba93260c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d0d7c),
	.w1(32'hbb99498c),
	.w2(32'h3c249707),
	.w3(32'h3884ad06),
	.w4(32'h3ab3e85e),
	.w5(32'h3d0d7345),
	.w6(32'hb9e651b4),
	.w7(32'hbb9e4634),
	.w8(32'h3caeaa0e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccaef47),
	.w1(32'h3c4deaa9),
	.w2(32'h3b7b27ea),
	.w3(32'h3d788686),
	.w4(32'h3d334a6b),
	.w5(32'h3b0853bc),
	.w6(32'h3d406905),
	.w7(32'h3cf87499),
	.w8(32'hbb401e0e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeafc1e),
	.w1(32'hb6ddca82),
	.w2(32'hba6ffa35),
	.w3(32'hbb75a50e),
	.w4(32'hbb29570d),
	.w5(32'h3b334235),
	.w6(32'hba0d2bba),
	.w7(32'hbaefc099),
	.w8(32'h38ee31d7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932a47),
	.w1(32'hbb9e94b8),
	.w2(32'hbb6eb19f),
	.w3(32'h3c081eb7),
	.w4(32'h3b61ea42),
	.w5(32'hba1b65bd),
	.w6(32'h3adf584c),
	.w7(32'h3b91a4a7),
	.w8(32'h3b7d10bf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c2336),
	.w1(32'hbb84c912),
	.w2(32'hbb0be44a),
	.w3(32'hb97bcaab),
	.w4(32'hba71df29),
	.w5(32'hb9d36e75),
	.w6(32'h3aa52b0f),
	.w7(32'hba3c6112),
	.w8(32'hba2a31e4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe382ee),
	.w1(32'h3ad9f3e7),
	.w2(32'hbcd3ff42),
	.w3(32'hbbe2af31),
	.w4(32'h3ac5e74c),
	.w5(32'hbbe8bb7a),
	.w6(32'h3a340cf4),
	.w7(32'hba51c7ec),
	.w8(32'hbc9fc94c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71f909),
	.w1(32'hbcc1b1e7),
	.w2(32'h3bbdda57),
	.w3(32'h3c221ea6),
	.w4(32'hbb8b00d3),
	.w5(32'hb9f7f079),
	.w6(32'hbb270eeb),
	.w7(32'hbc756d88),
	.w8(32'hb99ef4cf),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e3247),
	.w1(32'h3aa28509),
	.w2(32'hbb7171b2),
	.w3(32'h3a935df4),
	.w4(32'hb9a39bac),
	.w5(32'h386d9cfd),
	.w6(32'hba3fbcec),
	.w7(32'h3b00cd8f),
	.w8(32'hbba7a3ac),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0eab),
	.w1(32'hbbb28941),
	.w2(32'h3bbb72eb),
	.w3(32'hba1b6d98),
	.w4(32'hbc089841),
	.w5(32'hbacce38f),
	.w6(32'hbb9f6c9c),
	.w7(32'hbb5f8cf4),
	.w8(32'h3ad886aa),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06e366),
	.w1(32'h3ac3bd57),
	.w2(32'h3b1ce092),
	.w3(32'h3afcd780),
	.w4(32'hbb327177),
	.w5(32'h3b90ac03),
	.w6(32'hbb4f0004),
	.w7(32'hbb8affe4),
	.w8(32'h3a786741),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cef69f),
	.w1(32'h3a2b4f47),
	.w2(32'h3b1f9ce3),
	.w3(32'h3b92c4a5),
	.w4(32'h3b935619),
	.w5(32'h3b930e93),
	.w6(32'hbb1080c7),
	.w7(32'hbad94bca),
	.w8(32'h3b97dd77),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27649c),
	.w1(32'hb9bee068),
	.w2(32'hbb9b38d4),
	.w3(32'h3b0f0567),
	.w4(32'h3b5f3069),
	.w5(32'hbb3ca193),
	.w6(32'h3bb4ba41),
	.w7(32'h3ae90d7f),
	.w8(32'h3b1aaae6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b6647),
	.w1(32'hbb959e60),
	.w2(32'hbb41761f),
	.w3(32'hba7c2414),
	.w4(32'hbaf7c70e),
	.w5(32'hbb8d4ef1),
	.w6(32'h3a29ceb7),
	.w7(32'h3a9d0be1),
	.w8(32'hbb9f8d21),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb013fa0),
	.w1(32'hbbaca41f),
	.w2(32'hba4151aa),
	.w3(32'hbb14316c),
	.w4(32'hbb0cca61),
	.w5(32'hba3492bd),
	.w6(32'hbae4df8f),
	.w7(32'h38f550ca),
	.w8(32'hb7501afa),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb481f8e),
	.w1(32'h3a205a77),
	.w2(32'hbad69dbb),
	.w3(32'hba65f46f),
	.w4(32'hbb3a1c9f),
	.w5(32'hbac50353),
	.w6(32'h3b00acd4),
	.w7(32'hba24ece8),
	.w8(32'hbb3d3ae9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbcef7),
	.w1(32'hbbb262ad),
	.w2(32'hbb4c8237),
	.w3(32'hbb86f197),
	.w4(32'hbb235c40),
	.w5(32'hbba4bf35),
	.w6(32'hbac23fbb),
	.w7(32'h3b345563),
	.w8(32'hbbaaa887),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd00d42),
	.w1(32'hbaf24c8a),
	.w2(32'h3a9d820e),
	.w3(32'hbb16b409),
	.w4(32'h3ab0d2ba),
	.w5(32'h3b3ab410),
	.w6(32'h39797c6d),
	.w7(32'h3bfe42b8),
	.w8(32'h3b36c928),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4feee),
	.w1(32'hbb9238e9),
	.w2(32'h3b5c47c9),
	.w3(32'hba5d2f51),
	.w4(32'hbb0bc167),
	.w5(32'h3b65d292),
	.w6(32'h39a1bfca),
	.w7(32'h39cb5183),
	.w8(32'h3ba84978),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98002cf),
	.w1(32'hbb43047a),
	.w2(32'h3b9b0e81),
	.w3(32'h3ba13a07),
	.w4(32'h3ab9347b),
	.w5(32'h3b2ab982),
	.w6(32'h3a1fafdf),
	.w7(32'h39fc5e0d),
	.w8(32'h3ba81ec9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885d1a5),
	.w1(32'h3b13be02),
	.w2(32'h3b69cbc1),
	.w3(32'h3bb419a6),
	.w4(32'h3bc5575a),
	.w5(32'h3bb93d8f),
	.w6(32'h3b0c6355),
	.w7(32'h3a9ccb40),
	.w8(32'h3c25ce33),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3383e),
	.w1(32'h3bd7b0fd),
	.w2(32'h3a31b02a),
	.w3(32'h3a5e9a4e),
	.w4(32'h3b8b0d0b),
	.w5(32'h3b993307),
	.w6(32'h3b734e85),
	.w7(32'h3acfe8d1),
	.w8(32'h3af7a570),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5de930),
	.w1(32'h3ac117a4),
	.w2(32'hb98985d6),
	.w3(32'h3be947a5),
	.w4(32'h3b3565f4),
	.w5(32'h3b95b38d),
	.w6(32'h3b1c6971),
	.w7(32'h3b6ca76e),
	.w8(32'h3a87caba),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cdbaae),
	.w1(32'hbb528a17),
	.w2(32'h3b9a38b2),
	.w3(32'hbb937634),
	.w4(32'hbb690825),
	.w5(32'h3bcf4146),
	.w6(32'h39c662d8),
	.w7(32'hbb50aea5),
	.w8(32'h3b2728f1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52d5f4),
	.w1(32'h3b2d412c),
	.w2(32'h3c426816),
	.w3(32'h3b5f4ca6),
	.w4(32'h3b99895b),
	.w5(32'h3c5ce970),
	.w6(32'h3b049cdc),
	.w7(32'h3b9756aa),
	.w8(32'h3c6561e9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12cac5),
	.w1(32'h3c22ea4e),
	.w2(32'h3bd378c5),
	.w3(32'h3c8e936a),
	.w4(32'h3c86a3c4),
	.w5(32'h3b481d55),
	.w6(32'h3c9126c3),
	.w7(32'h3c8858c2),
	.w8(32'hbb829e6a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c801),
	.w1(32'h3abe6a39),
	.w2(32'h3bb2bbfb),
	.w3(32'h3b249adb),
	.w4(32'h3b4f0228),
	.w5(32'h3bb99c44),
	.w6(32'hbb6e27d1),
	.w7(32'hba7e2fcb),
	.w8(32'h3b4d50b4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a5221),
	.w1(32'h3b27e0ac),
	.w2(32'hba893f5d),
	.w3(32'h3b853410),
	.w4(32'h3af7844a),
	.w5(32'hba581006),
	.w6(32'h3b89bb77),
	.w7(32'h3bca4112),
	.w8(32'h39cc9db0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0786d2),
	.w1(32'h3a09cefe),
	.w2(32'h3a8d179a),
	.w3(32'h3bb761e8),
	.w4(32'h3b127b73),
	.w5(32'h3a482a67),
	.w6(32'h3bf2db43),
	.w7(32'h3b4a3023),
	.w8(32'h3ba47368),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfc443),
	.w1(32'h3b285d0e),
	.w2(32'hba8806dd),
	.w3(32'h3bf39548),
	.w4(32'h3b86b271),
	.w5(32'hbac32807),
	.w6(32'h3c17803c),
	.w7(32'h3b1ab828),
	.w8(32'hba5f52cf),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9478b6f),
	.w1(32'hba5fe834),
	.w2(32'hbba3e53a),
	.w3(32'hbba368a4),
	.w4(32'hbb3076f6),
	.w5(32'hbac12f7a),
	.w6(32'h3a3c552b),
	.w7(32'h3a90967e),
	.w8(32'hbac5270a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbfd46),
	.w1(32'h3b9a7ef1),
	.w2(32'hbb80af68),
	.w3(32'hbb69bade),
	.w4(32'h3a345b4c),
	.w5(32'hbb9bb337),
	.w6(32'hba5904bc),
	.w7(32'h3bcbdf8a),
	.w8(32'hbbe9ab06),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8c85e),
	.w1(32'h3b179a4c),
	.w2(32'hbc40f352),
	.w3(32'h3b63dc63),
	.w4(32'hbabefb42),
	.w5(32'h3c38df04),
	.w6(32'h3ba838ff),
	.w7(32'h3b5ad5af),
	.w8(32'hbb498595),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c805510),
	.w1(32'hbbee9e6f),
	.w2(32'h3b7a3d24),
	.w3(32'h3d44ce68),
	.w4(32'h3ca52af0),
	.w5(32'hbb55db03),
	.w6(32'h3d073200),
	.w7(32'h3bae819d),
	.w8(32'hb861eb66),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfcb5a),
	.w1(32'h3b3fda20),
	.w2(32'h3b467312),
	.w3(32'hbc00f5d7),
	.w4(32'hbb833c22),
	.w5(32'hbb34ae0f),
	.w6(32'hbbaf4475),
	.w7(32'hbb18567a),
	.w8(32'hbb2988d5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7aa202),
	.w1(32'h3bc4b9d6),
	.w2(32'hbaf79f8b),
	.w3(32'h3a026125),
	.w4(32'hbbc461dd),
	.w5(32'h3a81938a),
	.w6(32'hba18993d),
	.w7(32'h3b97d7ee),
	.w8(32'hbb4775c5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7885e8),
	.w1(32'hb9b0dbee),
	.w2(32'h3aac28b9),
	.w3(32'h3b2cce9c),
	.w4(32'hbb93ecd6),
	.w5(32'h3b0ed90b),
	.w6(32'h3b60c8da),
	.w7(32'h39d7b9b4),
	.w8(32'h3bf18c99),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c4ff1),
	.w1(32'hbb847dd1),
	.w2(32'hbb2b116b),
	.w3(32'hbb8d04cc),
	.w4(32'hbbc9979b),
	.w5(32'hbb925deb),
	.w6(32'h3b747ad1),
	.w7(32'hbbc67f2a),
	.w8(32'hba8eb537),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb97f4),
	.w1(32'hba8fd573),
	.w2(32'hbb45d312),
	.w3(32'h3c52f721),
	.w4(32'h3b48b478),
	.w5(32'hbb7aa0a4),
	.w6(32'h3bb7de64),
	.w7(32'hb88fafc9),
	.w8(32'hbbc0d3bb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb279c27),
	.w1(32'hbb00a5e3),
	.w2(32'hb9888e23),
	.w3(32'hbb9990be),
	.w4(32'hbaecf5f6),
	.w5(32'hba99b616),
	.w6(32'hba82b968),
	.w7(32'hbb1efcbd),
	.w8(32'h3b04eb8d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98d593),
	.w1(32'h3b22a24d),
	.w2(32'h3aa33042),
	.w3(32'h3c3ac3c4),
	.w4(32'h3c213e98),
	.w5(32'h3bd870d4),
	.w6(32'h3c714fe5),
	.w7(32'h3c0a9323),
	.w8(32'h38dcf8bc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62a067),
	.w1(32'h3b5990b8),
	.w2(32'hbac127fd),
	.w3(32'h3b93ec32),
	.w4(32'h3b17c3cb),
	.w5(32'hbb3ae139),
	.w6(32'h3b27129e),
	.w7(32'h3ab14276),
	.w8(32'hba5b648c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacde520),
	.w1(32'hb97a4996),
	.w2(32'hba4d44e8),
	.w3(32'hbb2f4bc4),
	.w4(32'h3939bca0),
	.w5(32'hbb51df96),
	.w6(32'h39ad017f),
	.w7(32'h3adaa749),
	.w8(32'h3bc7bb33),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b280b),
	.w1(32'h3aab08d0),
	.w2(32'h3b995390),
	.w3(32'hbb14aba6),
	.w4(32'h3a807b16),
	.w5(32'h3b7eef95),
	.w6(32'hbb3c4464),
	.w7(32'h3984f393),
	.w8(32'hbba2f8a9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa928fc),
	.w1(32'hbb284d81),
	.w2(32'h3b37a834),
	.w3(32'hbb1f6bb1),
	.w4(32'hbb54f01e),
	.w5(32'h3b83cf14),
	.w6(32'hb8474e76),
	.w7(32'h3b165d5e),
	.w8(32'h3b532553),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb1ebe),
	.w1(32'h38abb304),
	.w2(32'h3c41e52f),
	.w3(32'h3b3212fa),
	.w4(32'h3aa8f7c0),
	.w5(32'h3c8f12b0),
	.w6(32'h3be6683f),
	.w7(32'h3b6da6c2),
	.w8(32'h3c91aea0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a8fdd),
	.w1(32'h3c56d696),
	.w2(32'h3aa551e5),
	.w3(32'h3cb81141),
	.w4(32'h3ca9f2c4),
	.w5(32'hbaae303e),
	.w6(32'h3cbdf9af),
	.w7(32'h3cad2f0d),
	.w8(32'hbb090345),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad40ef),
	.w1(32'hbb0abe03),
	.w2(32'h3be28c7e),
	.w3(32'hbb3ef9ef),
	.w4(32'hbb9af2a5),
	.w5(32'h3af4ca02),
	.w6(32'hbbaa1d7c),
	.w7(32'h3b0c023e),
	.w8(32'hbb0d0cf9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3da185),
	.w1(32'h3979e6ca),
	.w2(32'h3b2327c0),
	.w3(32'hb81ceed8),
	.w4(32'h3b5d99f0),
	.w5(32'h3aedc5ed),
	.w6(32'h3b03c128),
	.w7(32'h3b56a1c9),
	.w8(32'hbb7ad5f4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8a3c4),
	.w1(32'h3996e4b7),
	.w2(32'h3b845544),
	.w3(32'h3b53e7d1),
	.w4(32'h3b2123ae),
	.w5(32'h3c243b10),
	.w6(32'hbaad4a5f),
	.w7(32'hbb6cd8d8),
	.w8(32'h3c070c5a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc44b4),
	.w1(32'hbab72867),
	.w2(32'hbb43d08e),
	.w3(32'h3bd926bf),
	.w4(32'h3bf0b4a1),
	.w5(32'hbba2eb5d),
	.w6(32'h3b5c2b0d),
	.w7(32'h3ba02488),
	.w8(32'hbb55a8df),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb146c2),
	.w1(32'hbbced2a1),
	.w2(32'h3c24db7f),
	.w3(32'hbbe4bbaa),
	.w4(32'hbbd3c442),
	.w5(32'h3caf34e3),
	.w6(32'hbba390bc),
	.w7(32'hbbab1ba5),
	.w8(32'h3c97daca),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85b7d7),
	.w1(32'h3c252ebd),
	.w2(32'h3bd88be0),
	.w3(32'h3d19f20b),
	.w4(32'h3ce5f549),
	.w5(32'h3b22999b),
	.w6(32'h3d015bc6),
	.w7(32'h3cbf2295),
	.w8(32'hb91af7f2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f2a7f),
	.w1(32'h39397916),
	.w2(32'h3adacb86),
	.w3(32'h3b0e335e),
	.w4(32'h3ab4a8a8),
	.w5(32'hbb943bcd),
	.w6(32'h3a86595e),
	.w7(32'hb958cc78),
	.w8(32'hbb3bfa9a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5e336),
	.w1(32'hbbe6d803),
	.w2(32'h3a9253ce),
	.w3(32'hbc2026ec),
	.w4(32'hbc4ed761),
	.w5(32'hbbcdd1c5),
	.w6(32'h3b3a12ff),
	.w7(32'hbb0538be),
	.w8(32'hbb80d523),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb152209),
	.w1(32'h3ab830f7),
	.w2(32'hbba2d754),
	.w3(32'hbbb4e13d),
	.w4(32'hbb8cb6f2),
	.w5(32'hbb5e186a),
	.w6(32'hbbb0949a),
	.w7(32'hba5b733a),
	.w8(32'h3b308254),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc45c0),
	.w1(32'hbb53370c),
	.w2(32'h3b33d464),
	.w3(32'hbbacec3c),
	.w4(32'hbb66c2b8),
	.w5(32'h3ad6bb00),
	.w6(32'hbb9e4fdb),
	.w7(32'hbb357152),
	.w8(32'hbb93352d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa962a5),
	.w1(32'hbb2874d8),
	.w2(32'hbbeebfb7),
	.w3(32'h3afe9b21),
	.w4(32'h38cd0e83),
	.w5(32'hbb936e7e),
	.w6(32'hba3c8262),
	.w7(32'hbb3c0b49),
	.w8(32'hbba33a9c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dd767),
	.w1(32'hbb458244),
	.w2(32'hbb374da1),
	.w3(32'hb90b9c05),
	.w4(32'h3b22b3d3),
	.w5(32'h3a1424d6),
	.w6(32'h3b1700f8),
	.w7(32'h39ec77d1),
	.w8(32'h3b0fe74c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aaacd),
	.w1(32'h38e23642),
	.w2(32'h3c0922fe),
	.w3(32'h3aab8fe3),
	.w4(32'h3ab9546b),
	.w5(32'h3aba50a9),
	.w6(32'h3b49fc61),
	.w7(32'hba908e17),
	.w8(32'hba6ad0c8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b265105),
	.w1(32'h3aabf4e2),
	.w2(32'hba39e127),
	.w3(32'h3ad2cd2d),
	.w4(32'hb9920654),
	.w5(32'hbb33481a),
	.w6(32'hbafe7eb7),
	.w7(32'h3ad12c4a),
	.w8(32'hbb9d9ee6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c8957),
	.w1(32'hb94a6f3e),
	.w2(32'hbb0c9475),
	.w3(32'h3b1c11d2),
	.w4(32'h3a3245c0),
	.w5(32'h3a5933af),
	.w6(32'h3b2f937f),
	.w7(32'hbb57890a),
	.w8(32'h3a2ceb68),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a3b90),
	.w1(32'h3af1274b),
	.w2(32'hba19b069),
	.w3(32'h3b808d87),
	.w4(32'h3ba4004b),
	.w5(32'h3b044bb0),
	.w6(32'h3b4c1155),
	.w7(32'hbb09aaa8),
	.w8(32'hbaabecaf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7faf66),
	.w1(32'hbb3e67d5),
	.w2(32'hb9672561),
	.w3(32'hbb3a4640),
	.w4(32'h3a55c864),
	.w5(32'hbb60a47e),
	.w6(32'hbb264d71),
	.w7(32'hbb0a45b9),
	.w8(32'h3a4a1412),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42f8ed),
	.w1(32'h3a15e9ac),
	.w2(32'h3b3bc7c1),
	.w3(32'hbb7f1cf1),
	.w4(32'hbb306a7b),
	.w5(32'h3aea1303),
	.w6(32'hbb0c4d6d),
	.w7(32'hb8f28c92),
	.w8(32'h3ba9b278),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a068a5),
	.w1(32'h3afe3a3a),
	.w2(32'h39ab3119),
	.w3(32'h3952e9ff),
	.w4(32'h3a9eb57d),
	.w5(32'h3b46fc3a),
	.w6(32'h3b0019c3),
	.w7(32'h3b9b1cd0),
	.w8(32'h3b9bbc55),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85dd01),
	.w1(32'h3afe4cf9),
	.w2(32'h3aa0cc85),
	.w3(32'h3b0940b0),
	.w4(32'h3b0b021b),
	.w5(32'hba2326b1),
	.w6(32'h3c024bbb),
	.w7(32'h3bfd2691),
	.w8(32'h3ba4f324),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02c61d),
	.w1(32'h3b2fb54e),
	.w2(32'h3b5f7a6a),
	.w3(32'h38cfa726),
	.w4(32'h3ba7cb14),
	.w5(32'h3ada9a3b),
	.w6(32'hba4bd96c),
	.w7(32'h3b6089c7),
	.w8(32'hba047540),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8461f),
	.w1(32'h3b77345a),
	.w2(32'h3a73a0f6),
	.w3(32'h3bdd9135),
	.w4(32'h3c0e4fca),
	.w5(32'h3948f2f1),
	.w6(32'h3b2fd0dd),
	.w7(32'h3b12bc7c),
	.w8(32'hbb0b1b13),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4336ac),
	.w1(32'hba7f645d),
	.w2(32'h3b5f070a),
	.w3(32'hbb2eed02),
	.w4(32'h3a5878e8),
	.w5(32'h3b8e3d17),
	.w6(32'h3b813bae),
	.w7(32'hbc137407),
	.w8(32'h3affcaa1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97087ae),
	.w1(32'h3b63a3b3),
	.w2(32'hbb1b7773),
	.w3(32'h3b9cf741),
	.w4(32'h3b70686b),
	.w5(32'hba8c3c0e),
	.w6(32'h3b4c88c4),
	.w7(32'h3a083241),
	.w8(32'hbbdbb711),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ab180),
	.w1(32'hbb21e7b4),
	.w2(32'hbb5ff906),
	.w3(32'hbad94498),
	.w4(32'h3b3d6092),
	.w5(32'hb9a42ea3),
	.w6(32'hbb1d521e),
	.w7(32'h3b4d93d0),
	.w8(32'hb97341a8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84b228),
	.w1(32'hbb6b7e6f),
	.w2(32'hbbad3cc4),
	.w3(32'hbb821a06),
	.w4(32'h39cf0127),
	.w5(32'hba1ccaa5),
	.w6(32'hbac735cd),
	.w7(32'hb977a87d),
	.w8(32'hba1dd82c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96efb55),
	.w1(32'hbaa832db),
	.w2(32'h3b27febf),
	.w3(32'h3b343932),
	.w4(32'hbaef2f12),
	.w5(32'h3a403c07),
	.w6(32'hbb00a0f0),
	.w7(32'hbb6b9299),
	.w8(32'h3b28e1fb),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bb8b9),
	.w1(32'hb7566b88),
	.w2(32'h3bdeffe3),
	.w3(32'h3a82e601),
	.w4(32'hba256c83),
	.w5(32'h3bdd5ded),
	.w6(32'h3bb05b74),
	.w7(32'h3b5dec49),
	.w8(32'h3bfa74aa),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe8794),
	.w1(32'h3b111b55),
	.w2(32'h3bc04dbf),
	.w3(32'h3bbc27f1),
	.w4(32'h3bb4d1b0),
	.w5(32'h3bb5a7d9),
	.w6(32'h3a87f0a4),
	.w7(32'h3a3e4b3e),
	.w8(32'h3b141172),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf57da),
	.w1(32'h3afcd6e9),
	.w2(32'hb9cc870b),
	.w3(32'h3b7682e0),
	.w4(32'h3b9d325e),
	.w5(32'hbb5a39aa),
	.w6(32'h3b2a8dd7),
	.w7(32'h3bc85254),
	.w8(32'hb9ec5683),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8867d5),
	.w1(32'h3a0af78e),
	.w2(32'h3a7e6cc0),
	.w3(32'h3a06c5d3),
	.w4(32'h3a737bdd),
	.w5(32'h3a8abcdf),
	.w6(32'hb9fd0843),
	.w7(32'h3ae9a3a9),
	.w8(32'hbb8aa1bd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9abf1a),
	.w1(32'h3ba6a81e),
	.w2(32'h3b40b22b),
	.w3(32'hb9f84b51),
	.w4(32'h3ab68ea6),
	.w5(32'h3b78d8a9),
	.w6(32'hba597f75),
	.w7(32'h3a7dbace),
	.w8(32'h3b634821),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf1991),
	.w1(32'h3bf542a3),
	.w2(32'h3c37abf3),
	.w3(32'h3b8122e4),
	.w4(32'h3bf291c9),
	.w5(32'h3c3da579),
	.w6(32'h3a9725d3),
	.w7(32'h3b82b7e6),
	.w8(32'h3c41c498),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c399db6),
	.w1(32'h3c2edf12),
	.w2(32'h3b19647c),
	.w3(32'h3c01432b),
	.w4(32'h3c052807),
	.w5(32'hbbcb2107),
	.w6(32'h3c212066),
	.w7(32'h3c10c5c8),
	.w8(32'h39a2251b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbec7b0),
	.w1(32'hbb3a1639),
	.w2(32'hb9f28942),
	.w3(32'hbc8642a6),
	.w4(32'hbc2cb25b),
	.w5(32'h3b99fe61),
	.w6(32'hbc1e82d1),
	.w7(32'hbbacfa46),
	.w8(32'h3b87facb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19c8b0),
	.w1(32'hbb02a592),
	.w2(32'h3ae1f878),
	.w3(32'hbb8ba3a3),
	.w4(32'h3b0352fe),
	.w5(32'h3a7a3e3b),
	.w6(32'hbb025232),
	.w7(32'h39ede85d),
	.w8(32'h3b58f7a1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977356a),
	.w1(32'h3b7e74f2),
	.w2(32'hb95debf8),
	.w3(32'h3ab41839),
	.w4(32'h3b83203c),
	.w5(32'hbb5f97bb),
	.w6(32'h3bb43f1e),
	.w7(32'h3bbb2a60),
	.w8(32'hbbb7d9f8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d211e),
	.w1(32'hbb9b63f7),
	.w2(32'h3b572e6f),
	.w3(32'hbb3ab16f),
	.w4(32'hbb66e382),
	.w5(32'h3b777ee8),
	.w6(32'hbabbc0dc),
	.w7(32'h3c04e979),
	.w8(32'h3b6e9521),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e2c95),
	.w1(32'h3b373ec6),
	.w2(32'h3b5d946a),
	.w3(32'h3a963aec),
	.w4(32'h3b5d07fc),
	.w5(32'h39cfc43f),
	.w6(32'h3b1260bf),
	.w7(32'h3b4c3b2c),
	.w8(32'h3ad7bab4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba985fb8),
	.w1(32'hba323296),
	.w2(32'hba067395),
	.w3(32'h3aa91982),
	.w4(32'hbb2ac8f4),
	.w5(32'h3b669c31),
	.w6(32'hb92c0c23),
	.w7(32'hb6b796de),
	.w8(32'h3c0276eb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba033503),
	.w1(32'hba7fbf88),
	.w2(32'h3a766a0d),
	.w3(32'hbb19d3f7),
	.w4(32'h3b86e3dd),
	.w5(32'h3b0c7cba),
	.w6(32'h3b6cdae0),
	.w7(32'h3a3ba367),
	.w8(32'h3bc853b9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaef6de),
	.w1(32'h3a3506ac),
	.w2(32'h3b6782fc),
	.w3(32'h3b0fafae),
	.w4(32'h3a4e9e85),
	.w5(32'h3a83a885),
	.w6(32'h3bc7d73d),
	.w7(32'h3b742196),
	.w8(32'h3a6954d0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc5469),
	.w1(32'hbb208242),
	.w2(32'h3b7e837f),
	.w3(32'hbb52733b),
	.w4(32'h3a738c4f),
	.w5(32'h3bce69cb),
	.w6(32'h3bb68953),
	.w7(32'hbbaa0389),
	.w8(32'h3a1bf0a8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4359b),
	.w1(32'h3b3ea3e6),
	.w2(32'h3bab73ae),
	.w3(32'hb872b4b8),
	.w4(32'h3b6a1fc0),
	.w5(32'hb8b5e347),
	.w6(32'h39ce1780),
	.w7(32'h3b12772a),
	.w8(32'h3af065b6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a5025),
	.w1(32'hb976b4c2),
	.w2(32'h3a92d20b),
	.w3(32'hbb888abe),
	.w4(32'h3b0da2f3),
	.w5(32'hbaf34952),
	.w6(32'hbaa3d781),
	.w7(32'hbb1b8f2d),
	.w8(32'hbac6c4c4),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c8096),
	.w1(32'h3b9ba01a),
	.w2(32'h3c839588),
	.w3(32'hbae0f513),
	.w4(32'hb9fb20b7),
	.w5(32'h3d502490),
	.w6(32'h3b1f898a),
	.w7(32'hba9ed68c),
	.w8(32'h3d0c6192),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4efe0c),
	.w1(32'h3ccb359d),
	.w2(32'h3b569549),
	.w3(32'h3dd6170f),
	.w4(32'h3d916adb),
	.w5(32'h39203e7f),
	.w6(32'h3daa1480),
	.w7(32'h3d49fafc),
	.w8(32'h3b5d6d5a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7e62f),
	.w1(32'h3ab96d9c),
	.w2(32'h3bb459a5),
	.w3(32'hbb38a791),
	.w4(32'h3a89c73f),
	.w5(32'h3bd6d1c7),
	.w6(32'h3b4d2803),
	.w7(32'h3ba829b4),
	.w8(32'h3beb206e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b2fe),
	.w1(32'h3b74d6ae),
	.w2(32'h3b8a08e6),
	.w3(32'h3ba06a43),
	.w4(32'h3b27d192),
	.w5(32'h3a8faa8c),
	.w6(32'h3b3dc8d3),
	.w7(32'h3b9db040),
	.w8(32'h3c02b182),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99f30d),
	.w1(32'h3aa6c75d),
	.w2(32'h3c127f09),
	.w3(32'hbb72f5b7),
	.w4(32'hba53ea07),
	.w5(32'h39df2a45),
	.w6(32'h3b1750d6),
	.w7(32'h3adf1b15),
	.w8(32'h3c051f61),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ddad7),
	.w1(32'h3bf4ba73),
	.w2(32'h3b8764aa),
	.w3(32'hbbfd1798),
	.w4(32'h3a477e80),
	.w5(32'hbab2c5c0),
	.w6(32'h38ca2213),
	.w7(32'h3bee34fd),
	.w8(32'h3b91430e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb0dcf),
	.w1(32'hb8965a54),
	.w2(32'hbb0347c4),
	.w3(32'hbad3c7fc),
	.w4(32'h3b476657),
	.w5(32'h3b49121b),
	.w6(32'h3b9984fc),
	.w7(32'h3b5c652e),
	.w8(32'h3ab13df1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8017e6),
	.w1(32'hb9229c91),
	.w2(32'h3b19b2ce),
	.w3(32'h3c404d2b),
	.w4(32'h3be799cc),
	.w5(32'hbb602a6a),
	.w6(32'h3c1f90f3),
	.w7(32'h3baaf1c1),
	.w8(32'h3a3167f1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfc883),
	.w1(32'h3a1a0166),
	.w2(32'h3ba93bbf),
	.w3(32'h3c57901c),
	.w4(32'hba66e8a5),
	.w5(32'h3b5dd6a4),
	.w6(32'h3bcec1e7),
	.w7(32'hbb1f9f79),
	.w8(32'h3b15f6fc),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b578045),
	.w1(32'h3aceb32c),
	.w2(32'h39e8b694),
	.w3(32'h39d6c920),
	.w4(32'h3b8be127),
	.w5(32'h3b437bed),
	.w6(32'h3a4d26a9),
	.w7(32'hbb32abdc),
	.w8(32'hbb0b702b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af826d1),
	.w1(32'hbaad9c8b),
	.w2(32'hbab78b9f),
	.w3(32'h388a5dcd),
	.w4(32'hba23656e),
	.w5(32'hbb8516ab),
	.w6(32'hbaa2ad4a),
	.w7(32'hba53afc2),
	.w8(32'h3a337c5c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2b69e),
	.w1(32'hba94e902),
	.w2(32'h3a3a1685),
	.w3(32'hbbd2952e),
	.w4(32'hba43e300),
	.w5(32'hb979cfc8),
	.w6(32'hbb3d6bd8),
	.w7(32'h3aca062d),
	.w8(32'hbb6fe37f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04856c),
	.w1(32'h3a8c5c78),
	.w2(32'hba2d6b8b),
	.w3(32'h3b705074),
	.w4(32'h3b302363),
	.w5(32'h3a9a9052),
	.w6(32'hba36db17),
	.w7(32'hbb2e1751),
	.w8(32'hbb4866b9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2712e7),
	.w1(32'h3a87aaf4),
	.w2(32'h37c49a57),
	.w3(32'h3aa89d28),
	.w4(32'h3b81a35d),
	.w5(32'h3af003d3),
	.w6(32'h39c5cf1c),
	.w7(32'h39011c42),
	.w8(32'h3b97fa16),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9099c8),
	.w1(32'h3aa59125),
	.w2(32'hbb6d7b2f),
	.w3(32'hbb521e7c),
	.w4(32'hbad1b56d),
	.w5(32'hba539ac8),
	.w6(32'h3b2c8caf),
	.w7(32'hbb6b122a),
	.w8(32'hba045577),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1731b),
	.w1(32'h3b42ce03),
	.w2(32'hbc10f7b5),
	.w3(32'h3b06596b),
	.w4(32'h3b3c3f63),
	.w5(32'hba253165),
	.w6(32'h3b446b18),
	.w7(32'h3afe9fe5),
	.w8(32'h3b87e1f3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e153df),
	.w1(32'hbb8b01c7),
	.w2(32'h387cd667),
	.w3(32'hbac19937),
	.w4(32'h3b13ef8d),
	.w5(32'hba68802d),
	.w6(32'hbbe5a281),
	.w7(32'hbb7797a9),
	.w8(32'hba1601f0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a764132),
	.w1(32'hba2152a7),
	.w2(32'h3bb4994d),
	.w3(32'hbb226a6c),
	.w4(32'h3b399d5f),
	.w5(32'hbba38fd8),
	.w6(32'hbbb0411f),
	.w7(32'h3aa69ac9),
	.w8(32'h3afb893d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca3d0),
	.w1(32'h3979aa8f),
	.w2(32'h37fef0f5),
	.w3(32'hbc85ce0d),
	.w4(32'hbc18ed86),
	.w5(32'h3bab98b0),
	.w6(32'hbc0d8f3b),
	.w7(32'hbb995867),
	.w8(32'hbb3abce9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16ed7e),
	.w1(32'hba6d912c),
	.w2(32'h3a1be5cf),
	.w3(32'h3b3873f7),
	.w4(32'h3b9e2713),
	.w5(32'hbaf4ea32),
	.w6(32'hb8919295),
	.w7(32'hbaa4a394),
	.w8(32'hba117d99),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a392865),
	.w1(32'h39edab95),
	.w2(32'h3b08c6cf),
	.w3(32'hbb47fd40),
	.w4(32'hbb277a53),
	.w5(32'h36b5186a),
	.w6(32'h3ab13425),
	.w7(32'hbbce2281),
	.w8(32'hbb5c3a18),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b745d),
	.w1(32'hb910786d),
	.w2(32'hb9d8046e),
	.w3(32'h3a25ca0e),
	.w4(32'hba7123fc),
	.w5(32'hba81a4e1),
	.w6(32'hb9f861b4),
	.w7(32'hba844f56),
	.w8(32'h3a012967),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67b4c1),
	.w1(32'hba235bdd),
	.w2(32'hbb193323),
	.w3(32'h3b03090a),
	.w4(32'hbac9ec75),
	.w5(32'hb90d37ff),
	.w6(32'h3b90b9f0),
	.w7(32'hb9c1171c),
	.w8(32'h3bae8b72),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b1cd5),
	.w1(32'h3c51918c),
	.w2(32'hbb016ecc),
	.w3(32'hbcc655a2),
	.w4(32'h3ad704a3),
	.w5(32'hbb9e02cb),
	.w6(32'hbcb5c96d),
	.w7(32'h3ac951ad),
	.w8(32'hbbfe5550),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4ee94),
	.w1(32'h3c21552d),
	.w2(32'h39418cba),
	.w3(32'hbc06833e),
	.w4(32'h3bd6fdf3),
	.w5(32'h3b4146f7),
	.w6(32'hbbd4f60b),
	.w7(32'h3c3650c1),
	.w8(32'h3b96dbf3),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef244b),
	.w1(32'hbbdea091),
	.w2(32'h3bef36b9),
	.w3(32'h3bd33099),
	.w4(32'hbc07413c),
	.w5(32'h3ac54eec),
	.w6(32'h3c44a153),
	.w7(32'hb9bcd037),
	.w8(32'hbb5e8c72),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd45d70),
	.w1(32'h3b873b6d),
	.w2(32'hbb1369cd),
	.w3(32'h3c25c91d),
	.w4(32'h3bb5881d),
	.w5(32'hbc0df653),
	.w6(32'h3c72ba11),
	.w7(32'h3bf69fcb),
	.w8(32'h3b5360ea),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a272b),
	.w1(32'h3c2bf9bb),
	.w2(32'h3a0ced1e),
	.w3(32'h3b82ef88),
	.w4(32'h3c4dbd22),
	.w5(32'h3aef4ed1),
	.w6(32'h38feac35),
	.w7(32'h3bfa99d9),
	.w8(32'h3bcb79ee),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b3b25),
	.w1(32'hba771388),
	.w2(32'h3c56484f),
	.w3(32'hbaf903a8),
	.w4(32'hbb33bc66),
	.w5(32'h3c5eb214),
	.w6(32'h3b595b3c),
	.w7(32'h37d277a7),
	.w8(32'h3c50e12f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c928d1b),
	.w1(32'hbab4c5be),
	.w2(32'hbb5de74b),
	.w3(32'h3d07edad),
	.w4(32'hbafcd70c),
	.w5(32'hbbac001b),
	.w6(32'h3d024c8a),
	.w7(32'hba507877),
	.w8(32'hbb0f2e67),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab2494),
	.w1(32'h3b4a63c9),
	.w2(32'hb9762325),
	.w3(32'hbb929ebf),
	.w4(32'h3b07224c),
	.w5(32'hbbaf1b18),
	.w6(32'hbc05125a),
	.w7(32'hb950284f),
	.w8(32'h3b3c4f4a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3877f),
	.w1(32'hbb697bbb),
	.w2(32'hbba668e8),
	.w3(32'hbbb762ac),
	.w4(32'h3ad467ca),
	.w5(32'hbc130988),
	.w6(32'h3b54c787),
	.w7(32'hbb68e844),
	.w8(32'hbb9834cf),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99443f),
	.w1(32'h3c3bd63b),
	.w2(32'h3b97696e),
	.w3(32'h3af6f9d5),
	.w4(32'h3c16782c),
	.w5(32'h3b14f456),
	.w6(32'h3b340f5d),
	.w7(32'h3c428326),
	.w8(32'hbba676ad),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2f9ad),
	.w1(32'hbb1ea9af),
	.w2(32'hbc9a8195),
	.w3(32'h3b6b478d),
	.w4(32'hbbd61313),
	.w5(32'hbc70ec33),
	.w6(32'hbb6800ba),
	.w7(32'hbbdb8cd1),
	.w8(32'hbc7a4522),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20f2cc),
	.w1(32'h3b4c7521),
	.w2(32'h3c0a6dc3),
	.w3(32'h3bd2c25d),
	.w4(32'h3c1b50ce),
	.w5(32'h3c2326a2),
	.w6(32'hbc55188e),
	.w7(32'h3bee858d),
	.w8(32'h3b3f38b5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87b49e),
	.w1(32'hbc030e1e),
	.w2(32'hbc1c5cf1),
	.w3(32'h3bdeb017),
	.w4(32'hbc2fd835),
	.w5(32'hbb4a6ff1),
	.w6(32'h3c900636),
	.w7(32'h39c99476),
	.w8(32'hbc287047),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43e5fc),
	.w1(32'hbb5c29ae),
	.w2(32'hbb8ffa7a),
	.w3(32'h3c3c3a48),
	.w4(32'h3b8ac164),
	.w5(32'hbbc83561),
	.w6(32'h3c6cc3f2),
	.w7(32'h3c575275),
	.w8(32'hbba1e6f3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3892eff2),
	.w1(32'h3a67f7bb),
	.w2(32'hbad0a131),
	.w3(32'hbbd24936),
	.w4(32'hbb368af6),
	.w5(32'hbb6df71b),
	.w6(32'hbbaa3b84),
	.w7(32'hbb9302fd),
	.w8(32'hbbf064ae),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb0b25),
	.w1(32'h3c252ec3),
	.w2(32'hbbd99307),
	.w3(32'hbb0fd1b6),
	.w4(32'h3c1222af),
	.w5(32'hbc45be2c),
	.w6(32'hbc25ad5c),
	.w7(32'h3b224d79),
	.w8(32'hbc5d4892),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f56c4),
	.w1(32'h3b65965e),
	.w2(32'h3b906d15),
	.w3(32'hbb003b05),
	.w4(32'h39cd513c),
	.w5(32'h3b5385be),
	.w6(32'hbbb05f1d),
	.w7(32'h3bf8371c),
	.w8(32'hbc20bec8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac33ca),
	.w1(32'hbc0d5306),
	.w2(32'hba89ce65),
	.w3(32'h3b525eca),
	.w4(32'hbbdd39aa),
	.w5(32'h3c42e58b),
	.w6(32'h3b803808),
	.w7(32'h3c296253),
	.w8(32'h3b48b154),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94ec02),
	.w1(32'h3b229f55),
	.w2(32'h3c432a02),
	.w3(32'hbc7360c2),
	.w4(32'h3a8f4371),
	.w5(32'h3c2407ac),
	.w6(32'hbc27e6c3),
	.w7(32'hbc2ee7c8),
	.w8(32'h3bc6c969),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfceaef),
	.w1(32'hbc850ef8),
	.w2(32'hb9e20de6),
	.w3(32'h3cbff8e3),
	.w4(32'hbc65d3cd),
	.w5(32'hbb683a67),
	.w6(32'h3d14261c),
	.w7(32'hb9dca462),
	.w8(32'hbbe5eea8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba23023),
	.w1(32'h3c231542),
	.w2(32'hbc00df96),
	.w3(32'hba76719b),
	.w4(32'h3c7247f4),
	.w5(32'hbc3a7e22),
	.w6(32'hbbd1619e),
	.w7(32'h3bc892a1),
	.w8(32'hbc182851),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefdbb5),
	.w1(32'h3b259098),
	.w2(32'hbb55fea4),
	.w3(32'hb6d07307),
	.w4(32'h3bba1034),
	.w5(32'h3ab72eac),
	.w6(32'hbc06beb9),
	.w7(32'h398b5612),
	.w8(32'h3ae10c53),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021505),
	.w1(32'hbaae270a),
	.w2(32'hbc2e941b),
	.w3(32'h3bffe73e),
	.w4(32'hbc2c017e),
	.w5(32'hbc2607fd),
	.w6(32'h3b82fb08),
	.w7(32'hbae8847d),
	.w8(32'hbb2874e6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc70e86),
	.w1(32'hb92c052e),
	.w2(32'hbbf3c51a),
	.w3(32'hbc825610),
	.w4(32'hbb1cf184),
	.w5(32'h3bbe2acd),
	.w6(32'hbb92496f),
	.w7(32'h3a324578),
	.w8(32'hbaab8237),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44ccbd),
	.w1(32'hbbda89d2),
	.w2(32'h3b4cb2fc),
	.w3(32'h3c0c7128),
	.w4(32'hbb5febfa),
	.w5(32'h3bb645ed),
	.w6(32'h3ae98ada),
	.w7(32'h39dfb1aa),
	.w8(32'h3b84c30f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec8018),
	.w1(32'hbb880144),
	.w2(32'hbabc5cc0),
	.w3(32'h3ba2494b),
	.w4(32'hbbe1986d),
	.w5(32'h3b4bcde6),
	.w6(32'h3bd0fc16),
	.w7(32'hbc2440e9),
	.w8(32'hbbb674d3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc687f5b),
	.w1(32'hbbfff01a),
	.w2(32'h3c4be11c),
	.w3(32'hbb054987),
	.w4(32'h3ba3ba0e),
	.w5(32'h3bba38ad),
	.w6(32'h3ab574e8),
	.w7(32'hbb7c09f3),
	.w8(32'h3b32b9fc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ccdc1),
	.w1(32'hbbc4ec80),
	.w2(32'hbbd1ba32),
	.w3(32'h3b09fc9b),
	.w4(32'hbbc1d037),
	.w5(32'h38fc88e2),
	.w6(32'h3bb825d9),
	.w7(32'hbbaf7bc1),
	.w8(32'hbc1ff7a1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c414743),
	.w1(32'h3ccb52dc),
	.w2(32'hbb499d73),
	.w3(32'hbc847aba),
	.w4(32'h3d182fa3),
	.w5(32'h3911c328),
	.w6(32'hbc72db81),
	.w7(32'h3cc1af1b),
	.w8(32'hbb87ae8b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38227a),
	.w1(32'hbbcbb04f),
	.w2(32'hbae37512),
	.w3(32'h3bb5ecd9),
	.w4(32'hbc2dd8dc),
	.w5(32'hb9fde070),
	.w6(32'h3c346f77),
	.w7(32'hbc46c0fa),
	.w8(32'hba97ee4a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51ee9b),
	.w1(32'h3c5e4b0f),
	.w2(32'hbc585684),
	.w3(32'h3ac1452e),
	.w4(32'h3c76c0bd),
	.w5(32'hbc01e677),
	.w6(32'h3bb5dfdc),
	.w7(32'h3c871929),
	.w8(32'hbb6aaf06),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd995dc),
	.w1(32'hbc0faaec),
	.w2(32'h3b86af20),
	.w3(32'h3b9f5876),
	.w4(32'hba8dee9b),
	.w5(32'h3c3961b5),
	.w6(32'h3b67e6b7),
	.w7(32'hb97af4bd),
	.w8(32'h3c0b7620),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8abf994),
	.w1(32'hbbdee54a),
	.w2(32'h39c9b5f4),
	.w3(32'h3c0fb953),
	.w4(32'hbc731485),
	.w5(32'h3ba7f571),
	.w6(32'h3ca904f6),
	.w7(32'hbbde3a3d),
	.w8(32'h3b8df0f8),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe63abb),
	.w1(32'hbb90602b),
	.w2(32'hbb89cfc4),
	.w3(32'hbc05d5d6),
	.w4(32'hbb8d177a),
	.w5(32'h3be604e6),
	.w6(32'hbbf2f550),
	.w7(32'hbbb9732a),
	.w8(32'h3bc28fb9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be906a6),
	.w1(32'h3c914e48),
	.w2(32'hbb95d5dd),
	.w3(32'h39cb7859),
	.w4(32'h3c012a0d),
	.w5(32'hba51012d),
	.w6(32'h3bfcabcc),
	.w7(32'hba81d81a),
	.w8(32'h3a966954),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedf938),
	.w1(32'h3adaedfa),
	.w2(32'hb9475e8d),
	.w3(32'hba233ca3),
	.w4(32'hba54d946),
	.w5(32'hbc09c172),
	.w6(32'h3aadb9cd),
	.w7(32'h3a79d7b3),
	.w8(32'hbbf1da4c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb9aac),
	.w1(32'hbc444de2),
	.w2(32'h3afc2443),
	.w3(32'hbc1e45c0),
	.w4(32'hbbab41b0),
	.w5(32'h3b269f88),
	.w6(32'h3b8999ad),
	.w7(32'hbbac831f),
	.w8(32'h3b8efe74),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa97778),
	.w1(32'h3b13d822),
	.w2(32'h3a1c2ca0),
	.w3(32'hbbfe94b3),
	.w4(32'hbb5a7dca),
	.w5(32'hbad0ae3c),
	.w6(32'hbbb259dd),
	.w7(32'hbbad9220),
	.w8(32'hbbbfd74c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac709e),
	.w1(32'h3c4d80a7),
	.w2(32'hbc6874eb),
	.w3(32'h3a73e0aa),
	.w4(32'h3c16bb0b),
	.w5(32'h3b09dfdc),
	.w6(32'hbbbcfa5e),
	.w7(32'h3bdc76d5),
	.w8(32'h3b1fb6e6),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe530f3),
	.w1(32'hbc583899),
	.w2(32'h3b0a51fc),
	.w3(32'hbc26e220),
	.w4(32'hbc84ed03),
	.w5(32'h3bb2abea),
	.w6(32'hbc82809b),
	.w7(32'hbc2829a1),
	.w8(32'hbb3890d4),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c252db3),
	.w1(32'h3b7bcd4c),
	.w2(32'h3a907d57),
	.w3(32'h3c1d3a3d),
	.w4(32'h3bac6aa7),
	.w5(32'h3aca279f),
	.w6(32'h3bc9b9c5),
	.w7(32'hbb0adaff),
	.w8(32'h3a1a27fe),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf64335),
	.w1(32'hb9d4dc51),
	.w2(32'hbca2a586),
	.w3(32'h3bc63417),
	.w4(32'hbac90bea),
	.w5(32'hbce30dbe),
	.w6(32'h3bb6e711),
	.w7(32'hba0589ef),
	.w8(32'hbcca3005),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9533449),
	.w1(32'h3c569f0d),
	.w2(32'hbbb45635),
	.w3(32'hba868d40),
	.w4(32'h3c15f74c),
	.w5(32'hba71c473),
	.w6(32'hbbae4e97),
	.w7(32'h3c15c495),
	.w8(32'h3bd0b6dd),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56b944),
	.w1(32'h3acea9f1),
	.w2(32'h3cbae925),
	.w3(32'hbccb43b0),
	.w4(32'hbbf5aa5e),
	.w5(32'h3cefc8ae),
	.w6(32'hbc719862),
	.w7(32'hbbdb2a25),
	.w8(32'h3cbbf6be),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabf601),
	.w1(32'hbbbf58c2),
	.w2(32'hbc90da80),
	.w3(32'hbb395393),
	.w4(32'hbc439801),
	.w5(32'hbcc39c46),
	.w6(32'h3b46d6d0),
	.w7(32'hbc785b76),
	.w8(32'hbcc27597),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c918676),
	.w1(32'h3c135943),
	.w2(32'hb9e3924a),
	.w3(32'h3c6a9867),
	.w4(32'h3c87ed03),
	.w5(32'hbbd7ca89),
	.w6(32'h3b025f25),
	.w7(32'h3c6a938d),
	.w8(32'hbbe206b6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1db7a3),
	.w1(32'h3a785395),
	.w2(32'h3b8bedd6),
	.w3(32'h3a612c2c),
	.w4(32'h3b8ece01),
	.w5(32'h3c28d492),
	.w6(32'hbb5caf4a),
	.w7(32'h3b087b14),
	.w8(32'h3c7843bf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb9528),
	.w1(32'hbb3c411f),
	.w2(32'hba75d92e),
	.w3(32'hbc395cd9),
	.w4(32'hbbd0af38),
	.w5(32'hbb543fac),
	.w6(32'h39985be3),
	.w7(32'hbc14b651),
	.w8(32'hbb91574a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aa577),
	.w1(32'h3c211934),
	.w2(32'h3ac6f050),
	.w3(32'h3a51c4e7),
	.w4(32'h3b334892),
	.w5(32'h3b7ddcdd),
	.w6(32'h3bf117ea),
	.w7(32'h390a0df6),
	.w8(32'h3ae42915),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90b11e),
	.w1(32'h3b9c7f72),
	.w2(32'h3c7231fe),
	.w3(32'h3c8af4e0),
	.w4(32'h3bd5dfa4),
	.w5(32'h3c4b746e),
	.w6(32'h3c95f0b9),
	.w7(32'h3c05776e),
	.w8(32'hbbbb8136),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8e23b),
	.w1(32'h3b32343a),
	.w2(32'hb94687ad),
	.w3(32'h3c8124a7),
	.w4(32'hbb89f4c4),
	.w5(32'hbbb8a0bf),
	.w6(32'h3cd2edf3),
	.w7(32'h3adf9b2b),
	.w8(32'h3a05efcd),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2f300),
	.w1(32'hb7707be8),
	.w2(32'hbaddf261),
	.w3(32'hba86afef),
	.w4(32'hbbfd3905),
	.w5(32'hbbeb091d),
	.w6(32'h3be7fea5),
	.w7(32'h3a364a71),
	.w8(32'hbc302884),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb10185),
	.w1(32'h3b58330a),
	.w2(32'hbac9c730),
	.w3(32'h3c0d2be8),
	.w4(32'h3c50e8e2),
	.w5(32'hba0c5a5d),
	.w6(32'h3bcd69f5),
	.w7(32'h3c0788d6),
	.w8(32'h3aba714e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1da4bd),
	.w1(32'hbbbd1912),
	.w2(32'h3ba2fc19),
	.w3(32'h3b1bcd3a),
	.w4(32'hbc32882f),
	.w5(32'h3c6cc717),
	.w6(32'h3bba3cab),
	.w7(32'hbba609e5),
	.w8(32'h3c66f14b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f433),
	.w1(32'hbc79110a),
	.w2(32'hbb6dd7b0),
	.w3(32'hbbf919fc),
	.w4(32'hbc97e6ae),
	.w5(32'hbc1ee7fb),
	.w6(32'h3b89e878),
	.w7(32'hbcc6cdc5),
	.w8(32'hbb58dd0b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b0960),
	.w1(32'hbbd11888),
	.w2(32'h3bdd6bae),
	.w3(32'hbc9b5e3f),
	.w4(32'hbc182d76),
	.w5(32'h3ca9bd8c),
	.w6(32'hbc9327e8),
	.w7(32'hbc86014a),
	.w8(32'h3baf98ac),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29cc3a),
	.w1(32'h3bf413b8),
	.w2(32'h3c04ecc8),
	.w3(32'hbc291b3c),
	.w4(32'hbb441007),
	.w5(32'h3ca9a518),
	.w6(32'h3b87bae1),
	.w7(32'hbc454b60),
	.w8(32'h3cfb89c1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd8a19),
	.w1(32'hbb50b05f),
	.w2(32'h38b83595),
	.w3(32'hbc89bd7d),
	.w4(32'h3983857a),
	.w5(32'h3bdbf66a),
	.w6(32'hbca21c2b),
	.w7(32'hbb5373f2),
	.w8(32'h3c577d05),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec9299),
	.w1(32'hbb574633),
	.w2(32'h3bb16d0e),
	.w3(32'hbc4945e4),
	.w4(32'hbbbc3c97),
	.w5(32'h3b418022),
	.w6(32'hbb91d195),
	.w7(32'hbc029adf),
	.w8(32'h3b0d39eb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad53e41),
	.w1(32'hba72cf55),
	.w2(32'h3a45bb97),
	.w3(32'h3a5abbf0),
	.w4(32'hbb4074ba),
	.w5(32'h399c79ef),
	.w6(32'h3af2b149),
	.w7(32'hb800e145),
	.w8(32'hbb35d19a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab47d8e),
	.w1(32'hbc36d0eb),
	.w2(32'hbb80bdb4),
	.w3(32'hbad7cdbb),
	.w4(32'hbc2fac9c),
	.w5(32'hbbb547e4),
	.w6(32'hbbca49c6),
	.w7(32'hbc202da8),
	.w8(32'h3b9234ec),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef4d1d),
	.w1(32'h3b501c49),
	.w2(32'hbb4ce9f9),
	.w3(32'hbc0812b5),
	.w4(32'hbc52e2d5),
	.w5(32'hbbc78e7d),
	.w6(32'hbc4f2ef7),
	.w7(32'hbca8e2d3),
	.w8(32'h3925e07c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b25a6b),
	.w1(32'h3b56ba05),
	.w2(32'h3c025a53),
	.w3(32'hbb18f512),
	.w4(32'h3a071526),
	.w5(32'hbb157985),
	.w6(32'hbb2480a8),
	.w7(32'hbb85abf6),
	.w8(32'hbbc3d269),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1eade),
	.w1(32'h3c0311e3),
	.w2(32'h3b0c7239),
	.w3(32'h3cbbc430),
	.w4(32'h3bd93ea1),
	.w5(32'h3b905956),
	.w6(32'h3caf42bb),
	.w7(32'h3c3bce6b),
	.w8(32'h3b99f0b7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4e1ad),
	.w1(32'hbc3b40c5),
	.w2(32'h3ad05d35),
	.w3(32'hbbb2bf04),
	.w4(32'hbc5983f0),
	.w5(32'h3b7b3e5b),
	.w6(32'h3a17f29a),
	.w7(32'hbb893ef8),
	.w8(32'h3b123f23),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaef5c),
	.w1(32'hbbb3f18a),
	.w2(32'h3c0647af),
	.w3(32'h3c0182e4),
	.w4(32'hbbe28747),
	.w5(32'h3b45bd10),
	.w6(32'h3c1d1457),
	.w7(32'h392b3e22),
	.w8(32'h3b5dd232),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c040b94),
	.w1(32'h3baba555),
	.w2(32'h3bd9fb16),
	.w3(32'h3bb1d19a),
	.w4(32'h3a3a3eb0),
	.w5(32'h3c576648),
	.w6(32'h3bf5fbbd),
	.w7(32'h3aebae33),
	.w8(32'h3bb51169),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebcdb2),
	.w1(32'h3bc83eee),
	.w2(32'h3a07b731),
	.w3(32'hba0b6847),
	.w4(32'h38d76c44),
	.w5(32'hbace47b8),
	.w6(32'hbc05c80f),
	.w7(32'hbc5d0d49),
	.w8(32'hbbc6c001),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc027986),
	.w1(32'h3b6c59b7),
	.w2(32'hbc33391b),
	.w3(32'hbc1a8d7b),
	.w4(32'h39fc6fcb),
	.w5(32'hbb319cda),
	.w6(32'hbc43601b),
	.w7(32'h3aa01c88),
	.w8(32'hbadb6837),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8588ab),
	.w1(32'h3bcf792a),
	.w2(32'h3b646ad4),
	.w3(32'hbce04ba1),
	.w4(32'hbac54f9f),
	.w5(32'hbb87dc38),
	.w6(32'hbbd4a0cc),
	.w7(32'hbc9546d2),
	.w8(32'hbbcbe8cc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81ddc4),
	.w1(32'hba2b55a2),
	.w2(32'hbb0956bb),
	.w3(32'h3c60223d),
	.w4(32'h3b7cfc14),
	.w5(32'hbc86a8cc),
	.w6(32'h3c133830),
	.w7(32'h3a97263c),
	.w8(32'hbc85ecc6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2a767),
	.w1(32'h3c4e6536),
	.w2(32'h3b294f2a),
	.w3(32'h3ca3d4a0),
	.w4(32'h3cbd6f97),
	.w5(32'hbc0e5cbf),
	.w6(32'h3bce06a3),
	.w7(32'h3cc44924),
	.w8(32'hbc6202b0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1884b),
	.w1(32'hbb477dd9),
	.w2(32'h3b969436),
	.w3(32'hbb216873),
	.w4(32'hbc21f054),
	.w5(32'h3aa858cc),
	.w6(32'hbbdb9952),
	.w7(32'h3c02e843),
	.w8(32'h3ab9e431),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8400be),
	.w1(32'hbbdb5002),
	.w2(32'hbaf8e5f8),
	.w3(32'h3c1c68ca),
	.w4(32'h3b418204),
	.w5(32'hbc057d11),
	.w6(32'h3bc8bbd4),
	.w7(32'h3b92a9b1),
	.w8(32'hbb2ea002),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a1f30),
	.w1(32'h3c030077),
	.w2(32'hbb2abd01),
	.w3(32'hbc9512da),
	.w4(32'h3ad90384),
	.w5(32'hbbbd8f40),
	.w6(32'hbc5ffffc),
	.w7(32'hb98aae5c),
	.w8(32'hbc1c813a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7da625),
	.w1(32'h3b828130),
	.w2(32'hba620d92),
	.w3(32'h3be0c364),
	.w4(32'h3c2b437c),
	.w5(32'h3bb7787d),
	.w6(32'h3b5ebaf6),
	.w7(32'h3bfb927c),
	.w8(32'h3a044043),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc147513),
	.w1(32'hb988e746),
	.w2(32'hbba20357),
	.w3(32'hbc2f0964),
	.w4(32'hbb7d67d5),
	.w5(32'hba9debe1),
	.w6(32'hbc7beb92),
	.w7(32'hbbb401d9),
	.w8(32'h3a26c2f7),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a08b1),
	.w1(32'h3b39d84e),
	.w2(32'hbba2429b),
	.w3(32'hbc5bc378),
	.w4(32'hbaade1bd),
	.w5(32'h39838df5),
	.w6(32'hbc229849),
	.w7(32'hbbf968d6),
	.w8(32'h3bba3e11),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55d76e),
	.w1(32'h3c07c6bc),
	.w2(32'hbbee1529),
	.w3(32'hbc83d2ae),
	.w4(32'h3b128264),
	.w5(32'h3be23f77),
	.w6(32'hbc48e037),
	.w7(32'hbb699da6),
	.w8(32'hb9a68a87),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b504c10),
	.w1(32'h3c8a73f5),
	.w2(32'hbc2ff6d8),
	.w3(32'h3b496969),
	.w4(32'h3cc77fba),
	.w5(32'hbb71d57f),
	.w6(32'hbc07610c),
	.w7(32'h3c0b4231),
	.w8(32'h3bf1cd01),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf2629),
	.w1(32'h3c2605d9),
	.w2(32'hbbb889cd),
	.w3(32'hbc80f304),
	.w4(32'h3ca2ab35),
	.w5(32'hbb4d28c3),
	.w6(32'hbc75c678),
	.w7(32'h3c8c291b),
	.w8(32'hbab33f7c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e860b),
	.w1(32'hbbbe0561),
	.w2(32'hbc88856c),
	.w3(32'h3b2c286c),
	.w4(32'hbbadf30e),
	.w5(32'hbb66f183),
	.w6(32'h3bec860a),
	.w7(32'hbb6f7add),
	.w8(32'hbb36ae99),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d21d9f),
	.w1(32'h3c117c9b),
	.w2(32'hbaeafcfc),
	.w3(32'hbcadc6a8),
	.w4(32'hbb3c0bf0),
	.w5(32'h3ba1e3d8),
	.w6(32'hbc20ca22),
	.w7(32'hbc449798),
	.w8(32'h3bbd1785),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67ef90),
	.w1(32'hbb983e33),
	.w2(32'hbc2e8ea2),
	.w3(32'h39f121af),
	.w4(32'hbb11c1de),
	.w5(32'hbc4251f3),
	.w6(32'hbb82437a),
	.w7(32'hbb5ba66a),
	.w8(32'hbc558294),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d6c59),
	.w1(32'hbafc5215),
	.w2(32'hbc54c32c),
	.w3(32'hbc407e8b),
	.w4(32'hbb5f4e9f),
	.w5(32'hbc539959),
	.w6(32'h3a71f51a),
	.w7(32'hba6a99b7),
	.w8(32'hbc304fd1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1d48a),
	.w1(32'hbb43b0a8),
	.w2(32'hbc51c511),
	.w3(32'hbbeca82e),
	.w4(32'hbc147ecf),
	.w5(32'hbca533a1),
	.w6(32'hbca68a33),
	.w7(32'hbc659f65),
	.w8(32'hbca18b81),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af60a79),
	.w1(32'h3c5a34d0),
	.w2(32'hbb6e2de7),
	.w3(32'hbb3e78dd),
	.w4(32'h3c38d7bb),
	.w5(32'hbb40380c),
	.w6(32'hbbf1e82c),
	.w7(32'h3c162ccc),
	.w8(32'hbc027d75),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b243d),
	.w1(32'h3be0433e),
	.w2(32'h3b17b065),
	.w3(32'h3bd9f74e),
	.w4(32'h3c17b034),
	.w5(32'hbbc9fe15),
	.w6(32'hb89e92b1),
	.w7(32'h3be1a636),
	.w8(32'hbbe5957c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd16552),
	.w1(32'h3b4abb01),
	.w2(32'hbbac70b9),
	.w3(32'hbaaa2b41),
	.w4(32'hbbb6c42a),
	.w5(32'h3ac3197d),
	.w6(32'h3b733e3f),
	.w7(32'hbab8aed5),
	.w8(32'hbb904aaa),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a506226),
	.w1(32'h3b582655),
	.w2(32'h3bd645f9),
	.w3(32'h3bea9d4a),
	.w4(32'h3bd5b36c),
	.w5(32'h3bf33773),
	.w6(32'h3b8189f1),
	.w7(32'h3ba1ab80),
	.w8(32'h3af3dfcd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba15dad),
	.w1(32'hb98a7675),
	.w2(32'h3b9a3590),
	.w3(32'h3cba1d9c),
	.w4(32'h3b35c338),
	.w5(32'hbb98282b),
	.w6(32'h3c89d91e),
	.w7(32'hb93b2364),
	.w8(32'hbc1c572a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21ecb6),
	.w1(32'hbbab1813),
	.w2(32'h3ac63a8f),
	.w3(32'h3b97298e),
	.w4(32'hbbb08ee8),
	.w5(32'hba62a224),
	.w6(32'h3bd953b6),
	.w7(32'h3c86687d),
	.w8(32'h3c0101b6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0b938),
	.w1(32'h3c430efe),
	.w2(32'h3b633c72),
	.w3(32'hbb9bf3ec),
	.w4(32'h3b9b27b9),
	.w5(32'h3acf9599),
	.w6(32'h3c057dec),
	.w7(32'h3bd5003c),
	.w8(32'h39f8ea98),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b306431),
	.w1(32'hbab21757),
	.w2(32'h3806e09c),
	.w3(32'h3bda6a22),
	.w4(32'h3b536591),
	.w5(32'h3b0a1d35),
	.w6(32'h3ba67406),
	.w7(32'h3b863684),
	.w8(32'h3af7fb46),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b0eac),
	.w1(32'hbbe028de),
	.w2(32'h3c9aff4d),
	.w3(32'h3a1ec9a1),
	.w4(32'hbc114c7e),
	.w5(32'h3cc2786a),
	.w6(32'h3bac206e),
	.w7(32'hbbba26c5),
	.w8(32'h3bb2701c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb93615),
	.w1(32'hbd08f8b7),
	.w2(32'hbbbb2c6b),
	.w3(32'h3bc51efc),
	.w4(32'hbd2b09f6),
	.w5(32'hbb0d884c),
	.w6(32'h3c80cbec),
	.w7(32'hbce3f064),
	.w8(32'hbb40f65d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf46220),
	.w1(32'h379eb935),
	.w2(32'hbc24901e),
	.w3(32'hbc041595),
	.w4(32'hbb50e27d),
	.w5(32'hbc11ba93),
	.w6(32'hbbcda19a),
	.w7(32'hbbb3bcdc),
	.w8(32'hbc3d1c86),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b8528),
	.w1(32'hbc5a7af7),
	.w2(32'hbb014372),
	.w3(32'hbcb15e68),
	.w4(32'hbc8fcc4e),
	.w5(32'h3c019add),
	.w6(32'hbc7d8960),
	.w7(32'hbc84c6e8),
	.w8(32'h3c07a965),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6622d7),
	.w1(32'hbc7fe7c2),
	.w2(32'h3b887e98),
	.w3(32'hbc901e1f),
	.w4(32'hbc953620),
	.w5(32'h3c23a209),
	.w6(32'hbc0b41d5),
	.w7(32'hbc91ae18),
	.w8(32'h3be8b8aa),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a8c10),
	.w1(32'hbbedc2a9),
	.w2(32'hbc298e39),
	.w3(32'hbcad347e),
	.w4(32'hbc3561bc),
	.w5(32'h3bad47a1),
	.w6(32'hbc83be5b),
	.w7(32'hbc471292),
	.w8(32'h3be7dc5e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule