module layer_8_featuremap_169(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3da39),
	.w1(32'hb9c5f3e7),
	.w2(32'h3b8c5993),
	.w3(32'h3c142143),
	.w4(32'h3a2b5352),
	.w5(32'hbb44b7a2),
	.w6(32'hba0bfb48),
	.w7(32'h3a86c272),
	.w8(32'h3ae20fc4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2c14),
	.w1(32'hbbb5aff2),
	.w2(32'hbb8d15d6),
	.w3(32'hba82228c),
	.w4(32'hbbb43861),
	.w5(32'hbbaf858d),
	.w6(32'hbbc31f05),
	.w7(32'hbafd6f28),
	.w8(32'h3a82be68),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebdb14),
	.w1(32'hbb2d818a),
	.w2(32'h3a4451c6),
	.w3(32'hbc166b70),
	.w4(32'hbbb592d8),
	.w5(32'hbb8a09f3),
	.w6(32'hbc36064b),
	.w7(32'hbb9f2991),
	.w8(32'hbb7e580b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eb797),
	.w1(32'hbb51e900),
	.w2(32'hbabbece8),
	.w3(32'h3aa26901),
	.w4(32'h3ac2c1cf),
	.w5(32'h3bc33673),
	.w6(32'h3b58fa8b),
	.w7(32'hbb80b431),
	.w8(32'hbba8f0f9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3084e),
	.w1(32'hbb307b08),
	.w2(32'hbb5405aa),
	.w3(32'h3bcd5bdd),
	.w4(32'hb9c0d790),
	.w5(32'hbaa5b2ea),
	.w6(32'hbb628301),
	.w7(32'hbae0fb40),
	.w8(32'hba3066a3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7246f4),
	.w1(32'h3b2c0d93),
	.w2(32'h3c4a2a0e),
	.w3(32'hbabb0983),
	.w4(32'h3c1b2e1d),
	.w5(32'h3c13960d),
	.w6(32'hbac07ff6),
	.w7(32'h3bd1fc4b),
	.w8(32'h3bb07721),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c198cb4),
	.w1(32'hba2d948a),
	.w2(32'hbaeaacf4),
	.w3(32'hb9e65808),
	.w4(32'hbb237ad0),
	.w5(32'h3803466d),
	.w6(32'hbab07900),
	.w7(32'hbb1e4d26),
	.w8(32'hbb33c77e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3f49f),
	.w1(32'h3b0a57c3),
	.w2(32'h3bb2359b),
	.w3(32'hbb8868de),
	.w4(32'h3aa66efc),
	.w5(32'h39b33036),
	.w6(32'h3b00c198),
	.w7(32'h3bc5f183),
	.w8(32'h3c05ee8e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb638f8b),
	.w1(32'hbbef4b3d),
	.w2(32'hbb3817e9),
	.w3(32'hbbc3df0a),
	.w4(32'hbbbb52a2),
	.w5(32'h3aadec42),
	.w6(32'hbc4aefce),
	.w7(32'hbbcb4cc1),
	.w8(32'hbbb927c8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83250e),
	.w1(32'h3c1628f2),
	.w2(32'h3c277d56),
	.w3(32'hbaee4e3a),
	.w4(32'h3c685093),
	.w5(32'h3ca36e43),
	.w6(32'hbbc9d945),
	.w7(32'h390233c2),
	.w8(32'hbab2d2b1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68357c),
	.w1(32'hbb4f2fc0),
	.w2(32'h3729cf09),
	.w3(32'h3cb83f0a),
	.w4(32'hbbd971c3),
	.w5(32'hbc11c625),
	.w6(32'h3bda4eb4),
	.w7(32'h3b2a2a03),
	.w8(32'hbb124377),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b154ffa),
	.w1(32'h39f96508),
	.w2(32'hba295a7d),
	.w3(32'hba796b2e),
	.w4(32'h3b587e26),
	.w5(32'h3b1fee05),
	.w6(32'hba27ade1),
	.w7(32'h3b15c61e),
	.w8(32'h3b524893),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0813a6),
	.w1(32'hbc410d80),
	.w2(32'hbc35f064),
	.w3(32'hbad035e0),
	.w4(32'h3c0c8788),
	.w5(32'h3c115e52),
	.w6(32'hbc60f280),
	.w7(32'hbc059c4f),
	.w8(32'hbbf4483d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a0d3f),
	.w1(32'hbb17c98f),
	.w2(32'hba0cc8a0),
	.w3(32'h39dc34be),
	.w4(32'hbac3fd17),
	.w5(32'hbbac0bbf),
	.w6(32'hbbbf0c1f),
	.w7(32'h3b66962e),
	.w8(32'hb98f7d0d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9af9a4),
	.w1(32'h3a999930),
	.w2(32'h3bb89840),
	.w3(32'hbb8322a9),
	.w4(32'h39e6a0a6),
	.w5(32'h3be7b282),
	.w6(32'h397c0dc7),
	.w7(32'h3af2fc89),
	.w8(32'h3b37304c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b835b52),
	.w1(32'hbae3286b),
	.w2(32'h3ac1396e),
	.w3(32'h3bc8c54e),
	.w4(32'hbb5153e0),
	.w5(32'hbbf5e8c9),
	.w6(32'h38b52fd8),
	.w7(32'hbae0d76d),
	.w8(32'hba81526a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7579d),
	.w1(32'h39d2c168),
	.w2(32'hbb014300),
	.w3(32'hbbc59b6d),
	.w4(32'h3ad9bb7e),
	.w5(32'h3b5f0300),
	.w6(32'h3b7b3256),
	.w7(32'hbb8f182b),
	.w8(32'hbb16a6d5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3db85d),
	.w1(32'hbadb10b7),
	.w2(32'hbb3549bf),
	.w3(32'hbb4d348b),
	.w4(32'h3b5c389d),
	.w5(32'h3b56e380),
	.w6(32'hbb7b11c4),
	.w7(32'h3bba115f),
	.w8(32'hbabf6010),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2165d6),
	.w1(32'hbc680d9d),
	.w2(32'hbc9c927f),
	.w3(32'hbb046235),
	.w4(32'hbb4b14f5),
	.w5(32'hbc75af6b),
	.w6(32'hba8dd411),
	.w7(32'h3a18eef2),
	.w8(32'hbc2f2939),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb90966),
	.w1(32'hbb08e636),
	.w2(32'hbbbfae66),
	.w3(32'h3b698143),
	.w4(32'h3b0df293),
	.w5(32'hbb983c12),
	.w6(32'h3aa4d0e1),
	.w7(32'h39ec172e),
	.w8(32'hbc03de1d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9996b2),
	.w1(32'hb73be2e7),
	.w2(32'hbb836619),
	.w3(32'h392539e1),
	.w4(32'hbb7c92a3),
	.w5(32'hbbaeb5ff),
	.w6(32'hbab238fe),
	.w7(32'hba26b438),
	.w8(32'h3a147f5c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a932f25),
	.w1(32'h3b4512ea),
	.w2(32'h3b951972),
	.w3(32'hbb3206dc),
	.w4(32'h3bb7e6de),
	.w5(32'h3a03dd53),
	.w6(32'hbb19432a),
	.w7(32'h3b51d8b7),
	.w8(32'h37877f0b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf8685),
	.w1(32'h38cb7241),
	.w2(32'hbb6c0d8f),
	.w3(32'h3c14cc09),
	.w4(32'h3b8734df),
	.w5(32'hbbbdf0c1),
	.w6(32'hbac70eac),
	.w7(32'h3b565588),
	.w8(32'hba700368),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac71b0d),
	.w1(32'h3b035afe),
	.w2(32'hba6b82e5),
	.w3(32'hba94812d),
	.w4(32'h3c0a127e),
	.w5(32'hb9cfa18c),
	.w6(32'h3bb991c3),
	.w7(32'h3baa68e0),
	.w8(32'h3902d26e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbae7e),
	.w1(32'h3b192573),
	.w2(32'h3c004285),
	.w3(32'h3a9219ea),
	.w4(32'hba1ec3e7),
	.w5(32'h381e77c7),
	.w6(32'hb7d5461a),
	.w7(32'hbabd2c27),
	.w8(32'h3b17e687),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7575d3),
	.w1(32'hbbf6e618),
	.w2(32'hbc28b805),
	.w3(32'h3b9f61de),
	.w4(32'hbbaec4fc),
	.w5(32'hbc3d6062),
	.w6(32'hbbbfb4aa),
	.w7(32'hbb661ee7),
	.w8(32'hbb1925e9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6da208),
	.w1(32'h3c748beb),
	.w2(32'h3ca6fedb),
	.w3(32'hbc3e42a7),
	.w4(32'h3bdb8fce),
	.w5(32'h3be568d4),
	.w6(32'h3c48f75d),
	.w7(32'h3bc54bf8),
	.w8(32'h3bbed75b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ce3dd),
	.w1(32'hbbb1b190),
	.w2(32'hbc17e993),
	.w3(32'h3c0b422e),
	.w4(32'hba42bb66),
	.w5(32'hbc5d0310),
	.w6(32'hbc187bd9),
	.w7(32'hbc429981),
	.w8(32'hbc33720a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ee14e),
	.w1(32'hbbf25089),
	.w2(32'hbbc7b330),
	.w3(32'h3ac1712c),
	.w4(32'hbba27bee),
	.w5(32'hbb3e86ba),
	.w6(32'hbb13e795),
	.w7(32'h3ab8e1b1),
	.w8(32'hbaf52b37),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56c0f),
	.w1(32'hba89dce0),
	.w2(32'hba1180fc),
	.w3(32'hbbac2daa),
	.w4(32'hbb404498),
	.w5(32'hba8d1ea1),
	.w6(32'hbabee6e2),
	.w7(32'h3943ea91),
	.w8(32'h3b6018e4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47e7ce),
	.w1(32'hbc0bbb33),
	.w2(32'hbc16ba73),
	.w3(32'hbbbeb0a0),
	.w4(32'h3af999d2),
	.w5(32'hb9dd9151),
	.w6(32'hbbdb98f8),
	.w7(32'hba8851a5),
	.w8(32'hb9173306),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb51a38),
	.w1(32'hbc1aec70),
	.w2(32'hbc1c0bcc),
	.w3(32'h3a2af7a8),
	.w4(32'hbb2a7a8b),
	.w5(32'hbbf21a52),
	.w6(32'h376fae74),
	.w7(32'h3c000d48),
	.w8(32'h3be566b5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a35ae),
	.w1(32'h3bcaf658),
	.w2(32'h3c0f4f7e),
	.w3(32'hbbb60428),
	.w4(32'hbac5b02f),
	.w5(32'h3bca6584),
	.w6(32'hbae1968b),
	.w7(32'hbb88a2f8),
	.w8(32'hbafa285c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c021d72),
	.w1(32'hba3da664),
	.w2(32'hba83d8df),
	.w3(32'h3bce2d74),
	.w4(32'hbae49e83),
	.w5(32'h3b92bf80),
	.w6(32'hba8111d1),
	.w7(32'h3b6b0e0a),
	.w8(32'h3ae2256b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cf75d),
	.w1(32'hba0f483f),
	.w2(32'hbb556c7d),
	.w3(32'hbba16b1e),
	.w4(32'h3b5d4603),
	.w5(32'h3b3464d3),
	.w6(32'hbb44e0a5),
	.w7(32'hb9a0f0eb),
	.w8(32'h3b519d87),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba760316),
	.w1(32'hbbf84c5b),
	.w2(32'hbc357e43),
	.w3(32'h3bb4ecdd),
	.w4(32'hbba71596),
	.w5(32'hbc3a9024),
	.w6(32'hb8f63acf),
	.w7(32'hbaf3a288),
	.w8(32'hb93f13ed),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9cfd9),
	.w1(32'h3bcedcb2),
	.w2(32'h3c1e581d),
	.w3(32'hbab1a120),
	.w4(32'h3ace5f06),
	.w5(32'h3b6bdb67),
	.w6(32'h3ba2c83f),
	.w7(32'h3ba98846),
	.w8(32'h3b5380f9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f1672),
	.w1(32'h3b019ad0),
	.w2(32'h3c25e1a7),
	.w3(32'h3a41b141),
	.w4(32'h3b4ccc94),
	.w5(32'h3c5cf185),
	.w6(32'hbb2a3a9d),
	.w7(32'h3b672943),
	.w8(32'h3b9ccb0e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4ba71),
	.w1(32'hb9affbf5),
	.w2(32'h3ae1e7cc),
	.w3(32'h3c1b41f2),
	.w4(32'h3be9529c),
	.w5(32'hbb89916f),
	.w6(32'h3baff715),
	.w7(32'hba1d56f8),
	.w8(32'hb8834398),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12d579),
	.w1(32'hb9a79816),
	.w2(32'h397ab056),
	.w3(32'h3a415a57),
	.w4(32'hbb2c5464),
	.w5(32'hbb18b49f),
	.w6(32'h3b46f3b7),
	.w7(32'h3b610110),
	.w8(32'h3b61fb4c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb082b2f),
	.w1(32'hbb125355),
	.w2(32'hba125a9e),
	.w3(32'hbb9fe464),
	.w4(32'h3b174356),
	.w5(32'h3b638216),
	.w6(32'hb9b3001e),
	.w7(32'h3b8c9d04),
	.w8(32'h3824736f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a265175),
	.w1(32'hbc022fb5),
	.w2(32'hbb9523ee),
	.w3(32'h3b76e602),
	.w4(32'hbac075f7),
	.w5(32'hbb8e300c),
	.w6(32'hbb914aca),
	.w7(32'h3b852a5e),
	.w8(32'h3b03fd28),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2efa79),
	.w1(32'hba316838),
	.w2(32'h3b56cb97),
	.w3(32'hbb98d7f1),
	.w4(32'hbb1128cf),
	.w5(32'hba9af150),
	.w6(32'h39335ee3),
	.w7(32'hba35432d),
	.w8(32'hbab5821e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10a984),
	.w1(32'hbb1912f4),
	.w2(32'hbb504ab7),
	.w3(32'h3b1b163f),
	.w4(32'hba2bd242),
	.w5(32'hba723146),
	.w6(32'h3b8adfa2),
	.w7(32'hba20762b),
	.w8(32'h3adf9450),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96d0cf),
	.w1(32'h3bf24f6b),
	.w2(32'h3ad56415),
	.w3(32'h3bb31dd4),
	.w4(32'h3c386503),
	.w5(32'h3c156b42),
	.w6(32'h3bf5a88b),
	.w7(32'h3c15827c),
	.w8(32'h3ac94cbd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b1327),
	.w1(32'hba5545da),
	.w2(32'hbbd69c9d),
	.w3(32'h3c3908bf),
	.w4(32'hbb1cd91e),
	.w5(32'hbbe5abee),
	.w6(32'hba1a2386),
	.w7(32'hbba8c6ed),
	.w8(32'hbb11442b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82aa0d),
	.w1(32'hbb3610f4),
	.w2(32'hba94a911),
	.w3(32'hbba1a3b0),
	.w4(32'hbb82e30f),
	.w5(32'hbb8a17f9),
	.w6(32'h3903f370),
	.w7(32'h3b82c7e9),
	.w8(32'h3b7a4d12),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f07474),
	.w1(32'hba8f24e3),
	.w2(32'hbbe13459),
	.w3(32'h3a496df3),
	.w4(32'hbc077b77),
	.w5(32'hbc06b62a),
	.w6(32'h3ab697f9),
	.w7(32'hbb204d49),
	.w8(32'hbbd3708a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bb796),
	.w1(32'hbbff6ae6),
	.w2(32'hbc583255),
	.w3(32'hbbebade0),
	.w4(32'hbc05eb2c),
	.w5(32'hbc955ed9),
	.w6(32'hbbf978c4),
	.w7(32'hbbaac76d),
	.w8(32'hbc46b29a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcff43),
	.w1(32'hbb560438),
	.w2(32'hbbca05c1),
	.w3(32'hbc3acbd6),
	.w4(32'hbbc7e9e3),
	.w5(32'hbb3e5764),
	.w6(32'hbb80ead7),
	.w7(32'hbb68015a),
	.w8(32'hbb8759a9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc350a66),
	.w1(32'hbb2f773c),
	.w2(32'h3a3b2ea7),
	.w3(32'hbc37f800),
	.w4(32'h3ac82c30),
	.w5(32'h3bacc951),
	.w6(32'hbaf51eab),
	.w7(32'h3b6b090c),
	.w8(32'h3b62bab7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95487c),
	.w1(32'hbc0ddef2),
	.w2(32'hbc82991b),
	.w3(32'h3b1c8d08),
	.w4(32'h3aec3274),
	.w5(32'hbc304fda),
	.w6(32'hba397fa6),
	.w7(32'hbb42916f),
	.w8(32'hbc6cda2e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc6e51),
	.w1(32'hbb616d16),
	.w2(32'hbbd2ea05),
	.w3(32'h3b7d73d2),
	.w4(32'hbac98b25),
	.w5(32'hbbbb02cb),
	.w6(32'h3b0ed4d9),
	.w7(32'h3ac0f22b),
	.w8(32'h39d8993d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a0f61),
	.w1(32'hbb93f0ec),
	.w2(32'hbb979b19),
	.w3(32'h39a39b00),
	.w4(32'hbb2203f2),
	.w5(32'hbb9e3d28),
	.w6(32'hbb560cdc),
	.w7(32'hbbe9e613),
	.w8(32'hbabac2f3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64f123),
	.w1(32'hbb247429),
	.w2(32'h3b123443),
	.w3(32'h3a949bb4),
	.w4(32'h3b1541a3),
	.w5(32'h3b0ca8bf),
	.w6(32'h3b137d5b),
	.w7(32'hba37f4ee),
	.w8(32'h3c15387a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947b5c3),
	.w1(32'hbae9048a),
	.w2(32'hb98f45ba),
	.w3(32'h394130d1),
	.w4(32'hba2a616c),
	.w5(32'h3ac8e4b8),
	.w6(32'h3aa0a427),
	.w7(32'hbb9b9586),
	.w8(32'hba984a5a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb11012),
	.w1(32'hbafa1ed7),
	.w2(32'hbbffe2c0),
	.w3(32'hbb22b9bb),
	.w4(32'hbbd23c4f),
	.w5(32'h3ab0145b),
	.w6(32'hbb857afe),
	.w7(32'hb99f569a),
	.w8(32'hbb76d25c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc175a57),
	.w1(32'hbb473269),
	.w2(32'hba971e08),
	.w3(32'hbb6dd5c9),
	.w4(32'hbb55e89d),
	.w5(32'hbaff285e),
	.w6(32'h39435ea5),
	.w7(32'h399eab11),
	.w8(32'hb99fbb4b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b091d),
	.w1(32'hbb1641b5),
	.w2(32'hbb64036a),
	.w3(32'hba4901af),
	.w4(32'hbb2a12eb),
	.w5(32'hbb509a1f),
	.w6(32'hba424810),
	.w7(32'h397f2fc2),
	.w8(32'hb9975c24),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0718b7),
	.w1(32'h3b2f4b0d),
	.w2(32'h3892b3e1),
	.w3(32'hbaf1652b),
	.w4(32'hba23bc23),
	.w5(32'hbafd7ba4),
	.w6(32'hbb87b040),
	.w7(32'h3b0b8970),
	.w8(32'hbb965ad5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc6b9b),
	.w1(32'h3c04dbab),
	.w2(32'h3c8bd919),
	.w3(32'h3b0d7508),
	.w4(32'hbb990263),
	.w5(32'h394e4e98),
	.w6(32'h3a3bec71),
	.w7(32'h38dd19b1),
	.w8(32'hb938d496),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c319921),
	.w1(32'h3c327b59),
	.w2(32'h3c9fe279),
	.w3(32'h3b48a2b7),
	.w4(32'h3b160621),
	.w5(32'h3b8d56b2),
	.w6(32'h3c1f96ed),
	.w7(32'h3c3ac7c6),
	.w8(32'h3c32d92b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c842d60),
	.w1(32'h3a909bcd),
	.w2(32'h3b253040),
	.w3(32'h3bf474fd),
	.w4(32'h3bcbff60),
	.w5(32'h3be3258f),
	.w6(32'h3ba594cc),
	.w7(32'h3c104906),
	.w8(32'h3b795c6a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8d185),
	.w1(32'hbabfda76),
	.w2(32'hba97e214),
	.w3(32'h3bbb9db6),
	.w4(32'hba1a810d),
	.w5(32'hb959b073),
	.w6(32'hbb6bc645),
	.w7(32'h3a173379),
	.w8(32'hbae20c41),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d11e2),
	.w1(32'hbb8114ce),
	.w2(32'hb9837d8b),
	.w3(32'h3aad8b98),
	.w4(32'hbb41f841),
	.w5(32'hba3ad201),
	.w6(32'h390185da),
	.w7(32'h3b8e7399),
	.w8(32'h3babaab5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e56ac),
	.w1(32'h3b81d401),
	.w2(32'hba805c66),
	.w3(32'hbafa486a),
	.w4(32'h3b1ca5ad),
	.w5(32'hbb399b52),
	.w6(32'h3bc94678),
	.w7(32'h3b571001),
	.w8(32'hbb8bf2e8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93b73c),
	.w1(32'h3bad6521),
	.w2(32'h3bf77869),
	.w3(32'hbb248feb),
	.w4(32'h3bcbf66b),
	.w5(32'h3c06af48),
	.w6(32'hba5cd565),
	.w7(32'hbbc992ea),
	.w8(32'hbb72fe22),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09f8f0),
	.w1(32'hbb933e52),
	.w2(32'hbc0a1226),
	.w3(32'h3bfcefe3),
	.w4(32'hbb86038b),
	.w5(32'hbbf182f8),
	.w6(32'hbb7006e8),
	.w7(32'h3a3d4a8c),
	.w8(32'h3af8b4f9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed296a),
	.w1(32'hbbe3c185),
	.w2(32'hbb8e9c11),
	.w3(32'hbbe98116),
	.w4(32'hbb401350),
	.w5(32'hbbd8612a),
	.w6(32'hbc27bd3e),
	.w7(32'hbba22a0a),
	.w8(32'hbb542cb6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27782a),
	.w1(32'hbbedb30d),
	.w2(32'hbbc1a69b),
	.w3(32'hbab2272e),
	.w4(32'hbb57d4f0),
	.w5(32'hbb0a6304),
	.w6(32'h3b46a934),
	.w7(32'hbb24cb88),
	.w8(32'h3b4571a2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5efa),
	.w1(32'hbbf6f75c),
	.w2(32'hbb4a29a5),
	.w3(32'h3a5f095b),
	.w4(32'hbb16a03e),
	.w5(32'h3b3b49af),
	.w6(32'hbc435ad9),
	.w7(32'hbbcac740),
	.w8(32'hbb1a15d0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc63e82),
	.w1(32'hbc32a6a3),
	.w2(32'hbc466e3c),
	.w3(32'h3a83c262),
	.w4(32'hbc064c9a),
	.w5(32'hbbf5a91b),
	.w6(32'hbb28c2c2),
	.w7(32'hbb5f5b25),
	.w8(32'h38abf1c0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf2ae0),
	.w1(32'hbbe30209),
	.w2(32'hbc111a54),
	.w3(32'hb984df5e),
	.w4(32'hbbb68648),
	.w5(32'hbbfa9afb),
	.w6(32'hbafbb579),
	.w7(32'hbb673e62),
	.w8(32'h3a101857),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e0a3f),
	.w1(32'hbb509987),
	.w2(32'hbb43b626),
	.w3(32'hbc10a251),
	.w4(32'h3bacaf1d),
	.w5(32'h3b743118),
	.w6(32'hbbd032ca),
	.w7(32'hbb89d288),
	.w8(32'hbb10ca03),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb72a0),
	.w1(32'hba8cf60c),
	.w2(32'h3acfeecb),
	.w3(32'hb9febe5a),
	.w4(32'hbbae92dd),
	.w5(32'hbbbca1b3),
	.w6(32'hba00a882),
	.w7(32'h3a3f9aaa),
	.w8(32'h3a13bd3c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedbc72),
	.w1(32'hbb75b644),
	.w2(32'hbbb9794e),
	.w3(32'hbbac1062),
	.w4(32'hba2094a2),
	.w5(32'hbb2a0991),
	.w6(32'hbaf24b5c),
	.w7(32'hbb91ea3b),
	.w8(32'hbb463cda),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ceaee),
	.w1(32'hba56ec72),
	.w2(32'hba752995),
	.w3(32'h3b8f0768),
	.w4(32'h3a244050),
	.w5(32'hbafc10bd),
	.w6(32'h3a392f17),
	.w7(32'hba4c3f0b),
	.w8(32'hbb240fbc),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb965fcd),
	.w1(32'hbb015477),
	.w2(32'hbb07727a),
	.w3(32'h39175981),
	.w4(32'hba568a22),
	.w5(32'hbb817ab0),
	.w6(32'h3b7c3f67),
	.w7(32'h3af3951b),
	.w8(32'hbb03b334),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0191dd),
	.w1(32'hbbbd6121),
	.w2(32'hbbd954fb),
	.w3(32'h3a599cb4),
	.w4(32'hba4cdba0),
	.w5(32'hbaccf7a8),
	.w6(32'hba515aba),
	.w7(32'hbae925a8),
	.w8(32'hbb8651fa),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef9448),
	.w1(32'h3a6a7b73),
	.w2(32'h3b8f1750),
	.w3(32'h3a135d4e),
	.w4(32'hbb46280a),
	.w5(32'hb9defbfe),
	.w6(32'hbb0734c1),
	.w7(32'hbb378315),
	.w8(32'h3b1df48c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395499dd),
	.w1(32'h3b2c2363),
	.w2(32'h3af2deaf),
	.w3(32'h3b01ee89),
	.w4(32'hbbb7f28b),
	.w5(32'hbb47a0f9),
	.w6(32'h3b24c103),
	.w7(32'hbaa3d37d),
	.w8(32'h3b8bc70a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28c41d),
	.w1(32'hbc48b6a6),
	.w2(32'hbc236995),
	.w3(32'hbb59f7a8),
	.w4(32'hbbf3694d),
	.w5(32'hbbcd4d9e),
	.w6(32'hbbc1a57a),
	.w7(32'hbba51eb9),
	.w8(32'hbbb69549),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97ad5b),
	.w1(32'h3b06c553),
	.w2(32'hbb3dfe8c),
	.w3(32'hbb122577),
	.w4(32'h3a52c93a),
	.w5(32'h3ac813b7),
	.w6(32'h3b13b059),
	.w7(32'hbb71606e),
	.w8(32'h3b1a55c0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2b4d1),
	.w1(32'hbc35cf10),
	.w2(32'hbbafefac),
	.w3(32'hba4bbf8d),
	.w4(32'hbb3f9839),
	.w5(32'h3913bba7),
	.w6(32'hbbfc1323),
	.w7(32'hbbd75557),
	.w8(32'hbbddd286),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb7dbb),
	.w1(32'hba868154),
	.w2(32'hbb9797f0),
	.w3(32'h3a856763),
	.w4(32'hba5f9cd8),
	.w5(32'hb9f5a3a0),
	.w6(32'h3b809f3d),
	.w7(32'h3be1a771),
	.w8(32'h3ab9106d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad299b),
	.w1(32'hbaa32ae9),
	.w2(32'hbb966329),
	.w3(32'h3bbb2ca1),
	.w4(32'hbb334960),
	.w5(32'hbc22807d),
	.w6(32'hb99caa2b),
	.w7(32'hbaa35598),
	.w8(32'hbaabca30),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba849fd2),
	.w1(32'hbb812ca1),
	.w2(32'hbba8d784),
	.w3(32'hbc9253d0),
	.w4(32'h39c41a50),
	.w5(32'h399138d4),
	.w6(32'hbbce83c4),
	.w7(32'hbbeaa911),
	.w8(32'hbbb1491d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb65bec),
	.w1(32'h3c1f4e73),
	.w2(32'h3c6f0ddb),
	.w3(32'h39d8a0c6),
	.w4(32'h3af5eb04),
	.w5(32'h3b81fc7e),
	.w6(32'h3c04cf50),
	.w7(32'h3c1962df),
	.w8(32'h3c22c165),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c770c61),
	.w1(32'hbb71860d),
	.w2(32'hbbb0893e),
	.w3(32'h3bd7f3b5),
	.w4(32'h3afcc2b4),
	.w5(32'h394217b4),
	.w6(32'hbb5e469f),
	.w7(32'hbb4a5fb3),
	.w8(32'hbaf958cf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb43803),
	.w1(32'h3b7b1072),
	.w2(32'hb9de03d4),
	.w3(32'h3adfa3af),
	.w4(32'hb96ad9f5),
	.w5(32'h3baa7538),
	.w6(32'h3bd0cfdd),
	.w7(32'h3b8eebb9),
	.w8(32'hb8ceb3e4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a0c4a),
	.w1(32'hbbbf95c4),
	.w2(32'hbbe27197),
	.w3(32'h3b5e1022),
	.w4(32'hbb943ae9),
	.w5(32'hbba2688e),
	.w6(32'h3a46e228),
	.w7(32'h3b1d2fc9),
	.w8(32'h3b6c56f3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5e06e),
	.w1(32'hbb7c3d01),
	.w2(32'hba8df235),
	.w3(32'hbb993fca),
	.w4(32'hbaa09cdf),
	.w5(32'hbb3f17a7),
	.w6(32'h3ad9dc3d),
	.w7(32'h3acb3f15),
	.w8(32'h3a66aed0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f6feac),
	.w1(32'h3a996769),
	.w2(32'hb7d873e9),
	.w3(32'hbbf31cf3),
	.w4(32'h3b795ab4),
	.w5(32'h3ae4e922),
	.w6(32'hba38a81b),
	.w7(32'h3a28d67e),
	.w8(32'h3a81f80a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b3fd0),
	.w1(32'hbb54be4c),
	.w2(32'hbbb1a0cf),
	.w3(32'hba7019a8),
	.w4(32'hbac13f07),
	.w5(32'hbb8ee380),
	.w6(32'hbb380d19),
	.w7(32'h39da45ad),
	.w8(32'hb898758f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d3aca),
	.w1(32'hbbced9a7),
	.w2(32'hbb15dbfc),
	.w3(32'hbbb52014),
	.w4(32'hbb53565b),
	.w5(32'hbb16f5df),
	.w6(32'hba5554b3),
	.w7(32'hbb6003a9),
	.w8(32'hba934249),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97cd85),
	.w1(32'hbc055c17),
	.w2(32'hbc150146),
	.w3(32'hb9cf290f),
	.w4(32'hbb70f8b1),
	.w5(32'hbb85edb8),
	.w6(32'hbbacc6a0),
	.w7(32'hbba81b3a),
	.w8(32'hbc1077ee),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4672d7),
	.w1(32'hbbff432d),
	.w2(32'hbc37a3a0),
	.w3(32'hbb819a33),
	.w4(32'hbb1788a9),
	.w5(32'hbbc02ca6),
	.w6(32'hbb394613),
	.w7(32'hba944523),
	.w8(32'hbc2e966c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b355f27),
	.w1(32'h3ba7ea3b),
	.w2(32'h3b6756df),
	.w3(32'h3a9fd1d2),
	.w4(32'h3ba1bd39),
	.w5(32'h3c1d97c1),
	.w6(32'h3b633f65),
	.w7(32'h3a7f1fdc),
	.w8(32'h3b709c1f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7ab96),
	.w1(32'h39b4bf6c),
	.w2(32'h3a8ab0cb),
	.w3(32'h3bfc68fa),
	.w4(32'h3b37e5b7),
	.w5(32'h3ae427ba),
	.w6(32'hbbcd4d3e),
	.w7(32'h3ab55189),
	.w8(32'hbad611ea),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbf214),
	.w1(32'h3bf87abd),
	.w2(32'h3c303519),
	.w3(32'h3ae41944),
	.w4(32'hbb00857c),
	.w5(32'h3bc4c14e),
	.w6(32'h3bc64e34),
	.w7(32'h3c271c35),
	.w8(32'h3bd320d4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b40f8),
	.w1(32'hba2cadb6),
	.w2(32'hbaa4f3c1),
	.w3(32'h3a8a6a34),
	.w4(32'h3a437936),
	.w5(32'h3af78901),
	.w6(32'hbc0b7590),
	.w7(32'hbc30d314),
	.w8(32'hbc0c3ae4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6701bd),
	.w1(32'hbb15a97d),
	.w2(32'hbb30e655),
	.w3(32'hbb1a4164),
	.w4(32'hb982cfbd),
	.w5(32'h3c179d16),
	.w6(32'hbc1510a3),
	.w7(32'hbc22681e),
	.w8(32'hbbb073a9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f3517),
	.w1(32'hbc16a55b),
	.w2(32'hbc1ddb16),
	.w3(32'h3b997287),
	.w4(32'hbb9e2115),
	.w5(32'hbc2091ed),
	.w6(32'hbacb16e7),
	.w7(32'hba4b4fb1),
	.w8(32'hb8d628fb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5580),
	.w1(32'hbbcdbbe8),
	.w2(32'hbbd44521),
	.w3(32'hbb68b158),
	.w4(32'hbbf06b45),
	.w5(32'hbb848b0f),
	.w6(32'hbac6e4f6),
	.w7(32'hbb455409),
	.w8(32'hbc1b32be),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba214917),
	.w1(32'hbc2f65cd),
	.w2(32'hbc24e7dd),
	.w3(32'hbb7e8686),
	.w4(32'hbbdb2ed3),
	.w5(32'hbbe6839c),
	.w6(32'hbc07f4e8),
	.w7(32'hbc1fa90a),
	.w8(32'hbba4aa64),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91c551),
	.w1(32'hbb500e81),
	.w2(32'hbbfcfa98),
	.w3(32'h3adcea8c),
	.w4(32'hbb1df4c1),
	.w5(32'hbbfeb67c),
	.w6(32'h3b862c49),
	.w7(32'h3b068072),
	.w8(32'h39876563),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a351b48),
	.w1(32'h3aade919),
	.w2(32'hba35dcb1),
	.w3(32'hbab1ed9d),
	.w4(32'h3bad62d9),
	.w5(32'h3b2086d5),
	.w6(32'hbc07bb24),
	.w7(32'hbbcd2e39),
	.w8(32'hbb91f2b6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd88450),
	.w1(32'h3adc4b65),
	.w2(32'h3bfd82cd),
	.w3(32'h39f01e4c),
	.w4(32'hbb600090),
	.w5(32'hbac04d1b),
	.w6(32'h3b9ac0b2),
	.w7(32'h3bf61704),
	.w8(32'h3c0a819f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe823b),
	.w1(32'hbb1da0b7),
	.w2(32'hba7d2bce),
	.w3(32'hba61cd35),
	.w4(32'hbbc75d0c),
	.w5(32'hbbb511ed),
	.w6(32'hbb49d4a7),
	.w7(32'h3ae656ff),
	.w8(32'h3aada74c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69bb2e),
	.w1(32'hbb23bde6),
	.w2(32'hba8e8ca6),
	.w3(32'hbbffaf5d),
	.w4(32'hbb48f004),
	.w5(32'hbb41d46f),
	.w6(32'hbb161f71),
	.w7(32'h3afdb553),
	.w8(32'h3b3cbdf5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02fe49),
	.w1(32'hbbdcb74d),
	.w2(32'hbae1118c),
	.w3(32'hbb99ddd0),
	.w4(32'hbbcf4fbd),
	.w5(32'hbb8b2979),
	.w6(32'h3a40bb64),
	.w7(32'hb9058e0d),
	.w8(32'h3b7549e7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1a0c8),
	.w1(32'hbb7028a4),
	.w2(32'hbba3f784),
	.w3(32'hbbd34ec4),
	.w4(32'hbb3075b3),
	.w5(32'hbbb4ba18),
	.w6(32'hbbc3c98b),
	.w7(32'h3aadffe9),
	.w8(32'h3ada3a5f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb294ac1),
	.w1(32'h3ad18b42),
	.w2(32'hbb593493),
	.w3(32'hbbba75b2),
	.w4(32'hbbbe70c5),
	.w5(32'hbc00dcb0),
	.w6(32'hbbe4490c),
	.w7(32'hbbf6e65b),
	.w8(32'hbbb6221d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cede6),
	.w1(32'hbc73045c),
	.w2(32'hbc586b8d),
	.w3(32'hbbf6cd1c),
	.w4(32'hbc159b12),
	.w5(32'hbc587125),
	.w6(32'hbbde7c76),
	.w7(32'hbc47efce),
	.w8(32'hbc1dcd4d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ae69c),
	.w1(32'hbbe543e6),
	.w2(32'hbbb7b903),
	.w3(32'hbc57c22e),
	.w4(32'h3b22ac70),
	.w5(32'hb9c02a80),
	.w6(32'hbbd279c4),
	.w7(32'hbbad90a6),
	.w8(32'hbbc47a89),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f0b74),
	.w1(32'hbb8ddb02),
	.w2(32'hbb2f85f7),
	.w3(32'hbb2cfb7a),
	.w4(32'hbb90b41d),
	.w5(32'hbb5edba3),
	.w6(32'hbb7969ea),
	.w7(32'hba239b01),
	.w8(32'hb9bfb2a6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e0376),
	.w1(32'h3b2c7b26),
	.w2(32'h3b9d1f7f),
	.w3(32'hbb919a2a),
	.w4(32'hbb9c4890),
	.w5(32'hbbcc4289),
	.w6(32'hba5d80c5),
	.w7(32'h3b8aa8db),
	.w8(32'h3b91a8cb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d46da),
	.w1(32'hbb64a91f),
	.w2(32'hbbb5299d),
	.w3(32'hbb224b34),
	.w4(32'hbb35a11e),
	.w5(32'hbb92ef92),
	.w6(32'hbaef4a06),
	.w7(32'hbb8c9489),
	.w8(32'hbb480c08),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ceb3f),
	.w1(32'hbb97803c),
	.w2(32'h3b31b066),
	.w3(32'hbb0ffc73),
	.w4(32'hbbcc5bf2),
	.w5(32'hbb57779f),
	.w6(32'h3bf99f8a),
	.w7(32'hb961d576),
	.w8(32'h3bccbb9e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3915a),
	.w1(32'h3b705a34),
	.w2(32'h3b9f1d87),
	.w3(32'h3b9403c4),
	.w4(32'h3a4d10ce),
	.w5(32'hba252f48),
	.w6(32'h3af7c80d),
	.w7(32'h3b1bd4dc),
	.w8(32'h3acc76ba),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1a10d),
	.w1(32'hbbe0c1ec),
	.w2(32'hbaee084f),
	.w3(32'hbb0f667d),
	.w4(32'hbaa597d2),
	.w5(32'hbb705bde),
	.w6(32'hbbb671ef),
	.w7(32'h39f88889),
	.w8(32'hbb13107a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961d960),
	.w1(32'hb89ab01c),
	.w2(32'hbac5715f),
	.w3(32'h3a788909),
	.w4(32'h3ace7a27),
	.w5(32'hbaf2e9c3),
	.w6(32'h3adebda4),
	.w7(32'h3c2a7140),
	.w8(32'h3b95fc8c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd3f3d),
	.w1(32'hbb1b8297),
	.w2(32'hbbbb075a),
	.w3(32'h3b97be56),
	.w4(32'hbb566d22),
	.w5(32'hbbbf9a04),
	.w6(32'hbb6aaaa4),
	.w7(32'hbb310452),
	.w8(32'hbb05a8f7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb2da6),
	.w1(32'hbbd716fd),
	.w2(32'hbc1cbf93),
	.w3(32'hbbf7abf4),
	.w4(32'hbb0374eb),
	.w5(32'hbbf44b27),
	.w6(32'hbbb9b7bc),
	.w7(32'hbbc7917b),
	.w8(32'hbbfd3a2c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5353f),
	.w1(32'hb93618fe),
	.w2(32'hbb2a0967),
	.w3(32'hbb850571),
	.w4(32'hbbc03323),
	.w5(32'hbbab897e),
	.w6(32'hbbd4811b),
	.w7(32'hbbbf57c6),
	.w8(32'hbb685be0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5b71),
	.w1(32'hbb48c656),
	.w2(32'hbbdc80de),
	.w3(32'hbbda3548),
	.w4(32'hbc01f139),
	.w5(32'hbbd2c730),
	.w6(32'hbbed169e),
	.w7(32'hbbfbe74e),
	.w8(32'hbc1ab790),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d172f),
	.w1(32'hba7efb2c),
	.w2(32'hbadacef8),
	.w3(32'hbb0a9ed1),
	.w4(32'hb9d3108e),
	.w5(32'hbabb8361),
	.w6(32'hb79aa16d),
	.w7(32'hba56d64d),
	.w8(32'h397c17d2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa06bb4),
	.w1(32'h38cd0f1b),
	.w2(32'hb930a26d),
	.w3(32'h3a1c567b),
	.w4(32'h3b00bd71),
	.w5(32'hbaa4cfce),
	.w6(32'h3ad43fee),
	.w7(32'hbb312b49),
	.w8(32'h3b140ac6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule