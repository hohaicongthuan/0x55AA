module layer_10_featuremap_227(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedb61f),
	.w1(32'h3aea2e99),
	.w2(32'hba6d5f33),
	.w3(32'hbb56f576),
	.w4(32'hbb12023b),
	.w5(32'h3c35f5d8),
	.w6(32'h3b6606b9),
	.w7(32'hbbfe186e),
	.w8(32'hbc19ca77),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6d48b8),
	.w1(32'hbc28c67b),
	.w2(32'h3b5f86f2),
	.w3(32'hb9bc326f),
	.w4(32'hbb4ef416),
	.w5(32'hbb385a06),
	.w6(32'hbb6152e4),
	.w7(32'h3b69db7b),
	.w8(32'h3b8761c1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d6232d),
	.w1(32'h3a8477d4),
	.w2(32'hbc25247c),
	.w3(32'hbb067f29),
	.w4(32'hbc1b50c8),
	.w5(32'h3a92f91b),
	.w6(32'hba9ac7cf),
	.w7(32'h3b3fcde6),
	.w8(32'hbc038cae),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9217af),
	.w1(32'hba91bf65),
	.w2(32'hbb9f77a9),
	.w3(32'h3b85b3bc),
	.w4(32'hbc444a09),
	.w5(32'hb727efe8),
	.w6(32'hbb102e51),
	.w7(32'hb9617723),
	.w8(32'hba147137),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cff1b),
	.w1(32'h3bfcac32),
	.w2(32'h3aca2ba8),
	.w3(32'hbba70ac0),
	.w4(32'hbb7544ba),
	.w5(32'h387b8d19),
	.w6(32'hbba4ce74),
	.w7(32'hba7bf756),
	.w8(32'hbbf36fd9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b137b50),
	.w1(32'hbba091a3),
	.w2(32'hbafa84f2),
	.w3(32'h3abec48e),
	.w4(32'hb7b9af6f),
	.w5(32'hbc0c4763),
	.w6(32'hbc040696),
	.w7(32'hba2664da),
	.w8(32'hbc1cee53),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec7916),
	.w1(32'hbb23104d),
	.w2(32'h3c024ee0),
	.w3(32'hbc02025c),
	.w4(32'hbcc85525),
	.w5(32'h3cad5d76),
	.w6(32'h3bb2357b),
	.w7(32'hbbfaec0d),
	.w8(32'h3c5e9b72),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a182),
	.w1(32'h3a1b1864),
	.w2(32'hbae3e4da),
	.w3(32'h3bc00b47),
	.w4(32'h3b969f57),
	.w5(32'hba0968be),
	.w6(32'hbc73705e),
	.w7(32'h3b473e33),
	.w8(32'h3c574513),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0ab18),
	.w1(32'h3c970e16),
	.w2(32'h3d1491d3),
	.w3(32'hbb83751e),
	.w4(32'hbb1932ee),
	.w5(32'h3ad9882b),
	.w6(32'hbc1dd4be),
	.w7(32'hbacab5b2),
	.w8(32'h3b2489ee),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a5b21),
	.w1(32'h3b2d0d0b),
	.w2(32'hbc5578d9),
	.w3(32'h3c02730a),
	.w4(32'hbad8fce0),
	.w5(32'h3ba10b30),
	.w6(32'hbbb31b01),
	.w7(32'h3ac310d4),
	.w8(32'hbb595d73),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae17d3),
	.w1(32'hbb9450d4),
	.w2(32'h3a500f2d),
	.w3(32'hbc19f733),
	.w4(32'h3b7b34bf),
	.w5(32'h3c31cb20),
	.w6(32'h39f6cba4),
	.w7(32'hbacf7bfe),
	.w8(32'h3b13101c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b803a45),
	.w1(32'h3b2d6707),
	.w2(32'hbc3a4e1c),
	.w3(32'h3b33a5d6),
	.w4(32'h3bf08252),
	.w5(32'hbbd08d21),
	.w6(32'h3b9941b9),
	.w7(32'h399bb74f),
	.w8(32'h3b8fc595),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc36a3),
	.w1(32'hbb5cd87c),
	.w2(32'h3bb857e9),
	.w3(32'h3ba9deaf),
	.w4(32'hbb80f77d),
	.w5(32'h3b1a88c7),
	.w6(32'h3c0859b7),
	.w7(32'h3b40a179),
	.w8(32'hbc354e62),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1074b),
	.w1(32'hbbfe2afa),
	.w2(32'h3c2c2daf),
	.w3(32'hbc0de641),
	.w4(32'hbd12a29a),
	.w5(32'h3be683a3),
	.w6(32'h3cda1633),
	.w7(32'hbb4dc6ea),
	.w8(32'h3ba5bc4c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc790b2d),
	.w1(32'h3c003f22),
	.w2(32'h3b93c7d1),
	.w3(32'h3b40fd83),
	.w4(32'hbb914693),
	.w5(32'h3b1f7446),
	.w6(32'hbbcf0d6e),
	.w7(32'hbb518eb4),
	.w8(32'h3a479dc9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3fa3d),
	.w1(32'h3a968532),
	.w2(32'h3bd617b0),
	.w3(32'h3a8585e1),
	.w4(32'hbb250d7a),
	.w5(32'hba8c2d25),
	.w6(32'hbb0f4d92),
	.w7(32'hbb384dec),
	.w8(32'h3cd4d398),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c359d),
	.w1(32'h3b7d11b2),
	.w2(32'h39a79f25),
	.w3(32'h3a9319f9),
	.w4(32'h37f61dc3),
	.w5(32'hbb3ccb8d),
	.w6(32'h3a8e32ba),
	.w7(32'hbb3757bf),
	.w8(32'h3ab4865c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc071cc),
	.w1(32'hbd4d5e48),
	.w2(32'hbbdc6943),
	.w3(32'h3c07645c),
	.w4(32'hbbdc5a98),
	.w5(32'h3a9005d6),
	.w6(32'hbc1932ad),
	.w7(32'hbb3ed793),
	.w8(32'hbb8754de),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28ad9c),
	.w1(32'hbba0eed3),
	.w2(32'h3bc97fe6),
	.w3(32'h3b944ed8),
	.w4(32'hbb516912),
	.w5(32'hbc22e4fe),
	.w6(32'h3b2c2e05),
	.w7(32'h3a9e8ab4),
	.w8(32'h3a95b5e5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd03357),
	.w1(32'h3a9c0023),
	.w2(32'hbc04dd8a),
	.w3(32'hbb58eaa5),
	.w4(32'hbb2b5043),
	.w5(32'hbb2ccbcc),
	.w6(32'h3b435b32),
	.w7(32'hba88d453),
	.w8(32'h3bbd4585),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f6100),
	.w1(32'hba9b87d9),
	.w2(32'hbcc9862f),
	.w3(32'hbb990602),
	.w4(32'h3ba14cd9),
	.w5(32'hb9a413c9),
	.w6(32'h3b36fca9),
	.w7(32'h3ac02c6d),
	.w8(32'hbbb20191),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bf1ee),
	.w1(32'h3bd1db69),
	.w2(32'hbab92ba2),
	.w3(32'hbb24effe),
	.w4(32'hbb58f126),
	.w5(32'hb9b77761),
	.w6(32'hbc232c45),
	.w7(32'hb9b2cf67),
	.w8(32'hbaf3f881),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac404b),
	.w1(32'h3b2d852c),
	.w2(32'h3d0b689d),
	.w3(32'h3b9e416d),
	.w4(32'hbb778cc8),
	.w5(32'hbc95f56a),
	.w6(32'h3ba0610d),
	.w7(32'hbb8ad3fb),
	.w8(32'h3c49f4ad),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92aa1c),
	.w1(32'hba433e74),
	.w2(32'h3c032037),
	.w3(32'h3bbadb2c),
	.w4(32'h3b8a5b37),
	.w5(32'h3bc573a4),
	.w6(32'h3b27dfb9),
	.w7(32'hbc8f90ae),
	.w8(32'h3b720b3c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeda75),
	.w1(32'h3c183001),
	.w2(32'h3aa5fa44),
	.w3(32'h3b3db6ea),
	.w4(32'h3c9257ed),
	.w5(32'hb82b8ba0),
	.w6(32'hbad26fc2),
	.w7(32'hbaea9c30),
	.w8(32'hbc9d60a8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b274b99),
	.w1(32'hbb777503),
	.w2(32'h3c243cdf),
	.w3(32'hbb57bce8),
	.w4(32'hbc27599b),
	.w5(32'h3b8d6f13),
	.w6(32'h3ab01a60),
	.w7(32'hbb26bc0c),
	.w8(32'h3b8481d3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89abda),
	.w1(32'hbb9fc8a1),
	.w2(32'hbb933a98),
	.w3(32'h3aa3f6c9),
	.w4(32'h3a5345ca),
	.w5(32'hbab9bd0d),
	.w6(32'hbb0aa6bf),
	.w7(32'h3bb63115),
	.w8(32'h3bb945ef),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dcfd2),
	.w1(32'hbc1faffd),
	.w2(32'hbba045a8),
	.w3(32'hba718e3d),
	.w4(32'hbb86f446),
	.w5(32'hbb791058),
	.w6(32'hbadfe122),
	.w7(32'h3aa56540),
	.w8(32'hbb00637c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bb714),
	.w1(32'h3bbf5fa6),
	.w2(32'h3abbcda6),
	.w3(32'hbbb3377e),
	.w4(32'h3b283809),
	.w5(32'h3b9a3b2a),
	.w6(32'hbc8efe66),
	.w7(32'hbab46eec),
	.w8(32'h3c8282d6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24aced),
	.w1(32'h3b99d0a6),
	.w2(32'h38c1c3f5),
	.w3(32'h3c1f5b77),
	.w4(32'h3b606ecb),
	.w5(32'h3c6034e3),
	.w6(32'hbb8b3978),
	.w7(32'hba4b20a5),
	.w8(32'h3abab3a8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb056f74),
	.w1(32'hbbe53538),
	.w2(32'h3baedd88),
	.w3(32'h3af5f647),
	.w4(32'hba9865b5),
	.w5(32'h3b7dbed3),
	.w6(32'h3ade0fc4),
	.w7(32'hbad72958),
	.w8(32'h3994d3f7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb28790),
	.w1(32'hbc36e19f),
	.w2(32'hbc35dc6a),
	.w3(32'h3b07f865),
	.w4(32'hbc244600),
	.w5(32'h3cf8d498),
	.w6(32'hbacc51dc),
	.w7(32'h3c24b4d8),
	.w8(32'hbaa9c4fb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a12bc),
	.w1(32'hbc620f05),
	.w2(32'h3c261fcd),
	.w3(32'h3b808123),
	.w4(32'h3a09ea21),
	.w5(32'h3c3d9ed1),
	.w6(32'h3b93f839),
	.w7(32'h3bad878f),
	.w8(32'h3b5dc1bb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9bcb9),
	.w1(32'h3ca73643),
	.w2(32'h3b61cd37),
	.w3(32'hbc0ebf1a),
	.w4(32'h3c98bd01),
	.w5(32'h3b0971e6),
	.w6(32'hbaca22c8),
	.w7(32'h3bf53a6f),
	.w8(32'h3afb1f5b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb939cbc),
	.w1(32'hbc36efb6),
	.w2(32'hbb92ccbe),
	.w3(32'h3bf50d27),
	.w4(32'hba9536b9),
	.w5(32'hbc6bb9cd),
	.w6(32'h3cabbeec),
	.w7(32'h3af574c7),
	.w8(32'h3bc602d6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b999f4),
	.w1(32'hbbf9c4a2),
	.w2(32'h3c58ae54),
	.w3(32'hbb64fe60),
	.w4(32'h3992dbc2),
	.w5(32'h3c4fbeed),
	.w6(32'h3b87525f),
	.w7(32'hbb687e50),
	.w8(32'h3c85c113),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cbedd),
	.w1(32'h39f4c083),
	.w2(32'h3b9355e2),
	.w3(32'h3c366153),
	.w4(32'h3ac9efa3),
	.w5(32'hbba4f8e3),
	.w6(32'h3b035cd5),
	.w7(32'h3c26acec),
	.w8(32'hbc562810),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fc4e7),
	.w1(32'hbaca500d),
	.w2(32'h3d00aa30),
	.w3(32'hbc6787dc),
	.w4(32'hbc227fb2),
	.w5(32'hbb84b822),
	.w6(32'hbbfba3a5),
	.w7(32'h3b1122cf),
	.w8(32'h3d1ba047),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42daa8),
	.w1(32'hbc0373fc),
	.w2(32'h3b51fec6),
	.w3(32'hbcc9b652),
	.w4(32'hbb66e4fd),
	.w5(32'hbbeaa58d),
	.w6(32'hbc73714e),
	.w7(32'hbbbeeee2),
	.w8(32'hbb734e93),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb093ba3),
	.w1(32'h3c022033),
	.w2(32'h3acfef18),
	.w3(32'h3b27a21b),
	.w4(32'hbb8405ce),
	.w5(32'hbc18efb2),
	.w6(32'h3aa27197),
	.w7(32'h3c20c056),
	.w8(32'h3c04208c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39113e67),
	.w1(32'h3c41eed8),
	.w2(32'h3bd463d5),
	.w3(32'h3c28bb75),
	.w4(32'h3b0dc561),
	.w5(32'h3be6e7c1),
	.w6(32'h3abf430a),
	.w7(32'h3b0aa1b5),
	.w8(32'hbbb33466),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55b267),
	.w1(32'h3a0d5ff0),
	.w2(32'h3c49759d),
	.w3(32'hbb088110),
	.w4(32'hb91c63c3),
	.w5(32'h3c14ca6b),
	.w6(32'h3b88cc42),
	.w7(32'hbac694c4),
	.w8(32'h3c17559b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bbbaa),
	.w1(32'hbb3f4205),
	.w2(32'hbb9227a7),
	.w3(32'hbc2c5008),
	.w4(32'h3c80587f),
	.w5(32'h3bbd9f84),
	.w6(32'hbc2335df),
	.w7(32'hbb6f9be5),
	.w8(32'hbb185da4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e114d0),
	.w1(32'h3b6bc2e3),
	.w2(32'h3c8158cb),
	.w3(32'h3bef08b8),
	.w4(32'h3b8bd817),
	.w5(32'hb81b46f7),
	.w6(32'hba923ab5),
	.w7(32'hbbdf30a9),
	.w8(32'h3b02d759),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b616f6a),
	.w1(32'hb83a89ed),
	.w2(32'h39ada597),
	.w3(32'hbba2652f),
	.w4(32'hbc0f793d),
	.w5(32'hbb24c1ab),
	.w6(32'hbbe1633a),
	.w7(32'h3b835eb2),
	.w8(32'h3b83d02b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e7efc),
	.w1(32'hb9e199c3),
	.w2(32'h3d1fc1f5),
	.w3(32'h3bb371b9),
	.w4(32'h3ca11429),
	.w5(32'h3beca268),
	.w6(32'h3ba7d35c),
	.w7(32'hbb9288bf),
	.w8(32'h3af1ec71),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a8e9d),
	.w1(32'hbb0cbe9e),
	.w2(32'h3a901e31),
	.w3(32'hbae3d42a),
	.w4(32'hbb24b1a6),
	.w5(32'hbc329b68),
	.w6(32'h3a645022),
	.w7(32'hbc5a4d0d),
	.w8(32'hbc03d8a4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3c4d6),
	.w1(32'h39810b63),
	.w2(32'h3a4739fa),
	.w3(32'hbbdb5bbe),
	.w4(32'h3bea664d),
	.w5(32'hbb672c90),
	.w6(32'h3c0a5c6b),
	.w7(32'h3be5d117),
	.w8(32'hbc1f43b3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb513cf9),
	.w1(32'h3bd0ed5c),
	.w2(32'hbb51551c),
	.w3(32'h3ad0419f),
	.w4(32'h3b04f8e9),
	.w5(32'h39ee5e0f),
	.w6(32'h397a3481),
	.w7(32'hbbefc028),
	.w8(32'h39ade46a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f10cb9),
	.w1(32'hba3af646),
	.w2(32'h3c90f7ef),
	.w3(32'hbc433d8d),
	.w4(32'hbb7cd0ed),
	.w5(32'hbc38dcf7),
	.w6(32'h3b9b3266),
	.w7(32'hb8d1567c),
	.w8(32'hb8c6ce2d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0ab90),
	.w1(32'h3b2e6fb6),
	.w2(32'hba8ec9ff),
	.w3(32'hba8f94dc),
	.w4(32'hba89b0b4),
	.w5(32'h3938db22),
	.w6(32'h3ad25f31),
	.w7(32'h3bd583f9),
	.w8(32'h3b23bbe9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2936c),
	.w1(32'h3c6e8dae),
	.w2(32'h3c214750),
	.w3(32'h3bc01875),
	.w4(32'hbad8b5ea),
	.w5(32'h3c9c71cd),
	.w6(32'h3bc3dbb9),
	.w7(32'hbbcae1ce),
	.w8(32'hbadf02f5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c739f84),
	.w1(32'hbb0fc829),
	.w2(32'hbb84dee1),
	.w3(32'hbaa9337a),
	.w4(32'hbc6752ab),
	.w5(32'hbc47e21e),
	.w6(32'h3bbca22d),
	.w7(32'h3b9d4484),
	.w8(32'hbbfbf84a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28a729),
	.w1(32'hbb8d0525),
	.w2(32'h3b1ef857),
	.w3(32'h3c103278),
	.w4(32'h3b690785),
	.w5(32'h3c130c47),
	.w6(32'h3bcd661c),
	.w7(32'h3c59954e),
	.w8(32'hbc61b067),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99238c),
	.w1(32'h3b0f05ee),
	.w2(32'hbb058697),
	.w3(32'hbba2767a),
	.w4(32'h3bee90dd),
	.w5(32'h3b2bcc6e),
	.w6(32'h3a9838e1),
	.w7(32'hbb59d6e2),
	.w8(32'h3a54b373),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd205bd),
	.w1(32'hbbc8c708),
	.w2(32'hbb543657),
	.w3(32'h3bb744c7),
	.w4(32'hbc727f35),
	.w5(32'hbc4d986b),
	.w6(32'hbb2e1708),
	.w7(32'hbb56263c),
	.w8(32'hbc1996c4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf29c8b),
	.w1(32'h3abc775a),
	.w2(32'hbaa0177b),
	.w3(32'hbbcd8fb4),
	.w4(32'h3a811443),
	.w5(32'h3ba30241),
	.w6(32'hbc231e2e),
	.w7(32'h3913eb18),
	.w8(32'hbaab0424),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1388b),
	.w1(32'h3a527136),
	.w2(32'hbb9c0e66),
	.w3(32'h3ad71052),
	.w4(32'h3c0a36ba),
	.w5(32'hb985c54a),
	.w6(32'h3b37eb3f),
	.w7(32'hbbf08995),
	.w8(32'h3c4d48bb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccb75f),
	.w1(32'hbb572f7a),
	.w2(32'h3ba86aad),
	.w3(32'hba4cb964),
	.w4(32'hbc433adc),
	.w5(32'h3b518641),
	.w6(32'hbc44542b),
	.w7(32'hbbb75ad2),
	.w8(32'hbb978120),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a200d),
	.w1(32'hbbf70649),
	.w2(32'hbb9ba47e),
	.w3(32'h3d0dc517),
	.w4(32'hbae0d519),
	.w5(32'hbbd08a81),
	.w6(32'hbab78879),
	.w7(32'h3a0c198d),
	.w8(32'hbb6de305),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be56781),
	.w1(32'hba8bf8cc),
	.w2(32'h3bb3c649),
	.w3(32'h3b4a62c4),
	.w4(32'hba5563c9),
	.w5(32'hbb3f7957),
	.w6(32'hbc631121),
	.w7(32'hbb82f32e),
	.w8(32'h3b7b8bbf),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09bae1),
	.w1(32'hbc1f48a0),
	.w2(32'h3a40c5f7),
	.w3(32'h3a77412f),
	.w4(32'hbaaba0e7),
	.w5(32'hbca50ae6),
	.w6(32'h3bf0db5b),
	.w7(32'hbba5f40c),
	.w8(32'h3b3ab0c0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28c43e),
	.w1(32'h3a49513b),
	.w2(32'hbbf368ad),
	.w3(32'h3c38878f),
	.w4(32'h3ac3a0fb),
	.w5(32'h3b5d6b09),
	.w6(32'hbca43c12),
	.w7(32'h3b4e97ff),
	.w8(32'hbc0404be),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eb410),
	.w1(32'hbc7c99d0),
	.w2(32'hbcda4424),
	.w3(32'hbb58f00d),
	.w4(32'h3b2e78f6),
	.w5(32'h3ab4885a),
	.w6(32'h3a59aa93),
	.w7(32'h3af4c0a5),
	.w8(32'hbbb12eff),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d6735),
	.w1(32'hbad1d4d1),
	.w2(32'hbaf77ba1),
	.w3(32'hbc49a60f),
	.w4(32'hbb781f55),
	.w5(32'hbb22781e),
	.w6(32'hbbb6c414),
	.w7(32'h3b1389fd),
	.w8(32'hbc211c99),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a285e37),
	.w1(32'h3aa21112),
	.w2(32'h3b02cd80),
	.w3(32'hbbc836e1),
	.w4(32'h3a184b7c),
	.w5(32'h3b3aa3f9),
	.w6(32'hbc36b5ce),
	.w7(32'h3a025784),
	.w8(32'hbd4b8ec4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e70c5),
	.w1(32'hbb27085f),
	.w2(32'h3a50816a),
	.w3(32'hbc2acce7),
	.w4(32'hbae1c102),
	.w5(32'hbb7754e3),
	.w6(32'hba85d6b5),
	.w7(32'hbba31ca1),
	.w8(32'hbb6958d5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99fb9b),
	.w1(32'hbc21bf96),
	.w2(32'hbd24e050),
	.w3(32'h3bb7d372),
	.w4(32'hba266464),
	.w5(32'hbb2dbbc1),
	.w6(32'hbc011f3e),
	.w7(32'hb882e123),
	.w8(32'h3c458f20),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42fc00),
	.w1(32'hbd26f5f6),
	.w2(32'hbb384db3),
	.w3(32'hbb2bccd2),
	.w4(32'hbb845df2),
	.w5(32'h3bb9b653),
	.w6(32'hbb7b77c5),
	.w7(32'hbd2d7f9f),
	.w8(32'hbb04d192),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0682fe),
	.w1(32'h3b7131bd),
	.w2(32'h3ac0e4aa),
	.w3(32'h3b6352cc),
	.w4(32'hbb580f0b),
	.w5(32'h3c254850),
	.w6(32'hbb862f1c),
	.w7(32'hbb9ac009),
	.w8(32'h3bc954a2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fad63),
	.w1(32'h3d8cbab7),
	.w2(32'h3a852f7f),
	.w3(32'hbb2a4487),
	.w4(32'hbb8aba40),
	.w5(32'h3c0cff26),
	.w6(32'hbc434e08),
	.w7(32'h3be0044e),
	.w8(32'h3ba7428c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e4fe9),
	.w1(32'h3b7fa3aa),
	.w2(32'hbad69a5c),
	.w3(32'hbab345f0),
	.w4(32'hbbcfb784),
	.w5(32'h3b89c468),
	.w6(32'hbbbd2e71),
	.w7(32'hbb63c931),
	.w8(32'h3bab27e1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6be91f),
	.w1(32'hbbadfeae),
	.w2(32'hba1ca92c),
	.w3(32'h3abf3d90),
	.w4(32'hbbb8276a),
	.w5(32'hbbdf695b),
	.w6(32'h3b4fc8fa),
	.w7(32'h3c0e7457),
	.w8(32'h39cbd8a7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98cc5f),
	.w1(32'hb9849d34),
	.w2(32'hb7e70057),
	.w3(32'h3be7b7d7),
	.w4(32'hbc2a73fc),
	.w5(32'hb99d4db8),
	.w6(32'hbb95000c),
	.w7(32'hb8980b01),
	.w8(32'hbbbbbc34),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0718e2),
	.w1(32'hbb78f7c5),
	.w2(32'h38adfd4a),
	.w3(32'h3ab5264f),
	.w4(32'hbcd5ddb9),
	.w5(32'hbb30d039),
	.w6(32'h3b87e6ec),
	.w7(32'hbb58edb8),
	.w8(32'hbb9e1134),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa992d6),
	.w1(32'hb8cefee2),
	.w2(32'hbb85df23),
	.w3(32'hbc1f3de0),
	.w4(32'hbae24974),
	.w5(32'h3ba3f604),
	.w6(32'h3ac9ef7f),
	.w7(32'h3bb8a95e),
	.w8(32'h3bbfaa0d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a14dc),
	.w1(32'hbcd51455),
	.w2(32'hbad9c56f),
	.w3(32'h3c52b30e),
	.w4(32'h3b7ab8b9),
	.w5(32'hbb8cc913),
	.w6(32'h3b898e00),
	.w7(32'hbc843554),
	.w8(32'hbc111ea2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb0792),
	.w1(32'hbb1979ac),
	.w2(32'h3bb6c0ea),
	.w3(32'h3c39e3b4),
	.w4(32'h3910a171),
	.w5(32'h3b608184),
	.w6(32'hbbb11d0c),
	.w7(32'hbb26defa),
	.w8(32'h3b9650c2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a953533),
	.w1(32'hba997e68),
	.w2(32'h3b120675),
	.w3(32'hbc8c8b3d),
	.w4(32'hb9bb253d),
	.w5(32'h3b5b115f),
	.w6(32'h393d5194),
	.w7(32'h3b03e2ce),
	.w8(32'hb9cc143c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bb2fa),
	.w1(32'h3b57cd79),
	.w2(32'h3c117e2a),
	.w3(32'h399c96ff),
	.w4(32'hbae98545),
	.w5(32'h3b70260d),
	.w6(32'h397edb0f),
	.w7(32'h3c52803c),
	.w8(32'hbc2f38bd),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ff061),
	.w1(32'hbc05f071),
	.w2(32'h3924bc45),
	.w3(32'hbb05570f),
	.w4(32'hbc8f8ffd),
	.w5(32'h3b830cf2),
	.w6(32'hbb63eff9),
	.w7(32'hbc359ada),
	.w8(32'hbac628c0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2cfe6),
	.w1(32'h3cad5821),
	.w2(32'h3be5190d),
	.w3(32'h3aa82bca),
	.w4(32'h3b7341a8),
	.w5(32'hbcd28539),
	.w6(32'h3bda2afb),
	.w7(32'hba55847d),
	.w8(32'hbc4e6893),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aa6ac),
	.w1(32'h398d8918),
	.w2(32'hbb1acb48),
	.w3(32'hbbd2e227),
	.w4(32'hbb5d220d),
	.w5(32'h3abd8cca),
	.w6(32'h39b63404),
	.w7(32'h3c0d3596),
	.w8(32'hbb6bc90b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e389a),
	.w1(32'h3a8adce0),
	.w2(32'hbb16389c),
	.w3(32'hbbc4d6bb),
	.w4(32'hba6d55e5),
	.w5(32'h3c02e6ae),
	.w6(32'h3a3b0f0e),
	.w7(32'h3bdde404),
	.w8(32'h3c117ce2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b699ace),
	.w1(32'h3b73952c),
	.w2(32'hbc56c1df),
	.w3(32'h3bbca56a),
	.w4(32'h3ba2983e),
	.w5(32'h3c0c183e),
	.w6(32'h3b15934d),
	.w7(32'h3b472830),
	.w8(32'h3baf8d16),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c237a7e),
	.w1(32'h3b876e26),
	.w2(32'h3c235288),
	.w3(32'hbc089126),
	.w4(32'h37298ea4),
	.w5(32'h3c5fb4c7),
	.w6(32'h3c39434b),
	.w7(32'h3b4a513d),
	.w8(32'h3b817a0d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccc94a),
	.w1(32'h3b4959cf),
	.w2(32'h3c2a1468),
	.w3(32'h3b874c88),
	.w4(32'hbc3e98ab),
	.w5(32'h3c468542),
	.w6(32'h3a9f6229),
	.w7(32'hbac44d6a),
	.w8(32'hb9f44dc1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7b16c),
	.w1(32'h3ad2f0e2),
	.w2(32'h3baa4d1d),
	.w3(32'h3c48bd37),
	.w4(32'h3b17b5d9),
	.w5(32'hbc891fce),
	.w6(32'hbac0694e),
	.w7(32'hbb7d6399),
	.w8(32'h3b8b44f7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaab2c5),
	.w1(32'hbaebb3b4),
	.w2(32'hbb76c332),
	.w3(32'h3bbedad6),
	.w4(32'hbad0544b),
	.w5(32'h3b812683),
	.w6(32'h3bd5dcaa),
	.w7(32'hbae0f29f),
	.w8(32'h3bdb0228),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a3585),
	.w1(32'h3c72c05d),
	.w2(32'h3bdb6064),
	.w3(32'h3ba5de33),
	.w4(32'h3bcc7268),
	.w5(32'hbb97f1eb),
	.w6(32'h3bab240e),
	.w7(32'h3bcb2447),
	.w8(32'hbbd95556),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e50a2),
	.w1(32'h3b8578a7),
	.w2(32'h3b1e140c),
	.w3(32'hbb0d24d1),
	.w4(32'h3b871102),
	.w5(32'h3b1777a8),
	.w6(32'hbb97ce11),
	.w7(32'hbb035a2d),
	.w8(32'h3bc9e543),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa2e83),
	.w1(32'h3a0abfaf),
	.w2(32'hbc8d5cfc),
	.w3(32'h3bfedffb),
	.w4(32'h3b261104),
	.w5(32'hbbc18486),
	.w6(32'hba057820),
	.w7(32'hbb310481),
	.w8(32'h3c4a02ee),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9990),
	.w1(32'h3c8aa8cd),
	.w2(32'h3c864e7a),
	.w3(32'hbbd6ac52),
	.w4(32'hbba6d5e5),
	.w5(32'hb77f57e0),
	.w6(32'hbaa69102),
	.w7(32'h3b8e21c3),
	.w8(32'h3c07f12c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d96d3),
	.w1(32'hbba91f47),
	.w2(32'h3ae0dc1f),
	.w3(32'h3bfca05e),
	.w4(32'h3c9cabea),
	.w5(32'hbc49327f),
	.w6(32'h3b95a2e0),
	.w7(32'h3b99d756),
	.w8(32'h3ba6e232),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc806b),
	.w1(32'h3bcdd3d9),
	.w2(32'h3a0fc56d),
	.w3(32'hbb885023),
	.w4(32'hbbbbd1a9),
	.w5(32'h3b4823a4),
	.w6(32'hba1295c1),
	.w7(32'h3a7c5343),
	.w8(32'h3a73ceaa),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66576b),
	.w1(32'h3c2e3098),
	.w2(32'h39bd7067),
	.w3(32'hbb39a6ee),
	.w4(32'h3cbb3431),
	.w5(32'hbb979275),
	.w6(32'h3c8923ff),
	.w7(32'hbc11b911),
	.w8(32'h3abf4a79),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914432),
	.w1(32'h3b995a95),
	.w2(32'h3b8c01fa),
	.w3(32'h3c2ad11c),
	.w4(32'h3bd18b22),
	.w5(32'hb9946c06),
	.w6(32'hbb2e49cf),
	.w7(32'h3a8ad5b4),
	.w8(32'h398d3d68),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b545231),
	.w1(32'hbc27c6ef),
	.w2(32'h3b8ba6cb),
	.w3(32'h3b0a4a63),
	.w4(32'h3bbe82d3),
	.w5(32'hb9844948),
	.w6(32'h3bd5882a),
	.w7(32'h3bca2eb8),
	.w8(32'h3bf91aa1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3937854b),
	.w1(32'hbc04e3b5),
	.w2(32'h3bbc55d3),
	.w3(32'h3bc2453a),
	.w4(32'h3a8d5479),
	.w5(32'hbb854519),
	.w6(32'hba478519),
	.w7(32'hbb50b272),
	.w8(32'h3bbf57c0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba329a71),
	.w1(32'hbbd290d4),
	.w2(32'hbc10cd30),
	.w3(32'h3c420377),
	.w4(32'h3bee2636),
	.w5(32'hba1ad854),
	.w6(32'h3c0f0b79),
	.w7(32'h39039b99),
	.w8(32'h3b83a733),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fd72c),
	.w1(32'h3c0897b0),
	.w2(32'hbb92e8ca),
	.w3(32'hbc10e1f1),
	.w4(32'hba8cd560),
	.w5(32'h3b0bec43),
	.w6(32'hbad43026),
	.w7(32'hbb5c6fc5),
	.w8(32'hbaf8852a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dab9a5),
	.w1(32'h3c0d3631),
	.w2(32'h3c316344),
	.w3(32'h3c6b77d3),
	.w4(32'hbac3f6c6),
	.w5(32'h3be08bca),
	.w6(32'hbc3aff8f),
	.w7(32'h3bd9a33f),
	.w8(32'h3cc6214e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6225c),
	.w1(32'h3a01afaf),
	.w2(32'hbb31d1fa),
	.w3(32'hbb4830cf),
	.w4(32'h3b268cfd),
	.w5(32'h3a5228f1),
	.w6(32'h3b9f324d),
	.w7(32'h3af71bee),
	.w8(32'hba4483fc),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00deaf),
	.w1(32'hb9bb1a8b),
	.w2(32'h3bf4a912),
	.w3(32'hb940e3c8),
	.w4(32'hbb4ad078),
	.w5(32'h3ba41558),
	.w6(32'h3bd7b32c),
	.w7(32'h3b186d47),
	.w8(32'h3be12877),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3be1d),
	.w1(32'h3ba6a3ba),
	.w2(32'h3b607332),
	.w3(32'hbac5fab6),
	.w4(32'h3b6bc597),
	.w5(32'hbbb62ef2),
	.w6(32'h3c52cc79),
	.w7(32'h3c28c8ab),
	.w8(32'h3b4b65bc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc27a6c),
	.w1(32'h3c557823),
	.w2(32'hbad4b74c),
	.w3(32'h3b972a26),
	.w4(32'h3b561fee),
	.w5(32'h3ade53da),
	.w6(32'h3a944309),
	.w7(32'hbb0a26b2),
	.w8(32'h3b8b87a5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd0f3d),
	.w1(32'hb9e580af),
	.w2(32'hbb32d3e5),
	.w3(32'hbb11de92),
	.w4(32'hbb19977d),
	.w5(32'h3bafa339),
	.w6(32'h3c1f3f8b),
	.w7(32'hbbcfc27a),
	.w8(32'hb922687b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0ccda),
	.w1(32'h3a2c9f6b),
	.w2(32'h3921e8dd),
	.w3(32'h3ab94181),
	.w4(32'h3a782628),
	.w5(32'h3ba4182b),
	.w6(32'h3af1769b),
	.w7(32'hb9a32886),
	.w8(32'h3af98fdf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd10031),
	.w1(32'hba24a4a8),
	.w2(32'h3c3fbecd),
	.w3(32'hb9d54b75),
	.w4(32'h3bc6d4de),
	.w5(32'h3b7dc2c6),
	.w6(32'h3c05552a),
	.w7(32'h3ac26bd6),
	.w8(32'hbb123882),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb192df),
	.w1(32'h3b31908c),
	.w2(32'hbadeb842),
	.w3(32'hbabce0b1),
	.w4(32'h3c8f70a9),
	.w5(32'hbb786a62),
	.w6(32'h3a0c09cf),
	.w7(32'hbbaf4ab4),
	.w8(32'h3c1d7983),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ce61c),
	.w1(32'hbc725f56),
	.w2(32'hbbc6deaa),
	.w3(32'h3c4d6ec7),
	.w4(32'hbaf7c602),
	.w5(32'hbca81445),
	.w6(32'hbbcb744e),
	.w7(32'h3bab0ce9),
	.w8(32'h3c499b6e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3c735),
	.w1(32'h3cfbddfd),
	.w2(32'hbc0fce93),
	.w3(32'h3c8a4a90),
	.w4(32'h3ad931ab),
	.w5(32'h3b5a45b7),
	.w6(32'h3a84d474),
	.w7(32'h3b988f4e),
	.w8(32'h3c1edbb2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc126712),
	.w1(32'hbc626fb4),
	.w2(32'hbc0b9adc),
	.w3(32'hbb243e46),
	.w4(32'h3b81989c),
	.w5(32'hbc63699f),
	.w6(32'h3b9c6803),
	.w7(32'h3c3a04ca),
	.w8(32'hba55462b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c352864),
	.w1(32'hbbb92df2),
	.w2(32'h39ea7aad),
	.w3(32'hba7c3b33),
	.w4(32'h39fe15d3),
	.w5(32'hbb98567d),
	.w6(32'hbb893c63),
	.w7(32'h3c0cac79),
	.w8(32'hbaafcc60),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc224663),
	.w1(32'hbbd254fe),
	.w2(32'h3af3d00c),
	.w3(32'hbc7419c9),
	.w4(32'hbb701cbd),
	.w5(32'hbbd12b14),
	.w6(32'h392d149d),
	.w7(32'h3c84811f),
	.w8(32'hbaa40eda),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc100080),
	.w1(32'hbb9e54ab),
	.w2(32'h3c85998a),
	.w3(32'hbbee9154),
	.w4(32'hbc0ff08f),
	.w5(32'h3c0ccf77),
	.w6(32'hbb27ff09),
	.w7(32'hbae29b12),
	.w8(32'hba81388c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81aa60),
	.w1(32'hbab4f36b),
	.w2(32'hbb4215de),
	.w3(32'h3b7b0ecf),
	.w4(32'h3a21cfbb),
	.w5(32'hbb4e8d68),
	.w6(32'hbac2dfaa),
	.w7(32'h3b2499f1),
	.w8(32'hbb04261f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc79a09),
	.w1(32'h3957bd38),
	.w2(32'h3c738e73),
	.w3(32'h3c844ba1),
	.w4(32'h3b061cb6),
	.w5(32'hba31b7d5),
	.w6(32'h3c46940b),
	.w7(32'hbc1f7b33),
	.w8(32'hbb0ce992),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabab72d),
	.w1(32'hbad0eb7f),
	.w2(32'h3a160cfe),
	.w3(32'h3b8bcb9d),
	.w4(32'hbaaa1dbc),
	.w5(32'hbc5e4500),
	.w6(32'hbada604b),
	.w7(32'h3b301c87),
	.w8(32'hbb2a608b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b5c66),
	.w1(32'h3a970c8d),
	.w2(32'h3b502c82),
	.w3(32'hbc1b06b9),
	.w4(32'hb947d25f),
	.w5(32'hb98ce6a3),
	.w6(32'hb9d18e95),
	.w7(32'h3cbad7b4),
	.w8(32'h3bf4c6dc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4de1de),
	.w1(32'hbc8f35e5),
	.w2(32'hbbb63770),
	.w3(32'hbab7ff85),
	.w4(32'hbc4bc8d8),
	.w5(32'hbc119927),
	.w6(32'h3c3ce12e),
	.w7(32'hbc57b73c),
	.w8(32'h3c26d21a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5520fc),
	.w1(32'hbc36ce3d),
	.w2(32'h3c1be9cf),
	.w3(32'h3c269054),
	.w4(32'hbc33178c),
	.w5(32'hbbab67b0),
	.w6(32'hbb747ae7),
	.w7(32'hbbd30597),
	.w8(32'h3c2d1432),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe9b06),
	.w1(32'h3c0abf37),
	.w2(32'h3b52bb24),
	.w3(32'hbbcf4aba),
	.w4(32'hbb77974f),
	.w5(32'hba9f9d37),
	.w6(32'h3b566a1a),
	.w7(32'hbb079ed0),
	.w8(32'h3b93cee9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43cc63),
	.w1(32'hbb87eea9),
	.w2(32'h3c772097),
	.w3(32'hb85de44b),
	.w4(32'hbc3edc2b),
	.w5(32'hbb9997ca),
	.w6(32'hbc6f21e6),
	.w7(32'hbc331a05),
	.w8(32'h3cba2d1d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d590),
	.w1(32'hba9caf80),
	.w2(32'h3a906433),
	.w3(32'hbb23caed),
	.w4(32'h3ba22ea6),
	.w5(32'hbb640783),
	.w6(32'hbc948cef),
	.w7(32'hbc4f4871),
	.w8(32'hbb466ec5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab12d3),
	.w1(32'hb69bce90),
	.w2(32'hbcca1c89),
	.w3(32'h3bba0f0a),
	.w4(32'hbaf86a1d),
	.w5(32'hbc2ea2dc),
	.w6(32'h3ba3fc4d),
	.w7(32'hba79fb29),
	.w8(32'h3a959ee2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc517f5e),
	.w1(32'h3c2b979b),
	.w2(32'h37d29161),
	.w3(32'hbba9d722),
	.w4(32'hbab69a6b),
	.w5(32'hbbe5d64e),
	.w6(32'h3aa9dfcb),
	.w7(32'h397315c8),
	.w8(32'hbb7a51cc),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c77dde),
	.w1(32'h3aa716e6),
	.w2(32'hbb388db2),
	.w3(32'h3c85e653),
	.w4(32'hbc50a41b),
	.w5(32'hbc040b80),
	.w6(32'h3b8560f8),
	.w7(32'hbbc095c5),
	.w8(32'h3ba74601),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bcae0),
	.w1(32'hbae95ef2),
	.w2(32'h3bd7a602),
	.w3(32'hbc2fc07f),
	.w4(32'h3cacd447),
	.w5(32'h3c670616),
	.w6(32'h3c14c07e),
	.w7(32'h3bc91748),
	.w8(32'hbc0cb9d7),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b951b42),
	.w1(32'hbb54c88c),
	.w2(32'h3a88ac8e),
	.w3(32'h3ba4ff30),
	.w4(32'h3a4be091),
	.w5(32'h3b3a2404),
	.w6(32'h3bd756c6),
	.w7(32'hbb89341f),
	.w8(32'h3b60533f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afefbe4),
	.w1(32'h3b120f97),
	.w2(32'hbc517bb1),
	.w3(32'hbc707cde),
	.w4(32'h3c563fa9),
	.w5(32'hbc4309f8),
	.w6(32'hb9bd3bf4),
	.w7(32'hbbe27bd8),
	.w8(32'h3b62b189),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80336a),
	.w1(32'h3ba6524b),
	.w2(32'hbb2801c7),
	.w3(32'hbc67b7b0),
	.w4(32'hba2e71ec),
	.w5(32'h3b058dbf),
	.w6(32'hbb6753de),
	.w7(32'h3b0faeaa),
	.w8(32'h3bde2c0d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5e782),
	.w1(32'hbc93e824),
	.w2(32'h3b239c0c),
	.w3(32'hbc41abe7),
	.w4(32'h3ba2203d),
	.w5(32'hbc1a4325),
	.w6(32'hbb0b0452),
	.w7(32'hbb182a09),
	.w8(32'hbb0bb929),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d8838),
	.w1(32'h3b149fdd),
	.w2(32'hbad9f65e),
	.w3(32'h3b312914),
	.w4(32'hbabfd4d0),
	.w5(32'hbaa434e9),
	.w6(32'h3b4ff88c),
	.w7(32'h3bd83c29),
	.w8(32'h39a27e11),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a9286),
	.w1(32'hbc036efb),
	.w2(32'h3ab3603a),
	.w3(32'h3bbd3c6d),
	.w4(32'hbc4e48ef),
	.w5(32'hbc9fda6f),
	.w6(32'h3c456a6f),
	.w7(32'hbbfc51e6),
	.w8(32'hb9199787),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d4a0),
	.w1(32'h3aa90678),
	.w2(32'h3c6a24a8),
	.w3(32'h3b5a4575),
	.w4(32'h3ae9d7c2),
	.w5(32'h3c9ead8b),
	.w6(32'h3bb6c4dc),
	.w7(32'hbb30a73b),
	.w8(32'hbb89edcc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f3a3e),
	.w1(32'hbaee2c6d),
	.w2(32'hbb2a8302),
	.w3(32'hb96d5234),
	.w4(32'hbb1e12e3),
	.w5(32'hbad1e767),
	.w6(32'h3b5ccde0),
	.w7(32'h3b8bc7f2),
	.w8(32'hba86fcba),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b252f8b),
	.w1(32'hbc0894e5),
	.w2(32'h3bf5e13d),
	.w3(32'h3bb6e0f7),
	.w4(32'hbc9ecb9d),
	.w5(32'h3b122390),
	.w6(32'h3bad02d0),
	.w7(32'h3bab0748),
	.w8(32'hbb8bf117),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba79ec4),
	.w1(32'h3bfe8dfd),
	.w2(32'h3c76b581),
	.w3(32'hbbdf454d),
	.w4(32'h3ad0b31a),
	.w5(32'h3bf5c475),
	.w6(32'h3bc9f561),
	.w7(32'h3b61e60e),
	.w8(32'hbc88c3e0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0f1cc),
	.w1(32'h3ae315bf),
	.w2(32'h3c04c346),
	.w3(32'h3c8a677b),
	.w4(32'h3c3a0dda),
	.w5(32'h3cd56f4a),
	.w6(32'hbd4fb942),
	.w7(32'h3bcaf602),
	.w8(32'h3c3588bd),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e134d),
	.w1(32'hbbe94ca1),
	.w2(32'hbb0c6b05),
	.w3(32'hbba72ac1),
	.w4(32'hbbb6f094),
	.w5(32'h3b8aa2c7),
	.w6(32'hbb9b163e),
	.w7(32'h3b9ec6a6),
	.w8(32'h3b33b9dc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c1b61),
	.w1(32'h3c04c126),
	.w2(32'h3c1a4263),
	.w3(32'h3c0a1fc4),
	.w4(32'h3a8738ff),
	.w5(32'hbc8de04a),
	.w6(32'h3ca3e5b3),
	.w7(32'h3a3703aa),
	.w8(32'h3cd88129),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc696804),
	.w1(32'h3ab4ead4),
	.w2(32'hbc74128b),
	.w3(32'hbc7fe756),
	.w4(32'h3b3a303b),
	.w5(32'hbba93d2c),
	.w6(32'h3b7be8b0),
	.w7(32'h3c83c87d),
	.w8(32'h3c840d5f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f3757),
	.w1(32'hbc47b9ff),
	.w2(32'h3cab15ad),
	.w3(32'hbc2bccbe),
	.w4(32'h3b938eff),
	.w5(32'hbcae2353),
	.w6(32'hb813e72e),
	.w7(32'h3c645f37),
	.w8(32'h3bf0f1a6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12b475),
	.w1(32'h3cc46618),
	.w2(32'h3cb3786e),
	.w3(32'h3b971c88),
	.w4(32'hba282480),
	.w5(32'hbb514076),
	.w6(32'h3bde2751),
	.w7(32'hbc871c2d),
	.w8(32'h3b1d658a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d22302),
	.w1(32'hbbc6bbba),
	.w2(32'hbc1d9bda),
	.w3(32'hbc2f76f1),
	.w4(32'hbb9e7033),
	.w5(32'h399a3d7b),
	.w6(32'hbb950826),
	.w7(32'hbbca2180),
	.w8(32'hba887dea),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc115ac5),
	.w1(32'hbb2f0d54),
	.w2(32'hbb564f5b),
	.w3(32'h3c25e38a),
	.w4(32'hbbbfeb98),
	.w5(32'h39b84e60),
	.w6(32'h3ca9442d),
	.w7(32'hbb71cc45),
	.w8(32'hbba15659),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0f911),
	.w1(32'hbc8e8bbe),
	.w2(32'h3bb0bd3b),
	.w3(32'hbaf9714c),
	.w4(32'h3c80a5c9),
	.w5(32'h3b802c34),
	.w6(32'hbbad86d8),
	.w7(32'h3cc58663),
	.w8(32'hbc43f63e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c975cc2),
	.w1(32'hbcd87bc5),
	.w2(32'h3c49b9b2),
	.w3(32'h3c1ac27c),
	.w4(32'h3ba33f69),
	.w5(32'h3c25d3c3),
	.w6(32'h3ad36dba),
	.w7(32'hbcb7dbca),
	.w8(32'h3bfa8b09),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5690b),
	.w1(32'hbc216781),
	.w2(32'h3b9e382f),
	.w3(32'hba66bba6),
	.w4(32'hbb8ebc1e),
	.w5(32'hbc95df11),
	.w6(32'h3d83c410),
	.w7(32'h3b921dc3),
	.w8(32'h3bb0a0bc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59e4b7),
	.w1(32'hbbfa989d),
	.w2(32'hbae3365d),
	.w3(32'hbc0d57f8),
	.w4(32'hbbff3a11),
	.w5(32'hbb5b0468),
	.w6(32'h3c7bc336),
	.w7(32'hbc51fcf4),
	.w8(32'hba88f53c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c287804),
	.w1(32'h3b44f01e),
	.w2(32'hbbd27dd0),
	.w3(32'h3bab26c5),
	.w4(32'h3c019d55),
	.w5(32'h3bc96720),
	.w6(32'hbbfcfa26),
	.w7(32'h3ad67b9a),
	.w8(32'h391289dc),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bd3ce),
	.w1(32'hb8835746),
	.w2(32'h3a2addee),
	.w3(32'h3a5c1dd7),
	.w4(32'hbc4d9449),
	.w5(32'hbaa86609),
	.w6(32'hbc95c6f3),
	.w7(32'hbaf39a85),
	.w8(32'h3873294c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb925184),
	.w1(32'hbc91de1b),
	.w2(32'h3b73ba59),
	.w3(32'hb9d8ab57),
	.w4(32'hbab30b96),
	.w5(32'hba4ef13d),
	.w6(32'hbc4a20f6),
	.w7(32'h3b073dfd),
	.w8(32'h3bcd1a08),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63fa11),
	.w1(32'hbb8f861a),
	.w2(32'hbb0e6549),
	.w3(32'hbc2807c1),
	.w4(32'h3c1bfbbb),
	.w5(32'hbc2eab27),
	.w6(32'hbc809187),
	.w7(32'h3b372f2d),
	.w8(32'hbcd0a234),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d8cef),
	.w1(32'hbc77ed50),
	.w2(32'h3b312afa),
	.w3(32'hbbad0846),
	.w4(32'h3bbb0560),
	.w5(32'h3c2679a8),
	.w6(32'h3b2cb5a6),
	.w7(32'hb8486f29),
	.w8(32'hb971afa7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6a531),
	.w1(32'h3bbc5e47),
	.w2(32'hbcb0d2d4),
	.w3(32'hbc03fc5b),
	.w4(32'hbb98544d),
	.w5(32'hbc7a8412),
	.w6(32'h3c69e361),
	.w7(32'hbbb8e0df),
	.w8(32'hbc3d457c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc22e3c),
	.w1(32'hbb78e4f7),
	.w2(32'h3a7767f1),
	.w3(32'hbb862589),
	.w4(32'h39e99cfa),
	.w5(32'h3b852699),
	.w6(32'hbca1b604),
	.w7(32'h3a4070ed),
	.w8(32'hbc24a44f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cab0c),
	.w1(32'hbb72f4de),
	.w2(32'hb981b627),
	.w3(32'h3c4258e9),
	.w4(32'hbca851fa),
	.w5(32'hbc135f7b),
	.w6(32'hbc1851ba),
	.w7(32'h3ba6f08a),
	.w8(32'h3b8a32b8),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb477bd4),
	.w1(32'hbbb3b4e1),
	.w2(32'h3c49e65b),
	.w3(32'hbaf8a8ef),
	.w4(32'hbc2d5d40),
	.w5(32'hbc151ae5),
	.w6(32'h3c96a3ff),
	.w7(32'h3bf714b5),
	.w8(32'hbbf9f683),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b077a),
	.w1(32'hbc18447b),
	.w2(32'h3ae5ec88),
	.w3(32'hbb05bfed),
	.w4(32'h3c86fc20),
	.w5(32'h3c7345f3),
	.w6(32'h3c9e2ab8),
	.w7(32'h3c6a82c9),
	.w8(32'hbc651a40),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba50efd),
	.w1(32'hbc8aae54),
	.w2(32'hbbef22d2),
	.w3(32'hbc845d1c),
	.w4(32'hbb448784),
	.w5(32'h3c2ef90a),
	.w6(32'h3b8d1f85),
	.w7(32'hbb8f64ff),
	.w8(32'h3c86bfb5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74dd31),
	.w1(32'h3cdf3601),
	.w2(32'h3b2f7659),
	.w3(32'hbbe4fbbc),
	.w4(32'h39dcfe2f),
	.w5(32'hbc020ed7),
	.w6(32'hbc3f48eb),
	.w7(32'hbbaf8b36),
	.w8(32'h3b174ee8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5b4b0),
	.w1(32'hbbbf81bf),
	.w2(32'hbbd262d1),
	.w3(32'hb9a4e699),
	.w4(32'h3b7b7e24),
	.w5(32'hba184a20),
	.w6(32'h3c25589d),
	.w7(32'hbc438bbd),
	.w8(32'hba87f32d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba712d42),
	.w1(32'hbb47f745),
	.w2(32'h3b9dc6fb),
	.w3(32'hbb92ae0f),
	.w4(32'hba9cbe4c),
	.w5(32'hbc6e387f),
	.w6(32'hbc71fbc1),
	.w7(32'hbaf5d59e),
	.w8(32'hbb29be1a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae19e2),
	.w1(32'h3bc1769c),
	.w2(32'h3bfe4ebc),
	.w3(32'hbbd7518d),
	.w4(32'h3b96ae39),
	.w5(32'h3ca14e48),
	.w6(32'h3bb6e86d),
	.w7(32'h3cae0b79),
	.w8(32'h3ce1f023),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ead49),
	.w1(32'h3c9c7848),
	.w2(32'hbb9fe725),
	.w3(32'hbc064ef9),
	.w4(32'h3c4ebb70),
	.w5(32'hbbab4765),
	.w6(32'h3bc1aec7),
	.w7(32'hbc85f4dd),
	.w8(32'h3cb5f85d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef9723),
	.w1(32'h3b3a7762),
	.w2(32'h3d3c1a59),
	.w3(32'h3c58d810),
	.w4(32'h3a5bb5d7),
	.w5(32'h3cf3f60e),
	.w6(32'hba66b5d9),
	.w7(32'h3ab1943c),
	.w8(32'h3bda916e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b627127),
	.w1(32'h3905baab),
	.w2(32'h3baeb3b2),
	.w3(32'hba3530f8),
	.w4(32'h3c30eedd),
	.w5(32'hbc5f52e3),
	.w6(32'h3d24e5d7),
	.w7(32'h3c1d1438),
	.w8(32'h3c337086),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eedda),
	.w1(32'h3b2340ed),
	.w2(32'h3aef5b87),
	.w3(32'hbb12834b),
	.w4(32'h3abb8f57),
	.w5(32'hbbbb42c9),
	.w6(32'h39f6dfb7),
	.w7(32'hbc081bd4),
	.w8(32'h3c577af7),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4fefae),
	.w1(32'h3b32ae36),
	.w2(32'h3c45b6eb),
	.w3(32'h3b60b3ba),
	.w4(32'hbc4d27ee),
	.w5(32'hbb115900),
	.w6(32'h3a60a2ea),
	.w7(32'hbc07c1ce),
	.w8(32'hbcffa216),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e850c),
	.w1(32'hbaff927d),
	.w2(32'hbd0df6d0),
	.w3(32'hbbdc0a02),
	.w4(32'h3c61614b),
	.w5(32'hbac73e9d),
	.w6(32'hbb1c691c),
	.w7(32'hbba26f6b),
	.w8(32'hbb472325),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc98ba0),
	.w1(32'h3b29ff8a),
	.w2(32'h3af86eb4),
	.w3(32'hbbe7d082),
	.w4(32'hbbc946e7),
	.w5(32'h3b96af61),
	.w6(32'hbb3ec981),
	.w7(32'h3b4fc2be),
	.w8(32'h3c6655c1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6f5f4),
	.w1(32'h3b705dc0),
	.w2(32'h39ee3e6f),
	.w3(32'hbca2b390),
	.w4(32'h3bbc3630),
	.w5(32'hbaa49e5b),
	.w6(32'h3bc297bb),
	.w7(32'hbbd9027a),
	.w8(32'hba40c005),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c375d),
	.w1(32'hbbeb5c12),
	.w2(32'h3b66b232),
	.w3(32'h3d07f22c),
	.w4(32'hbb00d446),
	.w5(32'h3bcbf7a2),
	.w6(32'hbaa6c779),
	.w7(32'hba75c8bd),
	.w8(32'h3c11ca8a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af02ce9),
	.w1(32'h3b880528),
	.w2(32'hb960728e),
	.w3(32'h3baaa960),
	.w4(32'h3a4a20a6),
	.w5(32'h3b81689a),
	.w6(32'h39ed5608),
	.w7(32'h3ca7fb26),
	.w8(32'hbbf94241),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc605879),
	.w1(32'hbbb679cf),
	.w2(32'h3b5e3960),
	.w3(32'hb9e42d0c),
	.w4(32'h3b36cc9d),
	.w5(32'h3b17bce9),
	.w6(32'hbb05c19b),
	.w7(32'hbbdd2e44),
	.w8(32'h3b207f15),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81cf7c),
	.w1(32'h39a1a725),
	.w2(32'h3b7045d7),
	.w3(32'hbccef6bc),
	.w4(32'hbc0b8bce),
	.w5(32'hbaba5470),
	.w6(32'hbc0499bc),
	.w7(32'h3c9d1ccb),
	.w8(32'hbc0b9492),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc428ba),
	.w1(32'h3c7f5955),
	.w2(32'h3c240b8e),
	.w3(32'h3b878b94),
	.w4(32'h3b4bb2a6),
	.w5(32'h3bc2e45b),
	.w6(32'hbbf6ef7d),
	.w7(32'h3ae67858),
	.w8(32'hbaa9adee),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4830a7),
	.w1(32'h3c0afba5),
	.w2(32'hbcb19f33),
	.w3(32'hbb8aded5),
	.w4(32'hbb01569d),
	.w5(32'hbab767bb),
	.w6(32'h3b7f8cf8),
	.w7(32'hb9ef5e35),
	.w8(32'h3cafb60e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08483f),
	.w1(32'hbc43e0de),
	.w2(32'h3ba61dc7),
	.w3(32'hbbbc2457),
	.w4(32'hbb6ee54e),
	.w5(32'hbc02d066),
	.w6(32'hbbafc3af),
	.w7(32'h39dbb8f0),
	.w8(32'h3a364dbb),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbea287),
	.w1(32'h3bfcc5ba),
	.w2(32'hb9bef557),
	.w3(32'h3c7066dd),
	.w4(32'hbab32adc),
	.w5(32'hb8b87db1),
	.w6(32'h3c0a820d),
	.w7(32'hbac50acd),
	.w8(32'hb9e893cd),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81e878),
	.w1(32'hbb914965),
	.w2(32'hbc0e4ef3),
	.w3(32'hbc10ebea),
	.w4(32'h3b5421d7),
	.w5(32'h3b3bde59),
	.w6(32'hb719040d),
	.w7(32'hbb32f9c4),
	.w8(32'hbb67fe68),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac94b6f),
	.w1(32'h3988f350),
	.w2(32'h3c81bd0b),
	.w3(32'hbbdb4ba1),
	.w4(32'h3b1ec738),
	.w5(32'hbc630a63),
	.w6(32'hba9dd8c9),
	.w7(32'h3bc59d8e),
	.w8(32'hbce6b202),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1c609),
	.w1(32'h3c391a61),
	.w2(32'hbbe76924),
	.w3(32'h3ce02b9d),
	.w4(32'hbca65953),
	.w5(32'hbbd19915),
	.w6(32'hbb8be8c1),
	.w7(32'hba540891),
	.w8(32'hbc5978c3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7533d),
	.w1(32'hbad3b347),
	.w2(32'hbc2ce975),
	.w3(32'hbc28d496),
	.w4(32'h3bd8443e),
	.w5(32'h3ab9c4bc),
	.w6(32'hbb288c98),
	.w7(32'hbab92771),
	.w8(32'hbb5d2ff5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e967f),
	.w1(32'hbad1d6c0),
	.w2(32'hbbc38618),
	.w3(32'hbb5607f1),
	.w4(32'h3bbc6ec7),
	.w5(32'hbb8cc87a),
	.w6(32'h3c3ad16d),
	.w7(32'hbd3d9e21),
	.w8(32'h3a373576),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c355357),
	.w1(32'hbb0d652d),
	.w2(32'h3bee8d83),
	.w3(32'h3bafe296),
	.w4(32'hb9e16756),
	.w5(32'h3c636038),
	.w6(32'hbaf8fa85),
	.w7(32'h3b8b0f37),
	.w8(32'h3b552c95),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0a4bc),
	.w1(32'hbc984c86),
	.w2(32'h3b8e9c00),
	.w3(32'h3b1983bc),
	.w4(32'hbb777cc2),
	.w5(32'hbc1b22e3),
	.w6(32'h3c9494dd),
	.w7(32'hbba1645b),
	.w8(32'h3b3e48ca),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba279b4d),
	.w1(32'hbb1ae178),
	.w2(32'h3d13dd83),
	.w3(32'hbb4748a8),
	.w4(32'h3ba3b4e7),
	.w5(32'h3a0ce943),
	.w6(32'hb866ce4a),
	.w7(32'h3aa77ca1),
	.w8(32'h3ba36a96),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9485b1c),
	.w1(32'h3c9cdba1),
	.w2(32'hbb807f50),
	.w3(32'hbc98edf5),
	.w4(32'h3b45bf13),
	.w5(32'hbbbd4dbb),
	.w6(32'hbb6fe6df),
	.w7(32'hbc00ce71),
	.w8(32'hbc2b6127),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1ad00),
	.w1(32'hbd19da82),
	.w2(32'hb9dbb934),
	.w3(32'h3b5a287e),
	.w4(32'hbbf08689),
	.w5(32'hb817a528),
	.w6(32'h3b039481),
	.w7(32'hbc8d5fc8),
	.w8(32'hbc9670a7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3ff0d),
	.w1(32'h3b86d137),
	.w2(32'h3a9a9855),
	.w3(32'h3a59394a),
	.w4(32'hbb4f96e2),
	.w5(32'h3b289a97),
	.w6(32'hb917ee90),
	.w7(32'h3b85fdb0),
	.w8(32'h3b2e3fe6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f3cfc),
	.w1(32'h3c83f8e1),
	.w2(32'h3cbd6160),
	.w3(32'h3afb3b40),
	.w4(32'hbc9b76f1),
	.w5(32'hbbad6bd6),
	.w6(32'h3b428ebc),
	.w7(32'hbc99ff59),
	.w8(32'hbb50e484),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be0e80),
	.w1(32'h3a4aed89),
	.w2(32'hbab7bf40),
	.w3(32'h3a9a8b30),
	.w4(32'hbbd439d0),
	.w5(32'h3b5c6b2d),
	.w6(32'h3ce13e1b),
	.w7(32'hbbce2afc),
	.w8(32'hba61e850),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe4be5),
	.w1(32'h3c0c555e),
	.w2(32'hbbb7fac8),
	.w3(32'hbd1e1f01),
	.w4(32'hbbf00d71),
	.w5(32'h3bb47c30),
	.w6(32'hbb620809),
	.w7(32'h3c9eee60),
	.w8(32'hb92e2feb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b3c26),
	.w1(32'h3c6c13cb),
	.w2(32'hbbba5df2),
	.w3(32'hbc9fa103),
	.w4(32'hbae53fe5),
	.w5(32'h3aad2af9),
	.w6(32'h3b156e69),
	.w7(32'h3bb3ad33),
	.w8(32'h3aa78bb6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13ca4c),
	.w1(32'h3a7dd93e),
	.w2(32'hbc511915),
	.w3(32'h3bab94bb),
	.w4(32'hbb46058a),
	.w5(32'h3a89ab00),
	.w6(32'hbb986f58),
	.w7(32'hbb96a39b),
	.w8(32'hb9c1b784),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb985958),
	.w1(32'h3d0cfd41),
	.w2(32'hbb74412e),
	.w3(32'h3bdfdfea),
	.w4(32'hbc0f9556),
	.w5(32'hba167a58),
	.w6(32'h3bdbe937),
	.w7(32'hb94ca496),
	.w8(32'h3b5a7592),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc133a05),
	.w1(32'h3bf1d3a6),
	.w2(32'hbc2401d2),
	.w3(32'h363b15dc),
	.w4(32'h3bed0d7c),
	.w5(32'hbbf20824),
	.w6(32'hbbb9c85f),
	.w7(32'h3b6399cc),
	.w8(32'h3b6d09bd),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb075b8e),
	.w1(32'h39e929d6),
	.w2(32'h3b048b29),
	.w3(32'h37e19bae),
	.w4(32'h3b4aaff2),
	.w5(32'hbb8d6dee),
	.w6(32'hbc1464a0),
	.w7(32'hbaa32bc5),
	.w8(32'hba34dd38),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed84ef),
	.w1(32'hbbaedcfc),
	.w2(32'h3c4b114f),
	.w3(32'hbbf5cffc),
	.w4(32'hbc01110c),
	.w5(32'h3b2a52de),
	.w6(32'hbbc15a7a),
	.w7(32'hba8d5f00),
	.w8(32'h3ac6b16f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ab8a5),
	.w1(32'hbb0be0cd),
	.w2(32'h3a9bdf4a),
	.w3(32'hbb0cd41b),
	.w4(32'hbbe30c3e),
	.w5(32'h390d846f),
	.w6(32'h37ebe126),
	.w7(32'h3cace3d5),
	.w8(32'hbba6c711),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f8b198),
	.w1(32'hbb97651c),
	.w2(32'h3baca46c),
	.w3(32'hbbd82700),
	.w4(32'hbc32b31e),
	.w5(32'hbad73518),
	.w6(32'hbc6dfeb0),
	.w7(32'h3b4be4d2),
	.w8(32'h39ad3f6b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb59257),
	.w1(32'hba691fa3),
	.w2(32'hba9ae968),
	.w3(32'hbb9fbdf3),
	.w4(32'h3ab487e9),
	.w5(32'hbb00f941),
	.w6(32'hbc451566),
	.w7(32'hba81c68f),
	.w8(32'h3bdb4543),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32f215),
	.w1(32'hbc17a145),
	.w2(32'hbba3777d),
	.w3(32'hbac8957f),
	.w4(32'hbc082322),
	.w5(32'h3b0aebf1),
	.w6(32'h3be398e1),
	.w7(32'hbb599920),
	.w8(32'h3c0b7411),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc95f8),
	.w1(32'hbc3c7903),
	.w2(32'h3bb45a14),
	.w3(32'hbaaf934f),
	.w4(32'hbbbd6ff0),
	.w5(32'h39031b1c),
	.w6(32'h3baebfc8),
	.w7(32'h3b914ff4),
	.w8(32'hbb4f41a9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820a3a),
	.w1(32'h3c850de7),
	.w2(32'h3beeb851),
	.w3(32'hbb619044),
	.w4(32'hbbe86df7),
	.w5(32'h3bf95fc8),
	.w6(32'h3bfd0ec1),
	.w7(32'hbb82271b),
	.w8(32'h3a6cb54f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b424d97),
	.w1(32'h3c076068),
	.w2(32'h3beffa87),
	.w3(32'hbabb199a),
	.w4(32'h3b29acc6),
	.w5(32'hbc71e17c),
	.w6(32'h3c0f2904),
	.w7(32'hba265b11),
	.w8(32'h3c0effb8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bc6c5),
	.w1(32'h3ace9044),
	.w2(32'hbc0545e2),
	.w3(32'h3c3d4443),
	.w4(32'hb978cc3a),
	.w5(32'hba64c32f),
	.w6(32'hbaab76fd),
	.w7(32'hbb7312d1),
	.w8(32'h3c11468d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8213e9),
	.w1(32'hba8b5a70),
	.w2(32'hb588583a),
	.w3(32'hb935bd46),
	.w4(32'hbb7323ff),
	.w5(32'h3a236a14),
	.w6(32'h3be47e50),
	.w7(32'h3b9d3e38),
	.w8(32'h3939bf59),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae70b),
	.w1(32'hbb0af1d9),
	.w2(32'hbb963555),
	.w3(32'h3b4925c6),
	.w4(32'hbb743ee9),
	.w5(32'h3b99f878),
	.w6(32'hbb73ef22),
	.w7(32'h3a541d99),
	.w8(32'hbc18d45e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f159c),
	.w1(32'hbc8953fb),
	.w2(32'h3b31a6ca),
	.w3(32'h3c36a99f),
	.w4(32'h3c1dbc87),
	.w5(32'h3b7e9aa2),
	.w6(32'h3b1e623d),
	.w7(32'hbbd009cc),
	.w8(32'h3b39b516),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38805543),
	.w1(32'hbb07ad50),
	.w2(32'h3a9e5289),
	.w3(32'h3b8fbb52),
	.w4(32'h3a74962f),
	.w5(32'h3c05dd81),
	.w6(32'hbbf06f8d),
	.w7(32'hbb764b62),
	.w8(32'hba7b4777),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabd7b3),
	.w1(32'hbbac40b2),
	.w2(32'hbbd80fcc),
	.w3(32'hbba9bafe),
	.w4(32'hbb5ee3a7),
	.w5(32'hbab6ddc8),
	.w6(32'h3bacfa3c),
	.w7(32'hbb0b8609),
	.w8(32'h38c9cb12),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0936dc),
	.w1(32'hbb9b96fd),
	.w2(32'hbbca827f),
	.w3(32'hbc3b9ad5),
	.w4(32'hba80db63),
	.w5(32'hbb7ad73b),
	.w6(32'hbb1aaaa9),
	.w7(32'hba061bd3),
	.w8(32'hba995a0f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef1c79),
	.w1(32'hbb268c08),
	.w2(32'hbbab4efe),
	.w3(32'hb9d58b74),
	.w4(32'hbbdc0d8f),
	.w5(32'h393ad4e9),
	.w6(32'hb88cb51f),
	.w7(32'h3a992dab),
	.w8(32'hba25ed4b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c4e4e),
	.w1(32'h3c387560),
	.w2(32'hbc1cdd97),
	.w3(32'hbb8fdf7e),
	.w4(32'hbbfa2633),
	.w5(32'h3bbc4129),
	.w6(32'h3b7afd4b),
	.w7(32'hba1747d8),
	.w8(32'hbc1a27a4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba537610),
	.w1(32'hbb39c727),
	.w2(32'hb9f2b002),
	.w3(32'h3ba579aa),
	.w4(32'hbb0d794c),
	.w5(32'h3be7fbf5),
	.w6(32'h3b9921c1),
	.w7(32'h3d06bd04),
	.w8(32'h3b6b4623),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7449c),
	.w1(32'hba40ea82),
	.w2(32'hba837058),
	.w3(32'h3a5a6589),
	.w4(32'h3ac5877b),
	.w5(32'hbbcfd3dd),
	.w6(32'hbb084cf2),
	.w7(32'hbb6d4ee4),
	.w8(32'hbc371bf5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d5888),
	.w1(32'h3c81d3cc),
	.w2(32'h390be7dc),
	.w3(32'hbb1a947c),
	.w4(32'h3bb43212),
	.w5(32'hbb250478),
	.w6(32'hbb11f8f1),
	.w7(32'hb9c3889f),
	.w8(32'hb9b3284c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3aec72),
	.w1(32'h3ae71ea2),
	.w2(32'hbb10f33f),
	.w3(32'hba64c3bb),
	.w4(32'hba385ac0),
	.w5(32'h3ba1e09c),
	.w6(32'hb9b0700d),
	.w7(32'hbb401602),
	.w8(32'h3c816758),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5af40),
	.w1(32'hbb7c7091),
	.w2(32'h3acc2d66),
	.w3(32'h3bbfa244),
	.w4(32'hbab09928),
	.w5(32'hbbaff59c),
	.w6(32'hbb0ab4d6),
	.w7(32'hbb4dba29),
	.w8(32'h3a1bdb55),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b921b31),
	.w1(32'hbb58f34b),
	.w2(32'h3b6b5925),
	.w3(32'hbaaa88a0),
	.w4(32'h3bd1c769),
	.w5(32'hb99ae8c2),
	.w6(32'h3adf951f),
	.w7(32'h3cb0ce72),
	.w8(32'hbc0d0ffc),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c933387),
	.w1(32'h395853d0),
	.w2(32'hbb97c4b7),
	.w3(32'hbc384db7),
	.w4(32'h3c1a4ef4),
	.w5(32'h3aff8176),
	.w6(32'h3ae9cd28),
	.w7(32'hbc0c37f8),
	.w8(32'hbb225088),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fa502),
	.w1(32'hbb2c6ef5),
	.w2(32'hbbce590e),
	.w3(32'h3ba9bc6a),
	.w4(32'hbbc879d5),
	.w5(32'hbbfc0284),
	.w6(32'h3b94f9ab),
	.w7(32'hbb45976d),
	.w8(32'hb9a36d03),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18b94f),
	.w1(32'hbb2a71bb),
	.w2(32'hbc9f78aa),
	.w3(32'h3bdce247),
	.w4(32'hbb883bd1),
	.w5(32'hbb6847e7),
	.w6(32'h3a8e1d06),
	.w7(32'hbb14ae04),
	.w8(32'hb9821be2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf57870),
	.w1(32'h3a575cdc),
	.w2(32'hb9eed20a),
	.w3(32'hbb8785f6),
	.w4(32'h3c0e3e36),
	.w5(32'h3b925aaf),
	.w6(32'h3b53bc68),
	.w7(32'h3bb85aaa),
	.w8(32'h39ff53fc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd49b7d),
	.w1(32'hbbaa86f3),
	.w2(32'hb935d496),
	.w3(32'hbb879fcc),
	.w4(32'hb91f2e7c),
	.w5(32'h3b06e2c1),
	.w6(32'h3c694dcf),
	.w7(32'h3baf8ba2),
	.w8(32'hbc0f6662),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caca52e),
	.w1(32'hbbfe0be1),
	.w2(32'hbaa3f33f),
	.w3(32'hbcdce2eb),
	.w4(32'hbb21efba),
	.w5(32'hbc994719),
	.w6(32'h3b89f56d),
	.w7(32'hbc00905a),
	.w8(32'hbbb0c389),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c948d77),
	.w1(32'h3bbc6768),
	.w2(32'hbaa3cce5),
	.w3(32'h3c447078),
	.w4(32'hbb70ad59),
	.w5(32'hbbf59704),
	.w6(32'h3d571925),
	.w7(32'hbbbee11c),
	.w8(32'h398eacc9),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4846a0),
	.w1(32'hbb2bd0fa),
	.w2(32'hb9e707f0),
	.w3(32'h3b4d2fb9),
	.w4(32'h39fc6cdb),
	.w5(32'h3c1692a3),
	.w6(32'hbbd619c8),
	.w7(32'h3b20f005),
	.w8(32'h3b203990),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1bc14),
	.w1(32'hb9a1a18e),
	.w2(32'hbc319c6d),
	.w3(32'h3c363436),
	.w4(32'hbbd0e800),
	.w5(32'h3c32f04b),
	.w6(32'hbc7b0dcc),
	.w7(32'h39a2c42c),
	.w8(32'h3cb686c4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5a856),
	.w1(32'h3ba5e431),
	.w2(32'hbbc81106),
	.w3(32'h3ba20ac7),
	.w4(32'hbb837ee4),
	.w5(32'hbc643b0d),
	.w6(32'hba7d6846),
	.w7(32'h3ac6731c),
	.w8(32'h3b770333),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fda0e),
	.w1(32'hbbbfa664),
	.w2(32'hbb911f91),
	.w3(32'h3b8c5193),
	.w4(32'hbc523be7),
	.w5(32'hbc0d6914),
	.w6(32'h3cc80202),
	.w7(32'hbb1b0c1f),
	.w8(32'hbc24a507),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64b40d),
	.w1(32'hbac9abca),
	.w2(32'hbbe9350a),
	.w3(32'hbc7a1426),
	.w4(32'hbcfcc582),
	.w5(32'hbba0a5d0),
	.w6(32'hbb09edd3),
	.w7(32'hba8febd0),
	.w8(32'h3c652b89),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48f2b8),
	.w1(32'h3be3706e),
	.w2(32'hbc97e585),
	.w3(32'hbc0a5d85),
	.w4(32'hbb4712e7),
	.w5(32'hbbd4a3ae),
	.w6(32'hbc0615b9),
	.w7(32'h3b969824),
	.w8(32'hb8455b2a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922a19),
	.w1(32'hbba1ca9b),
	.w2(32'h3ab316bd),
	.w3(32'h3b9c59cc),
	.w4(32'hbb364ab8),
	.w5(32'h3c380589),
	.w6(32'h3d04bb4d),
	.w7(32'hbc00d6f8),
	.w8(32'hba05967f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba40526),
	.w1(32'h3b8083e0),
	.w2(32'h3ca421c0),
	.w3(32'hbbd63a0f),
	.w4(32'hbbb8e2ee),
	.w5(32'hbbf3d2e7),
	.w6(32'hbbb503aa),
	.w7(32'h3b649691),
	.w8(32'h3a206468),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8833d7),
	.w1(32'hbabe5d2d),
	.w2(32'h3bb03e53),
	.w3(32'h3b56e8c5),
	.w4(32'h3ba77fc8),
	.w5(32'hbc763016),
	.w6(32'h3d129371),
	.w7(32'hbd5249dd),
	.w8(32'hbbd0723d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392336cb),
	.w1(32'hbc65c541),
	.w2(32'hbb934df1),
	.w3(32'hbba995ea),
	.w4(32'h3b99a6ad),
	.w5(32'h3c241de9),
	.w6(32'hbcebe594),
	.w7(32'h3cb92d67),
	.w8(32'h3d03d59d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7fdfd),
	.w1(32'h3a3a9f06),
	.w2(32'h3c0c2f2a),
	.w3(32'hbb159e72),
	.w4(32'hbc405467),
	.w5(32'h3c353125),
	.w6(32'h3c3f25cd),
	.w7(32'hbbf348b2),
	.w8(32'hbb63c26d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7a170),
	.w1(32'hbba159b0),
	.w2(32'hbc809e46),
	.w3(32'h3bb0c6d3),
	.w4(32'h3a48af3c),
	.w5(32'hbc29eef0),
	.w6(32'h3bfbfcb7),
	.w7(32'hbc830997),
	.w8(32'hbb5fb66f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb507dcb),
	.w1(32'hbc1d15f0),
	.w2(32'hbbf9aaed),
	.w3(32'h3bb6e260),
	.w4(32'hbc2faa27),
	.w5(32'h3a1c0d9b),
	.w6(32'h3c10778d),
	.w7(32'hbb95e604),
	.w8(32'h3af48a0d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37048017),
	.w1(32'h3a51969b),
	.w2(32'hbc02ca8f),
	.w3(32'h3bd0d589),
	.w4(32'h3ac53ffd),
	.w5(32'h3c8363f9),
	.w6(32'hba4ca819),
	.w7(32'hbc200dec),
	.w8(32'hba232e12),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2e97e),
	.w1(32'h39e7b538),
	.w2(32'h3c47f2d1),
	.w3(32'hbb8997b4),
	.w4(32'hb92c4847),
	.w5(32'hbaece8db),
	.w6(32'h3af676f4),
	.w7(32'h3b2eca5e),
	.w8(32'hbbe2f85c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3da43f),
	.w1(32'hbba1796a),
	.w2(32'hbc0cdc41),
	.w3(32'hbb953787),
	.w4(32'hbb5ab81c),
	.w5(32'hba49d480),
	.w6(32'h390dbcd2),
	.w7(32'hbb8e8061),
	.w8(32'h3b2f90ca),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb5d2b),
	.w1(32'hbc0fadec),
	.w2(32'hbb043f0b),
	.w3(32'h3ba382aa),
	.w4(32'hbbc4f755),
	.w5(32'h3a404993),
	.w6(32'hbbd9b914),
	.w7(32'h3ccb6867),
	.w8(32'hbad3daaf),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cba16),
	.w1(32'hbbcc54b7),
	.w2(32'hba277dd6),
	.w3(32'hbc40ede4),
	.w4(32'h3cb1dc23),
	.w5(32'hbb386750),
	.w6(32'hbb50b847),
	.w7(32'h39f3c717),
	.w8(32'h3b98bd8b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6718351),
	.w1(32'h3b793b54),
	.w2(32'hbbca2b33),
	.w3(32'hba9549de),
	.w4(32'h3aee99c8),
	.w5(32'hba602180),
	.w6(32'hbb387ca2),
	.w7(32'h3a489154),
	.w8(32'hba6bc524),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed666e),
	.w1(32'h3bf5fcd3),
	.w2(32'h3b86b815),
	.w3(32'hbbc132d1),
	.w4(32'hbc47ae89),
	.w5(32'h3bbe144a),
	.w6(32'h3af93a0a),
	.w7(32'hbbf9cfa3),
	.w8(32'h3cce2ce1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fcbcf),
	.w1(32'hbb528992),
	.w2(32'h3c79ee0b),
	.w3(32'h3bb0ecd2),
	.w4(32'hbc1fc4ac),
	.w5(32'h3b925fe8),
	.w6(32'h3ba853de),
	.w7(32'h3bd20535),
	.w8(32'hbcb8dd9d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c0289),
	.w1(32'h3bb01d48),
	.w2(32'hbc7946a2),
	.w3(32'hbcb2c18d),
	.w4(32'h3b38db55),
	.w5(32'h3a93b6f4),
	.w6(32'hbacca57a),
	.w7(32'h3c21bf33),
	.w8(32'hbc7879ca),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade1d0c),
	.w1(32'hbc318a7a),
	.w2(32'hbc24ef36),
	.w3(32'h3bf4b944),
	.w4(32'hbc4eeaf8),
	.w5(32'hbc9edfaf),
	.w6(32'h3c80ef95),
	.w7(32'hbc3fcbc9),
	.w8(32'hbc3cfcbc),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b124bc4),
	.w1(32'h3b3d146b),
	.w2(32'h39c3d6e4),
	.w3(32'h3bd849b7),
	.w4(32'hbc32f1db),
	.w5(32'h3b5b4e92),
	.w6(32'hbc8160b7),
	.w7(32'hbc7660cb),
	.w8(32'hbb7b31bf),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd3b77),
	.w1(32'hbc05aeec),
	.w2(32'h3c80b307),
	.w3(32'hbc9e4779),
	.w4(32'h3b8ab635),
	.w5(32'hbc8243bb),
	.w6(32'h3b730de2),
	.w7(32'hbbbb77d9),
	.w8(32'h3a8618da),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule