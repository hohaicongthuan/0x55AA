module layer_10_featuremap_111(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a9e29),
	.w1(32'h3c192adb),
	.w2(32'h3cf495d0),
	.w3(32'hbbe2bee7),
	.w4(32'hbbb637c3),
	.w5(32'hbcc86883),
	.w6(32'hbb3bc035),
	.w7(32'hbc14784d),
	.w8(32'hbc6e758a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab3a28),
	.w1(32'h3bea905a),
	.w2(32'hba620bf3),
	.w3(32'hbb8e9ce5),
	.w4(32'hb9e760f8),
	.w5(32'hbbc4cd00),
	.w6(32'h3ae40651),
	.w7(32'h3b492921),
	.w8(32'hbb38f30c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba400170),
	.w1(32'hbb28b239),
	.w2(32'hbb6a4327),
	.w3(32'hbaf51a69),
	.w4(32'h3b9d3c36),
	.w5(32'h3c2160db),
	.w6(32'h3bad9d62),
	.w7(32'hba64dc14),
	.w8(32'hba591a6e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb207ded),
	.w1(32'h3bd463a5),
	.w2(32'hbc06e986),
	.w3(32'h3bd5eb16),
	.w4(32'hbc302f32),
	.w5(32'hbb9f1b61),
	.w6(32'hbc024de1),
	.w7(32'hba0efeb6),
	.w8(32'hbba8751c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f6b90),
	.w1(32'hbb2c9c71),
	.w2(32'hbc337716),
	.w3(32'hbc07ba33),
	.w4(32'h3bb812b4),
	.w5(32'hbc0f7db1),
	.w6(32'hbba0e5a3),
	.w7(32'h3c00e7ba),
	.w8(32'h3c8c3a65),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3479e0),
	.w1(32'h3bb4920d),
	.w2(32'h3b35eb1c),
	.w3(32'hbcac76fc),
	.w4(32'hbbb2f979),
	.w5(32'hbc8bf8c0),
	.w6(32'h3c16f80d),
	.w7(32'h3c265e20),
	.w8(32'h3c2aa256),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08be6b),
	.w1(32'h3b0e9e2f),
	.w2(32'hb994c35f),
	.w3(32'hbc46188a),
	.w4(32'h3a4fd258),
	.w5(32'hbc59e907),
	.w6(32'h3a5acb0a),
	.w7(32'h3a848e8f),
	.w8(32'hbbcc83e8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49e3b4),
	.w1(32'hbc9be2de),
	.w2(32'hbc0ae16b),
	.w3(32'hbc000180),
	.w4(32'hbb313218),
	.w5(32'h3c11b3e7),
	.w6(32'hbc9d4084),
	.w7(32'hbb996faa),
	.w8(32'h3aab31fb),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b269b),
	.w1(32'h3b7b4a7a),
	.w2(32'h3a92b418),
	.w3(32'h3a501b3f),
	.w4(32'h3b844ce2),
	.w5(32'h3b046322),
	.w6(32'h3bf403b8),
	.w7(32'h3a9f1375),
	.w8(32'h3a8d10ff),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23ab9d),
	.w1(32'hbc1d6b37),
	.w2(32'hbc4aa0fc),
	.w3(32'h3acad268),
	.w4(32'hbbaa7766),
	.w5(32'hbc31ead5),
	.w6(32'hba364a54),
	.w7(32'h3c00d951),
	.w8(32'hbb96943c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bdd86),
	.w1(32'h3c632015),
	.w2(32'hbbacef76),
	.w3(32'hbb3bfe8a),
	.w4(32'h3ad4912c),
	.w5(32'h3b1d6112),
	.w6(32'h3c43ee92),
	.w7(32'h3c10d364),
	.w8(32'h3c06866c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0540e6),
	.w1(32'hbcb94daf),
	.w2(32'hbcbedf9b),
	.w3(32'h3c0e6e3b),
	.w4(32'hbc877c08),
	.w5(32'hbc77e53c),
	.w6(32'hbcbf6c19),
	.w7(32'hbcba032d),
	.w8(32'hbcdf6433),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1a0405),
	.w1(32'hbbf9224a),
	.w2(32'hba9e9b07),
	.w3(32'hbcbcaee0),
	.w4(32'h3b8c7571),
	.w5(32'hbab4597f),
	.w6(32'hbb44b0eb),
	.w7(32'hbba46d65),
	.w8(32'hbb8c0370),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6c09a),
	.w1(32'hbc731ad9),
	.w2(32'hb918cc89),
	.w3(32'hbadb179c),
	.w4(32'h3b8f12af),
	.w5(32'h3d21fd9d),
	.w6(32'hbce0f640),
	.w7(32'hbd165a47),
	.w8(32'hbc9dee53),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc22f33),
	.w1(32'hbb8d410c),
	.w2(32'hbd0daa8c),
	.w3(32'h3c780249),
	.w4(32'hbc4f91b0),
	.w5(32'h3a9ba125),
	.w6(32'hbc18031f),
	.w7(32'h3981d693),
	.w8(32'hbc288bab),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad11e7),
	.w1(32'h3b6f76ff),
	.w2(32'h3b84c1fa),
	.w3(32'hbcce9a72),
	.w4(32'hbb02c3d1),
	.w5(32'h3ae0e4b3),
	.w6(32'h3c397ea4),
	.w7(32'h3b51cef8),
	.w8(32'h3b3f5b64),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28c18c),
	.w1(32'hbb031141),
	.w2(32'h3a333268),
	.w3(32'hbb7aaea5),
	.w4(32'hbb4ad87d),
	.w5(32'hbb7132a6),
	.w6(32'h3bbafb44),
	.w7(32'h3acccac7),
	.w8(32'h3bcbefff),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda69dd),
	.w1(32'hbbcb86d0),
	.w2(32'hbb317c17),
	.w3(32'hbba9b03f),
	.w4(32'hbb7725a0),
	.w5(32'hbc0d4abf),
	.w6(32'h3b5a58fa),
	.w7(32'h3c4faa25),
	.w8(32'h39df204f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb511e4b),
	.w1(32'hbb03b12c),
	.w2(32'hba3e1a70),
	.w3(32'h3b867335),
	.w4(32'hbab72240),
	.w5(32'hbb0a076b),
	.w6(32'h3b9add22),
	.w7(32'h3b55cbc0),
	.w8(32'hb948825f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5276a),
	.w1(32'h3b2ad482),
	.w2(32'hba9a9bfc),
	.w3(32'hba7921e4),
	.w4(32'h3b312ede),
	.w5(32'hb9649a6c),
	.w6(32'h3b410935),
	.w7(32'h39903151),
	.w8(32'hb9de5525),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20584f),
	.w1(32'hbb01bbc7),
	.w2(32'hbb308695),
	.w3(32'hbb277daf),
	.w4(32'h3bbd031f),
	.w5(32'h3bfb0bd0),
	.w6(32'hbb9fe991),
	.w7(32'hbc0c8761),
	.w8(32'hbbb41149),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad01665),
	.w1(32'hbd0bb536),
	.w2(32'hbce3b88d),
	.w3(32'h3b4d5c78),
	.w4(32'hbbd1693b),
	.w5(32'hbc0403de),
	.w6(32'hbc757ae9),
	.w7(32'hbc7f4713),
	.w8(32'hbc68b902),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd973219),
	.w1(32'hbb86be0b),
	.w2(32'hbb71abc2),
	.w3(32'hbc79c72f),
	.w4(32'h3c7043ae),
	.w5(32'hbb2f353a),
	.w6(32'h3b9974d2),
	.w7(32'hbb2f2713),
	.w8(32'h3b26e7cf),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf74e5),
	.w1(32'hbb57bbe5),
	.w2(32'h399803b7),
	.w3(32'h3b0dc7e3),
	.w4(32'h3b58a6bd),
	.w5(32'h3be9e940),
	.w6(32'hb9d2c35f),
	.w7(32'hbbafb610),
	.w8(32'hb9c9942e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09d943),
	.w1(32'h3c7d8ca0),
	.w2(32'hbaa0052f),
	.w3(32'h3b46d4f3),
	.w4(32'hbc048544),
	.w5(32'hbc0ecf0b),
	.w6(32'hb9bf3da1),
	.w7(32'hbb05db3a),
	.w8(32'hbbc0e8dc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1e087),
	.w1(32'hbc46940d),
	.w2(32'hbcb1aa68),
	.w3(32'hbbb2fe47),
	.w4(32'hbb816d4e),
	.w5(32'hbb0d8650),
	.w6(32'hbb30c8eb),
	.w7(32'hbc169751),
	.w8(32'hbbf5d487),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5aefb6),
	.w1(32'h3b2062cb),
	.w2(32'h3a6fffc4),
	.w3(32'hbb80fadf),
	.w4(32'h3b859f88),
	.w5(32'h3b2558cf),
	.w6(32'h3a75f51c),
	.w7(32'hbaa2522f),
	.w8(32'h3a405251),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb10333),
	.w1(32'hbb26923f),
	.w2(32'hbbe1bb36),
	.w3(32'h3b316976),
	.w4(32'hbcb37e32),
	.w5(32'hbc798acf),
	.w6(32'h3c0d9be3),
	.w7(32'h3c37a8b1),
	.w8(32'h3b469e8e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba242d3c),
	.w1(32'h39f87a54),
	.w2(32'hbb1967b3),
	.w3(32'hbbe33ed1),
	.w4(32'h3ac89406),
	.w5(32'h3a26285e),
	.w6(32'h3c0ae4ab),
	.w7(32'h3bf6cfc2),
	.w8(32'h3b9e6411),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12ef20),
	.w1(32'h3c3b9071),
	.w2(32'h3a007437),
	.w3(32'h3b74f754),
	.w4(32'hbc08fb13),
	.w5(32'hbb977213),
	.w6(32'h3bb087b2),
	.w7(32'hbc1e8b45),
	.w8(32'hbbe3d7c7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7bf35),
	.w1(32'h3aad6fb1),
	.w2(32'h3b4ade82),
	.w3(32'hbadd8580),
	.w4(32'h3b8e919b),
	.w5(32'h3b84ad60),
	.w6(32'hbb070af6),
	.w7(32'hbb804280),
	.w8(32'hb9dfcaa3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b562a9b),
	.w1(32'hb94fb2d7),
	.w2(32'hbab83be7),
	.w3(32'h3b4027b2),
	.w4(32'h3b47abaa),
	.w5(32'h3a243ca3),
	.w6(32'hb7ff1d07),
	.w7(32'hbb747309),
	.w8(32'hba197997),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85ef6b),
	.w1(32'hbb0a6414),
	.w2(32'h3b90965a),
	.w3(32'h3b376a4f),
	.w4(32'h38550964),
	.w5(32'h3c59b9f9),
	.w6(32'hbb8ed3b9),
	.w7(32'h3bc72fff),
	.w8(32'h3b2b8929),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddee94),
	.w1(32'h3bcee6b3),
	.w2(32'hbbb60a24),
	.w3(32'h3c44af46),
	.w4(32'h3bb82449),
	.w5(32'hbb878723),
	.w6(32'h3b8b520a),
	.w7(32'hbb44e431),
	.w8(32'h3a918043),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad76510),
	.w1(32'h3a9cf7be),
	.w2(32'hbbe2dc26),
	.w3(32'hb9f3792c),
	.w4(32'hbbb904d8),
	.w5(32'hbc8e5519),
	.w6(32'h3ab4b2b2),
	.w7(32'h3c02cf8c),
	.w8(32'hbb8c98df),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb750c9f),
	.w1(32'hbbcac123),
	.w2(32'hbbb381af),
	.w3(32'hbc470e04),
	.w4(32'h3a1b18f9),
	.w5(32'hbb5eede7),
	.w6(32'hbb0f80c3),
	.w7(32'hbb05d0b2),
	.w8(32'h3a53dcd0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b416fe1),
	.w1(32'hbc465bd4),
	.w2(32'hbc79d065),
	.w3(32'hbbfc6af6),
	.w4(32'h3ba31da7),
	.w5(32'hba3ad77c),
	.w6(32'hbb77de75),
	.w7(32'h3ca344f2),
	.w8(32'h3b6507a5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c2708),
	.w1(32'h3bd66197),
	.w2(32'h3b17c881),
	.w3(32'hbc43b125),
	.w4(32'hbbd52ce5),
	.w5(32'h3a868e15),
	.w6(32'hbb80bfcf),
	.w7(32'hbbd10eff),
	.w8(32'h3b0b462c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083980),
	.w1(32'h3c39fd28),
	.w2(32'h3ad9cfe2),
	.w3(32'h3bd474f3),
	.w4(32'hbbb5e831),
	.w5(32'hbba6a52e),
	.w6(32'h3c33a1cd),
	.w7(32'hbbfcae0e),
	.w8(32'hbbc6ad25),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b2078),
	.w1(32'h3b5582eb),
	.w2(32'hbaa03bd0),
	.w3(32'hbb49dc4f),
	.w4(32'h3960fa9f),
	.w5(32'hbb0e556a),
	.w6(32'h3ad66887),
	.w7(32'h3b1e7b74),
	.w8(32'h3b397f13),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af45944),
	.w1(32'hbb5afd6d),
	.w2(32'hbb9bc8e0),
	.w3(32'hbb8474a0),
	.w4(32'h3a272e65),
	.w5(32'h391e0eea),
	.w6(32'hbb8db2f8),
	.w7(32'hbc1ba364),
	.w8(32'hbb4f7608),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75b236),
	.w1(32'hbb5d9659),
	.w2(32'hbbe239de),
	.w3(32'hbb14d8a4),
	.w4(32'hbb2df4c3),
	.w5(32'h3b0fdc00),
	.w6(32'hbbc0a592),
	.w7(32'hbb9da1e6),
	.w8(32'hbba05200),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb0773),
	.w1(32'hba8002f1),
	.w2(32'hb887ebae),
	.w3(32'hbb4542aa),
	.w4(32'h3baaedb5),
	.w5(32'h3ba36d09),
	.w6(32'hbb72df69),
	.w7(32'hbbb9bd05),
	.w8(32'hbb93785e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd6c7b0),
	.w1(32'hbb67f468),
	.w2(32'h3a802c3e),
	.w3(32'h3b0ab994),
	.w4(32'hba87f809),
	.w5(32'hbbffb180),
	.w6(32'h3c6a215f),
	.w7(32'h3c8ffc0f),
	.w8(32'h3bc49d1e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf39b1b),
	.w1(32'hb90e55e1),
	.w2(32'h3cd5a58d),
	.w3(32'h389f516f),
	.w4(32'h3aa0fe55),
	.w5(32'h3c9dd3d2),
	.w6(32'hbb8dd5c1),
	.w7(32'hbbd15d21),
	.w8(32'hba4cac20),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc75c2),
	.w1(32'hba14d5ce),
	.w2(32'h3c42e8b1),
	.w3(32'h3c8e60ef),
	.w4(32'h3c0639de),
	.w5(32'h3c1fafdf),
	.w6(32'hbba265d1),
	.w7(32'hbbe65f35),
	.w8(32'hbace8614),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccd8f3),
	.w1(32'hbc0bcd12),
	.w2(32'hbce471aa),
	.w3(32'h3aa5b863),
	.w4(32'hbc5c3d81),
	.w5(32'h3aa9cc1a),
	.w6(32'hbbf24f42),
	.w7(32'h3b5838c0),
	.w8(32'hbbf99305),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7d0e4),
	.w1(32'hbc027dca),
	.w2(32'h3a410a70),
	.w3(32'hbc684801),
	.w4(32'hb8588360),
	.w5(32'h3b1ec563),
	.w6(32'h3bb9fb0e),
	.w7(32'h3c215ad4),
	.w8(32'h3a6bea65),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7ea08),
	.w1(32'hbabf4545),
	.w2(32'hbb2cc9b7),
	.w3(32'h3968e58e),
	.w4(32'h3ac36cdd),
	.w5(32'hbae3a397),
	.w6(32'hbaa976e6),
	.w7(32'hbba0e702),
	.w8(32'hbb01b090),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bfa88),
	.w1(32'hbb58a589),
	.w2(32'h3b84875f),
	.w3(32'hb9e38279),
	.w4(32'h3b836b96),
	.w5(32'h3c771abd),
	.w6(32'hbbd08aff),
	.w7(32'hbc4cb47d),
	.w8(32'hbbb2cd3b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bf4e0),
	.w1(32'hbb9298a7),
	.w2(32'hbb2f059c),
	.w3(32'h3bbf8a49),
	.w4(32'h3bf48116),
	.w5(32'h3ce15046),
	.w6(32'hbc1bad38),
	.w7(32'hbc8935f1),
	.w8(32'hbc3ffd79),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70a3ee),
	.w1(32'h3af30685),
	.w2(32'hbcd6440e),
	.w3(32'h3b2416bc),
	.w4(32'hbc91ffaf),
	.w5(32'hbcd89d29),
	.w6(32'h3c4937b5),
	.w7(32'h3b8cb6d9),
	.w8(32'hbcae176c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd0633),
	.w1(32'h3c3bdfaf),
	.w2(32'h3c16f463),
	.w3(32'hbc2ffe98),
	.w4(32'h3b2c4765),
	.w5(32'hbc407763),
	.w6(32'h3c31e2f9),
	.w7(32'h3c6ddb58),
	.w8(32'h3ab84e85),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47367b),
	.w1(32'hbc57d941),
	.w2(32'hbc0b4963),
	.w3(32'hbc2eea06),
	.w4(32'hbc6914c5),
	.w5(32'hbcc45580),
	.w6(32'h3b397d7f),
	.w7(32'h3c89ca4d),
	.w8(32'h3bd50c6f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8995ce),
	.w1(32'hb83e2e77),
	.w2(32'hbb18b52e),
	.w3(32'hbc531027),
	.w4(32'hbb8bf8f2),
	.w5(32'hbc04df92),
	.w6(32'h3bc4c1f5),
	.w7(32'h3c143379),
	.w8(32'h3abc243b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9295a57),
	.w1(32'hbbe74a41),
	.w2(32'hbbf9b5d7),
	.w3(32'hbbc8f894),
	.w4(32'h3b126e05),
	.w5(32'h3b1b0d4c),
	.w6(32'hbb66f1d1),
	.w7(32'hbc16c673),
	.w8(32'hbb34bc58),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b8e46),
	.w1(32'hbae2a7d8),
	.w2(32'h3c049bf7),
	.w3(32'h3b31c4f7),
	.w4(32'h3c0b720e),
	.w5(32'h3cc159da),
	.w6(32'hbc095c46),
	.w7(32'hbc8c58e2),
	.w8(32'hbc339a3f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74316f9),
	.w1(32'hbae44bb0),
	.w2(32'hbc9c6ccf),
	.w3(32'h3c065a9e),
	.w4(32'hbae97ec5),
	.w5(32'h3b998803),
	.w6(32'hbc4af806),
	.w7(32'hbce329e6),
	.w8(32'hbbeac94c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba925b3),
	.w1(32'h3bb84334),
	.w2(32'hba53a751),
	.w3(32'hbc7e31e0),
	.w4(32'h3b189ffa),
	.w5(32'hbbd0753e),
	.w6(32'h3b7c28a1),
	.w7(32'h3b99818d),
	.w8(32'hbb02fbd2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da6551),
	.w1(32'h3a686334),
	.w2(32'h3b326444),
	.w3(32'h3a2a879e),
	.w4(32'h3abc8989),
	.w5(32'h3ac3e92c),
	.w6(32'h3ac9d8f0),
	.w7(32'hbbabac63),
	.w8(32'hbaa3f820),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bd44d),
	.w1(32'h3a62e1cd),
	.w2(32'h3aaa8291),
	.w3(32'hbace0615),
	.w4(32'h3b3b7ea2),
	.w5(32'hb9e4decd),
	.w6(32'h3bb04d38),
	.w7(32'h3bb68ff8),
	.w8(32'h3b05c6c5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68cf80),
	.w1(32'h3bbf75f7),
	.w2(32'h3cbfb115),
	.w3(32'hbaa21f7a),
	.w4(32'h3b4ed4ae),
	.w5(32'h3c1530bc),
	.w6(32'h3b9d516a),
	.w7(32'hbc0c0616),
	.w8(32'h39eb0bb1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0f149),
	.w1(32'h3b9f7dd3),
	.w2(32'h3b78ff45),
	.w3(32'h3bebab26),
	.w4(32'h3aa46f37),
	.w5(32'h3bca4a56),
	.w6(32'h3951b616),
	.w7(32'h3a15cf96),
	.w8(32'h3bae7ff4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7ef72),
	.w1(32'h3b156871),
	.w2(32'hbb06ef32),
	.w3(32'h3989b66f),
	.w4(32'hba62d801),
	.w5(32'hbc032d15),
	.w6(32'h3bcfd130),
	.w7(32'h3c52c43a),
	.w8(32'h3b5969fe),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23f4f5),
	.w1(32'h3bae678d),
	.w2(32'h3b901b60),
	.w3(32'hbb461bef),
	.w4(32'h3af7c47b),
	.w5(32'hba8d918a),
	.w6(32'h3c027749),
	.w7(32'h3bf95f52),
	.w8(32'h3a6bf8ad),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac69e70),
	.w1(32'h3a3a3290),
	.w2(32'hbbf98fc9),
	.w3(32'h39d7618d),
	.w4(32'h3b85b906),
	.w5(32'h3bf53bae),
	.w6(32'hbc300b00),
	.w7(32'hbca4a9c1),
	.w8(32'hbb9efe55),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc990729),
	.w1(32'hbc5648df),
	.w2(32'h3b5b93d7),
	.w3(32'hbc24811a),
	.w4(32'hbc2f7d43),
	.w5(32'h390cdafe),
	.w6(32'hbc2d4540),
	.w7(32'hbc24de69),
	.w8(32'hbc6a786f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f2aca),
	.w1(32'h3b2ec2ca),
	.w2(32'hbb43691a),
	.w3(32'hbb934603),
	.w4(32'h3be14939),
	.w5(32'h3b2a0225),
	.w6(32'hb98b816f),
	.w7(32'h3ab7e457),
	.w8(32'h3c07aaf6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2924c1),
	.w1(32'h3b68d19f),
	.w2(32'h3aee7f9a),
	.w3(32'hba991902),
	.w4(32'h3bb6122d),
	.w5(32'hbb9fd206),
	.w6(32'h3be717ff),
	.w7(32'h398ca841),
	.w8(32'hbacb1257),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf30795),
	.w1(32'h3c22a72a),
	.w2(32'hba5a6543),
	.w3(32'hbbbd7c1e),
	.w4(32'h3c4eedbb),
	.w5(32'h3d241f1f),
	.w6(32'hbcc410f5),
	.w7(32'hbd1809c0),
	.w8(32'hbc76950e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53ed42),
	.w1(32'h3b663ef4),
	.w2(32'hbaec4c71),
	.w3(32'h3b417f14),
	.w4(32'hbaa040f6),
	.w5(32'hbbeb5ea4),
	.w6(32'h3a5ce0a6),
	.w7(32'h3b8ddf6a),
	.w8(32'hba6d6002),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dfc606),
	.w1(32'h3ab278b7),
	.w2(32'h3b0dc251),
	.w3(32'h39f9b9f0),
	.w4(32'h3b25bd1e),
	.w5(32'h3b8970c1),
	.w6(32'hb985ac23),
	.w7(32'hbb5c9183),
	.w8(32'h3a929fd2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983c41a),
	.w1(32'h39b9fcb2),
	.w2(32'hbab1be60),
	.w3(32'hbba62624),
	.w4(32'h390bede9),
	.w5(32'h39ecc3f3),
	.w6(32'h3b0938b4),
	.w7(32'hbad89719),
	.w8(32'h38d10f34),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d164d),
	.w1(32'hbb38c715),
	.w2(32'hbb861307),
	.w3(32'hba54c574),
	.w4(32'h399161c2),
	.w5(32'hba1e57d0),
	.w6(32'hba0ce5bc),
	.w7(32'hbb841be8),
	.w8(32'hbb168ac2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d70da),
	.w1(32'h3bb556b2),
	.w2(32'hbad889b6),
	.w3(32'h3b5d2f76),
	.w4(32'hba53fa76),
	.w5(32'hbb987a2d),
	.w6(32'h3c023c4a),
	.w7(32'h3c206abb),
	.w8(32'hbb131fae),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e208a),
	.w1(32'hbc8c058e),
	.w2(32'hbc9647c8),
	.w3(32'hbae35a80),
	.w4(32'hbbf3ea9a),
	.w5(32'h3caed4c4),
	.w6(32'hbd05662a),
	.w7(32'hbc7d9910),
	.w8(32'hbc9e9aaa),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3ebaf),
	.w1(32'hbc63d1fc),
	.w2(32'h3af8c672),
	.w3(32'hbc8e28ac),
	.w4(32'h3bb1879c),
	.w5(32'h3c7e13db),
	.w6(32'hbc2464bc),
	.w7(32'hbbe16ea9),
	.w8(32'hb9ea5891),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86b88f),
	.w1(32'h3c079cc2),
	.w2(32'h3ba38414),
	.w3(32'h3b89b7fc),
	.w4(32'hbaac298a),
	.w5(32'h3be85d1c),
	.w6(32'h3bbeb846),
	.w7(32'hbad2fb10),
	.w8(32'h3a770f8e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56e99d),
	.w1(32'hbc0389e4),
	.w2(32'hbbd1b301),
	.w3(32'h3bb93d09),
	.w4(32'hbc05cffb),
	.w5(32'hbb8ff562),
	.w6(32'h3bd6bcea),
	.w7(32'h3b8bfda6),
	.w8(32'hb94b20b6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb894183),
	.w1(32'hbb9e508e),
	.w2(32'h3babc8e7),
	.w3(32'hba1b349d),
	.w4(32'h3baa6b50),
	.w5(32'h3bff1f74),
	.w6(32'hbb87962b),
	.w7(32'hbbeabbd2),
	.w8(32'hbb4e727b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1fe9f),
	.w1(32'hbb25e6ae),
	.w2(32'hbbadb326),
	.w3(32'h3b595de2),
	.w4(32'h39a0a857),
	.w5(32'hbb889abf),
	.w6(32'h3ae2b5a1),
	.w7(32'hbbc773ab),
	.w8(32'hbb12bb7f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896521),
	.w1(32'h3b2435e7),
	.w2(32'h3ad0797d),
	.w3(32'hba77f849),
	.w4(32'h3c0cac95),
	.w5(32'hbbcb33f4),
	.w6(32'h3acdcee3),
	.w7(32'h3bd6d43e),
	.w8(32'hbb161602),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79788a),
	.w1(32'h3b44bfe6),
	.w2(32'h378d0ac0),
	.w3(32'h3b04bd9e),
	.w4(32'hbb11161d),
	.w5(32'hbb81a24f),
	.w6(32'hba3711c4),
	.w7(32'hbaec594e),
	.w8(32'hbbd6a22e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e23144),
	.w1(32'h3bbd255d),
	.w2(32'h3bc03f4e),
	.w3(32'hbb876529),
	.w4(32'h3988527e),
	.w5(32'hbbb13982),
	.w6(32'h3b7c6f15),
	.w7(32'h3b5ecc14),
	.w8(32'hbb24ffa1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f34f7),
	.w1(32'h3bc42370),
	.w2(32'h39990055),
	.w3(32'h3b1ecfa9),
	.w4(32'hbc00fbdc),
	.w5(32'hbb95f258),
	.w6(32'h3ba78153),
	.w7(32'hb8d308a8),
	.w8(32'h391554ee),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79d52d),
	.w1(32'h3b4255ef),
	.w2(32'h3bbfb0bb),
	.w3(32'hbbeb6fa9),
	.w4(32'h3ae78608),
	.w5(32'h3b846bea),
	.w6(32'hb9a6a56f),
	.w7(32'hbb8bf3ba),
	.w8(32'hba9f1037),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc65ac),
	.w1(32'hbbf4e8e9),
	.w2(32'hbc5ab616),
	.w3(32'h3acc95a4),
	.w4(32'hbabce6ce),
	.w5(32'h3cc62ff0),
	.w6(32'hbcbce615),
	.w7(32'hbce24477),
	.w8(32'hbc86dc45),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc121be3),
	.w1(32'h3abcd947),
	.w2(32'h3b01ad7e),
	.w3(32'h3bedc3cb),
	.w4(32'h3b92725e),
	.w5(32'h3b77b84b),
	.w6(32'hbaff5908),
	.w7(32'hbb96c486),
	.w8(32'hba398f3e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83d0c9),
	.w1(32'h3b7e96c2),
	.w2(32'hb813db28),
	.w3(32'h3b1a6e3b),
	.w4(32'hbb1d3d5e),
	.w5(32'hbc01ad21),
	.w6(32'h3bc9cc09),
	.w7(32'h3c0ae2d3),
	.w8(32'h3b8554e8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd56822),
	.w1(32'hbbdb9aea),
	.w2(32'hbb15647a),
	.w3(32'hbc042950),
	.w4(32'h3bf2b5d3),
	.w5(32'h3b69747f),
	.w6(32'hbb5829f8),
	.w7(32'hbb9fb5e8),
	.w8(32'hbb809f3f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ca6b1),
	.w1(32'h3af24465),
	.w2(32'h3962b9ee),
	.w3(32'h3b704205),
	.w4(32'h3a80891e),
	.w5(32'h3a8fab1e),
	.w6(32'h3acddc2c),
	.w7(32'hbbc2b149),
	.w8(32'hbb991b18),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88f07d),
	.w1(32'hbb7e255e),
	.w2(32'h3bd94087),
	.w3(32'h3af321e4),
	.w4(32'h3c9f0b5e),
	.w5(32'h3c535cd7),
	.w6(32'h3b184c1c),
	.w7(32'h3b52a08a),
	.w8(32'hb8d212ff),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4068b),
	.w1(32'h3bb6e829),
	.w2(32'h3b944b60),
	.w3(32'h3c3c60f3),
	.w4(32'hbb38b75e),
	.w5(32'hbc797950),
	.w6(32'h3c04c762),
	.w7(32'h3c1a226c),
	.w8(32'h3a194ff2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc536230),
	.w1(32'hbc38bb39),
	.w2(32'hbc11486c),
	.w3(32'hbb8aeeab),
	.w4(32'h3a92024d),
	.w5(32'hbb717d8d),
	.w6(32'h3b1a6da1),
	.w7(32'hbbd940a9),
	.w8(32'h3859a999),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecdfae),
	.w1(32'hb9d4eb6f),
	.w2(32'hbb92b56c),
	.w3(32'h3a148b11),
	.w4(32'h3b0cb34d),
	.w5(32'h3bb588cf),
	.w6(32'h3b98a697),
	.w7(32'hba5a87a7),
	.w8(32'hbb5adf02),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a143ccb),
	.w1(32'hbafe5e62),
	.w2(32'h3c7d2deb),
	.w3(32'h3a79e987),
	.w4(32'hbc6c20ba),
	.w5(32'hbc8f8406),
	.w6(32'hb86f0a47),
	.w7(32'hbc42a0dc),
	.w8(32'hbb83350b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b710407),
	.w1(32'hb8410011),
	.w2(32'h398ba015),
	.w3(32'hbaca64dc),
	.w4(32'h3ae89503),
	.w5(32'h3b123e95),
	.w6(32'hbba1d4fc),
	.w7(32'hbba9bbcc),
	.w8(32'hbad7f672),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdd152),
	.w1(32'h3a11f942),
	.w2(32'h39dde0be),
	.w3(32'hba2c4326),
	.w4(32'hbb598725),
	.w5(32'hbca69fcf),
	.w6(32'h3c5be7cb),
	.w7(32'h3cf643c0),
	.w8(32'h3c38ebb1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe26b3),
	.w1(32'h3b659995),
	.w2(32'h3c85aeb6),
	.w3(32'h3b1fd1bb),
	.w4(32'h3c645758),
	.w5(32'h3b11af78),
	.w6(32'h3bfd701a),
	.w7(32'h3c7c3863),
	.w8(32'h3bb9c000),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cccb8),
	.w1(32'h3a589a66),
	.w2(32'hbc0286d5),
	.w3(32'hbc91f4fa),
	.w4(32'hbb03b62c),
	.w5(32'hbcae5b65),
	.w6(32'h3ba6b64e),
	.w7(32'h3c8be836),
	.w8(32'h3c1efd39),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b212),
	.w1(32'h3a8a77f3),
	.w2(32'hbc2ac530),
	.w3(32'hbcabbec8),
	.w4(32'h3c27505c),
	.w5(32'h3d045c79),
	.w6(32'hbb9f8957),
	.w7(32'hbc9ebba3),
	.w8(32'hbbc48740),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c43a6),
	.w1(32'hbb367937),
	.w2(32'h3c8a1ac0),
	.w3(32'h3ba94a4c),
	.w4(32'hbb81b88e),
	.w5(32'hbcd78947),
	.w6(32'hbbbd02b2),
	.w7(32'hbbfa055b),
	.w8(32'hbad4c081),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c0f6a),
	.w1(32'hbc88a880),
	.w2(32'h3c3befc9),
	.w3(32'hbcf9a352),
	.w4(32'h3ca99775),
	.w5(32'h3ce07291),
	.w6(32'hbbe10b99),
	.w7(32'hbbd76311),
	.w8(32'hbb665bab),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb121ea3),
	.w1(32'h3996b197),
	.w2(32'hba5ff549),
	.w3(32'h3c025b79),
	.w4(32'h3b116f05),
	.w5(32'h3bb7a4a6),
	.w6(32'h388259e2),
	.w7(32'hbb097436),
	.w8(32'h3b296291),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3aaaa8),
	.w1(32'hbc874805),
	.w2(32'hbc606b70),
	.w3(32'hbc89b022),
	.w4(32'h3bbb9749),
	.w5(32'h3c5adbed),
	.w6(32'hbc06b098),
	.w7(32'hbb2993ad),
	.w8(32'h3ae9a475),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7d77a),
	.w1(32'hbbc34438),
	.w2(32'hbbc0a859),
	.w3(32'h3b9fa215),
	.w4(32'h3b9f3a1f),
	.w5(32'h3aa7024a),
	.w6(32'hbafac0f1),
	.w7(32'hbaf0d8f4),
	.w8(32'hbae45343),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a871257),
	.w1(32'h3b1a8e98),
	.w2(32'h39b18512),
	.w3(32'h3b75c26c),
	.w4(32'h3ba59a0a),
	.w5(32'h3bbad400),
	.w6(32'h3bdae4f8),
	.w7(32'h3b83e234),
	.w8(32'h3aae2f85),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6a62e),
	.w1(32'h3b1fa56f),
	.w2(32'h3b342272),
	.w3(32'h3b0d0981),
	.w4(32'h3b907718),
	.w5(32'h3b86be5c),
	.w6(32'hbb9e5939),
	.w7(32'hbbf6e6cd),
	.w8(32'hbb286702),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84cbba),
	.w1(32'hbb8b4b59),
	.w2(32'h3be25a35),
	.w3(32'h3bd5ea91),
	.w4(32'h3be95d94),
	.w5(32'h3c5ac1fa),
	.w6(32'hb9af26fb),
	.w7(32'hbb8899bc),
	.w8(32'h3958a3f1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba051ef5),
	.w1(32'hbbe9c5fd),
	.w2(32'hbab1d337),
	.w3(32'h3b949662),
	.w4(32'hbb8686bb),
	.w5(32'h3c5d9212),
	.w6(32'hbbbb45f5),
	.w7(32'hbc5a1d43),
	.w8(32'hbbf1b699),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca4efe),
	.w1(32'hba31a68e),
	.w2(32'hbc372a1e),
	.w3(32'h3c24d18b),
	.w4(32'hbbf37540),
	.w5(32'hbc193b07),
	.w6(32'h3c230b6e),
	.w7(32'hba7f33bd),
	.w8(32'hbbdf611e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc101dbc),
	.w1(32'hb7a87656),
	.w2(32'hbbcf3ec4),
	.w3(32'hbbb060dc),
	.w4(32'hbc2024b9),
	.w5(32'h3a61fca0),
	.w6(32'hbc1b1c2f),
	.w7(32'hbcc8de89),
	.w8(32'hbcc526a5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b644b),
	.w1(32'h3c06e20d),
	.w2(32'hbb2878c6),
	.w3(32'hbb840402),
	.w4(32'hba169264),
	.w5(32'hbaef163f),
	.w6(32'h3b5aa202),
	.w7(32'h3c1552a4),
	.w8(32'h3c18dedc),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86c369),
	.w1(32'hbb3b8eb5),
	.w2(32'hbc11ab41),
	.w3(32'hbc70edae),
	.w4(32'h3a5e4b71),
	.w5(32'h3bddd521),
	.w6(32'hbba65ec6),
	.w7(32'hbc47f79b),
	.w8(32'hbb9cce4a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89beec),
	.w1(32'hbbf9172d),
	.w2(32'h3b01736e),
	.w3(32'h38f67d58),
	.w4(32'h3b3bf967),
	.w5(32'h3cb3a1a3),
	.w6(32'hbcac5283),
	.w7(32'hbcc619df),
	.w8(32'hbc85c80d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8affdc),
	.w1(32'hbb20d876),
	.w2(32'h3bfa1153),
	.w3(32'h3bfd90d4),
	.w4(32'h3bcb9af6),
	.w5(32'h3c9f78e2),
	.w6(32'hbb848a62),
	.w7(32'hbc1ef8a9),
	.w8(32'h3a193c56),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f85ec),
	.w1(32'h3b633e12),
	.w2(32'h3bef3040),
	.w3(32'h3bb2aac5),
	.w4(32'h3b71195a),
	.w5(32'h3bd3e703),
	.w6(32'h3b35a059),
	.w7(32'hb9191f17),
	.w8(32'h3b81dbac),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ade55),
	.w1(32'h3b761cb5),
	.w2(32'h3be7f3e2),
	.w3(32'h3a3348c8),
	.w4(32'h3b51b2dd),
	.w5(32'h3b23c506),
	.w6(32'h3ba3d294),
	.w7(32'h3b579c21),
	.w8(32'h3bd39e75),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6aacb7),
	.w1(32'hbc7ee23d),
	.w2(32'h3c09a176),
	.w3(32'hbad29f3d),
	.w4(32'hbba8e4eb),
	.w5(32'hbb847215),
	.w6(32'hbb2ecda0),
	.w7(32'hb8994657),
	.w8(32'hbc13851c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc849ef3),
	.w1(32'h3b6576f5),
	.w2(32'h3a727885),
	.w3(32'hbc0738b6),
	.w4(32'h3bee0a68),
	.w5(32'h3c4cbf88),
	.w6(32'h3b0afaf5),
	.w7(32'hbb7d534c),
	.w8(32'h3b3429b1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b17d5),
	.w1(32'h3af78707),
	.w2(32'h3b8cd8e4),
	.w3(32'h398e2876),
	.w4(32'hbb8d1e49),
	.w5(32'hbb6caf48),
	.w6(32'h3ad936a3),
	.w7(32'h3b9a3d6e),
	.w8(32'h3bfe5fb3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2e5f5),
	.w1(32'h3bf582e5),
	.w2(32'h3bd40487),
	.w3(32'hbb8aa140),
	.w4(32'h3b9a7564),
	.w5(32'hbbae043d),
	.w6(32'h3ba82bf3),
	.w7(32'h3bcd0c71),
	.w8(32'hbad1fe5b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88a6ef),
	.w1(32'h3bc70114),
	.w2(32'h3b996e85),
	.w3(32'hbc2503f8),
	.w4(32'hbb30b40e),
	.w5(32'h3b9a3cfe),
	.w6(32'hbb421c0d),
	.w7(32'hbc768e95),
	.w8(32'hbbacbd43),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7980e),
	.w1(32'hbc42cea5),
	.w2(32'h3ca2a77f),
	.w3(32'hba285ad5),
	.w4(32'hbc150528),
	.w5(32'hbc147995),
	.w6(32'hbc256c6d),
	.w7(32'hba940d90),
	.w8(32'hbbf22be8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a9255),
	.w1(32'h3c61a82e),
	.w2(32'h3cadd797),
	.w3(32'hbc5864dd),
	.w4(32'h3a846ec9),
	.w5(32'hbc944ccc),
	.w6(32'h3c372854),
	.w7(32'h3c874ec1),
	.w8(32'h3c275394),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65d4b5),
	.w1(32'h3b377178),
	.w2(32'h3a845af7),
	.w3(32'hbbcdad61),
	.w4(32'h3b9058e3),
	.w5(32'h3a66a2c8),
	.w6(32'hbab70e42),
	.w7(32'hbbc513ff),
	.w8(32'hbac77bd2),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab91afe),
	.w1(32'h3a0334fa),
	.w2(32'h38d79978),
	.w3(32'h3b3d131a),
	.w4(32'h3a519357),
	.w5(32'h398834b5),
	.w6(32'h3a667e6f),
	.w7(32'h3a33bb3f),
	.w8(32'h37091eaf),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5431e8),
	.w1(32'h3bf8d36b),
	.w2(32'h3accec89),
	.w3(32'h3a38d2a8),
	.w4(32'h3bacf4ac),
	.w5(32'hbba7710b),
	.w6(32'hbb34ab0d),
	.w7(32'hb7968463),
	.w8(32'h3b8c65da),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ccef0),
	.w1(32'hbbbda403),
	.w2(32'h3a8fd9f9),
	.w3(32'h3a460d01),
	.w4(32'hbb05ee56),
	.w5(32'hbab18163),
	.w6(32'h3a49fde0),
	.w7(32'h3ad8a120),
	.w8(32'hba2cc1ae),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d43b3),
	.w1(32'hbacf62d5),
	.w2(32'h3a0afd78),
	.w3(32'hba1cf494),
	.w4(32'h389593a5),
	.w5(32'hb8c5acfa),
	.w6(32'h39c6ee4f),
	.w7(32'h399f4f5d),
	.w8(32'hb9417196),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39338ae9),
	.w1(32'hba8121c5),
	.w2(32'hb987bdfb),
	.w3(32'hba5559f1),
	.w4(32'h37ab8052),
	.w5(32'h39c66b6a),
	.w6(32'hbaf76a3e),
	.w7(32'h3af8c523),
	.w8(32'h3ab36652),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3956fb17),
	.w1(32'h38a3a595),
	.w2(32'h3952f125),
	.w3(32'hb90da1d7),
	.w4(32'hb9d9352e),
	.w5(32'h3a5055ba),
	.w6(32'h3a5bd0e7),
	.w7(32'hb96ee4e9),
	.w8(32'h398728d7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e74a),
	.w1(32'hbaddf788),
	.w2(32'h3a2e0d6f),
	.w3(32'h3a64af00),
	.w4(32'hba07918a),
	.w5(32'h3a4b6a8b),
	.w6(32'h3abbf285),
	.w7(32'h3acfa480),
	.w8(32'h3a627c43),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb822639),
	.w1(32'h3b076367),
	.w2(32'hba1773c5),
	.w3(32'hbae3e4b9),
	.w4(32'hbad3375f),
	.w5(32'h3a2b90f6),
	.w6(32'h3b072282),
	.w7(32'hbb15b5d2),
	.w8(32'hbab0425a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc582e6a),
	.w1(32'hbc22678d),
	.w2(32'hba823fa9),
	.w3(32'hb8bb5422),
	.w4(32'h3889fb09),
	.w5(32'hbb894e4d),
	.w6(32'hbb2d6b19),
	.w7(32'h3b076bf2),
	.w8(32'hbb60eb96),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b231f07),
	.w1(32'h3b378dcc),
	.w2(32'h3a8002f0),
	.w3(32'hbad121d4),
	.w4(32'hbaf73f47),
	.w5(32'h39fe26d3),
	.w6(32'hba827761),
	.w7(32'hbb2e6501),
	.w8(32'hba4361b4),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0960a7),
	.w1(32'hba90c7d6),
	.w2(32'h3ac136c0),
	.w3(32'hbb4821ac),
	.w4(32'h3b0085e7),
	.w5(32'h3ad8667f),
	.w6(32'hb89424b1),
	.w7(32'hb9088180),
	.w8(32'h39e42f53),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaa181),
	.w1(32'hbbc368c4),
	.w2(32'hba894504),
	.w3(32'h3a14979f),
	.w4(32'h3b32a16e),
	.w5(32'hbafd57f5),
	.w6(32'h3a27048a),
	.w7(32'h3b4f7028),
	.w8(32'hba7a1cd1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83016d),
	.w1(32'h3ba01568),
	.w2(32'hb84df8e4),
	.w3(32'hb9fc0a0a),
	.w4(32'h3b4931c1),
	.w5(32'h3b78eaa4),
	.w6(32'hba571505),
	.w7(32'h3a966a41),
	.w8(32'h3bb337ef),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0f3ac),
	.w1(32'hbba9bfbd),
	.w2(32'h3a5c0cb0),
	.w3(32'hb9357cda),
	.w4(32'h3ac751ff),
	.w5(32'h3abb7981),
	.w6(32'h3aa70e14),
	.w7(32'h3b248d4e),
	.w8(32'hba312242),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e1902),
	.w1(32'hb9411325),
	.w2(32'hb8cede9a),
	.w3(32'h384983ee),
	.w4(32'h398f3022),
	.w5(32'h39743c46),
	.w6(32'h38bc72f4),
	.w7(32'h3973cc37),
	.w8(32'h39c992a0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb71d60),
	.w1(32'h3b7cd4de),
	.w2(32'h3b0940aa),
	.w3(32'h3aea7a02),
	.w4(32'hbbd083e4),
	.w5(32'hbb7acf93),
	.w6(32'h3b84ada1),
	.w7(32'hbb9d40e8),
	.w8(32'hbaef9324),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca532c),
	.w1(32'hb8c3550d),
	.w2(32'hba83e6e4),
	.w3(32'hb931d3c4),
	.w4(32'h39fbecb4),
	.w5(32'h3acbf67f),
	.w6(32'hba96450d),
	.w7(32'h39d73288),
	.w8(32'h3aae4d45),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b52eb),
	.w1(32'hb92e1a54),
	.w2(32'hb91df44a),
	.w3(32'hba046f3d),
	.w4(32'hb9748c67),
	.w5(32'hb96bdbc5),
	.w6(32'hb9313c77),
	.w7(32'hb78cf681),
	.w8(32'h38eaa2ca),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372aaaae),
	.w1(32'h38c59866),
	.w2(32'h39a71cba),
	.w3(32'h38cfc30c),
	.w4(32'h38071b85),
	.w5(32'h38831b92),
	.w6(32'h398ec70c),
	.w7(32'h38ea3274),
	.w8(32'h39864e53),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8cc07),
	.w1(32'hbaa95ddc),
	.w2(32'h36b1c605),
	.w3(32'hba341061),
	.w4(32'hb5824b98),
	.w5(32'h393b6e91),
	.w6(32'hb85476e6),
	.w7(32'h39983819),
	.w8(32'h3a718af8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb3c3),
	.w1(32'h3a9295a5),
	.w2(32'hbb15c024),
	.w3(32'hbb72cea4),
	.w4(32'hbb06d0b0),
	.w5(32'h39706b6b),
	.w6(32'hbb71003a),
	.w7(32'hbb5467df),
	.w8(32'hbb3fe889),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d02b8),
	.w1(32'hbb493d56),
	.w2(32'hbaac5b80),
	.w3(32'h398b9cc6),
	.w4(32'hbaa8698d),
	.w5(32'hbaf81bf5),
	.w6(32'h39224f64),
	.w7(32'h390bb82a),
	.w8(32'hb898058f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9229e95),
	.w1(32'h38e76ba3),
	.w2(32'h394c63eb),
	.w3(32'hb8c2085b),
	.w4(32'h392d752b),
	.w5(32'h39822e02),
	.w6(32'h3983b89d),
	.w7(32'h38e1e6ef),
	.w8(32'h393287ab),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe544c1),
	.w1(32'hbbc6b82f),
	.w2(32'h3a3c5d29),
	.w3(32'h3b00d3bc),
	.w4(32'hbad54f34),
	.w5(32'hb9e93a17),
	.w6(32'h3a521ef6),
	.w7(32'h3b15b16f),
	.w8(32'hba9f71e2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c662b),
	.w1(32'hb96ca39f),
	.w2(32'h3a0a4417),
	.w3(32'h3a80e013),
	.w4(32'hb944077c),
	.w5(32'hba0a1344),
	.w6(32'h3a841f2f),
	.w7(32'h399abb7f),
	.w8(32'hba93f2a1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3ea88),
	.w1(32'hbbe29fe3),
	.w2(32'hbacbd598),
	.w3(32'h3a9c0f8f),
	.w4(32'h3bd35b90),
	.w5(32'h3ae31cb0),
	.w6(32'hba869c2a),
	.w7(32'h3ad7ecc4),
	.w8(32'hbb656903),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46ba8b),
	.w1(32'h3b41b857),
	.w2(32'hbb1c23ac),
	.w3(32'h3bc93011),
	.w4(32'hbc03a595),
	.w5(32'hbae0cdc7),
	.w6(32'h3b0bbd84),
	.w7(32'hbbd67cb6),
	.w8(32'hbbaed9ad),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acefae0),
	.w1(32'h3adb49aa),
	.w2(32'h399d4d11),
	.w3(32'h38a4cb4c),
	.w4(32'hbacd448e),
	.w5(32'hb92a4c27),
	.w6(32'hb97ccff2),
	.w7(32'hbb13e6b5),
	.w8(32'hbadde1ae),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba643979),
	.w1(32'h38ba7749),
	.w2(32'h38b7339a),
	.w3(32'hb79eacd2),
	.w4(32'h3912d1fd),
	.w5(32'h3a5d1e79),
	.w6(32'h375a1c94),
	.w7(32'h39ff9dd0),
	.w8(32'h3a49fa89),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392bb7ca),
	.w1(32'h3b1711eb),
	.w2(32'h3add8eb8),
	.w3(32'h3996a59e),
	.w4(32'h390daac7),
	.w5(32'h3ab2ef28),
	.w6(32'h39d85f29),
	.w7(32'h3a858571),
	.w8(32'h3b20e211),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01b993),
	.w1(32'hba3c4983),
	.w2(32'hba057523),
	.w3(32'hbad6a156),
	.w4(32'hbb1bb853),
	.w5(32'h3a49a401),
	.w6(32'h3b22917c),
	.w7(32'hbb04cb94),
	.w8(32'h39d40d1a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9719ea),
	.w1(32'h3b78df80),
	.w2(32'h3b313430),
	.w3(32'h3a92cdd7),
	.w4(32'hb986e29f),
	.w5(32'h3b20838c),
	.w6(32'h39d907d4),
	.w7(32'hbadeee27),
	.w8(32'h391d6c9e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef5fe1),
	.w1(32'hbb2f4e33),
	.w2(32'h39fd095a),
	.w3(32'hb97e4d50),
	.w4(32'h3aa7e108),
	.w5(32'h38d30c84),
	.w6(32'hb9abc723),
	.w7(32'h3a321d99),
	.w8(32'hba33f329),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df57ae),
	.w1(32'h39860f74),
	.w2(32'h39a9dd48),
	.w3(32'h392ea0f1),
	.w4(32'h398b55d5),
	.w5(32'h39b82baa),
	.w6(32'h383a8d4a),
	.w7(32'hb809d0b3),
	.w8(32'hb905c4b9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc76ba),
	.w1(32'hbb6740a6),
	.w2(32'h3af5d5aa),
	.w3(32'hbb015213),
	.w4(32'h3a514190),
	.w5(32'h3a4ad853),
	.w6(32'hbaee0daa),
	.w7(32'h3accdf3c),
	.w8(32'h3a0bc093),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931a88a),
	.w1(32'hbab648f2),
	.w2(32'h39a740e4),
	.w3(32'h39ebf362),
	.w4(32'h3a0ada34),
	.w5(32'h3955e49e),
	.w6(32'hb7e19ba1),
	.w7(32'hba009f1c),
	.w8(32'hb9aa3899),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e1786),
	.w1(32'h3b692237),
	.w2(32'h3a7d7634),
	.w3(32'hba807e6d),
	.w4(32'hb9e9d773),
	.w5(32'hb91136b3),
	.w6(32'hb993d042),
	.w7(32'hbb093b90),
	.w8(32'h399a1480),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aee444),
	.w1(32'hb9157be0),
	.w2(32'hb9cd235b),
	.w3(32'hba1496f0),
	.w4(32'hb89092e5),
	.w5(32'hb968268e),
	.w6(32'hb97c9606),
	.w7(32'h38b96fa3),
	.w8(32'hb7b525d8),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b4041),
	.w1(32'h3b6f9343),
	.w2(32'h3ab22818),
	.w3(32'h3b463e6c),
	.w4(32'hbae663e5),
	.w5(32'hbb8eaf48),
	.w6(32'h3a713d3f),
	.w7(32'hba0763bb),
	.w8(32'hbace1afa),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f0f85d),
	.w1(32'hb9959fb1),
	.w2(32'hb9c40b8a),
	.w3(32'hba3e1e34),
	.w4(32'hb9bdece6),
	.w5(32'hba048304),
	.w6(32'hb9229e4b),
	.w7(32'hb934d715),
	.w8(32'hb9ff22cd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ffce5),
	.w1(32'hb8d94ba9),
	.w2(32'hb9cbd3a3),
	.w3(32'hb8e82750),
	.w4(32'hb94c61d2),
	.w5(32'hba2093dd),
	.w6(32'hb7356682),
	.w7(32'hb9c6c19c),
	.w8(32'hba4dd1b0),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae683f7),
	.w1(32'hba7a09be),
	.w2(32'hbb0a4c74),
	.w3(32'hba55fdec),
	.w4(32'hbad5931e),
	.w5(32'h3a51b812),
	.w6(32'hbad36cc1),
	.w7(32'hbacece08),
	.w8(32'h3aa2a3a6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074efc),
	.w1(32'hbb9b39da),
	.w2(32'hbb513243),
	.w3(32'hbb87a67a),
	.w4(32'h3b39de39),
	.w5(32'h389dfebb),
	.w6(32'hbbb691bd),
	.w7(32'h3b95823b),
	.w8(32'h3b68c25a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b5f89),
	.w1(32'h3ae2646e),
	.w2(32'h3a8181c7),
	.w3(32'h3a800b25),
	.w4(32'h3a1ce1d7),
	.w5(32'h39c96173),
	.w6(32'h3a404814),
	.w7(32'h39f1a126),
	.w8(32'h38217668),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37786d58),
	.w1(32'h3a72e21c),
	.w2(32'hbacee35d),
	.w3(32'hb9979440),
	.w4(32'hbb1696ab),
	.w5(32'hbb0fdcac),
	.w6(32'h3aadc6c1),
	.w7(32'hba356033),
	.w8(32'hbaf8f99d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad12c3e),
	.w1(32'hba73761b),
	.w2(32'hba95d564),
	.w3(32'h3ab5c1b9),
	.w4(32'hbb9809f5),
	.w5(32'hbb2b3eb5),
	.w6(32'h3ac4dbe6),
	.w7(32'hbb1fa70b),
	.w8(32'hbb250f9c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83e10d),
	.w1(32'hbb279524),
	.w2(32'h3a2402b4),
	.w3(32'h3a064be5),
	.w4(32'h3a2e3f2e),
	.w5(32'hba9c90ee),
	.w6(32'h3bf0b15c),
	.w7(32'hbb08598b),
	.w8(32'hba71f7a0),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e7950),
	.w1(32'hbb96641c),
	.w2(32'hbae1369f),
	.w3(32'h3a89680d),
	.w4(32'h3a2809c1),
	.w5(32'h3a94b750),
	.w6(32'hb9fb97c5),
	.w7(32'h3a7539a1),
	.w8(32'h3839241c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38f9e0),
	.w1(32'hbbae440a),
	.w2(32'hbaaa7c53),
	.w3(32'hba445915),
	.w4(32'h392905c3),
	.w5(32'hba2bea6b),
	.w6(32'h3a9ea2be),
	.w7(32'h3b597550),
	.w8(32'hb8eb2734),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df9682),
	.w1(32'h3909cbce),
	.w2(32'hb84ae2e7),
	.w3(32'hb8d2e7cc),
	.w4(32'h3991e48a),
	.w5(32'h3893a709),
	.w6(32'hb87539a2),
	.w7(32'h3a5845af),
	.w8(32'h3a5788dc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7a1f8),
	.w1(32'hbac612d5),
	.w2(32'h3b0a6dd0),
	.w3(32'hb97cf17b),
	.w4(32'hbb002eaf),
	.w5(32'h3a5d4fdc),
	.w6(32'h3aa35bd2),
	.w7(32'hba07dce3),
	.w8(32'hba75d7cc),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3752c8fb),
	.w1(32'h39734f3a),
	.w2(32'h399b6d6e),
	.w3(32'h38076eed),
	.w4(32'h3960a046),
	.w5(32'h39600873),
	.w6(32'h39841c38),
	.w7(32'h397bbe40),
	.w8(32'h3979c52a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27dccb),
	.w1(32'h39bbec28),
	.w2(32'h3a708613),
	.w3(32'h3995c183),
	.w4(32'h3a5daa4b),
	.w5(32'h3a7b0ce5),
	.w6(32'h38058601),
	.w7(32'h3a4924b6),
	.w8(32'h399ab6e1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1b5ee),
	.w1(32'h3996a30f),
	.w2(32'h38628615),
	.w3(32'h3982d6a4),
	.w4(32'hbad8efd4),
	.w5(32'hb9ba6f0c),
	.w6(32'hba6d5966),
	.w7(32'hbabf449b),
	.w8(32'hba77dc61),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe2da7),
	.w1(32'hb8c5728a),
	.w2(32'h3b3f84a4),
	.w3(32'hbaca2579),
	.w4(32'hba5b2fae),
	.w5(32'h3b3489fa),
	.w6(32'h3ab75f17),
	.w7(32'hbb0a136a),
	.w8(32'hb977832c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bf3d9e),
	.w1(32'h3703dee1),
	.w2(32'hb8f47e99),
	.w3(32'hb7443095),
	.w4(32'hb7a11068),
	.w5(32'hb92360fa),
	.w6(32'hb8d143f2),
	.w7(32'hb954b1ac),
	.w8(32'hb96c1d5c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1095a5),
	.w1(32'hb96cd8a0),
	.w2(32'h383f4178),
	.w3(32'hb9ff2493),
	.w4(32'hb8864e41),
	.w5(32'h38e24224),
	.w6(32'hb9353df0),
	.w7(32'hb7986a54),
	.w8(32'h36976d23),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c7d1a),
	.w1(32'h3b5c9988),
	.w2(32'h3a26563f),
	.w3(32'h3a0eb20d),
	.w4(32'hba390efb),
	.w5(32'hb9aa1391),
	.w6(32'hba2b43da),
	.w7(32'hba93f94c),
	.w8(32'h394cc316),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb307cb2),
	.w1(32'hbaf59403),
	.w2(32'h39b4fd1b),
	.w3(32'h3b84a370),
	.w4(32'h3bb4a07a),
	.w5(32'hba3ecfb0),
	.w6(32'h3bc4d690),
	.w7(32'h3afed9de),
	.w8(32'hbb69ece7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a5f7e),
	.w1(32'hbbd9c2aa),
	.w2(32'hbc0d6f84),
	.w3(32'hbc043b46),
	.w4(32'h38b351f8),
	.w5(32'hbb00644c),
	.w6(32'hbbf55ecd),
	.w7(32'h3986aa35),
	.w8(32'hba37653f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a800a6),
	.w1(32'hb9ed3897),
	.w2(32'hbaaadd95),
	.w3(32'h38da5116),
	.w4(32'hb955f362),
	.w5(32'hbaa5ad48),
	.w6(32'h39f92d0c),
	.w7(32'hb9eb40d3),
	.w8(32'hba58a789),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc788965),
	.w1(32'hbb946d55),
	.w2(32'hbb6cb09f),
	.w3(32'hba846b03),
	.w4(32'h3b263a37),
	.w5(32'hbbbb53e9),
	.w6(32'h3b2b8add),
	.w7(32'h3b23fc05),
	.w8(32'h38cf7a63),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb76ff),
	.w1(32'h3b13dabe),
	.w2(32'h3b592fab),
	.w3(32'h3b6f083b),
	.w4(32'hbba3a914),
	.w5(32'h3ba34226),
	.w6(32'h3bd2c253),
	.w7(32'hbb6fb68e),
	.w8(32'hbb064ff6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f951cd),
	.w1(32'hbb8c3285),
	.w2(32'hb972828c),
	.w3(32'h3a332abf),
	.w4(32'h39a0b9d8),
	.w5(32'hb9b374d5),
	.w6(32'hbad13626),
	.w7(32'hb9966a2e),
	.w8(32'hbb1fdf2a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb810e01e),
	.w1(32'hb9a71089),
	.w2(32'hba021cd6),
	.w3(32'h37bdfd44),
	.w4(32'hba07aca8),
	.w5(32'hba3e0ff2),
	.w6(32'hba095ae0),
	.w7(32'hb9e5a088),
	.w8(32'hb988dd7e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39995b),
	.w1(32'hb8d43b3c),
	.w2(32'hb950b460),
	.w3(32'hb9ea2ef1),
	.w4(32'h3807cf4b),
	.w5(32'hb946c8df),
	.w6(32'h3a1a6139),
	.w7(32'h39cb4df1),
	.w8(32'h38e60990),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb792ba3f),
	.w1(32'hb80f69b6),
	.w2(32'h37e5b59c),
	.w3(32'hb7f250ac),
	.w4(32'hb8d3bc3b),
	.w5(32'hb8f58a35),
	.w6(32'hb8461b22),
	.w7(32'hb8a61570),
	.w8(32'hb818a99f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bb547),
	.w1(32'hbb5617e5),
	.w2(32'hba773dc6),
	.w3(32'hb9801092),
	.w4(32'h39ec4728),
	.w5(32'hbb6d484f),
	.w6(32'hbae83ab8),
	.w7(32'h395b77bc),
	.w8(32'hbb06fb94),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c6c6d),
	.w1(32'hba9cfb8c),
	.w2(32'hb9d44b57),
	.w3(32'hb89e2e88),
	.w4(32'h3a648a28),
	.w5(32'h3a554f20),
	.w6(32'h3a10d698),
	.w7(32'h3a404e0f),
	.w8(32'h3a2e052f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ca5b0),
	.w1(32'h3b7d5541),
	.w2(32'h3933507a),
	.w3(32'hba018727),
	.w4(32'hba997ce5),
	.w5(32'h3a6f19d8),
	.w6(32'hbb141063),
	.w7(32'hbb0f67c9),
	.w8(32'hb905e696),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c14064),
	.w1(32'h3a846373),
	.w2(32'h3a2a4c92),
	.w3(32'h37bd5f6b),
	.w4(32'h39f74daa),
	.w5(32'h3a88903d),
	.w6(32'h3925467c),
	.w7(32'h38c95cb9),
	.w8(32'h3a3a783f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba0c00),
	.w1(32'hbb4b22c8),
	.w2(32'hbb00f08e),
	.w3(32'h3a484dd0),
	.w4(32'h3ad526c8),
	.w5(32'hbb8a742c),
	.w6(32'h3b0b9861),
	.w7(32'h3b404168),
	.w8(32'hba57b6d4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a74a9),
	.w1(32'hbb07ec40),
	.w2(32'hbb2973de),
	.w3(32'hbab698a7),
	.w4(32'h3aa185da),
	.w5(32'hb9ea16fe),
	.w6(32'hba99b82d),
	.w7(32'h39dcb131),
	.w8(32'h3a9f5784),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97fb9a2),
	.w1(32'h38b436b6),
	.w2(32'h392b0e58),
	.w3(32'hb98108e9),
	.w4(32'h38bd09d5),
	.w5(32'h392f10d5),
	.w6(32'h379a7818),
	.w7(32'h38a8d51a),
	.w8(32'h390011a1),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8968d),
	.w1(32'hba13035d),
	.w2(32'hbac144a0),
	.w3(32'hbaa8a420),
	.w4(32'h3b216718),
	.w5(32'hba0f60f8),
	.w6(32'h38ef351e),
	.w7(32'h3b0cd8a6),
	.w8(32'h3a5fb6a2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c6383),
	.w1(32'hb7fe7231),
	.w2(32'h38a6e020),
	.w3(32'h38973653),
	.w4(32'hb59f0417),
	.w5(32'h391669a5),
	.w6(32'h3890e4ef),
	.w7(32'h36856fbe),
	.w8(32'h38a86571),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f13d9),
	.w1(32'hba7eb4a9),
	.w2(32'hba8a9fa8),
	.w3(32'h396208a4),
	.w4(32'h3a2a7392),
	.w5(32'hba6e3327),
	.w6(32'h3a2cedf9),
	.w7(32'h3a9f3cc0),
	.w8(32'h3930a347),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b950b),
	.w1(32'h3b65b0e2),
	.w2(32'h3a6303cd),
	.w3(32'hb9986017),
	.w4(32'hba8d3689),
	.w5(32'h3b85504e),
	.w6(32'hba1a50f7),
	.w7(32'hbb80352d),
	.w8(32'hb9c0a84d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a55575),
	.w1(32'h3ac4861e),
	.w2(32'hba02f70f),
	.w3(32'h3a8db4a7),
	.w4(32'h38c8c056),
	.w5(32'h3a810006),
	.w6(32'h3a6be366),
	.w7(32'hb82a2181),
	.w8(32'h3a2f55a9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab29979),
	.w1(32'h3a1f1b5c),
	.w2(32'h391b519d),
	.w3(32'h3a1daad9),
	.w4(32'hb90f0fa2),
	.w5(32'hba2b5ba1),
	.w6(32'h38be999e),
	.w7(32'hb9136b11),
	.w8(32'hba2508e9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81f63b),
	.w1(32'h3b42b147),
	.w2(32'h39598277),
	.w3(32'h39836cc8),
	.w4(32'hbb17ea7a),
	.w5(32'h39fc747e),
	.w6(32'h3a8e64e2),
	.w7(32'hbac166b5),
	.w8(32'hb9858bbc),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb1cca),
	.w1(32'hbb82d355),
	.w2(32'h3a28152c),
	.w3(32'hbaaf6bc8),
	.w4(32'hba1943ba),
	.w5(32'h3aa835d1),
	.w6(32'hba1527c6),
	.w7(32'h3ae82a6e),
	.w8(32'h3a6aa587),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29df01),
	.w1(32'hbadc1c16),
	.w2(32'hba4b057c),
	.w3(32'hba224749),
	.w4(32'h39bf9c43),
	.w5(32'hba7f5f86),
	.w6(32'hba2d16aa),
	.w7(32'h3a0a7e23),
	.w8(32'hb9be9bf4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb859785a),
	.w1(32'hb7b2bf20),
	.w2(32'h36170c06),
	.w3(32'h37763550),
	.w4(32'hb8a1378e),
	.w5(32'hb8d6789d),
	.w6(32'h38a0e262),
	.w7(32'hb7883a14),
	.w8(32'hb940afa2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7200efa),
	.w1(32'hb9291803),
	.w2(32'hb901318e),
	.w3(32'hb91b2ac4),
	.w4(32'hb9c16b4b),
	.w5(32'hb9b1c24f),
	.w6(32'h39cdb2fa),
	.w7(32'hb9926822),
	.w8(32'hb98a08d7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c032704),
	.w1(32'hbb530da9),
	.w2(32'hbac277fe),
	.w3(32'h39fd8cc4),
	.w4(32'h3b80eef7),
	.w5(32'h3b0fb930),
	.w6(32'hbb3770ce),
	.w7(32'h3bb4a849),
	.w8(32'h3c05807e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcdb8c),
	.w1(32'hba0f7a17),
	.w2(32'hbac21933),
	.w3(32'hbaa8ab17),
	.w4(32'h3b8ba234),
	.w5(32'h3aa71c58),
	.w6(32'h3ab8fd71),
	.w7(32'h3b98603b),
	.w8(32'h3b4ffad5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83e5dd),
	.w1(32'h3b495fb1),
	.w2(32'h3ac28120),
	.w3(32'h3aeb4bad),
	.w4(32'h3abaeb20),
	.w5(32'h3b64a70f),
	.w6(32'h3a3344f3),
	.w7(32'h3a6b6df8),
	.w8(32'h3b3681bb),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7b6a3),
	.w1(32'hbb80ba72),
	.w2(32'h3c372691),
	.w3(32'h3b0aaafb),
	.w4(32'h3b16efa1),
	.w5(32'h3b884e81),
	.w6(32'h39a14a72),
	.w7(32'h3b227f7d),
	.w8(32'hbbadb8cc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c9a53),
	.w1(32'h3a86c252),
	.w2(32'hb9532526),
	.w3(32'hba0e213e),
	.w4(32'hb92b386e),
	.w5(32'hb9ee5f89),
	.w6(32'hba06cf02),
	.w7(32'hba6c1350),
	.w8(32'h3959df37),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2dd20e),
	.w1(32'hba80a8d4),
	.w2(32'h393f7338),
	.w3(32'hba6968e2),
	.w4(32'h38d95664),
	.w5(32'h3a4b6fcc),
	.w6(32'hba88d397),
	.w7(32'hba39ffc7),
	.w8(32'h38c6e5ce),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbf2be),
	.w1(32'hbb69021f),
	.w2(32'hbbc55ce6),
	.w3(32'hbb297a11),
	.w4(32'h3b474cdc),
	.w5(32'hbbb708de),
	.w6(32'hbbea47de),
	.w7(32'h3a2f6876),
	.w8(32'h3b674dd3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cf8bd),
	.w1(32'hbbaf3a62),
	.w2(32'hba29be5e),
	.w3(32'hbb077952),
	.w4(32'hba05bd23),
	.w5(32'hbb8dbfa6),
	.w6(32'hba08c124),
	.w7(32'h3a4ad177),
	.w8(32'hba838c52),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bcab8),
	.w1(32'hbbd1ee41),
	.w2(32'hbaccbab8),
	.w3(32'hbb8b2fc6),
	.w4(32'h3bcbccb2),
	.w5(32'hba90fedf),
	.w6(32'hbb9e36d1),
	.w7(32'h3b40d645),
	.w8(32'h3a5e7092),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b642d26),
	.w1(32'h3b8ac03f),
	.w2(32'h3b11b5c6),
	.w3(32'hb9c97110),
	.w4(32'hbb09d132),
	.w5(32'h3aac2dec),
	.w6(32'hba94e02b),
	.w7(32'hbb683797),
	.w8(32'hb8a52afd),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00444c),
	.w1(32'h3b0628fd),
	.w2(32'hba33ef42),
	.w3(32'hbb544c1b),
	.w4(32'hbb8510a1),
	.w5(32'h39c568b9),
	.w6(32'hbad13169),
	.w7(32'hbbbcd168),
	.w8(32'hbaf86a6e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb721a393),
	.w1(32'h3893a712),
	.w2(32'h38e6b4dd),
	.w3(32'hb78811de),
	.w4(32'hb7a8f5df),
	.w5(32'hb76eb708),
	.w6(32'h37bb80c5),
	.w7(32'h3881314a),
	.w8(32'hb7e82168),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8144076),
	.w1(32'hb8279fc4),
	.w2(32'h378f5fb5),
	.w3(32'hb91e388e),
	.w4(32'h3741bdb3),
	.w5(32'hb81226ec),
	.w6(32'h38586b66),
	.w7(32'hb83918f3),
	.w8(32'hb8c1e726),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bd7e3),
	.w1(32'h3b8487a3),
	.w2(32'h3b650d07),
	.w3(32'hba599c31),
	.w4(32'h38e1155a),
	.w5(32'hb8b3ed3d),
	.w6(32'hb9b85e97),
	.w7(32'hb9a9e622),
	.w8(32'h39db1eaf),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a5aeed),
	.w1(32'hb9a87d8d),
	.w2(32'hb9922b03),
	.w3(32'hb72c3f5e),
	.w4(32'hb9d06eb4),
	.w5(32'hb9d1e348),
	.w6(32'hb9b3682d),
	.w7(32'hb9c51c4e),
	.w8(32'hb94e238f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c2f78),
	.w1(32'hbb348d63),
	.w2(32'hbb6b3c66),
	.w3(32'hba1040ec),
	.w4(32'hbb107357),
	.w5(32'hbb8764d4),
	.w6(32'hbadf8d39),
	.w7(32'hba79dc0f),
	.w8(32'hbb695b70),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbee3f7),
	.w1(32'hba1a5c00),
	.w2(32'h3a4f50e6),
	.w3(32'hbb324447),
	.w4(32'h3b92ed12),
	.w5(32'hb9b13ea1),
	.w6(32'hb93b19f2),
	.w7(32'hb93e5156),
	.w8(32'h3b8b010c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73a9427),
	.w1(32'h39bb7885),
	.w2(32'hb8780737),
	.w3(32'h3a382bbc),
	.w4(32'h3a70ed94),
	.w5(32'h3a885082),
	.w6(32'h39751a1d),
	.w7(32'hb893168a),
	.w8(32'h39d29ee7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c3aed),
	.w1(32'h38963855),
	.w2(32'hb92c9f99),
	.w3(32'hb9fab207),
	.w4(32'hb9147729),
	.w5(32'hb9897dc6),
	.w6(32'h388642c8),
	.w7(32'hb99abcb1),
	.w8(32'hb9b4fbd5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7ae9d),
	.w1(32'hbc633ec3),
	.w2(32'hbb5e1b04),
	.w3(32'hbc07e217),
	.w4(32'h3b7f5ea2),
	.w5(32'hbb8c5d29),
	.w6(32'hbc1d969a),
	.w7(32'h3b686dec),
	.w8(32'hb98d4d96),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb878bbc),
	.w1(32'hbaa4fd3e),
	.w2(32'h3aaf3402),
	.w3(32'h389bf4fa),
	.w4(32'h3a98743e),
	.w5(32'h3969c6b4),
	.w6(32'h3a110299),
	.w7(32'h3b1dc5cb),
	.w8(32'h3a34a557),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9332ed4),
	.w1(32'h38ef3b1c),
	.w2(32'h391e6931),
	.w3(32'hb8cf0ea4),
	.w4(32'h39142f25),
	.w5(32'h370d0746),
	.w6(32'h387aa9bb),
	.w7(32'h37bd23bd),
	.w8(32'h39298a7e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6e74),
	.w1(32'hbb8c6c0b),
	.w2(32'hba290238),
	.w3(32'hba6a70ee),
	.w4(32'h39b41ebf),
	.w5(32'hbacdfeee),
	.w6(32'hbaa6b55c),
	.w7(32'h3a89c1cb),
	.w8(32'h37c2de25),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a14556),
	.w1(32'h396ce26e),
	.w2(32'h39a2c841),
	.w3(32'h397d7787),
	.w4(32'h393a2810),
	.w5(32'h392d52e1),
	.w6(32'h39a2f9d0),
	.w7(32'h39a8a676),
	.w8(32'h39295477),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70fa88b),
	.w1(32'h399c807d),
	.w2(32'h39d7a948),
	.w3(32'h395c01bd),
	.w4(32'h3a101875),
	.w5(32'h3a60986f),
	.w6(32'hb95dde92),
	.w7(32'h399b0795),
	.w8(32'h3a150187),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39232e12),
	.w1(32'h394c4ed8),
	.w2(32'h394af333),
	.w3(32'h3967bfc2),
	.w4(32'h399a4d98),
	.w5(32'h397a4315),
	.w6(32'h396d2b95),
	.w7(32'h399d184c),
	.w8(32'h39acd874),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3382f),
	.w1(32'h398f04c8),
	.w2(32'h399043b1),
	.w3(32'h39cd905c),
	.w4(32'h392bdd1a),
	.w5(32'h38e7bbbd),
	.w6(32'h390492c8),
	.w7(32'h394c0222),
	.w8(32'h391fc643),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07fa94),
	.w1(32'h3b159462),
	.w2(32'h3a8416bc),
	.w3(32'hb9803763),
	.w4(32'hba5eac12),
	.w5(32'h3964f522),
	.w6(32'hbadacdfe),
	.w7(32'hbadfe4be),
	.w8(32'h3995f2ed),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc472a6b),
	.w1(32'hbb884abe),
	.w2(32'h3b2a48a9),
	.w3(32'h3aeee6f0),
	.w4(32'hba4b362e),
	.w5(32'hb6eac3f0),
	.w6(32'h3b384dec),
	.w7(32'hbae9eba4),
	.w8(32'hbb69f32d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0febfc),
	.w1(32'hbbcf1e96),
	.w2(32'hb9de6551),
	.w3(32'hba546d90),
	.w4(32'h3867deb5),
	.w5(32'h35e9b90c),
	.w6(32'h39188166),
	.w7(32'h3b5a47c2),
	.w8(32'h3aa04065),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42e287),
	.w1(32'hbbb5a2e7),
	.w2(32'h3894ee5f),
	.w3(32'hba76fe1c),
	.w4(32'hbb05d09e),
	.w5(32'hbb22b10d),
	.w6(32'h3a198696),
	.w7(32'h386b5827),
	.w8(32'hbb0d7675),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0dd24f),
	.w1(32'h3a370a89),
	.w2(32'h3a0a6658),
	.w3(32'h3990babb),
	.w4(32'h39ee94f3),
	.w5(32'h39aa6455),
	.w6(32'h38df85b8),
	.w7(32'h39cc0c86),
	.w8(32'h394cc47d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb7ebe),
	.w1(32'h3a312724),
	.w2(32'h38811ae1),
	.w3(32'hb84ee1dc),
	.w4(32'h39382106),
	.w5(32'h3895c974),
	.w6(32'h398d9702),
	.w7(32'h39c61427),
	.w8(32'h395cf60d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e15772),
	.w1(32'h380cdd64),
	.w2(32'h38fc07a2),
	.w3(32'h3985e613),
	.w4(32'h37fbd489),
	.w5(32'h38c71d8c),
	.w6(32'h379a5cb0),
	.w7(32'h387b7772),
	.w8(32'h3929a940),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389e86d3),
	.w1(32'hb7758e7d),
	.w2(32'hb87fd6a3),
	.w3(32'h3915192d),
	.w4(32'h38f4bd00),
	.w5(32'h388f837c),
	.w6(32'h38b09390),
	.w7(32'h38c1f230),
	.w8(32'h38f64666),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3895),
	.w1(32'hbaf50a51),
	.w2(32'h3a8f2ab2),
	.w3(32'hba8f2da1),
	.w4(32'hbb04a209),
	.w5(32'hba945d90),
	.w6(32'h3b3653b4),
	.w7(32'h3a84cf90),
	.w8(32'h39089d66),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2382d1),
	.w1(32'hb8b67830),
	.w2(32'h37831b91),
	.w3(32'hb9e2af3c),
	.w4(32'hb93fb2e2),
	.w5(32'hb9b16cba),
	.w6(32'hb8e6e9b2),
	.w7(32'hb99293c1),
	.w8(32'hba2da522),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dabeb),
	.w1(32'h3a9532d2),
	.w2(32'h3a8c0d57),
	.w3(32'h3aac2348),
	.w4(32'h3abc4d01),
	.w5(32'h39e7b8d1),
	.w6(32'h3a34d516),
	.w7(32'h3a25193a),
	.w8(32'hb9528b79),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e22ad),
	.w1(32'hbadbe2a5),
	.w2(32'hbada1d5a),
	.w3(32'hbb09646f),
	.w4(32'h38e54561),
	.w5(32'hba61f815),
	.w6(32'h391abc11),
	.w7(32'hba9ef1d6),
	.w8(32'hba0455bc),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b0c9c),
	.w1(32'h38cefc13),
	.w2(32'h3912696c),
	.w3(32'h38646c0e),
	.w4(32'h3988f97c),
	.w5(32'h38e4d808),
	.w6(32'h39a730af),
	.w7(32'h398bebac),
	.w8(32'h34ded388),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c672e),
	.w1(32'hba099784),
	.w2(32'h3810f10e),
	.w3(32'h3a55ed8f),
	.w4(32'h3917c966),
	.w5(32'hba69e538),
	.w6(32'h39513a49),
	.w7(32'h3a09f63d),
	.w8(32'hb9ccf840),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7737904),
	.w1(32'hb9969880),
	.w2(32'hb9fc1964),
	.w3(32'hb8c58657),
	.w4(32'hb9cf6072),
	.w5(32'hba279733),
	.w6(32'h38e14c28),
	.w7(32'hb93961c0),
	.w8(32'hba47a64f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cdfa6),
	.w1(32'hbaef4bef),
	.w2(32'h3b0fdd21),
	.w3(32'hbb006918),
	.w4(32'hbb6dece8),
	.w5(32'h3a2a5176),
	.w6(32'h3b8fb109),
	.w7(32'hbb4978cf),
	.w8(32'hbb2e49fd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392eabaf),
	.w1(32'hbaabcfbb),
	.w2(32'hbae18cfb),
	.w3(32'h3974c175),
	.w4(32'hbaa94666),
	.w5(32'hbae0aa04),
	.w6(32'hba90b1df),
	.w7(32'hbaea1148),
	.w8(32'hb9bc48fa),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28169a),
	.w1(32'h3b0f7f48),
	.w2(32'hbb1ab658),
	.w3(32'hbaf9b885),
	.w4(32'hba6476f2),
	.w5(32'h38a96008),
	.w6(32'hba7a8225),
	.w7(32'h3b0d7db8),
	.w8(32'h3b8c3125),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule