module layer_10_featuremap_265(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad24e44),
	.w1(32'hbaf235ea),
	.w2(32'hba89a680),
	.w3(32'hbb01a30d),
	.w4(32'hbb001485),
	.w5(32'h38b73ce8),
	.w6(32'hbafb84ae),
	.w7(32'hbaf44939),
	.w8(32'hb99bc26e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba747a),
	.w1(32'h3b42fa2c),
	.w2(32'h3b8e366d),
	.w3(32'h391ef3f8),
	.w4(32'h3ad20b25),
	.w5(32'h3aa86459),
	.w6(32'hb99e84bd),
	.w7(32'hb9059d45),
	.w8(32'hba407474),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a440f),
	.w1(32'hb93cf7d8),
	.w2(32'hb924baf9),
	.w3(32'hbb065896),
	.w4(32'hba26fca2),
	.w5(32'h3a0e8ffc),
	.w6(32'hba8adcef),
	.w7(32'hb9e2ecac),
	.w8(32'hba46dadd),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d262f),
	.w1(32'h3a5d6917),
	.w2(32'hb7ff714a),
	.w3(32'hba0f86fa),
	.w4(32'h39ee7985),
	.w5(32'hba831606),
	.w6(32'hbb05f7a9),
	.w7(32'hba7468d8),
	.w8(32'hbae8a3d9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab36574),
	.w1(32'hbb7d5e5a),
	.w2(32'hbb9c605d),
	.w3(32'hbade3640),
	.w4(32'hbb07196c),
	.w5(32'hb99700f0),
	.w6(32'hbaf0b529),
	.w7(32'hbb0ad81f),
	.w8(32'h3a01abcf),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bfa89),
	.w1(32'h3a9ae190),
	.w2(32'h3a863610),
	.w3(32'h393e3eeb),
	.w4(32'h398ac15e),
	.w5(32'h3a630671),
	.w6(32'h39fed1ed),
	.w7(32'h3a06e4c7),
	.w8(32'hb7b11d80),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f80d8),
	.w1(32'hb9635159),
	.w2(32'h3aa164de),
	.w3(32'hbb5b6a37),
	.w4(32'h3b2530f4),
	.w5(32'hbb6e792c),
	.w6(32'hba6f06fb),
	.w7(32'h3aa1bd97),
	.w8(32'hbc54705c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1efdb),
	.w1(32'hbc0cb1bf),
	.w2(32'hbc674051),
	.w3(32'h3b7a8d11),
	.w4(32'hbbb70be7),
	.w5(32'hbc347be5),
	.w6(32'h3c08da97),
	.w7(32'h3afe437d),
	.w8(32'h39d44e26),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b5c9a),
	.w1(32'h3a7e9304),
	.w2(32'hba6d1a35),
	.w3(32'h3aebf572),
	.w4(32'h39af7e55),
	.w5(32'hba9ebab9),
	.w6(32'h3a1bc23d),
	.w7(32'hb9b86596),
	.w8(32'hba7d01d4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be94aca),
	.w1(32'h3ae58278),
	.w2(32'h3ad32191),
	.w3(32'h3966bb40),
	.w4(32'hbb3416c7),
	.w5(32'hbabfad8a),
	.w6(32'hbbcbdbf6),
	.w7(32'hbc045c0e),
	.w8(32'hbc2064d5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab16038),
	.w1(32'hba97cbed),
	.w2(32'hbb254cae),
	.w3(32'hbb0afd79),
	.w4(32'hbaf9fbbc),
	.w5(32'hbb04e924),
	.w6(32'h39fbc0a3),
	.w7(32'h3a329c4c),
	.w8(32'h3a96e76c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2eeb17),
	.w1(32'hbb48cf27),
	.w2(32'hba9cffc8),
	.w3(32'h3a990a42),
	.w4(32'h3b3c90ca),
	.w5(32'hba5b9bd6),
	.w6(32'h3b39ea1e),
	.w7(32'h3b961f85),
	.w8(32'hbae05d06),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b911998),
	.w1(32'hbb546377),
	.w2(32'hbbcdc397),
	.w3(32'h3bac93c3),
	.w4(32'hba93604a),
	.w5(32'hbbd19ceb),
	.w6(32'h3aad8fd8),
	.w7(32'hbb4a898b),
	.w8(32'hbc3f774f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9c620),
	.w1(32'h3a3538dc),
	.w2(32'hbab559ef),
	.w3(32'h3b39516d),
	.w4(32'h385569ca),
	.w5(32'hbb4719b1),
	.w6(32'h3b334cf5),
	.w7(32'hba3a8365),
	.w8(32'hbb3aac33),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0e9ed),
	.w1(32'h3c004b1c),
	.w2(32'h3be4ac8c),
	.w3(32'h3afc6ce3),
	.w4(32'h3b6f1789),
	.w5(32'h3b4ba045),
	.w6(32'hbb6b63a2),
	.w7(32'hbb2cf210),
	.w8(32'hba8d84f8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbba956),
	.w1(32'h3baefe78),
	.w2(32'h3ad25223),
	.w3(32'h3c0dcc8d),
	.w4(32'h3ab77cf1),
	.w5(32'hbb23a724),
	.w6(32'hba4c9393),
	.w7(32'hbb9a9de7),
	.w8(32'hbbdb6d85),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b5603),
	.w1(32'h3a24e5b8),
	.w2(32'h39d96db7),
	.w3(32'h3a304459),
	.w4(32'h3ad658bc),
	.w5(32'h3a339af0),
	.w6(32'h3a816d08),
	.w7(32'h3a8373ed),
	.w8(32'h3a2a657b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac29024),
	.w1(32'hbc224960),
	.w2(32'hbc42ef23),
	.w3(32'h3ac13990),
	.w4(32'hbc00e622),
	.w5(32'hbc412f4d),
	.w6(32'h3b3fc231),
	.w7(32'hbb145dfb),
	.w8(32'hbc6c98bc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b018371),
	.w1(32'hbb4206f4),
	.w2(32'hbbbafda2),
	.w3(32'h3a78b85a),
	.w4(32'hbb6eff82),
	.w5(32'hbbc6de51),
	.w6(32'h3ab2f311),
	.w7(32'hbb704a54),
	.w8(32'hbbf6e743),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4620e4),
	.w1(32'hbac3df0a),
	.w2(32'hba80a1a8),
	.w3(32'h3992b100),
	.w4(32'h3aa62549),
	.w5(32'h38a1f0dd),
	.w6(32'hba000cef),
	.w7(32'h392e1545),
	.w8(32'hba8cfc69),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09a390),
	.w1(32'h38bb499a),
	.w2(32'hb9b10c5e),
	.w3(32'hb8a45c45),
	.w4(32'hb9208f34),
	.w5(32'h3a45b980),
	.w6(32'h384f326c),
	.w7(32'h36c46515),
	.w8(32'h3acd3703),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22e621),
	.w1(32'h3b89aa6f),
	.w2(32'h3b9f4bb2),
	.w3(32'h3ad78247),
	.w4(32'h3b517530),
	.w5(32'h3b355ab2),
	.w6(32'h3b16a014),
	.w7(32'h3b5b8eff),
	.w8(32'h3b407391),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c520098),
	.w1(32'h3bdf8833),
	.w2(32'hbb475099),
	.w3(32'h3c8ba738),
	.w4(32'h3be9720d),
	.w5(32'hbb685d26),
	.w6(32'h3c06c80a),
	.w7(32'h3bb10ee0),
	.w8(32'hbbe6b296),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b999fda),
	.w1(32'h3b3f456f),
	.w2(32'h3b516c1e),
	.w3(32'hba8d09aa),
	.w4(32'hba79d11d),
	.w5(32'hbb728e88),
	.w6(32'hbbaf272a),
	.w7(32'hbbb0daf2),
	.w8(32'hbbd9628e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15b062),
	.w1(32'h3bea11b4),
	.w2(32'h3c0e5a61),
	.w3(32'hbbd4c95c),
	.w4(32'hb99e94b9),
	.w5(32'h3b92fbf5),
	.w6(32'hbbf1345d),
	.w7(32'hbb7b21d9),
	.w8(32'h3b15b2c9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08ab20),
	.w1(32'h3b29a317),
	.w2(32'h3b2a67bd),
	.w3(32'h3b213dac),
	.w4(32'h3b14b4f1),
	.w5(32'h3a8c86c8),
	.w6(32'h3acdbac3),
	.w7(32'h39a6366a),
	.w8(32'h3a072a32),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fdfd9),
	.w1(32'h3acb988f),
	.w2(32'h3a0ae3b5),
	.w3(32'hb9d8bd18),
	.w4(32'hba67a533),
	.w5(32'hbaef4e83),
	.w6(32'hb9358f2b),
	.w7(32'hba1f22e2),
	.w8(32'hbaba9362),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a721e4a),
	.w1(32'hbc5d19ba),
	.w2(32'h3b0711ee),
	.w3(32'h38797710),
	.w4(32'hbca04df2),
	.w5(32'h3aaafcde),
	.w6(32'hbbba132c),
	.w7(32'hbc916b34),
	.w8(32'hbb7c1e2a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d71ff),
	.w1(32'h39bb4feb),
	.w2(32'h3a9efe83),
	.w3(32'hba287f9d),
	.w4(32'h3b17ef2d),
	.w5(32'h3a5a3298),
	.w6(32'hba1ffd43),
	.w7(32'h3b285f02),
	.w8(32'h3ace4cfe),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd0708),
	.w1(32'h3bd38e28),
	.w2(32'h3c452378),
	.w3(32'hbb4d6e62),
	.w4(32'hbbd6132f),
	.w5(32'h3aa363e5),
	.w6(32'hbc041d07),
	.w7(32'hbc458246),
	.w8(32'hbb41c2a2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd04ff),
	.w1(32'h369b2606),
	.w2(32'hba1b5db6),
	.w3(32'hbb2ed120),
	.w4(32'hbb284704),
	.w5(32'hba6cc822),
	.w6(32'hbac86e84),
	.w7(32'hbb659584),
	.w8(32'hba25eacf),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba2fc5),
	.w1(32'hbb3b3824),
	.w2(32'hba13dd71),
	.w3(32'hb9071266),
	.w4(32'h3993c551),
	.w5(32'hbac503f1),
	.w6(32'h3a36df46),
	.w7(32'h3ade28de),
	.w8(32'h3a5f04f2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b966da4),
	.w1(32'h3b19633c),
	.w2(32'h39576e46),
	.w3(32'h3b46e138),
	.w4(32'hba315980),
	.w5(32'hbb3d6669),
	.w6(32'h3a90a9be),
	.w7(32'hbb193c88),
	.w8(32'hbbb59d5c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac210e5),
	.w1(32'h3b2f5c13),
	.w2(32'h3b788b2d),
	.w3(32'hbaa55154),
	.w4(32'h3b13fd27),
	.w5(32'h398de504),
	.w6(32'hbb6c83ac),
	.w7(32'hba3d6a7c),
	.w8(32'h38dad40b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1bf9d),
	.w1(32'h3971a8f3),
	.w2(32'h399a91aa),
	.w3(32'hb92fb1a4),
	.w4(32'hba96b789),
	.w5(32'hba8c3197),
	.w6(32'h3a42b0b2),
	.w7(32'hbab55022),
	.w8(32'hbb25f21d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e54ef9),
	.w1(32'hbb0506a2),
	.w2(32'hbb3c3200),
	.w3(32'hba8c905c),
	.w4(32'hba51d45f),
	.w5(32'hbb69a5e1),
	.w6(32'h3aa2d139),
	.w7(32'h3aae84de),
	.w8(32'hbaa11881),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa13aad),
	.w1(32'h3b68dbf0),
	.w2(32'hb9d2d04f),
	.w3(32'h3c07adee),
	.w4(32'h3c7a1517),
	.w5(32'h3c05d6ca),
	.w6(32'h3b40583d),
	.w7(32'h3c70e598),
	.w8(32'h3c8b02c6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7af55),
	.w1(32'h3bc5845b),
	.w2(32'h3c5175db),
	.w3(32'hbc113dff),
	.w4(32'h3aed279f),
	.w5(32'h3c0a0736),
	.w6(32'hbc29a45b),
	.w7(32'hb80997ee),
	.w8(32'h3be3a7f2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc51aa),
	.w1(32'hbbfc0620),
	.w2(32'h3b3e646f),
	.w3(32'hbc1e9861),
	.w4(32'hbc24c4bb),
	.w5(32'h39b60016),
	.w6(32'hbbe65fe7),
	.w7(32'hbc38ef70),
	.w8(32'hbbe3c02b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2bada),
	.w1(32'h3b467d17),
	.w2(32'h3b31209d),
	.w3(32'hbaca6794),
	.w4(32'h3aa25569),
	.w5(32'h3af7a1e9),
	.w6(32'hbaac1f08),
	.w7(32'h3aadd26d),
	.w8(32'h3ace5b43),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a667c),
	.w1(32'hbac6d4c9),
	.w2(32'hbafbe64c),
	.w3(32'hba3b2e24),
	.w4(32'hba8b68d4),
	.w5(32'h3a31d5d0),
	.w6(32'hb9e7a554),
	.w7(32'hb987af22),
	.w8(32'h3acdeab5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dcb103),
	.w1(32'h3a1ce916),
	.w2(32'h39be59d9),
	.w3(32'h3a86b27e),
	.w4(32'h3a857095),
	.w5(32'hbb10b00f),
	.w6(32'h3b11ac08),
	.w7(32'h3a8d871e),
	.w8(32'hbb1afb46),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf64923),
	.w1(32'hbb08669e),
	.w2(32'hbacd223c),
	.w3(32'hbb907a20),
	.w4(32'hbb3fece2),
	.w5(32'h3a1a620f),
	.w6(32'hbb9c0b58),
	.w7(32'hbb2e469a),
	.w8(32'hba876585),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd0a31),
	.w1(32'hbac43a4f),
	.w2(32'h3a53e217),
	.w3(32'hbbdb3a97),
	.w4(32'hbbe6c6c4),
	.w5(32'hbc49b119),
	.w6(32'hbbe4574d),
	.w7(32'hbc4e36f2),
	.w8(32'hbc863b79),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0feba),
	.w1(32'h3bb5aaff),
	.w2(32'h3bf94003),
	.w3(32'hbb2fd891),
	.w4(32'h3abaef72),
	.w5(32'h3b7d0e74),
	.w6(32'hbbed7606),
	.w7(32'hbb3fe8d4),
	.w8(32'h3a7dd912),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19f378),
	.w1(32'h3b939e71),
	.w2(32'h3b6b50bb),
	.w3(32'h3a0f1e30),
	.w4(32'h3b570f6c),
	.w5(32'hbb18a66f),
	.w6(32'h3a1e6303),
	.w7(32'h3b40adf4),
	.w8(32'hbb9eef74),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc660a),
	.w1(32'h3b8f224d),
	.w2(32'h3bad3abe),
	.w3(32'h3b51a6c7),
	.w4(32'h3b93fe1c),
	.w5(32'h3b7825d1),
	.w6(32'hb8ef7604),
	.w7(32'h3a30bd43),
	.w8(32'hbaceed9e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c460d11),
	.w1(32'hbbefc9c4),
	.w2(32'hbc7ce6af),
	.w3(32'h3c6c2374),
	.w4(32'h39c5d59f),
	.w5(32'hbc12a910),
	.w6(32'h3c88b6db),
	.w7(32'h3b9d2b65),
	.w8(32'hbc04964c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba145c2c),
	.w1(32'hba48839b),
	.w2(32'hb9f7ca62),
	.w3(32'hb8f39145),
	.w4(32'h3a4a9190),
	.w5(32'h3a8aaf56),
	.w6(32'h386296d3),
	.w7(32'h3aaf86de),
	.w8(32'h3a4e6efa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fa463),
	.w1(32'h3b90cc2a),
	.w2(32'h3b9fe578),
	.w3(32'h3b4befc9),
	.w4(32'h3b66cdc0),
	.w5(32'hbac67388),
	.w6(32'h3b402826),
	.w7(32'h39d41983),
	.w8(32'hbb45aa93),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b3c1a),
	.w1(32'h3a37e264),
	.w2(32'hb8f699da),
	.w3(32'h3ad90814),
	.w4(32'h3ab52739),
	.w5(32'h3a97971c),
	.w6(32'h3abb3389),
	.w7(32'h3abe717b),
	.w8(32'h3a122745),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ffca4),
	.w1(32'hb959a708),
	.w2(32'hb99bc817),
	.w3(32'hba5d31ed),
	.w4(32'hba4c6d3a),
	.w5(32'h38b2c301),
	.w6(32'h3ab2f177),
	.w7(32'h3aaea02d),
	.w8(32'hba00f2b5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ff03f),
	.w1(32'hba1698e4),
	.w2(32'hbb0df733),
	.w3(32'h3b2215e6),
	.w4(32'hba2a0e52),
	.w5(32'hbb0a82ee),
	.w6(32'h3ac4f553),
	.w7(32'hba20a874),
	.w8(32'hba85ac2b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7f6e5),
	.w1(32'hbba9deb0),
	.w2(32'hbc2d1aa0),
	.w3(32'h3bc208a6),
	.w4(32'hbb80d6b5),
	.w5(32'hbc0fd3cf),
	.w6(32'h3ae9807a),
	.w7(32'hbb9a574c),
	.w8(32'hbc4c260c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47084a),
	.w1(32'hbb52554a),
	.w2(32'hbb19ba00),
	.w3(32'hba83bed1),
	.w4(32'hbb143332),
	.w5(32'hbb72a68e),
	.w6(32'h394eacdc),
	.w7(32'hb8411456),
	.w8(32'hbb1db528),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d64ed),
	.w1(32'hb9a7d6b2),
	.w2(32'h3a9ba836),
	.w3(32'hb94b2906),
	.w4(32'h3a1e69ac),
	.w5(32'hba1d088b),
	.w6(32'h39192583),
	.w7(32'h3a6ea8af),
	.w8(32'h39502d2e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996c5c4),
	.w1(32'hb8912824),
	.w2(32'hb9251289),
	.w3(32'hb94ed6bf),
	.w4(32'hb910e97e),
	.w5(32'hba9a950c),
	.w6(32'h389a61ac),
	.w7(32'h39d07bf7),
	.w8(32'hbad4cf66),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab80cca),
	.w1(32'hbadabd4d),
	.w2(32'hba304d14),
	.w3(32'hbb18e87b),
	.w4(32'hbb09144e),
	.w5(32'h3aa6f5ab),
	.w6(32'hbad62bd7),
	.w7(32'hba887231),
	.w8(32'h3aaae11d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4cecd),
	.w1(32'h3af498d9),
	.w2(32'h3ad26891),
	.w3(32'h3abe5fb0),
	.w4(32'h3ad15a27),
	.w5(32'h3a89074d),
	.w6(32'h3b26d677),
	.w7(32'h3af4c67a),
	.w8(32'h3b12fb4a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392fd934),
	.w1(32'h397d4e2a),
	.w2(32'h3a9ab956),
	.w3(32'hbaa983ab),
	.w4(32'h3983262b),
	.w5(32'hbae35cea),
	.w6(32'h3a8fe520),
	.w7(32'h3b2218d2),
	.w8(32'hbaeb8083),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a5e1b),
	.w1(32'hba3cdd10),
	.w2(32'hbaf07714),
	.w3(32'h3a71a288),
	.w4(32'hbaee6ae8),
	.w5(32'hbb831bfd),
	.w6(32'h3b337048),
	.w7(32'hbb1a90e7),
	.w8(32'hbb95f67d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb775cd),
	.w1(32'hbbac09b1),
	.w2(32'h3a640bdd),
	.w3(32'hba08775a),
	.w4(32'hbbcfbe0a),
	.w5(32'hba1e417a),
	.w6(32'h3710289f),
	.w7(32'hbbdda3ea),
	.w8(32'hbab3f4b4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938fdc3),
	.w1(32'h39516c08),
	.w2(32'h399a2a00),
	.w3(32'hbad78296),
	.w4(32'hbb0d02d8),
	.w5(32'hb987ad7d),
	.w6(32'h3ab4c145),
	.w7(32'hb9b1de1b),
	.w8(32'h3a5435e8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38849c8c),
	.w1(32'h3a680151),
	.w2(32'h3a23920e),
	.w3(32'hb97c616e),
	.w4(32'h39aa7d47),
	.w5(32'hba6dee2c),
	.w6(32'h3a46ed91),
	.w7(32'h3a4f6ff8),
	.w8(32'hba22f3ed),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56b47f),
	.w1(32'h39cc092e),
	.w2(32'h3ab90f47),
	.w3(32'h39c11465),
	.w4(32'h3a3eedb5),
	.w5(32'hb9fcfb42),
	.w6(32'h3a6cd007),
	.w7(32'h3a882203),
	.w8(32'h39e7f1df),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87ab49),
	.w1(32'hbab6b392),
	.w2(32'hba8460ec),
	.w3(32'hba8549ef),
	.w4(32'hbab44c5b),
	.w5(32'h3a14e1b2),
	.w6(32'h3a1d2ba9),
	.w7(32'hba5d770a),
	.w8(32'hb9545e1a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa28d95),
	.w1(32'hbbf04e47),
	.w2(32'hbc1f151b),
	.w3(32'h3c088ce1),
	.w4(32'hbb83d808),
	.w5(32'hbaddf713),
	.w6(32'h3b9fe895),
	.w7(32'hbc3c61cd),
	.w8(32'hbc736750),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48e696),
	.w1(32'h3aece94b),
	.w2(32'hbc079950),
	.w3(32'h3c048d97),
	.w4(32'hbac88fcb),
	.w5(32'hbc75e48d),
	.w6(32'h3c2593b5),
	.w7(32'h3b92a22b),
	.w8(32'hbbf02532),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba952d8),
	.w1(32'hbb385b72),
	.w2(32'hbbe70259),
	.w3(32'h3932030f),
	.w4(32'hbaba8ab8),
	.w5(32'hbb92765f),
	.w6(32'h3b4ee3fc),
	.w7(32'h3aff4608),
	.w8(32'hbbf7618d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c321a0),
	.w1(32'h3c0ce13c),
	.w2(32'h3c38f77f),
	.w3(32'hbbf03da3),
	.w4(32'hbb1a392a),
	.w5(32'h3b2bb938),
	.w6(32'hbc4e0ba7),
	.w7(32'hbbd61d0f),
	.w8(32'h399468f7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac37b6),
	.w1(32'hba120672),
	.w2(32'hb9a46cea),
	.w3(32'hbaa0b97e),
	.w4(32'hba8d9d6e),
	.w5(32'h39047a49),
	.w6(32'hbaf983e0),
	.w7(32'hbabb1f49),
	.w8(32'h3912ae23),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990192d),
	.w1(32'h3901e05c),
	.w2(32'h3ae8431c),
	.w3(32'h3a46dd26),
	.w4(32'hb642675a),
	.w5(32'h3a2bd0ea),
	.w6(32'h3ade3052),
	.w7(32'h3aa0042a),
	.w8(32'hb81d5d28),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984e426),
	.w1(32'hba4cac05),
	.w2(32'h367c0876),
	.w3(32'h39529097),
	.w4(32'h3a01c731),
	.w5(32'hbac5e56a),
	.w6(32'h39907c87),
	.w7(32'h3a21493d),
	.w8(32'hba09a4a6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37a713),
	.w1(32'hbabbd169),
	.w2(32'hbb165e03),
	.w3(32'h3a84726e),
	.w4(32'hbaaed555),
	.w5(32'hbae242cf),
	.w6(32'h3af3d144),
	.w7(32'h388acc80),
	.w8(32'hbaa620b3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a878766),
	.w1(32'h3a8fba76),
	.w2(32'h39becb8d),
	.w3(32'h39f3bfab),
	.w4(32'hb92ddf75),
	.w5(32'hbad70614),
	.w6(32'h3a6a3e81),
	.w7(32'h3a1e8d07),
	.w8(32'hbad5d0eb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d59d1),
	.w1(32'hbbd1350f),
	.w2(32'hbbdcbca0),
	.w3(32'h3a8bdea1),
	.w4(32'hb932b8b3),
	.w5(32'hbb6ac133),
	.w6(32'h3b029179),
	.w7(32'h39861816),
	.w8(32'hbb0f4de6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c378a8a),
	.w1(32'h3b0e7905),
	.w2(32'hbbfbb197),
	.w3(32'h3c1358c2),
	.w4(32'hba656a42),
	.w5(32'hbbe32728),
	.w6(32'h3c1c3c59),
	.w7(32'h3b0b256d),
	.w8(32'hbba5cb2b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ebd0a),
	.w1(32'h3b03cea2),
	.w2(32'h3b8000c2),
	.w3(32'hbb60c8b1),
	.w4(32'h3a9c0cc6),
	.w5(32'h3af10ac9),
	.w6(32'hbb6012c5),
	.w7(32'hbb26edf1),
	.w8(32'hbadd3970),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bcbc9),
	.w1(32'hbbb01907),
	.w2(32'hbbabb958),
	.w3(32'hbaacd5d0),
	.w4(32'hbb8541f3),
	.w5(32'hbb853153),
	.w6(32'hbb38d4b2),
	.w7(32'hbb6a1e3f),
	.w8(32'hbbc1bbc3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b822ca2),
	.w1(32'hbb4836f3),
	.w2(32'hbb5f1d01),
	.w3(32'h3b3a1441),
	.w4(32'h3b3871e0),
	.w5(32'hbb8addd1),
	.w6(32'h3acb2d08),
	.w7(32'h37cc69fc),
	.w8(32'hbc2618d2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cc8e1),
	.w1(32'hbb9e87b3),
	.w2(32'hbaa892cf),
	.w3(32'hbbc1de01),
	.w4(32'hbbef0cb3),
	.w5(32'hbabcb4f7),
	.w6(32'hbc295c17),
	.w7(32'hbc015324),
	.w8(32'hbb5a5c6e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a706ea0),
	.w1(32'hbb898024),
	.w2(32'hbbaa79b7),
	.w3(32'h3aa1fb5b),
	.w4(32'hbaea3e7d),
	.w5(32'hbb6f774a),
	.w6(32'h3ac03b7f),
	.w7(32'hbaed67a9),
	.w8(32'hbbac08e6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f41c0),
	.w1(32'hb9dfd8f8),
	.w2(32'hb9bcf3d5),
	.w3(32'hba550e5a),
	.w4(32'hba61b47d),
	.w5(32'h39b7a500),
	.w6(32'hba5843eb),
	.w7(32'hb9f30c43),
	.w8(32'h3a0b8d8a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1db83e),
	.w1(32'h3aa52d71),
	.w2(32'hbabb80b6),
	.w3(32'h39bbd0ec),
	.w4(32'hba9efffd),
	.w5(32'h39d757fc),
	.w6(32'h3a23cf55),
	.w7(32'hbaa98e16),
	.w8(32'h39eb1c53),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390726cf),
	.w1(32'hba3f7666),
	.w2(32'hb9e6ae90),
	.w3(32'hb9d2c070),
	.w4(32'hb9cf85f4),
	.w5(32'hba845e3c),
	.w6(32'h3805e57d),
	.w7(32'h37bcc20b),
	.w8(32'hba90788b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9ca99),
	.w1(32'hb972cd8c),
	.w2(32'h3adb9a30),
	.w3(32'hbb30afe9),
	.w4(32'hba02e57b),
	.w5(32'h3a1fa4d9),
	.w6(32'hb9d632d4),
	.w7(32'h3996c741),
	.w8(32'h394d487f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ba38c),
	.w1(32'h3b5656f0),
	.w2(32'h3b24ad4d),
	.w3(32'hbb6954e3),
	.w4(32'h3a6bb4e3),
	.w5(32'h3b0aca4e),
	.w6(32'hbb84b2ab),
	.w7(32'hbade6902),
	.w8(32'h3b4d9eab),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f90e2),
	.w1(32'hbac220f0),
	.w2(32'hba92bcaf),
	.w3(32'hba056083),
	.w4(32'h3a03d4dc),
	.w5(32'h3a54a29f),
	.w6(32'hba4e49a4),
	.w7(32'hba868843),
	.w8(32'hb98cbe00),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d89f9),
	.w1(32'h3b97126c),
	.w2(32'h3b638b5b),
	.w3(32'h3b29b092),
	.w4(32'h3a5a9c62),
	.w5(32'hbb744f15),
	.w6(32'h39f48f8b),
	.w7(32'h3b45d86b),
	.w8(32'h39e8a541),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc156e2),
	.w1(32'hbabe4888),
	.w2(32'hbbf4cfed),
	.w3(32'h3b8a0993),
	.w4(32'hbb2df6f0),
	.w5(32'hbbf2663e),
	.w6(32'h3bb7a296),
	.w7(32'hbb4e3bd2),
	.w8(32'hbbfae7de),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0186f),
	.w1(32'hbb55a74a),
	.w2(32'hb9b3e268),
	.w3(32'hbb852263),
	.w4(32'hbb308d42),
	.w5(32'h3a67e3cd),
	.w6(32'hbb09ffb4),
	.w7(32'hbb0c41ae),
	.w8(32'hb9f18760),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba30ac3),
	.w1(32'hbb92a488),
	.w2(32'hbca4193d),
	.w3(32'h3c3da677),
	.w4(32'h3bc41069),
	.w5(32'hbc06007d),
	.w6(32'h3c543f11),
	.w7(32'h3bb36e87),
	.w8(32'hbc18e1bb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a5a21),
	.w1(32'hbae86ccd),
	.w2(32'h3a78da77),
	.w3(32'hbb9b1e5a),
	.w4(32'hbab4d77d),
	.w5(32'h3acac71f),
	.w6(32'hbbd4b6d7),
	.w7(32'hbb59434e),
	.w8(32'h3a04d06d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3718a),
	.w1(32'hbb9fc251),
	.w2(32'hbbaea8a2),
	.w3(32'h3b7d560a),
	.w4(32'hbb97a281),
	.w5(32'hbc2572c4),
	.w6(32'h3b32b4de),
	.w7(32'hbc074fb4),
	.w8(32'hbc676c9b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae45864),
	.w1(32'h3a64bb68),
	.w2(32'h3b446a65),
	.w3(32'h3a263f30),
	.w4(32'h3a8231da),
	.w5(32'h3aa0ff94),
	.w6(32'hbb1c38c3),
	.w7(32'hbb422042),
	.w8(32'h391af645),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80dfc0),
	.w1(32'h3a641af0),
	.w2(32'h3b50c7da),
	.w3(32'hbb88f434),
	.w4(32'hbac49c0d),
	.w5(32'h3b4acb71),
	.w6(32'hbb8a28df),
	.w7(32'hbb85ec9f),
	.w8(32'hba973c32),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29f160),
	.w1(32'hbb1d3f24),
	.w2(32'hbb16469d),
	.w3(32'hba6b114d),
	.w4(32'h39d239ab),
	.w5(32'hbba08148),
	.w6(32'hbaadab8d),
	.w7(32'hba8a2a32),
	.w8(32'hbbbc7759),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8144ef),
	.w1(32'h3b3affa9),
	.w2(32'hb9f83883),
	.w3(32'h3be8e07c),
	.w4(32'h3b0bcb77),
	.w5(32'hbbc5cfbb),
	.w6(32'h3abf0ccb),
	.w7(32'hbb684d50),
	.w8(32'hbc53f809),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab86ebe),
	.w1(32'hbbe4d191),
	.w2(32'hbb8e5b72),
	.w3(32'h3b2bdf81),
	.w4(32'h3b42d09f),
	.w5(32'h3b574306),
	.w6(32'h3b46968a),
	.w7(32'hb8b85218),
	.w8(32'hbc1cf3f1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd02e2),
	.w1(32'hba3cdbf5),
	.w2(32'hbc1fff9a),
	.w3(32'h3c1f9617),
	.w4(32'h3ba3de31),
	.w5(32'hbbae54dc),
	.w6(32'h3c249e1e),
	.w7(32'h3c8df2b5),
	.w8(32'h3c97793b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7c2a5),
	.w1(32'h3bafae15),
	.w2(32'h3b1c9e98),
	.w3(32'hbb849d37),
	.w4(32'h3c5c5317),
	.w5(32'h3c1da14d),
	.w6(32'hbb6dfa36),
	.w7(32'h3bafe828),
	.w8(32'h3b8af640),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3d550),
	.w1(32'h3c21e57c),
	.w2(32'h3c31212f),
	.w3(32'h39a1582d),
	.w4(32'h3ba25164),
	.w5(32'h3b0e7463),
	.w6(32'hbbb06870),
	.w7(32'hbad2bedf),
	.w8(32'hbab66dbc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba947a5b),
	.w1(32'hbc2a2bf0),
	.w2(32'hbc0b7622),
	.w3(32'h3bc2e994),
	.w4(32'h3bacdcbf),
	.w5(32'hbba35fcb),
	.w6(32'h3bb81d0d),
	.w7(32'h3b8cc7ad),
	.w8(32'hbc0bb1b3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fcc62),
	.w1(32'hba5e3168),
	.w2(32'hbb45ec52),
	.w3(32'hba2234c7),
	.w4(32'hb9720a78),
	.w5(32'hba9a55e9),
	.w6(32'h3a8c5644),
	.w7(32'h39e9aa97),
	.w8(32'hbb4edcd8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd283b5),
	.w1(32'hbb581174),
	.w2(32'hbba376d5),
	.w3(32'h3aaa5f4a),
	.w4(32'h3bb891a8),
	.w5(32'h3b16b6ab),
	.w6(32'h3bb7f52e),
	.w7(32'h3c14e391),
	.w8(32'h3c8b69f4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a50d9),
	.w1(32'hbb275fa8),
	.w2(32'hbb680103),
	.w3(32'hba8811f0),
	.w4(32'hbbdb3b1f),
	.w5(32'hba6fa884),
	.w6(32'h3a3856f4),
	.w7(32'hbbecb1e8),
	.w8(32'hbaf2ba00),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa52fa0),
	.w1(32'h395982ae),
	.w2(32'hb9e4bf2b),
	.w3(32'h3a95f629),
	.w4(32'h3a19b6f0),
	.w5(32'hba9907b5),
	.w6(32'hb9b2058b),
	.w7(32'hba26c2e5),
	.w8(32'hbad4bf57),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad59e17),
	.w1(32'hb71f103f),
	.w2(32'hbb14f0ae),
	.w3(32'h3aa7ec95),
	.w4(32'h3a41eaca),
	.w5(32'h39012c92),
	.w6(32'h3a932a00),
	.w7(32'hb99f375e),
	.w8(32'hba34e933),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd76718),
	.w1(32'h3a72bc4f),
	.w2(32'hbaac1309),
	.w3(32'h3b628acf),
	.w4(32'hba40afff),
	.w5(32'hbbc7c71f),
	.w6(32'h396cbe89),
	.w7(32'hbbaffafe),
	.w8(32'hbc37fe1a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae57e52),
	.w1(32'h3b96b976),
	.w2(32'h3bd45cc4),
	.w3(32'hbb97e027),
	.w4(32'h3a481c2b),
	.w5(32'h3b111764),
	.w6(32'hbbdf4f5f),
	.w7(32'hbb9401a1),
	.w8(32'hba7911d0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7743af),
	.w1(32'hbbb0d5ad),
	.w2(32'h3a79910b),
	.w3(32'hbb372954),
	.w4(32'hbbc843b4),
	.w5(32'h3b02c3ff),
	.w6(32'hbbc86d22),
	.w7(32'hbc25b3c3),
	.w8(32'hbb82db6a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9716c1),
	.w1(32'h3ae8b57c),
	.w2(32'h3b32c1e6),
	.w3(32'hba9ae35a),
	.w4(32'h39cd1f42),
	.w5(32'hba19f7f6),
	.w6(32'hbb666a2a),
	.w7(32'hbb184597),
	.w8(32'hbb62f9de),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2fd71),
	.w1(32'h3b4c0e56),
	.w2(32'h39dcd44d),
	.w3(32'hbba32533),
	.w4(32'hbb0a390f),
	.w5(32'hbaf5203a),
	.w6(32'hb9f198a5),
	.w7(32'h3be3a151),
	.w8(32'h3c2fd1e8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9437a),
	.w1(32'h3ae1327e),
	.w2(32'h3ac8dc1d),
	.w3(32'h3b67cf3e),
	.w4(32'hb8b7c9c0),
	.w5(32'hbb963628),
	.w6(32'hb9df4436),
	.w7(32'hbb727fac),
	.w8(32'hbb82b1af),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bfd56),
	.w1(32'h3b1b2191),
	.w2(32'h3ae48026),
	.w3(32'h39810e7a),
	.w4(32'hba33c80c),
	.w5(32'h382219cf),
	.w6(32'hb9ee80c7),
	.w7(32'hbaca2882),
	.w8(32'hba5d05a2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39990eac),
	.w1(32'h3a941df5),
	.w2(32'h38ed6bbb),
	.w3(32'h3a6187b3),
	.w4(32'h3aaff3fb),
	.w5(32'hb9770bd2),
	.w6(32'h3aabbb86),
	.w7(32'h3a919d07),
	.w8(32'hb9c562d4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89acd00),
	.w1(32'hba33fec1),
	.w2(32'hbad1a5c9),
	.w3(32'h39883a31),
	.w4(32'hbaa1e3c8),
	.w5(32'h39f2ea2f),
	.w6(32'hb9c341e6),
	.w7(32'hbac67b5d),
	.w8(32'h37f47dc1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b9501),
	.w1(32'hb91510cb),
	.w2(32'h3a2775c1),
	.w3(32'h3a2b01e0),
	.w4(32'h3b031d4e),
	.w5(32'hb9dcaa87),
	.w6(32'hb909ea5a),
	.w7(32'h3a8e68a4),
	.w8(32'hba15a9f2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df02e5),
	.w1(32'h3a9ced47),
	.w2(32'h3b125328),
	.w3(32'h3ac2b290),
	.w4(32'h3b225925),
	.w5(32'h3ab6801d),
	.w6(32'h3a67cc43),
	.w7(32'h3aa10b7e),
	.w8(32'hbaa6038a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad495f5),
	.w1(32'h3b372fe3),
	.w2(32'h3b7dfc1f),
	.w3(32'hbb2230b1),
	.w4(32'h3a528548),
	.w5(32'h3aeb5489),
	.w6(32'hbc070a60),
	.w7(32'hbba96942),
	.w8(32'hbb12beff),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8975328),
	.w1(32'hbb0c5750),
	.w2(32'hbb897387),
	.w3(32'hba03aafb),
	.w4(32'hba2a69b5),
	.w5(32'hba99f357),
	.w6(32'h3a54f61a),
	.w7(32'h3abebd59),
	.w8(32'hb986f389),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50a1c0),
	.w1(32'hba1698e5),
	.w2(32'hba082815),
	.w3(32'h3b4bbc90),
	.w4(32'h3a998fd9),
	.w5(32'h3a37c66c),
	.w6(32'h3acdf8fb),
	.w7(32'h3adc9c49),
	.w8(32'hba461867),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba0d78),
	.w1(32'h3b9e58f8),
	.w2(32'h3c15795c),
	.w3(32'hbaf830af),
	.w4(32'hbacd2fb9),
	.w5(32'h3b9b3b2c),
	.w6(32'hbb5bb7db),
	.w7(32'hbb6ce963),
	.w8(32'h3add46e6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86d712f),
	.w1(32'h3a86e37a),
	.w2(32'h3a7e2867),
	.w3(32'h3a629407),
	.w4(32'h3a8b42c3),
	.w5(32'hba2cb63e),
	.w6(32'h3aa50928),
	.w7(32'h3aaad3aa),
	.w8(32'h38ad7a21),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9456e4c),
	.w1(32'h3a0e2fa0),
	.w2(32'hb93880d0),
	.w3(32'hb9f8ed2b),
	.w4(32'hba64dc58),
	.w5(32'h3ab26471),
	.w6(32'hb9fb65bb),
	.w7(32'hb9fbe8e1),
	.w8(32'h3abab99c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad57160),
	.w1(32'h3ae4177c),
	.w2(32'h3aaa42a0),
	.w3(32'h3afb402b),
	.w4(32'h3ae0798a),
	.w5(32'hb999c94b),
	.w6(32'h3b33b094),
	.w7(32'h3acb3c97),
	.w8(32'hba7bbc32),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d29b5c),
	.w1(32'h39dad3b2),
	.w2(32'h3a417152),
	.w3(32'h36809386),
	.w4(32'hb9d6fc43),
	.w5(32'h3a6a4d77),
	.w6(32'hb95fbfac),
	.w7(32'hba09aeb2),
	.w8(32'h3a64ac2d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3daef3),
	.w1(32'h3b20ad64),
	.w2(32'h3a349adc),
	.w3(32'h3b063aad),
	.w4(32'hbb37226e),
	.w5(32'hbc535ac7),
	.w6(32'h3b8f8f5b),
	.w7(32'h3b11aa88),
	.w8(32'hbbeea9f0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dbda2),
	.w1(32'hbad2f0d7),
	.w2(32'hbb03f9c3),
	.w3(32'h3b3feca2),
	.w4(32'hbba166b7),
	.w5(32'hbae604ed),
	.w6(32'hba9e92da),
	.w7(32'hbbf51d09),
	.w8(32'hbc0556f0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393afbbb),
	.w1(32'hbaa5159a),
	.w2(32'hba2ee837),
	.w3(32'h3aa0e2b9),
	.w4(32'h39dd9d0a),
	.w5(32'hbae48029),
	.w6(32'hb806af1e),
	.w7(32'h388f3540),
	.w8(32'hbac33344),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5f6ee),
	.w1(32'hba047dec),
	.w2(32'hbb0b208e),
	.w3(32'h39cc34a2),
	.w4(32'hba185142),
	.w5(32'hbb4ba01c),
	.w6(32'h393ede6a),
	.w7(32'h3a3bab03),
	.w8(32'hba86aa87),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba143bdb),
	.w1(32'h3a088c0a),
	.w2(32'h3a0b8d05),
	.w3(32'hba5f69b2),
	.w4(32'h390f3c10),
	.w5(32'hb9f27a17),
	.w6(32'hba0b3c25),
	.w7(32'hb8839032),
	.w8(32'hba095da1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad1eec),
	.w1(32'hba3a2a0f),
	.w2(32'hba46299b),
	.w3(32'h3aea7cc5),
	.w4(32'hba2ef204),
	.w5(32'hbb368a61),
	.w6(32'h3aec3e93),
	.w7(32'hbaedb90c),
	.w8(32'hbb8a871f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57763d),
	.w1(32'h39591654),
	.w2(32'h3a140660),
	.w3(32'hba94a0ec),
	.w4(32'hbb233a09),
	.w5(32'h3a0fad29),
	.w6(32'h38b74e25),
	.w7(32'hbb86e7d3),
	.w8(32'hbab2fd98),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc18b25),
	.w1(32'hbb873040),
	.w2(32'hbb9f7a16),
	.w3(32'h3bd5fda4),
	.w4(32'hb9efa0bd),
	.w5(32'hbbb2cb2b),
	.w6(32'h3afac2ac),
	.w7(32'hbb96fd8c),
	.w8(32'hbc6c19ef),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944e188),
	.w1(32'h3b3e25c6),
	.w2(32'h3b5fee98),
	.w3(32'hbaf80e1a),
	.w4(32'hb96a0ed5),
	.w5(32'h3a09482f),
	.w6(32'hbb64b373),
	.w7(32'hbb704b60),
	.w8(32'hbafce5bb),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab56257),
	.w1(32'hba798a22),
	.w2(32'hbb19efc3),
	.w3(32'h3b06923c),
	.w4(32'h397177bd),
	.w5(32'hbb177713),
	.w6(32'hbb6a4663),
	.w7(32'hbb92a39c),
	.w8(32'hbbfe271c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6040e),
	.w1(32'hbbe18ba1),
	.w2(32'hbc0e86cc),
	.w3(32'h3b9a5951),
	.w4(32'h39e0ab08),
	.w5(32'hbbc1c38e),
	.w6(32'h3b7a2139),
	.w7(32'h3ae23422),
	.w8(32'hbba44bbf),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a455220),
	.w1(32'h3ab7fe70),
	.w2(32'hbb054997),
	.w3(32'h3add25b2),
	.w4(32'h3b1e74a7),
	.w5(32'hb8395b56),
	.w6(32'h3b3a3510),
	.w7(32'h3b69cf5d),
	.w8(32'h3b9ecc45),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b5e7e),
	.w1(32'h3b8e2f7b),
	.w2(32'h3b154c43),
	.w3(32'h3bae1ace),
	.w4(32'h3b2649ae),
	.w5(32'hba2de66b),
	.w6(32'hb9c39bcd),
	.w7(32'hbb12cd37),
	.w8(32'hbbceaa63),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f3d75),
	.w1(32'h3ac4c18f),
	.w2(32'hb8d2858d),
	.w3(32'h392afba3),
	.w4(32'hba6698ba),
	.w5(32'hb9e3f20a),
	.w6(32'hb9d1a2ad),
	.w7(32'hbacd1eef),
	.w8(32'hba73eab5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3edb05),
	.w1(32'h3c057295),
	.w2(32'h3c2c8faf),
	.w3(32'h3bed7392),
	.w4(32'hbb3e345c),
	.w5(32'h39cbd7fa),
	.w6(32'h3b929e3c),
	.w7(32'hbbefaeb8),
	.w8(32'hbb86939e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea53a),
	.w1(32'h3b3d9bef),
	.w2(32'h3b15dccd),
	.w3(32'hb921101b),
	.w4(32'hbaced399),
	.w5(32'h3b4423d4),
	.w6(32'hbb6186b3),
	.w7(32'hbb6c009d),
	.w8(32'h3a4a5658),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b21f94),
	.w1(32'hb9f89c70),
	.w2(32'hb8d6fb8d),
	.w3(32'hb79d0be5),
	.w4(32'hb9f1159b),
	.w5(32'hba7bbf9e),
	.w6(32'h391e2fc6),
	.w7(32'h394f6fd6),
	.w8(32'hba71318a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba588764),
	.w1(32'hba40239f),
	.w2(32'hba1dabc1),
	.w3(32'hba6e5a7b),
	.w4(32'hba9e8cec),
	.w5(32'hb8c39177),
	.w6(32'hba8e11e6),
	.w7(32'hbaaa9a48),
	.w8(32'hb9260208),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f976f0),
	.w1(32'h39c495d8),
	.w2(32'h38287751),
	.w3(32'hb95a6fdd),
	.w4(32'hb97de3a1),
	.w5(32'hb843a0b0),
	.w6(32'hba66af77),
	.w7(32'hbb19f344),
	.w8(32'h39c1ef78),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3680056f),
	.w1(32'h3bc963fb),
	.w2(32'h3ba7314b),
	.w3(32'hbb85adf0),
	.w4(32'h3b1b9a79),
	.w5(32'h3b0f3ba8),
	.w6(32'hbbd737d0),
	.w7(32'hbb8bed24),
	.w8(32'h39c9bc82),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b165477),
	.w1(32'h3a470560),
	.w2(32'h3a03cfab),
	.w3(32'h3a9f0844),
	.w4(32'hbaa0c1b8),
	.w5(32'hbaf6681d),
	.w6(32'h39cfe269),
	.w7(32'hbb3cd43b),
	.w8(32'hbb76edd1),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b3652),
	.w1(32'h3a478f37),
	.w2(32'h3a6f41eb),
	.w3(32'h39a73d8f),
	.w4(32'hb8cc085e),
	.w5(32'h39f10033),
	.w6(32'h3a947e8e),
	.w7(32'h3a51f920),
	.w8(32'h39a1f016),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd535e0),
	.w1(32'h3b200d0a),
	.w2(32'h3ae46a26),
	.w3(32'h3b8571af),
	.w4(32'hbac86452),
	.w5(32'hba95450b),
	.w6(32'hba80eda0),
	.w7(32'hbbe7cdd4),
	.w8(32'hbc05a9fd),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd2118),
	.w1(32'h3bd5fdaa),
	.w2(32'h3bd61cfe),
	.w3(32'h3b52068e),
	.w4(32'h3b20294b),
	.w5(32'h39a9af6e),
	.w6(32'hbb0aa26b),
	.w7(32'hbb654375),
	.w8(32'hbb4f5986),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b33ad),
	.w1(32'hbb20d326),
	.w2(32'hbbb1f93d),
	.w3(32'h3c39d581),
	.w4(32'h3b4781a9),
	.w5(32'hba8b79bc),
	.w6(32'h3c0943db),
	.w7(32'h3ab0f3da),
	.w8(32'hbbc5cc31),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2633a),
	.w1(32'hbbd61197),
	.w2(32'h3ba76452),
	.w3(32'h3b5b46bd),
	.w4(32'hbc23eaec),
	.w5(32'h36b89740),
	.w6(32'hbc0596ea),
	.w7(32'hbc84db27),
	.w8(32'hbbe2c24f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9843801),
	.w1(32'h3ae193a0),
	.w2(32'h3a6e6d2d),
	.w3(32'hba9aa0c7),
	.w4(32'hb9488e7e),
	.w5(32'h3a8eeb2b),
	.w6(32'hbad9a419),
	.w7(32'hbb72580a),
	.w8(32'hbae261c8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada6b8b),
	.w1(32'hbb86f60c),
	.w2(32'hbb5c89a1),
	.w3(32'h39485f2b),
	.w4(32'hba6343db),
	.w5(32'hbb30172a),
	.w6(32'h3997b2a7),
	.w7(32'hbaefd148),
	.w8(32'hbb91c669),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61bde6),
	.w1(32'h3a2aa148),
	.w2(32'h3b4a99ed),
	.w3(32'hbb7de383),
	.w4(32'hba8d0dd7),
	.w5(32'h3b81e3f9),
	.w6(32'hbbb41f4b),
	.w7(32'hbb4b1ac2),
	.w8(32'h3b210599),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13aa38),
	.w1(32'hba5835ed),
	.w2(32'h3b325d2d),
	.w3(32'hbaa6116a),
	.w4(32'hba4162d9),
	.w5(32'h3b8b9b64),
	.w6(32'hbb683944),
	.w7(32'hbb55df37),
	.w8(32'h38e6dd8e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb880f269),
	.w1(32'h3bb40cc0),
	.w2(32'h3be3b76b),
	.w3(32'hb99f5a8c),
	.w4(32'h3b6d67e3),
	.w5(32'h3bc2a6bc),
	.w6(32'hb89e1fc6),
	.w7(32'h3b484ca6),
	.w8(32'h3b89cc16),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65ad4e),
	.w1(32'hbb43a7a0),
	.w2(32'hbaf78a5a),
	.w3(32'h3b6fdb6f),
	.w4(32'h3a9daf2a),
	.w5(32'h3a5d0e53),
	.w6(32'h3a981ff5),
	.w7(32'h39a5ea35),
	.w8(32'h3ad58d47),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b273db7),
	.w1(32'h3b5d4dc1),
	.w2(32'h3b16264f),
	.w3(32'h3a8238df),
	.w4(32'h3a709353),
	.w5(32'h3b18ad52),
	.w6(32'h3ac73a58),
	.w7(32'h3ac59430),
	.w8(32'h3b00d3ae),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfc55c),
	.w1(32'h3a800bac),
	.w2(32'h3a8a6727),
	.w3(32'h3b9aee69),
	.w4(32'h39996f87),
	.w5(32'hbb09f305),
	.w6(32'h3b39cf06),
	.w7(32'hbabb4a6c),
	.w8(32'hbbc6c906),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ad916),
	.w1(32'hbae2dc4a),
	.w2(32'hb88c3b13),
	.w3(32'hbab1f753),
	.w4(32'hbac4e896),
	.w5(32'hba91a75e),
	.w6(32'hb9d44600),
	.w7(32'hba4a2544),
	.w8(32'hb9993fe6),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ba4be),
	.w1(32'h3a891cc3),
	.w2(32'h3b5007e1),
	.w3(32'hbb2b0c7b),
	.w4(32'hbb2c3574),
	.w5(32'h3a13f0dc),
	.w6(32'hbb4a9ed1),
	.w7(32'hbae0fffb),
	.w8(32'h3add6cf4),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909fefb),
	.w1(32'h38b16b89),
	.w2(32'hbaa5a4a2),
	.w3(32'h38789d1f),
	.w4(32'hba21b43c),
	.w5(32'h3a9a7f25),
	.w6(32'h3986f326),
	.w7(32'h39dda46a),
	.w8(32'h3a919e2a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16aeed),
	.w1(32'h3b18e181),
	.w2(32'h3a1224a1),
	.w3(32'h3b9bffee),
	.w4(32'h3a9932c4),
	.w5(32'hbaeff506),
	.w6(32'h3b6f9308),
	.w7(32'hb99481ee),
	.w8(32'hbb7b921f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bbdb9),
	.w1(32'hba9cae81),
	.w2(32'hba6b917c),
	.w3(32'hbab14de1),
	.w4(32'hba943c11),
	.w5(32'h3a0dead1),
	.w6(32'hba96d33c),
	.w7(32'hba977b10),
	.w8(32'h3949de3b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36df4ca5),
	.w1(32'hba002022),
	.w2(32'hbaa3bbe3),
	.w3(32'h3aaf4bbc),
	.w4(32'h3a10418a),
	.w5(32'h3a990675),
	.w6(32'h3a5fd5f7),
	.w7(32'h393bf382),
	.w8(32'h3b1c94c7),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46f7aa),
	.w1(32'h3b7a1d18),
	.w2(32'h3bdbf046),
	.w3(32'hb9e53ea9),
	.w4(32'h3b3f16aa),
	.w5(32'h3b240b70),
	.w6(32'hbb353fd7),
	.w7(32'h3a051a68),
	.w8(32'hbad843ba),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d72a1),
	.w1(32'h3c13f91f),
	.w2(32'h3bd86e82),
	.w3(32'h3c095278),
	.w4(32'h3b3ed760),
	.w5(32'hba9bb49e),
	.w6(32'h3a1ce7db),
	.w7(32'hba066c07),
	.w8(32'hbb86485e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8565c),
	.w1(32'h398b2b24),
	.w2(32'hba7835d1),
	.w3(32'hb93d8379),
	.w4(32'h3a22082a),
	.w5(32'h39fffde7),
	.w6(32'h3a5a840d),
	.w7(32'h3a94002f),
	.w8(32'h3a4acd5e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c3754),
	.w1(32'hbb679a53),
	.w2(32'hbb440d0c),
	.w3(32'hbac8b98d),
	.w4(32'hbabcd706),
	.w5(32'hba435458),
	.w6(32'hbb41adb3),
	.w7(32'hbb89f68b),
	.w8(32'hbbd30a0e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bcdc7b),
	.w1(32'hbb71020f),
	.w2(32'hbb0f718a),
	.w3(32'h3a91aefd),
	.w4(32'hbb3d7a28),
	.w5(32'hbad4b7e9),
	.w6(32'hbb9460dc),
	.w7(32'hbba0a98f),
	.w8(32'hbb806f7b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ed817),
	.w1(32'hbb3efc32),
	.w2(32'hbb3fd106),
	.w3(32'h3b1dd67d),
	.w4(32'hbba7c7d3),
	.w5(32'h3a1527c1),
	.w6(32'hbb38374f),
	.w7(32'hbb28bc2e),
	.w8(32'hbbdd7147),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a186fba),
	.w1(32'hbb1c0e46),
	.w2(32'hbba16ab5),
	.w3(32'h3b761f60),
	.w4(32'h3a2cb978),
	.w5(32'hbb712f5d),
	.w6(32'h3b28e0f7),
	.w7(32'hbadd01f4),
	.w8(32'hbbab6efe),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f4f3),
	.w1(32'h3b17acf6),
	.w2(32'h3b466234),
	.w3(32'h3b3ad040),
	.w4(32'h3b1ad952),
	.w5(32'hbb90dfa6),
	.w6(32'hbb1808d7),
	.w7(32'hbb90b7d5),
	.w8(32'hbc4bc2a2),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999f0fc),
	.w1(32'hba2e4559),
	.w2(32'hb9ba99f3),
	.w3(32'hbabb46de),
	.w4(32'hba39344d),
	.w5(32'h3a979dc2),
	.w6(32'hbb0f8b27),
	.w7(32'hbab25a3b),
	.w8(32'h3ab5993e),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab74dcc),
	.w1(32'hb9a8fb4b),
	.w2(32'h3a140689),
	.w3(32'h3b30010d),
	.w4(32'hbad397f7),
	.w5(32'hb91e5423),
	.w6(32'hba8dc16a),
	.w7(32'hbb5d588d),
	.w8(32'hbb2db0cc),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00ec8d),
	.w1(32'hb9d9543e),
	.w2(32'hb99fea46),
	.w3(32'hb9dc5fa7),
	.w4(32'hb9f25745),
	.w5(32'hba9842d5),
	.w6(32'hb9fb6a18),
	.w7(32'hba390cc6),
	.w8(32'hba2ffaa5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a138e80),
	.w1(32'h399b9dc3),
	.w2(32'hba2f76b6),
	.w3(32'h39ef7151),
	.w4(32'h3a26bae8),
	.w5(32'hba222c80),
	.w6(32'h3a551b76),
	.w7(32'h3a11a06b),
	.w8(32'hba3d32f2),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928c464),
	.w1(32'h39f1f0f4),
	.w2(32'h3a3fc681),
	.w3(32'h39adc78c),
	.w4(32'hb93b0685),
	.w5(32'h39aac6fe),
	.w6(32'hb96275f2),
	.w7(32'hba0db900),
	.w8(32'h3a8b6888),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19f634),
	.w1(32'hbab4f1f7),
	.w2(32'hbb889ea2),
	.w3(32'h3b6383f3),
	.w4(32'hba86a0d3),
	.w5(32'hbb0d86a3),
	.w6(32'h3b40fcf2),
	.w7(32'hbacec8f3),
	.w8(32'hbb7859bb),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90b23e),
	.w1(32'hba72e1f4),
	.w2(32'h39ac87d1),
	.w3(32'h39e5d7cc),
	.w4(32'h3a81d255),
	.w5(32'h3a71e6cf),
	.w6(32'hba32f8f0),
	.w7(32'h39f29ca3),
	.w8(32'h3af00b90),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f0c20),
	.w1(32'h3b01fde9),
	.w2(32'h3add8aed),
	.w3(32'h3a4b4bcd),
	.w4(32'h3a9cefcb),
	.w5(32'hb77f08f1),
	.w6(32'h3ade3427),
	.w7(32'h3ab2a4fe),
	.w8(32'hba17eb0f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3810bde8),
	.w1(32'hb9b7e9a0),
	.w2(32'h3ae3858b),
	.w3(32'h3a685141),
	.w4(32'h3948d439),
	.w5(32'h3aacd841),
	.w6(32'h3a330898),
	.w7(32'hb9b84614),
	.w8(32'hb5b2f3fa),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0cea4),
	.w1(32'hbbd5853b),
	.w2(32'hbc14d6c7),
	.w3(32'h3b09888e),
	.w4(32'h3a02cde9),
	.w5(32'hba7b6c68),
	.w6(32'h3a7eb5c4),
	.w7(32'h3b9a7a53),
	.w8(32'hbbd092b8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba014423),
	.w1(32'hbac578bc),
	.w2(32'hbb70e55f),
	.w3(32'h3909fada),
	.w4(32'h3ab9a1b9),
	.w5(32'h39e6c218),
	.w6(32'h3ab15dfb),
	.w7(32'h3b201910),
	.w8(32'h3bcefc08),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a939f),
	.w1(32'hbafaccbe),
	.w2(32'hbb54ff86),
	.w3(32'hba085ce6),
	.w4(32'hbaa0ef36),
	.w5(32'h39e6ee22),
	.w6(32'hb968418c),
	.w7(32'hba838012),
	.w8(32'h3ab55de6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c537784),
	.w1(32'h3c046187),
	.w2(32'h3a42d128),
	.w3(32'h3c1e664b),
	.w4(32'h3ac1ae5a),
	.w5(32'hbb7ae442),
	.w6(32'h3c18013d),
	.w7(32'hb758e2c0),
	.w8(32'hbc4d9225),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a8c7),
	.w1(32'hbba4e0da),
	.w2(32'h3be0c0be),
	.w3(32'h3aa2a05a),
	.w4(32'hbbeff504),
	.w5(32'h3b822493),
	.w6(32'hbb01b121),
	.w7(32'hbc42a951),
	.w8(32'hbb57ba0c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90b80b),
	.w1(32'hbad70068),
	.w2(32'hbb0b3b7c),
	.w3(32'h3a5934fa),
	.w4(32'hb7a47c54),
	.w5(32'hbb136e40),
	.w6(32'h3aa37ea0),
	.w7(32'hb910c72a),
	.w8(32'hbae69478),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba398028),
	.w1(32'hba60dc2f),
	.w2(32'hb9dd2210),
	.w3(32'hb94a0efb),
	.w4(32'h3a2e4be8),
	.w5(32'h39a6047c),
	.w6(32'hb9087b0f),
	.w7(32'h38fbc31f),
	.w8(32'hb94e8b42),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba111b90),
	.w1(32'hb9ac4a4c),
	.w2(32'h3a8e74cd),
	.w3(32'h3ab63a21),
	.w4(32'h3b0c926e),
	.w5(32'h3a0a1938),
	.w6(32'h3ac7a994),
	.w7(32'h3b310431),
	.w8(32'h3a364637),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd379f),
	.w1(32'h38985b23),
	.w2(32'h3a649ac5),
	.w3(32'h3a63dec9),
	.w4(32'h3acd665a),
	.w5(32'h3aa04c17),
	.w6(32'h3a9cca44),
	.w7(32'h3acc0e59),
	.w8(32'h3b05d180),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1b6cb),
	.w1(32'h3b0ead72),
	.w2(32'h3b24c47d),
	.w3(32'h3b25b1bb),
	.w4(32'h3b62ca57),
	.w5(32'hbaceb4f3),
	.w6(32'h3b28e1a9),
	.w7(32'h3b113b12),
	.w8(32'hbb9ef66a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad702c2),
	.w1(32'hbb5c484a),
	.w2(32'hbb94407f),
	.w3(32'h3a91cacb),
	.w4(32'hbb6cb30f),
	.w5(32'hbb692445),
	.w6(32'h391e4528),
	.w7(32'hbaff7059),
	.w8(32'hbb23cc93),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2d15b),
	.w1(32'h3ba961ff),
	.w2(32'h3b8375dd),
	.w3(32'hbb3929cf),
	.w4(32'h3b1e3414),
	.w5(32'h3b5d60ae),
	.w6(32'hbb957624),
	.w7(32'h38fcdfdb),
	.w8(32'h3b6ff8b4),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54faad),
	.w1(32'h3a42f3c6),
	.w2(32'h3997de90),
	.w3(32'h3a24a045),
	.w4(32'h3a5b6302),
	.w5(32'h3af7bae6),
	.w6(32'h3a4dc583),
	.w7(32'h3a27674e),
	.w8(32'h3a7b460f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b860086),
	.w1(32'hbb3f9db9),
	.w2(32'hbbc0f26b),
	.w3(32'h3b9552ea),
	.w4(32'hba8c1b47),
	.w5(32'hbba3cce7),
	.w6(32'h3b72d410),
	.w7(32'h39244a74),
	.w8(32'hbbcb856e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64b530),
	.w1(32'hbb463072),
	.w2(32'hbb6e1bdc),
	.w3(32'hbb235087),
	.w4(32'hb8d5cf16),
	.w5(32'hbb226c55),
	.w6(32'hbb405c5e),
	.w7(32'h3a2cc4c2),
	.w8(32'h3a5a2708),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c577b5),
	.w1(32'h39937c23),
	.w2(32'hb9f9189d),
	.w3(32'hb9b1b970),
	.w4(32'hb9637121),
	.w5(32'hb8b53a22),
	.w6(32'h399f2ac5),
	.w7(32'hba701053),
	.w8(32'h39f4a73c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3139d3),
	.w1(32'hba098332),
	.w2(32'hbb628632),
	.w3(32'hba612cd2),
	.w4(32'hbb2c922a),
	.w5(32'hbb00e212),
	.w6(32'h3621e0e0),
	.w7(32'hba9dd3c3),
	.w8(32'h3ae96629),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3795f1c8),
	.w1(32'h3964f795),
	.w2(32'h3a1189b0),
	.w3(32'h391828d8),
	.w4(32'h38e90f5a),
	.w5(32'hba552072),
	.w6(32'h3a41a0c3),
	.w7(32'h39b562d5),
	.w8(32'hb988d0f5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e5a3c0),
	.w1(32'hbabd1c47),
	.w2(32'hbb533de6),
	.w3(32'hba42ef4c),
	.w4(32'hbb107884),
	.w5(32'hbb62a3f3),
	.w6(32'hba7723da),
	.w7(32'hbb1a6d97),
	.w8(32'hbb48bbf8),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c1c5c),
	.w1(32'h3b80536b),
	.w2(32'h3bc3998e),
	.w3(32'hb9df8384),
	.w4(32'h37b477df),
	.w5(32'h3b82aa2a),
	.w6(32'hbba02454),
	.w7(32'hbbae6b7e),
	.w8(32'h3a3e4a4e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa898f3),
	.w1(32'h39ce7af2),
	.w2(32'hb9da58f1),
	.w3(32'hb9d3695d),
	.w4(32'h396b6c8a),
	.w5(32'hba76e4a1),
	.w6(32'hbb4dc81b),
	.w7(32'hbafc5807),
	.w8(32'hbab4e544),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952bccc),
	.w1(32'hbae01ac5),
	.w2(32'hbb491cfe),
	.w3(32'h3a1b4bba),
	.w4(32'hb96a5dd1),
	.w5(32'hbb130a55),
	.w6(32'h39c952fe),
	.w7(32'h39abcdd2),
	.w8(32'hba870e1b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f149ac),
	.w1(32'h3b101595),
	.w2(32'h3b577b86),
	.w3(32'hbab8f758),
	.w4(32'hba65519a),
	.w5(32'hb9c9bb3d),
	.w6(32'hbae2b0ff),
	.w7(32'hbb67d17f),
	.w8(32'hbb40e6e7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ec17e),
	.w1(32'h3a5da4c5),
	.w2(32'hb94c8081),
	.w3(32'h3b18dc0f),
	.w4(32'hba2d066f),
	.w5(32'h39b26a31),
	.w6(32'hb9b511b9),
	.w7(32'hbb8a0e3a),
	.w8(32'hbb1e8886),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4847f3),
	.w1(32'h3b419e28),
	.w2(32'h3b37c157),
	.w3(32'h39f45072),
	.w4(32'hba09d04e),
	.w5(32'hb939c927),
	.w6(32'hbaeee05c),
	.w7(32'hbb827999),
	.w8(32'hbb879b3a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906e39f),
	.w1(32'hb95f46a2),
	.w2(32'hba2f3cac),
	.w3(32'hb8c1e0b2),
	.w4(32'hba679183),
	.w5(32'hb9e3324a),
	.w6(32'h39e73e13),
	.w7(32'hb9e4bb63),
	.w8(32'hb9700930),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8383072),
	.w1(32'hba59121c),
	.w2(32'hba637b3d),
	.w3(32'hb9740f00),
	.w4(32'h38284b49),
	.w5(32'h3a9392f2),
	.w6(32'hb9c150c3),
	.w7(32'hb99232bd),
	.w8(32'h3ab78339),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75e3fb),
	.w1(32'hbb91375c),
	.w2(32'hbbedc17f),
	.w3(32'h3aa2ebee),
	.w4(32'hbb572166),
	.w5(32'hbc2ba4d5),
	.w6(32'h3b9cee15),
	.w7(32'h3ae3c312),
	.w8(32'hbb9cd075),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b42c2),
	.w1(32'h3bc5b5c3),
	.w2(32'h3ad8edd2),
	.w3(32'h3b1ee3d5),
	.w4(32'h3af5f684),
	.w5(32'hbb82a499),
	.w6(32'hbab8c650),
	.w7(32'hbabeb7cd),
	.w8(32'hbbd2e1a1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0af599),
	.w1(32'h3b9a1a33),
	.w2(32'h3b3accd2),
	.w3(32'h3a80d81e),
	.w4(32'h3b3636c6),
	.w5(32'h3ab11d91),
	.w6(32'hb9b4441f),
	.w7(32'h395a4990),
	.w8(32'hba7985ea),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9569b),
	.w1(32'hbbc14ff8),
	.w2(32'hbb149727),
	.w3(32'h3b226d75),
	.w4(32'h3b9cb038),
	.w5(32'h3b914f32),
	.w6(32'h399627db),
	.w7(32'hb8d4c24c),
	.w8(32'hbbc3c47a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bd262),
	.w1(32'h3a45e8b5),
	.w2(32'h3648c3bf),
	.w3(32'h3ab40ab2),
	.w4(32'h3adaed92),
	.w5(32'hbac10968),
	.w6(32'h3aa88f0f),
	.w7(32'h3a318573),
	.w8(32'hbb16dedb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a9afc),
	.w1(32'hbacfc91d),
	.w2(32'hbae4c049),
	.w3(32'hbabc6082),
	.w4(32'hbb2f58d5),
	.w5(32'hbb1b7473),
	.w6(32'hbadce1d3),
	.w7(32'hbb44d536),
	.w8(32'hbab5685d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88832be),
	.w1(32'hb9b2a050),
	.w2(32'hbb85a58c),
	.w3(32'h39fcfeb1),
	.w4(32'hbb5d920c),
	.w5(32'hbbebc190),
	.w6(32'h3b29eeaf),
	.w7(32'h3b9a06c4),
	.w8(32'h3ae0fdeb),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b848ee2),
	.w1(32'hbb07e969),
	.w2(32'hbbd27888),
	.w3(32'h3bbfe28b),
	.w4(32'hbb89f1f4),
	.w5(32'hbbe449df),
	.w6(32'h3be2ff4b),
	.w7(32'hb8a46132),
	.w8(32'hbc07e826),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4625b),
	.w1(32'hba95b4fa),
	.w2(32'hbb0c95e5),
	.w3(32'h3c120bdd),
	.w4(32'h3b9f25f3),
	.w5(32'h3786c11c),
	.w6(32'h3bf98176),
	.w7(32'h3bbcad11),
	.w8(32'h3ac19c37),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38464ba5),
	.w1(32'h3b60c951),
	.w2(32'h3bbb07e3),
	.w3(32'hbb4e505a),
	.w4(32'hbae2cd75),
	.w5(32'h3ac94180),
	.w6(32'hbba13ff4),
	.w7(32'hbb3db25c),
	.w8(32'h39217a17),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6ab2),
	.w1(32'h39a05274),
	.w2(32'h3bcd54b4),
	.w3(32'hbb7dbf7e),
	.w4(32'hbad1e6cb),
	.w5(32'h3b3afcdc),
	.w6(32'hbbf334b6),
	.w7(32'hbbc41c64),
	.w8(32'hba241f83),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb834c),
	.w1(32'hb98c425d),
	.w2(32'hba1561e4),
	.w3(32'hb9e08b02),
	.w4(32'hba2700ef),
	.w5(32'h3adb8222),
	.w6(32'h393e3b40),
	.w7(32'hb999237a),
	.w8(32'h3b20ab17),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5bfa2),
	.w1(32'h3adc5e76),
	.w2(32'h3a5b8558),
	.w3(32'h3a18b0f2),
	.w4(32'h3a1d7159),
	.w5(32'hba9cac31),
	.w6(32'h3a13f615),
	.w7(32'h39a36019),
	.w8(32'hba4b4512),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa6ebe),
	.w1(32'hba6235c9),
	.w2(32'hb91630d8),
	.w3(32'hbb102e41),
	.w4(32'hbb430fc1),
	.w5(32'h3a1ea5fc),
	.w6(32'hba24f213),
	.w7(32'hbae31a03),
	.w8(32'hb9273090),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d297a),
	.w1(32'hba75fc4b),
	.w2(32'hbacaeb40),
	.w3(32'h3aa98a75),
	.w4(32'hba003e96),
	.w5(32'hb9cecaac),
	.w6(32'hb92863a9),
	.w7(32'hba92f506),
	.w8(32'hb954c212),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11464f),
	.w1(32'hbad308c1),
	.w2(32'hbc0975ae),
	.w3(32'hbb6d4dda),
	.w4(32'hbbf850bf),
	.w5(32'hbc19cc35),
	.w6(32'hbb38fbe2),
	.w7(32'hbb8e5e8b),
	.w8(32'hbc054292),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66dcbc),
	.w1(32'h3c15147e),
	.w2(32'h3c113439),
	.w3(32'h3c172c02),
	.w4(32'h3b1e6bea),
	.w5(32'h3abe2988),
	.w6(32'h3c37fcaa),
	.w7(32'h3bb1ca76),
	.w8(32'hbb22ee37),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c113207),
	.w1(32'h3b0767ac),
	.w2(32'h3bc215f4),
	.w3(32'hbbad294e),
	.w4(32'h3b25c15e),
	.w5(32'hba862ed7),
	.w6(32'hbc70a564),
	.w7(32'h3bc1162a),
	.w8(32'h3b8db11a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b7436),
	.w1(32'hbbd15d9e),
	.w2(32'hbbe6ea39),
	.w3(32'hbbb0861d),
	.w4(32'hbbfef3ac),
	.w5(32'hbc06738b),
	.w6(32'h3b78ae13),
	.w7(32'hbbff114d),
	.w8(32'hbbb214bb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf80fd6),
	.w1(32'hbc7c5338),
	.w2(32'hbbe6122e),
	.w3(32'hbb20d35a),
	.w4(32'hbb8ab002),
	.w5(32'hbc7a0d27),
	.w6(32'h3b0e252e),
	.w7(32'h3b68dded),
	.w8(32'hbc91573a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc70dd2),
	.w1(32'hba774f1b),
	.w2(32'h378a74ed),
	.w3(32'h3b208235),
	.w4(32'h3b82bbd6),
	.w5(32'h3b8a14bc),
	.w6(32'h3b6163e2),
	.w7(32'h3be9750b),
	.w8(32'hbb172ce0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1be61c),
	.w1(32'hbbc0e5bd),
	.w2(32'h3a1b95f2),
	.w3(32'hbba3e74a),
	.w4(32'hba9c48a2),
	.w5(32'hbb4015d6),
	.w6(32'h3b05eff3),
	.w7(32'h3bbcd2c9),
	.w8(32'hbbb0f3a5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11de68),
	.w1(32'hbbc1b2b8),
	.w2(32'hbb3e00c7),
	.w3(32'hb96936b7),
	.w4(32'hbaf8df78),
	.w5(32'hbc7fcf58),
	.w6(32'hbb0c26d6),
	.w7(32'h3ba71161),
	.w8(32'hbada7cca),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98aa667),
	.w1(32'h39cd9efa),
	.w2(32'hbb5693a3),
	.w3(32'hbb1d65ae),
	.w4(32'hbbed1b29),
	.w5(32'hba792e5c),
	.w6(32'h3b883112),
	.w7(32'h3b652589),
	.w8(32'h3b2c7f5a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6b572),
	.w1(32'hbc3d5dca),
	.w2(32'h3b9f8ffa),
	.w3(32'hbc3a4f97),
	.w4(32'h3bcf3d8f),
	.w5(32'hbb3346ad),
	.w6(32'hbc3e3f9e),
	.w7(32'h3b1234ee),
	.w8(32'hbb7f0cb5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad0eb4),
	.w1(32'h3b933263),
	.w2(32'hbba8ea5e),
	.w3(32'h3b15211c),
	.w4(32'hbb8b9fd9),
	.w5(32'h3a078b8f),
	.w6(32'h3953bc8a),
	.w7(32'hbb46bea6),
	.w8(32'h39de1b0d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab806e9),
	.w1(32'hbb42c4cf),
	.w2(32'h389bc21c),
	.w3(32'h39428d92),
	.w4(32'h3abce898),
	.w5(32'hbbd5235d),
	.w6(32'hbb41a8fa),
	.w7(32'h3a886575),
	.w8(32'hbbd03a6e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2da1ff),
	.w1(32'hb949af56),
	.w2(32'h3b315665),
	.w3(32'hbc122b57),
	.w4(32'hbba5946d),
	.w5(32'h3be224ef),
	.w6(32'hbbfc3e85),
	.w7(32'hbb636c93),
	.w8(32'h3c1d92ef),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3ed75),
	.w1(32'h3a07aab5),
	.w2(32'h3bab6b36),
	.w3(32'hba543d0a),
	.w4(32'h3b8b8012),
	.w5(32'hb98d9c7e),
	.w6(32'hbc00bf8f),
	.w7(32'h3b2f3eca),
	.w8(32'hbc1d9594),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77417d),
	.w1(32'hbbafd5cd),
	.w2(32'hbbf84051),
	.w3(32'h3b3e4f6b),
	.w4(32'hbb4a03ac),
	.w5(32'hbb4247cc),
	.w6(32'h3b472f30),
	.w7(32'hbb82fbdb),
	.w8(32'h3b99fe0a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf7194),
	.w1(32'h3c250125),
	.w2(32'h3bb8bf4b),
	.w3(32'h3a35cf26),
	.w4(32'hbb1e125a),
	.w5(32'hb9ad1cb6),
	.w6(32'hb97c4799),
	.w7(32'hbba2c61b),
	.w8(32'hbc1ea3e1),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb00627),
	.w1(32'h3bfd1bed),
	.w2(32'h3bcfbb23),
	.w3(32'h3b22a722),
	.w4(32'h3bd97d74),
	.w5(32'h3a4bd226),
	.w6(32'h3c4fa746),
	.w7(32'h3b375985),
	.w8(32'h3baf635b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c852587),
	.w1(32'h3c1e34c1),
	.w2(32'hbbc237f0),
	.w3(32'h3b982268),
	.w4(32'hbaa4804a),
	.w5(32'h39dc1215),
	.w6(32'h3bf9503e),
	.w7(32'hba2bea0d),
	.w8(32'hba8ab6c3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e12aae),
	.w1(32'hbb6a6ff6),
	.w2(32'hbaa60f79),
	.w3(32'hbba36994),
	.w4(32'hba81d8f5),
	.w5(32'h3b50008e),
	.w6(32'hbb6f8ce4),
	.w7(32'hbb1f5f61),
	.w8(32'hbbc948b1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a2d17),
	.w1(32'hbc075441),
	.w2(32'h3ac199c6),
	.w3(32'hbad8760a),
	.w4(32'hbbc2942e),
	.w5(32'h3b9c54d9),
	.w6(32'h3a9385ba),
	.w7(32'hbb54f9ae),
	.w8(32'h3b37d34b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00d600),
	.w1(32'hbba25e15),
	.w2(32'hbb765ae0),
	.w3(32'hbb87ff32),
	.w4(32'hbbaf16c1),
	.w5(32'hbc577d24),
	.w6(32'hbad56ffd),
	.w7(32'hbb1b15c1),
	.w8(32'hbc52b794),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e7deb),
	.w1(32'h3b37bbe9),
	.w2(32'hba687444),
	.w3(32'h3bdcb053),
	.w4(32'h3b870223),
	.w5(32'hbb9d82f7),
	.w6(32'h3b981d04),
	.w7(32'h3b386b26),
	.w8(32'hbb9f585c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0091d0),
	.w1(32'hbc4cf3ef),
	.w2(32'hbb2954ff),
	.w3(32'hbbfe80ea),
	.w4(32'hbba68a77),
	.w5(32'hbbad1533),
	.w6(32'hbc1fb6c5),
	.w7(32'h3b331e35),
	.w8(32'hbc0c9e2c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dd735),
	.w1(32'h3b87c7ce),
	.w2(32'hbb60d045),
	.w3(32'hbacdde59),
	.w4(32'hbc0f29e2),
	.w5(32'hbc91be44),
	.w6(32'h3c2704f8),
	.w7(32'hbb091bef),
	.w8(32'hbc9c5af2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc310611),
	.w1(32'hbb8d6d5f),
	.w2(32'hbbbfc70e),
	.w3(32'hbc10a2bb),
	.w4(32'hbbaf50f8),
	.w5(32'hbb3dacad),
	.w6(32'hbbbb0bdf),
	.w7(32'hbbfaeb44),
	.w8(32'hbbd21d46),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc030a),
	.w1(32'h3a8482c3),
	.w2(32'hbb49259c),
	.w3(32'h3b4ba184),
	.w4(32'h37dd0cd0),
	.w5(32'hbc1d5413),
	.w6(32'h3b26ef7a),
	.w7(32'h3a8a46e2),
	.w8(32'hbc30b0f0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe37c5),
	.w1(32'hbb59aebb),
	.w2(32'hbb81e063),
	.w3(32'hbb139718),
	.w4(32'hbb7fb58a),
	.w5(32'hbc13ec04),
	.w6(32'hbba6bbe1),
	.w7(32'hbba896e1),
	.w8(32'hbbe02180),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62fd16),
	.w1(32'hbc89da78),
	.w2(32'hbc1b388c),
	.w3(32'hbb2ff52a),
	.w4(32'hba15a92a),
	.w5(32'h38b558d6),
	.w6(32'h3b84245f),
	.w7(32'hbc08738e),
	.w8(32'hbc1e012b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48ec35),
	.w1(32'hbae6a5ff),
	.w2(32'hbab82335),
	.w3(32'h3b2ea700),
	.w4(32'h3b9db660),
	.w5(32'h3b259870),
	.w6(32'hbb070e18),
	.w7(32'hb9876cd5),
	.w8(32'h3c9de5ae),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf27cdf),
	.w1(32'hba8bf371),
	.w2(32'h3beedc03),
	.w3(32'hbc2d1a65),
	.w4(32'h3af46d49),
	.w5(32'hbad86610),
	.w6(32'hbc43d864),
	.w7(32'h3b90dae1),
	.w8(32'h3bfc7a4b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule